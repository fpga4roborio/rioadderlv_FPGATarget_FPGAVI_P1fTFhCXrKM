`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
ddtXksX2+yylW5zu6QL2Lhnb2d1sD00763mmSITNX595NcHTEkwn0zB1Dry37fOW
FufOhVzEJp80NC5qZ/+F0Vk7Ik02dIR0elf3clrjeJRK85K4e3Hoo4xn7YbFUIms
l/8VZSb14+JVGURjfswrIyCUotIzlzVYZ6gzoZwDXIi5gQIBf/gI+KxNXPaKV+PQ
Ufys/12rjO6aI/pPlqSm0hCvftmBcnezN2hk1UeXgOIuKZnogjOsf0iJVX2aOOWE
6pD/psybjbnsNB6kH5uFTA5frkzIzkzl5d9+YDm9OyC+k84E83I/7/j+rk4L2dah
QJOvksSIzN867/4Qt8qYTQ==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="MvBXkzurAa5VTw+1JJ70nePUfoQXBvZOku/SMmg4TwQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
oRtzZL4VJ4iwysPsC8SXYCzXS8Fw2gtZTOskLcDV+1B9Nzn1zTyNtlo6lNICRmmK
ZRVu2BmCc2G+fmzynYlNTnSa7C0Cuel6FYpxCBlOuk3OF2tzAmLAuDyOH3Z1Yjzk
a0aHuoCdIRKv7BrZCdALt03JeUmXKPdOmIlkVGFl8yw=
`protect rights_digest_method = "sha256"
`protect end_toolblock="Jn9CQpRhJt4rnzZPRk+dOpzAubz7omckX1MrFd4p81o="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 22400 )
`protect data_block
gD6l00tciPUa6pDNTk/+t0OO0nC/UTtBwLB41d4inuAUA3i/ALrNyoJVcBnAmEQW
ptbcNp5fxEUJjnOxnedyZEuEBxWRieZFQnkRdF269oObrzpRPNh/F2Ut0wuRVj5L
s3Nsal7K6IYnBp069YNI7x5LWUJEBPkDtt1ZeyUN1xYXajl6CYKooesz38MofdCE
J92xTwib1J95LBvF8oHwmYa1yxmoCkPtX/u924tC9kRo5SUIN8Q/rihHyylHOmq1
GkdlCMlnfmQr7il46zdqr55SCUQHQOlBl2++FW1/FL8xoDsHPFFNEQDfv53Rq+3Q
dp5HAUwgu/VS0vQuSlty03LB0ky3vl6VIGGarwAcYs+riQT+7G7oE1W2eRVAYani
/Cpjn4msVBcBv3sgM4A0OnAHb80TiVyU5Gfruz/Z5E/Uy1nSUNuGLDSxxdSRlBb+
vnxdTsajUSOO79wuPN58XWIGeky5kjSQFHy1ryweEG75KF8NbeMAQuT5L/TyzRUP
SXx1eMNaFUqshHUDpZUQKPBhD4yJgTJI5VdFdoNJyD4quzNeTm2ppFLzJsgK7rGH
GbkkG7PP0NwKMBmTZcdxg8k5vWJvF56W8dsTF/AdA4ORoYj5TUi+tr4AvvCNlH2O
J7GNlRumQTBrbIo4AdzbRkoTL4CHEGcgMat8E8Zb57Osluiv196QiI//6AXd58vd
Imowj9oPSM7wL5OqgIlMXHrpFsJw6UPFY2pUPhwpS2OSIaGaev7f4zOmwlbgrB1/
WEbwG8l2cBp2NJXQieeOgiaqXsX7OWbdlVVItBrDvBYH/Euo23CD/wufogzyilrp
7sYshojxKxxGfGq64PU0eFM6c0BSxVn1kxYLPy1iu4ajwDz7WQtX8OKV1eSdk9Xc
Dw3FypUxxyzY8obHmTHBY/9MXLS4Vi5ZxUKcTQX81krlzsEaX9lhE8Zjcun2707l
zb6FeGWSZYsuCD9W/wZ5JdDwkQz+rDUmbepr4e9T500pnQrDObGsHW8kjwMg8r+w
IbZ4iKgofyDjuRReJBJFARo/ICF2XG/hFB3ile0UdlhrJ7Z3s/ESbZqIZCGuTmwx
qlbDoJlK2c39eEV7K0hLn8naO2uC9Ay9Biokwm5BqECxTMI3TKv1GDFMLPo0W23a
qmeRT7Xd824PGxGPE9NMIBoa/siB0/Fhh+r3EmP0UEVkr5TPVadzRh/5gP0S+wcj
3BvLv1Ojl76D42nSBkjcm0niy3trpKexzQd8EHLc7jQMulQ/DQOKNlFpTRAK0YdR
CsNWGEK7R3MIJfwONOwYSVA2bHZldSBFcX3l9/GSgyDVUi7T2jkow4MqntqN8twl
tfs04s2RQUINb8f1tl+ZfZ8uVZR1rf+NnJ+lw0hKnnhtDXDAKcDF2QlkMiDnAZNM
sxE+1yVheu4qYjRHb++opOiUj1CzSxXRTls1u40jq6kShQVT7acdEJOyq2EkRsO+
u/XPBtCt47cwRzkKT4HjiRic1OHXEEISp0TDv/EZLpH5EoeOCgoTG12XSJ4m2YJQ
TLOcmMD2kplqzw8tNeuvTZeHmzHClDQjVOF6zISYOur3Pq5Im9FPmOP8o2vXOraR
C2MrxNgoi0qLcubTEd2ga/ZYoIx+JlbrB2QuNi3XB0r6VrVJyDOXk1XO0nPHRk53
7hYcztug8wXD9bZjRozmN1wCSDlOEAzMADXytl+/oClCBPq8wv9RsWFKYJj2AZr2
pXfu0bIo420ZpSyynf4TNwqUOb1vsM4e6PMa1PiOJFP2WIy4X8LW3LEBMUS0CSdV
7dSYVHoIAR3N6zU7Apy66ddK6yEZGCI/yIC0cl3sWjIJmP+aT1wVg1yHIwh5PQ33
ty3Ks7g6hRlVUoSbOHnTggGJQzeteiCW7GUOJTUD0HgxKDwVaDs1pwFT2QsxQT8E
PYxaU/ImtFJ4Qi/ENomi8+VmH2DOmYVFento0g7QE24p0Nd5pU9OYAZEB9gT0Hdp
fgpVZmG28A7w9rOfDWT//Ic8neqc7mdlsZv2HImvCXM9UYyQjepBIqZ9d4ionAMF
ebVFs/XYz3vGuL5viBqXiDFOdH30lQO2IuL1FHqo7gyrzD/Tx/0xy7yT+moJwuLK
/lWovx1YQVY7jdFklJ6EGC5mRXhkb1vH7yX9edV3VozObmmyBMameH5/2frJv3bv
HZ58IJUBQBGGME+om/s5wpVGM+LNEu4gme3jS9bZoOupeoLtbk4AznfrPpZH/wC2
FZpiMK3msPntuGKK/OmqhmyxVHIKxuK9KG1t+Yktek9dOZJiUiNQ7BC5lxrhXWj0
WygUB7MkzDmoowjLlGyI81xhwq4fsKV9IGNzRr8pxN/SPbf56evUJY06ASisxOXm
5MHEVYPJi3j7WCiIu9RyaZHU3i0HgpPQuCUfvwLe3VO6DYonT8wsjMRxjM0mqAuw
xOPgt2Dq7gcpDxx+rTot3XURALXQpA47DDI6hAdfixULsopcaw4+BFNoW5FIqf5b
7Oxz6rXcsoxxBQ4Gn7QKV4/KMPl612OJEE+WWpY5anZK9xJLVAHtcRgDbQXoPHYf
8FyY5+3orea513v/TZGMB+JN8x/mdLXqjXC4rGO0BILbTPzahBcVJEntFc2rvUuY
7F14r6EbpHp+ZBkwCwdlEYOtl0vnyrE6YMFnUdJafuka5I0dluWcbWbcLepYhi27
r1+gXvD/0jfyz9MkdxICHr803LcUoDiuFr51bVi6kg2c6Cad9VI0vOPRtUGfeqhY
YKKa8rCEqWq09CyRudt2qbP2lEvurgjASZwXnkYfyrA9xUBrC7yfRK9FVgg9g08u
eoG5R+8p3tX/+q41hk/hpWpl9kbxWFJGgqFeSXUn2gI3/onLCuj3/76c5h34ySYV
Fm54HiCfxgoPY94sJ6uFs8guXrA+qPJIS2iqH5eYjXW7+gIifhADPAIdFspgzMnY
qsSO50CQCzNgvdEOGTjxCNLFH/+MXRBPHSnF5bk3f7w1lKl4R23Kv0FGGM2pE+Kw
C116/S867NR9dYKGxzE8pBpUgOcD0aHCceGbgHYWLClg8mjWdKcJY9NvBkXw0Got
6IQ7leQK1Q03FTWyafCSxxRMcTh7ZpzUNGnshXwDpbg/f17HzEUBaS+cOqqzz1Wq
92hSIgTLji/idFJ49Z1HJ/uvfGAWZ93IKAEn3yx8/my/WC3TDhsdtOBp6T6l0ZT4
+R/AqvCBqG8Hlos1rG1xnAyPpHWHoF4FStiCgUPpMsRONfWCX/wYhboDz6P7NBV4
mijUXh2icjsr42TCVhPKTfSnIgh7tQYjNkApfsNaUt7vvZDQwL1KXTTpNY4yvUC8
q/iA8wWUpCWGfKy3+Nai6BgwUmxvCLiETWe8ZG+bED7ARX1Dt7vod7p7s1JpYAw3
8nCW50gDC0oScxMIWlH5BQ6yJ71v5i9bhMtU1RFpEBFRBpvNx1x2sPtHmpJ/d7ox
iMXHnErkE9waH2Nj8anaJufcnnEnTe6uDr7EdCqHN76HYQ6vVdXs58cc4IfCeyQv
zHLJvIYXNnJtAwkWJBgwjB+M6Yigy+TW1JeJxAUthQJ12jCIQpJSHlpLXcFR7fzq
BXueQKc6Hl1Yzq+SNxv+Pv6xK9PNqnXQNMrRRbSM33C8MyL5zrB70Bz9nh6knMJh
/RQvcQ6toDZ/EXruiPTr1y9rdCHqDj0gewl+yKkFYVvVR4L10Kj7AYNAuTq7Lbos
fRQxzKhUwi0dY/SBJCosRd+8gByFjYgRuSfq8lI/WhKkC8XlpACUc//RoiZ6f22Y
iXtWZjKUfehpr8cIXl3cPU9ItUNMr45zFSVoIja4tdEXtFwq8lBo7SBTgvJgJ3J7
nlSO6b9Uo1BJQu3AfuxlpNGMD3h+nss1Ps4n9vaCt+2cOpdLvsLyicC8fwE07ftH
C8nh6fVAEAFjogC0D12xL1khZYVazTXUWl8EjWmItOB8Eg2SQ4jRqBXZYza0LJGC
XnCKZNibxuaM66u7d0EQO9SZpW6OXro4rnhFmyvMTyYFNU6soye/vxqOjg9KJOHF
57CmE6G/Pp1YZbPN5Z/OBLD+LEr64LApqYidJfW0oRbOWzPv7PBDL0F7aamY10IY
lsAsP6AlIDSUXiAAaRoxZpkGgMT1Nv1bEgSVgoFokdJYhXJOQsO7UWpFY+ggB+g6
DkqzKoo80ubNsnBfQf3zVcghNv8xhLc8yse/O5i0JOC2W6Tpt7pHP8VtIcrCBgFg
7D7xjob/cItXbWMh53IlMmoX+oXgezQvZDt3fqx9QaJY7NFPnDdNN9MmoJWwGZmJ
yimod56Qavjl+/hbqabiZqVERj/j/3s9328bdQZTENbkk8IV4RD4ef+ZZ2pN4etE
8J9dcEAK3lMvhjharew+FrpZXrAgQ9cWr9VDhAF0rMX4Dm6tNotYWorUlF3T+vec
7Q+XGEP9xe0EjQF8rfPI4eK3wE14nWl/Kq7/dYvTQGs7I/CjJB4KQonaAkbweMTj
QFnzufjMcuJHL51j/rhbU6lWtdre2kfMO4YJujT+HSl78YZIZZJeTcfL9blLwc+J
mzshVt2t/eXa2SenyEFIyVBq5gjxZGAee2xCfoimb7QLUQjg/7W2Du2zmdD2V0ol
kQWkUSJJJw8EJcaxO/EafNRVOVTY6lWaypmwcFahctoaIPP1Yfy5OwqtXhUyz9XK
VvhWaQv7MQd64hl0SjbamaQ+AVuC4XVy6grvgCz7j89aE90lvt30cItVN3nKNMyX
ycw9uUft+wXVmVdjKdBIcosEMpWybTq7rUHUUCDvTu4KwVN4RYxOyz4tnVLUhRcY
OV6FE2thtnS5sK4xrJuwTQJOeo9ANwVNgICMk4eP9OWiu7ps6xp0ypZzV41kNJTe
rmxlMUu8zoh7GsdO+MhASyK88zvC2pKpKz7Pid9WDZlDm1hkv9ifnwqZAJmDkuAv
C93W3hZDy5VPYQmAhRlnL23qYXKcv6HyQo2WlonBe3KFmi9lhglMX2JqZOZaTnY6
bDCdzK4uPPXbO/6DOXF2K/eltWb6KqiS2+/PP2t011f6r2J8NpDnoFzwTme6bJ1U
1fHuqSlK8dfYj2TNPwbM8R/iapA+NjwucrpEKg6U1YDd5p6xhvvULzDMfkUiLSVw
E9zXFwa802SoW2VLCMqwsviDO8dPwEhMmpDl80eM52+UwZFQ8+UEm6MDIYT6Qwsm
dF65NjA5Dvcsqq5KPrO1mxuUtKIYwBTisiRVyi/zIm8SsCJpHe5m9vDzcZOiHjef
VYFrfoIjXeFkMePshM8Konl4XprLL+O7Pv6qMuxDVBacAPe59MNPj+IvGOvGHTaN
D9tRvAO/jWVoLTaLqH3OqOBc4xBWslZoHMeHe93NU1XMGAfK8DE9bQBQPwiRDv7G
tzUmARjJoM4FGHkZyDNbJ66JaonW8eBmC2Rtp6j+P7m86ygYIpp9m9XVO5BjlSFA
Bv+rPXgYEcZvou3GESmct6MuFFYiukiJd27w5S36Z5UkCn2lZM9ld2DOmYC0ygWZ
qQSREjzIEFONDs18hl3miq4F1vxnY00LOPyAX9NAfF9baQQ57ktv7lMGhDxdSVMG
XGM1KBCQXgFR+jITUNVq0wISL6SI90hnYXn8pCCdGGz4banZi8bHljle0ZKdybVR
1zdjEmCU8VzLRGi0m2dK1iB1FQCDGVASJTbjQ1ssPz2IWJtdxkQOCg+QOBnTHbT/
wrhBTOtqN2iocHY8jv6PHUPHUwwicU5As35NMRcwhsLPO23g5gUjCmcNNJHVvox5
4xF3mpXI7zt5D0HwYYMNg5ybu7cD7a3iv1AvacJTKVhVCK5nGt6NNkNtQ6iebfFb
Kcex0NlKN1MBp7rpFQsA3Sy9izM6y5YWd44ZuDa8ARBP1oz652MY4tBzNC1v4+Vp
iAJEjZHsdD+SPwIvKFeInDA1X0Hs4VnxrbozMV6eXjw1Ypk1Qui5dhWYCyYbMG0A
DPNZsVAG8wwbjSRTwpa3WDGDLtbDw899BGhfW3fs8G3c/T3Tj3tvqKd7u31ZPRe9
r94fHHR+Xb1WTs0I8xTmzC7MJtgVBYQx4CjPbLvOpJRqQmiqVPQXDK9OQRC77Ara
osbuOBhdgyCifApw5Jh2mqwbFy5aHtUtJzNrjyK1px5mU+drCAdmfeSB1H+M/lhq
L0uO0J0sdQrV+oVwLeCUKXcH/Ru7/F0q58SCPMDh8N+WX+JXyGGOPtKCKLs2c1cL
7Rk59Zxi0SIHyBSwQH+NC8Qo79HHLPFIK9HUhvZxO9Wl8WkASUg8jlwcnUVvEOSK
uQxMkxXzKeDOlhZrKmZekbWC+N3e6A3HLiM3LGMbLo6D2lJuek92oMCyHvMLJ3ed
aXSE1JewS4q7X3v04MMnIM+/mY1RAkXjXEqct+fdFmN/p7IL6GX0/c0L6898UnAI
HLPKyHHSuPsOgESLebEjnKpOtRlU5vvZ0l8JGTuojn9fpWdAYNCsr+sSIgMel1MQ
Ydz8265VWPdIFqT2czTnufAXx2uqvYV3v8KBDT0kOCM5W5Xbso0bGnEIWBDzjQUB
PPSk4XOVtNVxpET/td/1/aboktPmdHGJH9MFEIn5k5FIlPp1gfEgFZcADWxkWFI1
VQcJ6K1o8ygFQIBsnu6R8t3iFgJOtQyVadtOqEvvh3FEmoVz0zZvp3WzpP2Jegfm
gPQWGenbtclmWTdTLXiUcUXTpezCNTuiRc+HeJ/VUGHKzE2L13CCPP7zSdroyVRt
Tb/9bByDsG+SbLccknqUgShRVD8s8RhEsZkdvli9IkrMEwuti3j/28osrisGmfB6
bksf0bFkTFpHcCZbB3SCkHl1h1HVi315ObNZterZZN4kI1ZRvyddHjLtdky/veIO
NSecSEATIZ1Ka8q7pYmwKSo6xsDriAqeB/gX/8aW5Z0v+L1BUhhndQs4NfkEKC1F
gQApvMKggBVUcOuruQ1guJF25m37d42ArvKVO7KJAkGqJKH3ZOoN+QtbsY7TWaKh
S7QVTv7cNsoQbapanatrm8Dw0X7zP47g//KqMaHGmR6yvzRa6kmfoU58jMtFHsCG
f3wCSvSP9hek0daz2oFF3QnnkfVCBm/Q8JGt/HjVCPoY6XEt3+npzJoJUHfkP+84
iucGB8iLJc2L+6HCt/17fSWBiYMrdDtFYpYp+gMqfyBa/gpLhIoFZYNIAt2TC4+a
Kb66+mm01buDtN8FFd5D7isPhi1gl34Y9yD9t4re8lT1hkBTMJU8NHYHz/EYOYm8
DP/WyFgMYdtMZMspIZdMoHH3RsuJEhKOEyrj+RbIle/cO/S8VynNZAqDX9j7Xscs
77Z/NXYSGBYQ0r95ivLYoYeFPUqepWj+kuMZPPmwfm/MA2ju4cdlyA2SvqPJ90JK
3wwEBtWd/G+SLYQqJeGcum7zn5VUxT+fdGzTVVjNVpD9QvfcoVqY3eXN0U9HNWI4
rMd3RV1Hn9ehs5NAzg5nLXRlUik/Ibw/ytWrbAUZkMI2d0tRgvpjXu70MtuwshFq
vxe1QOIHsMnJ8baoFbL/fR1V3t5v4ztLTQYSREjI44ucroudQmasY2SU1iO1GzON
BNYucDmcflow2x6cpIf6rdEAs2Fk8G//HzDNg8V9OB1vCT1z1nguy5axexvkBxhU
/MnjGNQDsZMjgeJlzL32CaOuTYFMoWSaCD9sC1t7PBJ+hsGGZX2SZoaHFX9oMwfa
XRFnEf25Arbh1riyAtDz4seb7KysLIqrKhyu5z1mpvkg35sU/YWk43jjAGBgY/u2
zoU1WiykRGPG54LpoB0H91kNMcKdZFB8M5Oais7B/AbJsKauMZ5DT0AODw2Mwho0
s3seZGCdQJNaGRj8RVX60cY0FO9NdZWkirSiC/S30FBHhWzBJPGnCsr7Yip2mZY4
rgPQ4pZdAUMYmWpeugJ1y2O6cIdetXRr1vquA/2kPefnxHejAzq6yFQd9u5bzVLV
iki1dLw7bNrCgYoy8U0UqjNoCuuP6SwnQ6Qt5r/BqQ5R1GPjXlvpieEBQxdhW3LW
gd332DxtI6Uvaqud/Tv6BXmbxg3cKbZuW2Z3H/m+JravtI9fIARPqd9fWsQYQ4Uw
Nd5p3Am7rxWFt0cLqlAIb5nAbHaQ7swTzTxa1hbzorBO4vL4qrKoaMq3T38Uo5C3
jwXruYjlcuNBA/ImlMMKfFqv3XDFPahoXCRei9M4NuwpQJzZ0xJS1HGjoNwBDR/p
9qlcSc2sOZ8fJ7mfpar73K6WWQ77k6ZtrVS/W7NHaLubkdNOEXAOFhC552O1uhYy
qlynzA+93LnkERxb5dm7fN8Ytgl9ORwzKmpJGcdAFqTnMEmsQRrhgLxxVgXiRUAy
B5UjQ/6GixWe+fYywk2jE3KY/OUQy5d9lXcOnZYyegvFvSV86kebSMqNBSN6rWQJ
CTgIyKpgKHQBhU4oeXpuA6gYC/jCWaynVA6Lgttp5G1+fu2KSNdidvj/qrCnB5qk
hnt50Cx1r8phHwA9PsuMVp0wOgcSOoKUslkZLicibAjp38qaXCVFTKZtM3U2ebwW
3S0Kcb+k36aFg+I1I7uVlImZNuYJjkB3ZfhEw3cR5MXnFxZvK0H8Uof09CLsq+Rx
OsqF/XWVYLtJql3kP98gcd+i6rLaz2G2t3V/7uvq8twdKnqicKM4TLyVK6Jm7vrs
jwQ6x4o5+3Mjy+QxxTDrBMSj7RfbFhsTh4Xi5P5leNvYIyPPJxFFcfxJIKkgxlmG
lld9fVPJ6OEWNpV+kKUCoMTKdDJEnKk5hlD9JWztvLf4SymXtBRMrWv7sjUHh4Jg
mTDDR5L4gn4kHI5gQjDAHkKqzQLOf3AMGyOllyc6ftbVJIV35VcgKnvR6+vpRlYE
fFXqda7vPz8CGc0Ee99jK5qXcJTZPsX7Lk44HCxLqDB3X9fC89jAlbRu3LD1BkM5
a5YNC7PRHlpfCCnqgzEfEPZ2YJS+55I7gfdxBJ0rp4B40FLb8MWyMt4Uok7Q7ltW
CeuAFANzK7EGHlSxu3wW9DBggtVDwqdLN7oPggJ2Okioxc4mabL4W3+jrK1wVEgs
k/5F0eLjLGUZ7YRuriKbZ6yx38+LPnKdh6WZT296wvluGPxa1y5PFtR23FjqU/wa
FhImVppZG2TnTVgkT8nBuz5IXbELh2UX7ww0I1D0Y+2CznH1QbZ50jaCAkV/rBs8
IVyk+Apex9cbNIHoc69Qjz/QZTSLbYudd8t87sNiYO6u8wYdKNPjf0HHpXor1PeN
C86kNbHbnewXOMlcOsml/IrJra0y/Eze3na8UhK+Ds1oozEF2vgfVFfZ2E5wt5c8
KKtFPvc7HknEAIrw3HXsjfpv0JDpbv5z6695BpJGuttjQ5D0FrClIbg9hDYaKAdv
LCll1QzHBp+SK1Wd3J+Jvid62eSZDRW9wCbZ6KR+/aXtBGqLmKdrUjVrUtJSXzD8
nNxC2aZNFn5aa5GWxBQNeV/0RL6jx3fEdgD3ANG+FWw9pD04u85XpIEXhOjjINFu
v39xM9+SuE3f8Cn6BZv4HkBsav6yCdxyUTdmF2N3yrm+RLdsOVk7qTvgmvzVXB9F
FpuAZ14KANtu/gcJk68GX1m8l2eIQoMLAmUuqQrqLlJAxXy3c9NLmTMJsvryEjqX
PflWdHXUHZqro1IQ5BPpOEjzyOdx8/ftfTpLhfH3PeGYhrUg6j6trh7CNDe5netk
KHWWNJPiBYWCytl5+qFEVO9SZddnvQbnNzhbU3uGc51PgNX+GOgnJ2Nvp0zMuJTZ
i9HyEN7tRtLrFbs0fkX1j8w+Y8LH/YBeUBiGg6Tqas0/yL+kLcIrfpRYAkLWuKnn
YY/po1FGTawLgClKRsmXs11zKgBnRvJmcRiPNVMJwETqm8hK/l5mmOC7iRWIk4uj
aUKykFonJl5m87AcuhqUG21U6CtJkfvuBf5eNAeL8YcGTZfbImlmky1ECiXTrFj4
WwNbONhB4/NIX1rkWGSfkd8lkSybhDU76wPo8HYZT5L+K/rBdQCnrxAXCOgDNfQQ
gLTYV0Z6A3Q632If3INZRUKeiLmP/nw5x8ydDWR+X9BevzsYCc7xX4evE2omrPIh
wClAvlBoEqu+5RR+/cFzy0bll7HpDJoi9hl4nkDqsNGo8/5UBGd+lk8q6bMJUQAq
ZaebyAnHQU/zsVZGxeuLJmGQp6I92q2U9zeDrXj+idcg+g7OvWHmIrRfFZuf0FFo
157uNnmF1dpFDIfltmkHWcnSeTc0jEncGqYmTMKBdQMRUSIK62d860SkhU4BbyOH
TotQ4OPROaHCcwg2stTv9przeshptMIsa9eZMjhg709scfhR3d/9NGuIvDn/j8il
22hDjgcvW2J6dgBtydTwrwFNXKTJ4DUX4Cgu8MW5Q02vuyT1/tHz0FVsRPS/ziao
Y2goCtEuyZmXEpJYgPAXCciVGA3MPAp4/OlA+YYRWbp9Vujov1/3gVBwjJPVsrUL
iKtxwC/9M+9loi1IT4xXOK46NnJEEJv0kxYvU+di9cIz0u6q1vlzEEhNOEAbZa/1
n1NwSGyQDIVoc6MjxSD1B74JN08JXg61zZ8w8TTfqCgvwhjKKwprvk7FCU+WDZR7
Y6V9CjaRN5lS6KMI08DRrjHWXL17EejndAzRgo1XFreTLCvCVDO3VEuKtdnOCYJs
rOLZ9Yd2zkUtf9yZLf6KFokP+mRQ/qcmMGCz0G5qZ8caHvd/W3xqy5BcljwNa8G3
Er1NDdb/eRIGS5z4a/STLnt9CYbgV2z337uAeA9ZpUoGSv6I6n6YQLeWYuA23od/
2dHs+zh0TgAyjCHpTns9oXDGANnQtfbnFkqPBRb4+mAPlA7UkO0MM+udNknoIUu5
gM2HhMtsjUvpAxwtfduMC7qtliD3p6FxC1ilZ5xqdRRPLM5IQD8ngl2/1JiUVJV0
MvUMudXN9bJzU7BCpj1+odgz4DMbAu6w5OTdXPexyX55d/xp7ozMuqQcbBRHXmfh
87btoD+xfiHhN7YCULk6jxWPZa8XEyNwFruhWxSxIXBkC+w8FdH9nk2lHHDYq1oV
b6eWKAv6HHzRmp6FUj2ymQjUoprDQnH9NgY67kodsU39mQzW+FQiCm7r4nHIVdqE
pR4/4RM2PFs/Kxnjel+yHITi7ipGbL5PDZkkmAalmBLXWtuZrAREb6bQ3ReVPp3J
BLOB5vHZ8sl7zhVIHWyFBO8OemfTrx7+Bu7eS5atOuXcxYYFD39xjVu9TDVSGCC0
nxTkej+YS+tS3w9vwMdP0KoxlYsNpZiB0fDcbID7dum16tLpYG5WwHMMfvl66Whi
IBwyuSuSOPnzeZAElYSmt9den10Ox/c4MYFkFNY6vMgxocejNZ7JMLxK11Q8PTgR
kV/8ea7Gd4zJjY685iHsXICdMx0v6aI2J8/UaGVAYi4+WBCpRhyZQXOm6zzdjrXS
+4XCOhqgk12LVx4AB8Ms1ZuetEN2HeBha0PjlhYZyNMRf9eNQyxR8FdL8pbBxOtT
EJk5NsWUmcCnrBDd/S2VXvsnL0AhGj/UdYCxl3IfCInhwbeDLlsBKgpP0UbpQ++m
d1K1LW5Rp1xt4+ty7PvgY1ewzM72mezYE1XWwsJnVK3Nncwg1Vpy2pUsHJGzKqrt
Wa5bxE3BLVQeROMJfaGPJKgBG8/WmVxFHEB8FqVTMrIMLF2d9Zgvw26yQU6o38I7
zL4DoAUJKZp3ykCL7C1dVVlCwcMX6SiDJPxKQfjC8pPdOU8iGCjzH0ykVl0wC7YY
1km5LFrtMOkRi3nRQC2SVV0ieKAmy/NA4aULdFxMgTDs4u+pRnyfe2bNE1jAymaO
bxjL0bZSTCU2Y63TWqPzgH69AudTFM1ibFkmS8/r3sC08CM5yS9CW1OMCyf+hO5j
djSpCNzMye26WBpHQza+8+Ah8sotzDYbZ3wgRv7iDqada6W4hEYfHR6ynUto24cs
bRp7HISdOGdWDy8nZQKqxxNKTy4osiI2AlOdp78KyYvveJQLmRsA4NWAklK66l66
lb/9ZfBioTFOEps1+dTEcz44iAv+kIL4Kf786NJm86di5cZYJZ5VE8dMcqp1ZEIL
kVQyyQ+MAjDkllP3zlWoJ2pX1Ie1bPt6uPQyCL9kqFPZBuPH6lbHwfcbj4BrHwK2
/MeWBZbPSxl8kWcHKx5+ck+77OB63HutMZIE1IXxdwcDCRuMnowxlyTuwKzTszaY
TA+k9VtKdkVWyvmgNa7cJYwmwP0M0QvfD4ybPs4aajyNFifaCpq5MNImlKvA33m2
zD65PDAI8uGK0Y/M5CM7T2girnl6kN4O6am8yJQCO7uTMVCfCZfywitjgW1L0qPD
r79+oGps28T4J+FGh54oHfZkk16nUs69FfdIq9JyYrhOBHx7EclEmHgphFypwofb
9IQKbl6VWivUrmbi/RY2J+dJOAqz0eQAa+S3tKd9kvsF5EqKYfhwtJEH+1jJoSc1
jl5zqKmKlrudru8wqAMPXLWysjnhdmcdB9w6BPYDvAP9/ASGYMFH0OGUDwWoT1xi
NvJfCNlxbJxBfE35C46T2HlSkfMoaJM8D7aDrXYeki72XbZV8a8+p5Pvb90TLUR1
dXsLOcyZU5SGcqRsOf6PCEelzkbKjGAbaiTRqwCd/QMUWkUzbqeBVzjdxgyXfyO1
7rgGpxwKtNz1lRxE09D/8mDw1qFnm7eDrQqw+fMwwdDPDIK6oOUpE2HdgW+BC+/I
fl39vN+Q6UfyziiPrquTMWQhMOuO+cKImHP/C4gmhbBhR1oRd9G1mW/B9Dw9zq9v
coDnUgAZxjU6Y0z3E9gUS9JmEJmAmK8B8kPKEw1WCnmIkZk7iCeYn9SGJM52wnwf
lw1XPQN94nDwXf61SYGd0/29+punwdFiRM48zJPlKqltxhBCaKohXa9Ccr/r8YBJ
bDAZfor5pCjudQwvIs4s6KmX9g0gheYF75+qea54EO0+GJrk/3v3P5UOWYRjClsM
P0aed+wzZzBSdhbtA78MDLxgKduaa49R101cXG0hElnfd51d7uTfJ/BRwVSeaFR7
F5XYcH870WC2cJqAMITJK19suGZqtw74XwmOqjlDSv2SkFDyCdcrreayXyYrZqjs
GYxLdWOwAyaowjNATibac25vkBq+DTRKCyod2bmjlDJmiWgvVKFiTDo8NbDnfCGC
IVjpWQJYPHwZUykau2m0emId7j8nVxhdskzn14sFp/EvPbrd/lfjLUylVcNL890h
NRaXkZOIzMdIVS5kL3Xvk3nmHHVi0LBciVL3EhNOLbgb7A1AIYPoNTqZvp4yStmU
MyrLzdnOOB7j9Mgt1Cu4lOFwAb1ZbQAZMCT95L3PGLWfKVN9QpHzcLrTuHoe3vJN
puwYBcQQBGzvnE+bAkwxv+YjcaozRWOrAoDpmeMM2Tb/BPwv1EeQJwXmVTv4cfA5
kgPPRiRXhJX7oVV/YU7+wk6bjjWRUuxeGhsZdVBlv4eQlHa8nAEA3ViWaFZdvWb1
jBrQfaytC969KMfSNZ29+n2EUEkMUrfDn7KFGmx+t1mFXS9c2KYzfBcQfualcBEN
yOk0A+QFqQLUl/AQiw9yEhfTUVK4GSEQCLp0IQLze+DP20i09+gy/k8eAUSWQrBe
XwizrJYnPxtx8GVgYFG7sY0VK2zf0mJVC0ZMqUpGW3PSQ4S96SJYIjVj1Xh5zFQS
I6ov3ZUdqNpaVlWA1HRVv+g/bQbEDkP8vbfLTRJOs895xpeB7RCew5mghb4fMqe4
2eYuGpi9biG1cD4FZAbl0qFUxrBruOjn7hXLw1I5pNpWTiHe0VuYIqk3tfLZg3o2
vqlWiBeLWXNdSjKzPABkdi7VyUenxolwdZ/wY+wmbKfnEEpEeEHD0SJ4yjeywrjQ
MhQtRqvKOesWP+TaAPXIfnlH7KxDINR4/PagVule++REB+Vfx4CWNAsBMo4GZl+O
ckkt1gsJsETCRVh2KN+pKiDGgR2njd+PCjUv21U3xDjMtrdKKZm+GK7o4hq/zmKp
qmMVfENPHYyyq7hARBkr5Tlxh2CG3lFcRAVhPcVVVUJe2mMDXgTHCjIC7xQjcut/
fXqxuvqVCvLte+5WuuRtLvgLlGGFgKvtDAkJdtUh7TbOt6EhO1uTGZGXbuL8S9Lv
E7tSveKIZ7vhHtueA65O4D4r40Z2qTUh3N7KFmUmykUN5vR5qj7SDNavceOwqWEp
KdujWoPJiCqTV7a5m3GaXSiWNdhnV5l6iJ/Eibw/NW0nPT/mTMMO6lwtc+am0MKy
yuqsu6bUq0Qfuamla3s/cg5a0upOblBMlMRX/h6XinZKTaiUdydPVRDysbZhIXQ4
ZtHgurRNDeYi0kc8YhRYQAFetHj4Lk5tHhHmCUXj1ocjmqxQQ8jYb6i/3MGSHjY7
YmTAIzQz/UH6/pBgO4N704UGS8Noe5QumsKx4X8U4XhBiOkdsjoTsIT9Jss1Riuy
Clwyj1mnvpWrlWTh8bbNllHVMAvaeTklZCblF4ITLMcmO0MOglHG9dzurnY59Qgc
i7HFyGB14B3bpmia4b1Er0YsO0TU2cuDewQZTLjBaULtIfz3RuXTa2bKO+BIgLDx
QKu+hI++ZT/mBvYwmeEmeJnrn9u/vZpzs3Zod/5tu4drV9RoJZGTtk1O+8WrKKk4
3/lzHmI23xCgbzWgizU96RN26Rp+pWuSccr7JmWB7b76TfldodyZmnS0Pc1zJh0P
4rGJjLuoRryomY2DQ24eM7FD+ILPFG4VX/0VnK03DpbB/CuOGjXlnLo7pPuAcEhV
LBOSt8KK//t+o2BzO0mp7/+HaJiWge4U3Bm+IlYUFl1/FETeZpBlRMnpp3UWPfMn
hUVBy4EJIsUjUkn80LRPFgBKR2b3OkMzHFbrgYfnFSowL7PL3X/BIVOQME/RT11n
m9hKP6vaLu5iajXRSrYFQXqOZTF2+C6N5/+DU4X7bjabHP4ahm3aO7Oy8GyRspL4
WnkI+t3g8oEOGOlAlJ29NQQ6pDestsBcaE4bHcKIJLHavWsaewdoJDGtqa4CFu0g
d6qKxwJcvl3U4hMiWxiTMR3jeVH2ENELm6SP7YTz19R7fxDCbSSncpVrXC7ppIZ1
SerPSrhr5YuZTrg9rrfYn3cAkb4ZotWpiwzz0DJFMM5bKJCMljh06dUxRdDlovIb
ex8R/YOe4gEok+6GyKgI615C2MdRAkHrGleE5Za4KxoGhU+hlj82/4PK+BX2Ppgg
G6mOkYgmeW6SZhQwrlMBXazlIfKgGA22nj1afxdlVPz47FnjwOePhjgn1RM0sQZk
ner+AtfFBZbMM/ng5zmJJGQNG0NSSLG03MzmxD2oCNCHd4V/ftz6UmF+TvJQl6m+
XGlnRolxS2o7Sw9xJdBilGIERwsm9jZ1WMOB60mp1UWxAIwbcYY4EjLtRmwyjrV4
gX6WAaAcXnT+Cm9/CqDmfl8EUH2XuXmZTg5emeJob18oxwi/qJZORiA0eYURm7hA
FLb425IwwE7FxZI4Q2MnETzGEBua3DGxPBgRh78jPedC0fWUg36qtEoevCjq9C/J
3MBP8mypzo0V2+fSy0qWUgrwvduq5w3H+nymo7FLJBapgK1gu56hCbdWg0to/4Sk
ZkODdMKmFMmiTydWdp5eJXVN31nSF3VRwZl6Xe0hWUl1x+/r6RBho+ZiWOKLWJC8
qrNoDkmKReD0/SWX3g9qQp59RSms9DC02Oav4ja/hUMdJk7Coe5Nr+n/h7Cx6sxU
KscBxLL/4HIiIurovWs09d6AIhHuXVMbvF8FMNJ5isBTWCdunY+qp2syHBEQ9+2y
yOPH/tNvvWlfY/FRK7hvbkLyavpV9LpdH8FhuI3OgnSp4mf5DaM2KN/b808nluaM
AoUxoqQihdtboWS6xm2CmKvKw5BkbKpp9TkvxWdap6ej7qkOpJFZNd4y3lYQ3s+i
YbqgZZtf3MDBUZuxhkEJiQvahKAFPgbvBsLpVu/JIP1vfekuQaMymc5BoNmgpqLq
hgWCAzLN4QyFfrCRNopGIQYapOLP8oW4MMmJoC/HMMcnl3ryrohh3MLgLn3W66c8
pay8jGbVYoVRhiq2hkUw50nUnkEQ1IPPWMiE/83TEE0EYgwTg5nwOKdcn5ghokBe
Zi/ZqGgO8pJLuMe05tQsp16BFEZewjIlVqo1xwnkjam83LnPNbXlOR1lAM9Jwe0o
cMplG01EguYfiALrVAQg9hvASLXbVAdIYPYPBQ3tA+MTYAfPc560HVWv5xfinRCy
RINDtlKOUdI3tOFjXxc6TsLb9eyRKUikzrdhDfhWpe4hH3B3gradpftyAbJUExu1
w5gwQ9vevpgCMyjc9f4WCY+Je+u/wMs7/og1+T4uKmJrZ7JH8luk+j9aOrwVlPOl
GPTC2OKnoZZ72AOtsmI8479ZU3hLuMabxoJ+BPcY/LKbWn08iXkBLthlK89tqdXR
OMTbXG1x1vh6GMF7rpjkn0nUJkQegZj/8eScBhMxpbkWQjhA8DcDF52xQRIX8Qu/
bJ0hPu4x/LT4PvVGa7xlX9gL+ju50LzRkzhYOjhZ3ha0Zgpn09JqEJNxYa6ezzuF
8VG1iA7Hb0vIakI0zzRozSZIF9qMzO5MAVzKCBxofxz2akeF9XY3ltMitE5d941w
2UXeVQmeCdTpbHwH7bw9b7Rm7kvhiUs/I/ivFOllqVNoIEAl6SVSTPiO/4X/QhME
GZ/EaxQJbvI3OPwIv9BLVO6scDuGA5qD77f9a2yHHMwcLM5UdM8PgTt4vEr/+uAo
G+dl6OtodO8arC2iFUCDAH1YvxdpRcF5+slKr9pe4hC7/i4u4jf1zS6miY+TdoHs
ADqG3rtUDMHv/xPJY0DKMlCTAZT5I4+ulkkMYZijh7e/20gy5lh2pTICPh81EsfI
HApojzmT5XOGq9k1iKUvSX9VE4Xvi/LA0rrUSSjp+UjX61eX6uzCarEHLNv+6UK1
RKs4HOkWerUQ87iTN+xY05u8edkVJHYNwjhYZs3+7mNV8kWVe/yELZCA1G791Lp5
PGBCdhKaf95ANPyFz0sVCg2OibThMRq6RJxjwKOplam0/CnQzFOC6Fx5yIrog552
xhDU9m2NZIZXrSOXYHBN4UxB25jXDagd/HAqGYmPbaC826QTcm3VV8LUfWnrtfUb
Gl3+Uqyj3BE5Ea2A8FgF10Ix9+Ke6CwWluneljpUNJatKgbB1tlXiTiutLn3xguL
rqWC/0/mOBsYxVc5nTF+FA8qsGPbuRQiErSnn5Rod9TdhEm7Rd6WlbEKHcy440Fl
4s81u9xFXj2C1vcZTdI5JFQ0yJ+bRYHQys4bAZvtQDpjyqE1O1yt31doqZSrV8Fb
Mg+DCn6ixFlLEI4NrkRahJ6FPmC0fr9HjaRvEu39fXg/QqRWRqD9nqvk6Bw+0uLV
mJsQqyF4AOiMLXKUPw5FGs9sQiwkJnPspDvYIg5EKF1npnbgYXLB4nhCV0OJgvaw
hlcOQNlTgIyR6KNbMUB6DGmxb/oU6J1vFx7i/owHSS6ZWBfGh5KGtVclPIzDLpl+
QNQSdiiWyiEkIK2xHKVRa4362aBgXW5+FHafuPhIaoslzoQyE7n5KVDXZHULtVRq
pJD7lYdom/EbXjWvWVyoxXo7ElXMnC9YW3q2Y3CI304u/+f/y9c8uGJaKDuptbsa
ArxjKN9LiPPZH0jyTeRxhQX0o1NHAxh8MowNhJXvH4UGkHNwOtPd4CjJiXlgjbC1
xFvzK8xpkeuwCWDfkA5yMK4HUvCL4Ak/tge9UNhdG/0bQPIHuJd0Dc8CoK5W2U6W
Kqf0K4RefKYJA9euzjePreZuuiQ2J9yGSM8UzL4f1si4ZqoeRYTPl/QVd1uGYHZS
NMwYOVsbSk0TLEv44GIJeLq3yDwuQAFHkYQ1Zcsxwz4JBuj5VhaQC8c7PdaKdfNi
+HPB3J0Yd7VahEj5EO+0QR1sDlsP6EPfuL7uu5pxWBaEQrkFRMvGSmtLnjBbhMGv
VyU5NRputq1xqMOqnLpVSsG20CtpDy2o17eO5ejpCcenoE3AFr46yzIdX1M7vCBR
848hOMV45M8TBiJLOmkDkXzcDtB8pcF6YIfmtzUtjb6RPuSU1K21BZ82jIGHngNl
vTVlYWzf0TyRZbW2mSC08JqOR5ZT+FpcRWHxmFd5BfwzYc017sbtq6sjwPh1Y6qc
ywejQyBDc9TT5OPILiuRB2t8uK5lN7hOnUu9QhreIs0hjRYonJ9Ik2m5rqSXvMPo
+7whpAWSB6T04ZeJXMr3Gh9IueLNLhXBCreoLLetvT2apzRahG1HdcgH8gaQm5q4
ZkHk7/nqU+HYs3X0nzJgkkrRug0KJMyp4Ec02cDXaKGP7LGbROiaaUb5RxGInKOj
itIKY0VN6LvZk3YnQ0K2VC2wYtL5oBAJ0et2reYPBbh1wvjdbzMWwiLaaiYrce56
jnO3MtwpmBCPkAuazqxCwM8Oat8BSmZ3vl7wbezPETcB2BXcEVoF3PEfHXXBPwKo
7rORgM/pqpLuuk9wZu4Ka60oThDbSEZCFvh1+4iyJM6Y5FggBEfbwMmzFcM+1Xrg
KLrBVa11VSKdCWMWc2xdxA2Yw1XGQvtYELbpvG7d181p0vVMZg6d4Q2O1Y4Vtg/L
dLZmpqYJsWPr06lt+KFvjJJV8mzHEgbb7/ez9H68dkAwQZSXijgradXvXbprbXzv
tjlCBy2NGzE83gsbuDo80L/DPk5x79F86HCxAQfgH+e62CULOQCZ3XUs39gv1yMz
ji5qyYRXhx8LVEwRg8ZT73TDTnWikcRbNDSzKj74HnWd32LxILsseRW3w+VeXc7J
gQyvPu4WjW6VJDB9Y7bfoRnDygKjGZUSc41vnlfZb4noaBic4T47WtRnJA06hRkw
E+WPHIN/vIAX6ZG3Pb2gUBq2hbY97YqKsGtOVbenPNahRkRBzrXWibcypjlzbcbc
Nt9ojHFyMT0vUZjLvSqe3PBSotGvWc+lkoQ83axnnrGxw14EHDjqhyp0lAL3YOVK
Do3Ve7E7/J0UxQdZ2vmzHJCISYKZsL78IT2OOSg5Wnq1XLyaRAkw93FzRf4rtNjT
qxMjtoidggAsv04FRVXOtIb3TuDSz1q9Ktx6QKowcfyAb3y81BlJfjU9MueB36Iw
UdkhrNcjkUwc8o2g20KmwJ95EaN6wwFKqIxhuLPXYISOxppWg4+cSOZ7J6z94+Y9
cdRwrlRnuhtByIlHc7tDN51+n2zV0q/QS6WMVtbrGAWp5Q14r6fLZnd50rW69Llr
hI5VYZuO7RWbnL9/1bv7h2ZurWqkxPSWReSlgwZyamG8vFGedyp/izkGiYUB9Psw
PHmmoDIkEmNDqyfrg49oi0c8hSJ8Hv/LH0+Fac/oh55REBVmWMtiUS+QUvQxvXFH
lUJX4HiF/Og3T42fA/9+TkNMVtX+ub3fz6dcKKPFSzdwbQC2mBNe75FztKu7+hO4
+d39MG59d36T71z48RJhmBuzc/aWveyDSH8bSfUxvilqmrz68a2XsKA7JeS5orWC
pKuGvm1OgsreIwG++OpYdZpscJcgatpfJyZAeLpexxaYNTJfR+7WX2PcOQWKEdZP
srMOlP1gEdT6HLfeSko/zj7ixPypHOiECCQt0slF29fmhHKsi3a1r26AQQPjkjbX
inuaweU5cgGDc1n1InTHB68ZIa3zIwmGQQNILyF0U7W7QLbHtx1b0hc20vzyiCcc
YsxuSPRWU5urKJ/HVE2JGkRYmW5xZBANqPlSUkndOC6N/vePMfk4vkNsm8ThqqLX
troGepX+E7rrdo0IudYzQrkd45RHOR1SeM1QZH/7MAfwEkuRP48DLsnQToHYT3GY
pCsNQaPGYJoctPFDPe5xOdJpS2IqSUhZTBikagS9VlM4wRd8TwKNxHf/XeCFnfWv
fmtufM6b90KP1OXl4gQX7NRTBobD6zGW3h3yJNg6tNtIhr6Ta78HuK1oKrQNF0XE
C2A0m8+Y6ftc0ZpPhMMLw/fRlbTk+V5k1i8ngdaZ2HEuFgBBS56/FRh5rSfzAaN3
8fluuQrRejQyAA4HKl5e5lbTVeU8KVpE29dxeuVEsr2Aw1F59AorKzzWXvN4+0b3
hsDvusxFkKjOATLXE/PrWq7j5qcrwQcfMfWEn+SfpX9SuomFgfNoKfX1guG9GX1L
ufoHKHvfcf/9Gz/huoZ1dfRAULyeXR/DbaKrXQGBUVT7VCbtAH/3sZlOFqmWZiqQ
dpuLVHC9LQFXMBGMJikZ+fpW4k/+SJ5/lT/NjImxGpnaM9Z9+9eflnbbp26um28q
pOjoAIuiC3dP7jGU6BETNR8TT7Ee4d5K3ojKmsIXT58PVA4Nl+cdkjjrb3WF6rCj
NK/kENia5tmVDwLnmKQjA6/BdJ7Q+/UN30hQF+wG5T1Tymsp2/e8Zg8FMMNe6Y2b
Yp2N/i5Ov8nEYSZPQz2KrYqh6EGLLnbrfo4xW4U9+17Ad1RvWK+FVt7sUHV4G82v
nyFdKtGVOSAA3dKLkXQUdxO86F0r1Atnxv7jZe4VMCOKPTUskKuVPPqEjNn9lZus
/RoxnYWDvIqLiVx1WN9cM6dAjV7P3tfKPc5z+KGsIb3g1T2mDKXTybTX+fcsqBIZ
UKbXIk1Ikm7YreoNbvFxiAHGHS6kkIYkp/x1Wvdyyz0ftzN+wllt1Qa8sqjLS0ri
oJNt4JIdwwk0OlEis1Icwig7PUMC42Kqk9qlOQOz0G5lsvYQxZfCmcuhg9iddjFN
kTFqFNvblvPyafImvp6vw5pjHb4pEf8e5VcTELaCjvwOzVBPFZTey+56x9WdoUwg
43O0KdVMAd1yE+v1/aMPf00uVZk576xhFYYKSHqADdLPlkum7eILDRwbnJfGEx5C
Q/e9rWgdOzzBuXiVYQbYA9Mg9ARhFZLsjABrqNm8TrqOYMOhf/qb/DBIjj2Pitr1
c6n/Xmm/V9qBfdPzsEIJCDC8mmGnPSS7oiyunLDi7f3yZ28Si51bu04kMA3EqoPe
swZk52avmd06L+QEPeEN3LlmA9OAGVDkO/dLbf9g8Y2hQZMdcSwBmZMp4v/TcovB
mTFOubl51f3SRW6GnYT1ZFxGF1LwU9JMdOJeWvb+lW5ZqlrNI+XnYZNnbLoSGr3U
hZitU/Shpi9LblL0yhLcTO4sWmmg6dayKr4wbh27ek5t293W2VXTOMEiw+AWNIsa
cYwDQNltl5oCPPmTQ0BBvk3O6LlvOsc+VepYk+izxaJq/7hLBR7BRk4hEEHejuZ1
24+2CdDxIXQV8qgYMHqlveTQnhrZRa8kdi4v/SZV6h/Bg949TgPOAE7+kkqFkSk1
NdXtfDXPBiMzPceIOMn1elx9MFwj2QpLX9X2vbsQbxQHIHxu0lvDiB/bQDos30aT
w9eT1zStEuMDGSMtSw3jv8pqO4FkXHHLu4i5q5bqqSXS38/KV3hYrylB9reoUmem
g5O8EmI4aacM5EYi5wPw3twtGm71qW6qfBuLdpZl8H4q6WFREvl7X22s02xn3t7v
vSPMa5vV4bgkMFcIcrwaEfbvvJYMnnvaB8mlYlcTAuBTS9X1TB6SIvEkhMFpGu6B
rKCjQ9XWboW9UI9e0PS+x22KeiBPuqtuVHl9jQMI44WVR3XwAjQYNnBCauNmXUJM
XrmWY0pIwZuci/wQf2ITrxAdN5Q+QOXuy2aOjL533C3YXeDgLsuQ6B2ai3M4osfv
dO+/K7Kf3069abJnfDStr/yy+wEYT5tHJ1ada1aTPR/P3BhIu7f3LccAYsVNbB9h
cN7lL3fmkYVC/IfPKNL7lVn5QZHtWeYDdE+aGb0tV9piNsc6UGaQrbt9CS9mLUJA
RZ03zsWOLck5loPGS1KzsLY1Fx/1Kz3ElbjRaVqwS3UZ1MHgrMaG1WNsrQNq/fZk
HDCOqCY1LlQevyVwd1QwGx/fEDg0sxlmsLDSxgIrRajPd0Hau8uvPeSEvQ94N5x+
/X68o1kP2ePbKcHYtMT/djQrwDBEMLfT9mM/7TrhQJ0D5zu+e6FOJSTOe0yp5U28
ke0Kqs8VY+OcnGUVaB5OxCsbhtwDFyG19ioqhEyw0hzAsxXGNlH6ZYTQtUB1aVou
fZ17wtZictoYpW0VAqRLwtV+m6Ys52HaauVpS+3GYEiQ69enk627+12kpGf3cIXC
KNYk3pzkqK0fCZ4Drx2gE1/A8Vmi0AEyXz5AqHHgVSaxQPFLbboiDd4ka7HbdZ5R
wlM6oIUvHil58YOMQOvBAuR7B48762tbtRgPwLK8uRNgGr2L0lEYL28F2WncXMew
bbaX5FF5WMImTBvCOuPZVZGGeKni1MNOIo3wE5ro1e/70YiLUwCfwXjpuY91NrLW
QqND8/SvGVvAO1MA/rEx6eaOXYWMikcdLqtenCfkvnthap3G1owp/kmyJ+MeZIcv
pgw6nthuQtPlFny6lujGRtyKIVkZQK7cw48HIdJ8ndo7dhONG5TmUoJ9KHPMh83I
yhEhsAf7CamQBovEYEvSekC8B+ifID54PNCUIeHiOeHExRzRCt0uugeevv82+B3Q
WFNfdUPE804bnm9nl/vYTsFq5lLFJ741kZeNLQCtHFqdmut6Lj5KfK+q1yXDAmnt
o9H7v/Dxb4DQzsvH7GvJOwLcGHq0+DrTUuI8Ce1o0fyJSkxkAhBhbcdpSIaw+Dwn
Q+pm2gWXU6S8C5vRCo0MknBbvUzr34+X2tWTVA3IhXs7Sr4dyK2I9IKyItaCDwM9
2DmlHjKDf8MTZiJI0vz6dXYibldX//4rXEDo1Lc+LE8q9xxw8uZO1RejmV+j0RJQ
16d/UD4gD86kYA8rDMnpaAuaIIMeytQPAcNgetbGTjkffaTG2Vqe9Qdq+RZXIWd3
YfCn1UY0cw43RBpgB8o6A+TGpd5IVMG1JRjZpS+3nCk6zWcUQ5RrW+m2i0I9ehAd
oNgEFVkFR9guDSGisujqPOv5IF4m/KmJbFMr+7XgtEo5CiDDnoCX8sjfeIXJEJ8i
NlSy7qXc/WF4Jy8Dgj5SgqqZC5rSKRvEesQWnIwTkfM8A1yjxgAeRUxMXqa9O34U
V9ZWXqKQQH4B07YiR/KRsQnpI16UzTMHiO9mtC58293NTP+3HQsKF8tZjmjmnQqN
CUl/vdEel+pxxNTOWIGWGjlDZltIGWpP5vlsM+QfzIPeCAF1FCpZrQ0SaQeW11fM
zhCx0ZqhWXC6l9djvDy++9TyDpgcICsIDNFuvw5vyf/AKfmfDURqeFxu7XKZrSRP
lVIOHA+OTvjulqhkV0c41l7hYpbr9C0raciYS12dJmsmNz22wdUbUSzV0wZNOmaF
0HybSjKwZC93Linbw4EqbACAwnF+1BhmBz9xGpKk804A+BvZtcRaX1k/VNbymlwA
H7KvIrha4dmICnfRp9djlP/CyKPnQWJRb0ZXXkXEFWLYq/eI7xf8heEKQ/xW+A+W
zeEDggrzLLv2uM73VxT1WLTxYKb13GJJxRtmu4JCMU1jYJAeAz2BcRCyKNGMrVzq
2Z9hxBlIhPlLbacK1gAgG8lYVqmJJbn+ATW9x4uLqsz0aFEYhC6sMQ4lNlz25jfM
y+D/RN28+BueRj7mmpg/Sy4ZdWsHtropoM11Db8w9s9oq5s9QUb4yiskptOIgPjn
7FdMUeg9TycnW+snccAWQTm7uMevVjI9A8azy0/+AadXq4LsFDLQsSSX/8pU8MWm
rOBHp1P3vEWvzw5jSszrsh6ZAJZh3KilirUL3L0zNsAd8R2VMgaiVqi5aoNfb6ZU
FnzN2bJqWuzWSgqm9sgzIJsG4VNphvmC00Dzum8tvY0NvsMF0jzwOp9loU1pMSH8
SOVVqJ3l08TWZiIQ5jybMTwu8bGSu7h+DpbAy7BuWepGaHjFj0XwzwLIgBuqck+H
atyABbzVHH28OLStPR96h4dcKvExrtIjM+MvouieXlboPqs1gawi5rEKqn7KPGXG
+SzFRbUi7CxtjboDD8e5No4rnO6wwnJcd13TlqvmFpTdqGwOUsQagPAIvpBxBV7P
v3G9hMGnB8wTzu+ivELZqfs0QM054mJ/D4kR1X66wZR62t61FxDyVUPXDemBD8u7
n3vuC1VSKSVCRERmw/KB8AhSYKlrKWOzKSRIgEiHGUiUDaAFYPRNCdS1DwBDpt5G
c1EqxTkDjXoSAXEzRxCKUmvJ22u5qIlmu5jDjXdyWxRpJ3nXaORc7IlssgiKew+K
JImVXuZsHsdmynLhxjJf9krte58z7L/ih+qwtCIqzqGpVl2nkh3hYq27DgVc3oad
8cQj18l2fU2SL8XoUKe5DE+7/8OKgYQy78Fs/56gx/7GSlhc7SF4ARW1BT7UBREU
X433aOe8QdO2Vf2MyX8jlo89IDeVyPPLaDZei6Lol2sAocXbIDoYwaPCLeY2d/Xi
zTyIklI3+vfq+tokeA2A03LN7mjE9pn7+vtBLLp4CErKXP1KkFr5lILLKEBM/Srp
mfOwWNZzG0GxDNTqmytwU5WGtJgTIifCAemCEYtHh/UsGLLd/WOuQDH1lVbzb2Ac
R2O3JO4yQNWRq6CTqBrGbQ8o5GW2waW5z7c0qcN4gxngb9CKlZhLcUTsRVubQeiD
XVXadgR1JIRmAev+5v9KdUB5YMc3G4u7G8LVFhcLzizdvDbWhDcNMFT4gXBKHGk3
QxYDlQ6UXdImd/cWgmxa2gmz/nUG2bZDUGUKWRi2HDVIAPEjL4ZGuIyZVR5hKPyo
IFuCl/tRRtsvZgyUTgEu0YAIqPl5Tm/zRnWypOvAiYmVA3Vs8Gi5vyADYhSps0Z2
5B/tWK1xjd/V2CqSIxLrJC60p1MahzCi8iptBVZg20P5xix/NkcCZkLxQ9mEHiYS
yeAFgor+3mdsyN+vAhuGQTjiC1k56VDNwYq5h8btE9EyVZnLulLI/5GUwdFk8beT
5teIY7ymn60C8jqhcFBQHS1DFe4EV8FoXAgolATquj/GYhbB4ujSdcjCNkVttNwy
eWEnBwUNtSfq1lG22i7RN6LJ1qOhCkjlekgD9WbVqIICkbLWPKdFeYGNwOD5Zq/F
QLMzUSxbW3LR4p1UphYnSAgwtFrfBc3mm7mS4AE1feSNqqjR65UgDDlkqk7EJOOk
NKsrDaXDH9fESlZzWRXhcWa5Ul6UFAWaNJBjUSxsqZR6/MP8EOy5w+lS05rlt14O
wJ+5mnnQbIR8OVHgmMCyGMlnA93u+M4SAGstMcqBVhLFexh5gIzdVgwz/OApxhzL
o+WFJNYxUsGAccYU8VF58op39/TrfTogmG7llcKslAHHyaxk6rwCQjUX18wIVW6Z
g3dPrTl7Nmqa6bwHHYJVQrbxxzXvQjP/KJDqFDHaAzlVmFH4LtlojVuSQnjttqWr
CARTdqX5ri+Q8gM71Vxvh6sIySWNiibVRKEcHx/glSdUvPxXQVsIw0uqrk0FQkSf
OT1fMMyL96UJbwRmDaIh6oV128+XtZ2joWpSZ0onE38us/jIsMwH3nLVJLwEEA7x
8qs4eGnBj6GnF8tqTuhcWb8IbQ5PoRbA7eK9LHJlXqZhuE6ugn8rMW7aw4R4dt8c
VSvFYZK+5Zi9jRjxJV5k9jCxd3m3uCAarTuHQFZKS2fy5i2AuN96PIAPnbD2Islm
Yx3MKn9QkMTTUGphy0NoG+cxKkPJlbKqAlbb52tt/xZth3XR7ZAW6i+LrzrzwYYH
Ez04H8BF8BqJM8VspEYHytFLNjOxJOaGrT5PDLoOasKGvCqe79KZigXOubSFPP9F
93HH8zJw8+Vps4lp6sEXazwKjFYekJbPeHwpRgXtHknZ9JD4Uxd52wMwLXxCbtif
LcfdpGWa+XlJ69Ya51+PLm0Lxrl4Adv+zO9+72TR/Afs5OkAlbGKBQ1U7CL9EVxT
wuSWWPxYBbmflZbJDYQqX2ObRrfRN2j4TURvDorz92tzeW3V/vCxerFeg1bCwO1s
JyTcZFkRN2TWpQpozE9ILr66wQErkfKjSKkF9s+TlYtdjadgOV9jUGhm8Ia7JQs+
Tlg1x+E9Kerqfm2PWQe8x7hGzeiEwHfhLO6KvISeMfQP07Uhq371nIfb2nvxWke+
Zqs1RpSE+HJST1afI2IyW/QtbeMvbyvYRSEDZxCEfrKAtIsJlLRQ6EZTR3z9nhNi
p+Ijc2oFRmoCDss9LcEdy5+MR2W8e0+U/rHN4mInPpcmEsKGU6kjPWIDQPS/3Qyz
muyKWTVQ8bUDlc5Yv+rJztzni1ZimCAXbJg1ApSngLMeLCQUL7NmPI/AVGbyoUYq
vRcwd8+EDkPYtrGBjZGwbDObe4lFkNM82ZvjqZV/6NKUOe/DxPSPtoGyGbyf45o0
LRB9ZYNVrFq4ZRnq5CFhgu/I1shThIAMDWjCyZ1abn57u40XG/MsJcCw2rqEsBYi
58kgJcVLtTNaIXkELNKXM0DIWoTwKeNruh0KVhxvArQQYn4NN01WHIjkgYWuRC6X
ms4nDESm0ayzwQYudfcJpTlamuzfT5e26g/mk5AvyCxE658JnI4nHrcZz3V6Hn3d
wSQFVaNBoXMfDfcg5/TJ7xcE0TVJc6+fH9mRa6cuWXYjrUtmYePm0Laj723iJRnm
4pCRpkCucRM+QiGIAL4cu8ZKukU8YMZ0CwLrZU+pFdWx1hJcJsUqIxAFnoWXwKj9
eLTlUQTr0keoChTzkU+EejRjcA3VCRikmuklzS/4fWzRnmfd2B6wNn0pQJ6XxLuv
Ekzg14G1+WA1w9nTa+z6MTPSjORgfLPGuqCrqiB/762gLvspiONWWaD8UQcezddg
4+IIxZOl/QEZ8PBHCNfFsshOTPc2KUEVqMUyMc1qRH0uJO1ERVTAt+gAZOEf0oiS
8wTqns0/ZEPkYrcvXffoyIuPWIrtoY0b/4/iWXeisMJRownDHio0f0O0bifdaVKq
cyHihaBtDTsKYFLXHil68+rikJp0auVoqdi5ne72GdmGLOzeMPOWqnz26uqxqhQF
WkFCufHXYFaHnTr4IY3TtEYd68i405ww4uH+XbEGGMMduqz4Dn5WDFlU7SYlO3l+
GtLa8xEmGn0zZNlnnLljEkYBkGr7hLpwnUJU+cpsbqqHuBv5dHBmB+HOQpyMRdvs
Mojmzzjq3zsDZsWtZLztLdSYKc1N41HffwmusXD6jh+MzoZlTbv13FHbchGZ0lEM
zlWfANMFZqydni3F4jMds4CIr4q1t9fL1MPWwnF5Im4DPWeR5Voap+v+mChiD7dT
2ANpP4KdyHMdza/QKBpyFXRvkk4RGpU9QR5VIxGhkGPYVlqvWkAYdjv9KcyiVUT1
w5uEUISokVIjY/q+BgAcw0MhGGR8P4UKyzC72tvUgjK8V7pki94d2dtK6PgME/4s
AcKxgTyg0qeLMXazNPTPhEeBMDc6Aajkv3tlYw1TGA9gW9MJZJEHdnwDgcJe4o4k
MUagdDOH7yZ7k8WpotyM7TqpYYBP3sRx0asetYP6fwLYdI0fIIy8Gp7dNweqsyV3
xhH/DGnqFOBlRvCvu2kWaN81lAOIGlYU478oquUvPySnI0kR+arXpG/L30zgqB0l
ilw41TuZj7/hslXUXuatze9FHfAGp0WY5JumpzxcbZuNMEmxoO8R+j4tv8DSdgl8
OSMJr5zV2ggAe9DVmd5ti3g9MCwx1nrEyfVyUlvx/cBEP+icWHpjc0/QsWipgjQv
mS2mLnJBeNQaq3hBhZpgvzXnVpM12KmKABnUVa4j2/T8J9LZXeY0BKbD7BishWpH
31Ngu+pfFLTHmCr3r9ArDJ4ToZmwjZCsyMxXRbnBiQhwEx/0gNi55GChfAYJYFxq
9gZvpuvgl76zTSAlx7E55JjPkip0ssifvP0JSzP6A1S6Zt3nk5w83guBo3qzGV1f
kmY+y2p3ORkD5ecgLEO9OvPHrjWfXK/ScY0rz8f1vG7nhBPGjmu+NwI3LsJZPB+b
sPZokkrIx9gxPdO4nFi3cheT8+ZG2Jwbh6F6GYSB1MO6R8GWzLxlysGpZMPhyuE4
M/ANXN1/u5X9IrRuMuVrr9vNyEnsYI8RPfCzYhLblG3AOLn50H5olsDPCUUatDcv
l4kkSnSFV/zJGDndPp3Qrhap+4Snppyt5Dq6Z2V3CNrDrOhfxN+lxrnTZRsQlJko
OGgXYMh1FQmsUhBdR9X0lQ45aUM2wjHI6AjYTQ8JcUNvRUUwIPGQfwTqCV0E/fGG
WfxAnrKJ/OBskBXhXF/wMTm8PqRJW+EKlO5d+z6Ios6u6lReeuu7/V7QMbNagyD8
wXPSKql1yeTMT0RrpYWZoQdDJVkX3vWm0bsxT6HmslMYFrpyGN3jjGy6ikIfeh52
Q9MUhZTDm7++EXp+tANEPvrEn/8AZvoaRaajqsEbZYcSj4p/a4abnQ7Nj3I7/odR
tZ9hVxcPrsDjpnO9hOWNvE73ojvI02eqx6RtK9dhPo7jLMBhOO9nFqWqVMVDBj9Y
tAYBoWbWLQ/REPm5Qg9QCqylhy14ColNL7Y9HvkcBSm9rMrkYTRMuuaszqvsnYe8
fZjNU8Wcj3fhwZKPy0RjSnM48kU/IZcsGxuK95XhcfDuxXimUKIHx8DKkGXWRj03
CuNuDmPG7H5+cTMtLgp/CTU2rj40aI9UftbED2exHRbNGJT6s6GfUVgE3zpBj+ob
msm0roIWlDmiizehoJx4QGlQuH2TJCM9ESs+z3hAUb8nW1r71ZzNeIEFl3iXzBKk
b9WdHxatz39nYVmpKrkYkUYGUWHzcF+l3wIdGQs962uOXlZk4QkXn6ZxWsh15D8E
g8MF8pr7MSIB1S5WoqMXfH+M8N6WJ8F6xZ+ppsmCu2w6/UUtfLUyVN+cHE9ZmsCy
2HiQke+xsEF1nsFG3o6luRz2F82vMg/hSwvF+KFol3pBFliyWmRI1NqmmDcxS2zA
ZGt+dj8Fq9B8B5fxVJoKM2KgARbuYq/7F/0+THaXUgKVPHRJ5vXnS2byz3b/nDIp
HKfsKaEDycrnCzfcVZ7b8OETIyg9NWPU7XCwcaI6dgen/dUTsgUdcQlcXt2F7vdZ
g15KEFzMEJK6DOhiD2f0WuN9guvCTJdP3zhtDGYnMgTdLh9XEqRPvyxyNuwuNB9G
rZF/i1WJqNoNWM5//wNhD5V3eh+301m9hklARdnmc/KDPgzWYZo8R9uh6mpoA5iD
GjGJjISk3mgYzv/OxjdzafbHkJ8c/Sy9oWenWlHZwzmoogIaLcanbbcU/mG3oHGC
E9I8scLDxn8/ImM738iIak3whn5NVTQvqzM4uC4OVrAkjQoPSVpy9hNQb7hNQrtm
x3gYclQU1hiGMN6ohD6aivgKN8mUlnxFjUdUH85dMIhBnqeXHtMU/v/YSjD1O22T
bp/PgtXqmvdqnKA9eAV3AjeEQkhcIZMpWwz1ChI7ZKHngpaIsuPdvRYot0f5SpVH
iXRK/HHsXkoJjp4ZWxOA1SgN67qAoUxqLHKZu3rZDfJp86gyZ/ViDCZuPKhjR2/O
F/Tr3Gdpntq1ASEOP97t8mIV8OnKPdjL5z9nmm44jy2JG192CUKLr/4pKsmZ9Spf
Yjnu2dVmio9xkFitM2eutYd83plAugMFd2M2GncRpE22l4ApW/KC5xH/70yKJiru
4ob4ozaChXDltN0Ot32K7rcLpF6Zwv/3buuFMiRCLWI0kUS+W8QMLJs+bxD8obQy
/RTtmv4UPq4IPkNd2ELROd3M2hTFuTXkzStRKDGj2ZpW9m0zPOGqCV7L/jk+VHPA
+kZtDArg+NN28TVF1jl3oZqzFj9X5MmZy2kzWMlPUoSQk/9DnExuHmnWSa4EE3rG
3zcyyi/O/WRDtWi7EQnFZrVjs04j3oZtdHUQ49eYq6NOCAR4mRmFOSPs9aKbega+
tTdWdUrkqk8hfLV2HsjBByfYuseEu0k3vCA6uP9VvJoCoDBrP76X3TpY7BwMtiBf
KXeslFS4kDaKL3ur14luFG/M08F4IfNvC+uQEw48F3A=
`protect end_protected