`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
ddtXksX2+yylW5zu6QL2Lhnb2d1sD00763mmSITNX595NcHTEkwn0zB1Dry37fOW
FufOhVzEJp80NC5qZ/+F0Vk7Ik02dIR0elf3clrjeJRK85K4e3Hoo4xn7YbFUIms
l/8VZSb14+JVGURjfswrIyCUotIzlzVYZ6gzoZwDXIi5gQIBf/gI+KxNXPaKV+PQ
Ufys/12rjO6aI/pPlqSm0hCvftmBcnezN2hk1UeXgOIuKZnogjOsf0iJVX2aOOWE
6pD/psybjbnsNB6kH5uFTA5frkzIzkzl5d9+YDm9OyC+k84E83I/7/j+rk4L2dah
QJOvksSIzN867/4Qt8qYTQ==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="MvBXkzurAa5VTw+1JJ70nePUfoQXBvZOku/SMmg4TwQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
oRtzZL4VJ4iwysPsC8SXYCzXS8Fw2gtZTOskLcDV+1B9Nzn1zTyNtlo6lNICRmmK
ZRVu2BmCc2G+fmzynYlNTnSa7C0Cuel6FYpxCBlOuk3OF2tzAmLAuDyOH3Z1Yjzk
a0aHuoCdIRKv7BrZCdALt03JeUmXKPdOmIlkVGFl8yw=
`protect rights_digest_method = "sha256"
`protect end_toolblock="Jn9CQpRhJt4rnzZPRk+dOpzAubz7omckX1MrFd4p81o="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 27648 )
`protect data_block
gD6l00tciPUa6pDNTk/+t0OO0nC/UTtBwLB41d4inuAUA3i/ALrNyoJVcBnAmEQW
ptbcNp5fxEUJjnOxnedyZEuEBxWRieZFQnkRdF269oOe719cio1HQ+6376a10o8e
GCdRs8f1Vn+bdYPfGagiCUmfLoMUTDDghIpV/zyjE3Y2rEMGhwHl9+cQuBc8GnJT
D5A4vSVbHeL3IGgiYt/KgZNhRo1BVJDuOPVfNXl9qw2vz5w8qlmIUR9JUnWiBFhs
JQOaBTZNtCPKraNmfs47prBTHYnu6IYFvF6xch7geaWRfYcnBkrGTcdEbrj+rULf
9ZV3PLiGDJj7mUDXFmzvmLJ4WwzEUN3p21X/zzoUgBLbjjDBonlAFzeFCU5FFkN1
92V9N0YXSWkxKKxWptQXy0CRds8a0JwHDfPeR0iLSfdXkaHX+fNOXkL03F2LsqNl
0RuUKbDuwo9nBmn3/E4Di6/aULDbAtsA12k/EzHLC/0InY7UNOR7TQ5HpTDZyB9M
AfP/sLrzilv01IZ/feNnw5C+R32mlPuxYxqNpd2km2Ei3ma0yfTaskkn6zQ9cZsm
NBFuMLOpn62xZOTM9bJi9UU3BeMqsCe0iNlBnLebJRbig0kLBOOBkpnhfIs6wPGQ
mwDWS0X5kmVBCDNDqaUxnbYx1HubpkGG9dcaXU7yYTT2kL99x48vYoYI/AgwdxQ/
mge6p2oSS3VAZfYWsuAk9Erlb28hGJMq7s8rHdVWq2yn5CowQ3XGwuWmdedu9AxM
VFENZLgDn/ltGbRYiK/xQnv0raxBqsoOJaKudzlTj7c2lZYm7Z4h2npjOFz9pLNj
srE7HjraL9KbHwiYKCC6uo6KYcmchKcgV8jUG969usDFDRDB2saZtzF20XrqrGrO
ILQSTYG336QcvFAFCzVhuk6NX15J5MshIaQj2QqjVVssgxbEb1LSkIbRDQBy6GnB
1NKo4mDHMPXw7xbCwVYRDxOP6PEWkHhI0GowID2ClIfacoxA4PWixBqIk0MCPQsR
4EE3kmSDDt+yZ9eyJ1Bqcs6SSLCkK3M1bcK2Yx9eB/yUrOX7d4r2TITKzJ1PwcE3
XCrkYYp7h3ggrEhLuVJ22IMo8inRBkKpVbB3IfXvZ6ySHka5eXvkKjY/MG8Ka0e7
k+kF4+YgZJABLp8FfEnB3ti1J+lIxSSsepYzJA3ghVClh+mnAUEGXIekuXdwFn5+
xhJ69C8fDwejy/3S/50Br3q3L4WGTJPZJtvt4x8Ov4rkSS0BuBb4VcNOrBP4M48A
g+FXPfR6vfbqvlLYVRZoxZ3y51nXO67RmUxU0eEWjc8yTlK2fyrmQfRMpu0v2PVB
GBmFFm1IlGCD+UutInlauJudD2u2GL7md2YmVS7AL/bKYojVtp/MfnvOWdonzUgZ
v7pTIgmJq/EgIGmCZLHPOSNk6F6RoSRMIry/U3V5368P3i9kkiX3wdKlItxQzZwU
9EVIziaTh/eT48QGXK58JO6Z5BaxJz5KZG1YSOvpVhJmPv4jbV15V8efH7dHC+ZO
9nqkivqW6oy8yOhMAnSGnG62LGD9twCMD7C144aARHNQ+S+GjbqGkQ0KZFnzb3lk
tVn6rZbvIalpwzlK8U9vn0Tpq1KIxmnd13lYVds4hHUeVCCE4JA9NsRjo5+Dshqf
WzZOX4cN8OA9jIyB3jumqFnZA5o/u8Y39MMPaRF9RS/9O+aRQFGkBeVY3fvi4xZy
hrxUoMDjcFnLtz+xdCGHcMgbnLC4pbEkHeXZuP0SGnV5Pz1RuQGw2gcwzigD/Mgg
XG+FY+Up674t94/scb+hgB2UkRGnUcQ97do+emASSJr2+nP1LVTtP/NtX3rGd2l8
4XmwgAlYhLDNJMoHpwHXhZ6hBGoynIJp0UgWV9MbN5kYUQCoJH1kNHJ4zg7cqWgr
GSgPyukcJS2RtSHyTvCqF5AJWqXDKJU717n/gJi6xY3owJxN7+IzZQVR7xJKaYTY
ISIP7rwuOmROXRA6eBF2CiaXfpvyOk+nv1Nt8HHT+jsoR5u+BHbxu/wMBjWXUBgq
lYNQWF2cpsww4xDhjuTzJlxMjm/8fpZ1yoxdovBmJWt8RAUVfxuCv4Yfy1cE1ZiI
GjplgwDsNnzIJp+wq+oXJpFsC4kKq471cVX7u7hA0kn75moWsnFGdMkh61YxlmuU
H6FBgBo6DmyGx7M/+hj3DCscg16dVsD64yU6yOR5jVNkiseVdIY/9ASdLwiz/KBm
P+Zf63OYUXbtMdwnCrj9mUmGrjzi6Mpts6RBz26DPLnkx2uzSJhS3hliZUh8Hrn7
lth/QyC+vRH11Xpd6gde01S98Py4PXqdVKBpc00p0zB6sXpyDjBIz+t6bTuenGIA
Dft+WxjxCvZQQDfqYMega38xSzz0fCVh+7T4bbr0YdAatFiy2dVy7xhucPuKdOyA
Xr6wCtSSfM1SwRSO8ZpkrABqbu7h51ppPXxK01euaJHp9ay+AZ6iLrwkb2lJWbST
qKgV3BtXrvgtTJnr/ur90fi5pt3tazoSfURhtpejDp4wg+dPGESYeRib8fVMJDkH
1/lyKRnNRrO3wlL0uEEp45M/2WxZFEoS4gajbVa4mrUVmLNxyCMGUIwjg92o+dcg
5AnhPYO/3l4PC7GmngT+Aunbii0cPOoYlcZxRuyBLkAeAUlBu5PqkIVpoax541M5
oScl2KUsd+kv93dWqWOAl5F6k0E4TzrYOkGTjhJnHPWjNB0Iw4yLld/ZQSfBZdk/
ywkiV8Jrc9b9u4NvIcb9OSFpbeXEyx2V7Utq664oWHJrWwBxCcwa0yGf3TqhqlST
Dm+w2HlkzNVlFeRiARhswYvXbkl8VBFx9iQ/j/PdiqY5ibeg5rFQYqNc5455lu6g
4HktMLP2WJl7TK/EtJy+OL5vkFUCkjt7YCc8taZOx4Tq5RhiI58g62RFN/Df5IIx
2B1+sHOeghT9nX+pMG0Ax4abn3wB8mpCYmpF3hFYJ6fsBhi8oiShkw4VTUoZhazJ
uhpvR3QYQZ96JJ3oDrFhxadbyIw1L7hu+/1I9db3qTsJvfSkjQXQa7HUMu7xAOgR
RVx1ELz3MMyL58d9krDMj+bjyIREnR92HdQMLREHvMW7bLIu6ZVB+5mgjJXJ4Vcd
vvGfOJ0j7G1UUA3iLJT+bvvc6g6HPxw7g99mguyunX8YrpEzcnGOB+NuLU72j8zD
qfgNDM+TZx8N4kNsLUXnaInAEy/OHHd3uu5O9j+MuIfGyn2dbjLCYbfbxeJDgttb
3N+Ya5J0EkkfuHEsI9Npl/9rjAgWB0aWiYEkyJpC4ED2B9TJQLqXaC3ZVAwOkAjE
TQR7cYRl2J2BINasjwm1eH6/EJ3B5uWjVZkLcKksjb3/c9gl3XeZH9P2k9OELGc5
Tkbr6dOjMzsrChdyvy54yo0F+orWFeCMFN75/D22aWUw85Xh1YphmY3zCElp0DMH
3BLEN5vGIjhhKbnS5OtxrIwHclMGSebsKKPDenQ0xxun5O+Rp3Z9M4zmD1R+sVYH
cb5q1i5BQcAqIELHnLkHsVhtUHOt6uIshWRyCDN+ONh1F2PSICRN4ZQLBrhW78+z
Ww41LPiBnCgIUEOtvrL3JBdmZH8Sa2pokL0L9sLnK1WU79Wclnu62eezjXTX+xKa
mimp03kbcwm1VDrNXyX86e/NYQr75siZnqTlFfZe/hvXcu22LG5QSOaxhs4v403r
KANzAdE5rmBdnX0CRtlBA6IWeT22Uq23aLE5HHHXic4bfSd++/T1jAIzgPj3SiNc
Ed3po4731WUWossrxVoJfEswteZXJDSm0q31FnYipke2A3fyPGbWjRR60UTQLj0Q
CvZwm5eziXfevW035AWZ6nDptt9/qCev+wfU6vuj6E8eloLicEXFD7xssaDXrZOJ
z0hdahWvdkroef7pSE3j4rPmjdzShxwoyk/XxV1tXtaEX0PZ5nGLVGz4bqLuF+wJ
PIQiQteaYxmh6dSqRpxxI6w8J7hdE2OWAhm9/rIvSeybLyCAjgOXQvflMWEJPUxy
PUcteZbtk8V6k9Xqjj+ghpGmNyDwBTEGE6advCBi0NL0+lpvTdERXLIz2UtL6aYf
zwI6BBd1xRXN8RDra1k6aGOa+S9IwCM19v/87/eiw9oYd/DJRm/HcLu1LU+EX43h
8JxOVPLdt8O14bktO5GCLo2s9dajFzag9loSosMnZmSDnSu1cwfPO8c2ueEuAUHA
ak8HBjt7hl3ZHa0B8OJBzP/Rc6rvw03Fmz29OzcmhNK2S3itQyp4JnFuVJEKtSel
GghY9lBG+B5w95J0dTzBWP9u2rZ9abXJuVJozXaAlFTPnCOT5cR1M5a/x89tV4PW
xepEQeysDVHckVo7TeMN+VztxkwwK8LrutmSCqsAFzkqzOLGeHvkawjvobYNmT8P
rEUbjsO/B9z0Ot1Zvuub64ah2Q0r5hCbN3vwO6T5qKG3B4jgk6LwbpuRWejCyVpG
hEYf+U+ANOfiRmU04IbiR9ZpFIDoRHUiDSXaWxwFrEXTSoPD2M1hHTazdC2FHox8
Dw/OlVe/wbPFeOJXHcqymMfpVfnm2t82k1KY0eq2V+kb+buL21thuUIoF37584TC
d7WbxBXceJeq6v+FLYKM6QB0zMSjN1fPTOJ5sHnDXxBOvxLSFf8c+b6mxl1B6SQb
vsjooi2RuaMXLw4BFGOw/xMUUTeFac8gOJWhYHeXYJHvqQafCyUGdIM++4Q3j///
P/p/gJs6Wc3dpA8XKJmgaemPw98gA+CzS87Pt1goAZ7dvrXg14Xuig2a0U6sXZwy
7ptZdhoOSO6hlIvj4A9cUn3rsgI/c4vE0tPAFayjtH/GjghRQS+wMrE7w2yY0j7I
jIjj0vsd6iALQ6KIvtJdFiKNXFrkiC5/OuTwgBCR35NO8aMZrrxBNO3KNKImMQVA
m2M5q+I9tVphqZZFdcWuM0d1n5u+b05wjXmugusNqnz3lWGnVC1RrwgDRQdJLEDT
lbUBKO0b+Abot48kTOzMde4Od+wLid33CCnWwupVLWEhO5n9Af9TYgZm/QSJKNaB
jqIVV33awONom3/1LSGBv5kaJgdaQhIr1EMLEjidzQY3/06aLacRifbAbuCLVSUa
8SrDdv/csWoKNEpmvZLFD10IhTCnRHGyhaMPCCH8wPMwFBEgX/YfBEGaqwptEgoI
LMOmyjSdA0cOHn52eDvmMXMih0p66Mu6pUIS0Flpn5Cicu9ktoXnS+CqEsKodTjW
KAcajdnIU4NMRvN4CB4m19NGBmQyZU+liyHGbrMuJSRMT9NP8+VQ7MtZ6tsiEF2D
2Asb1ki4rtMCPSze/jeso8TKaayzRsWNJ9BlIdsSZRjV9KzEsc0WhwmVgqlbBGIn
aiiDPvB7FlNp2c3F9syzBE5Fj0RlUw6vzx6NU27+PB+W6hSjgk/3uY821GF+SnNI
a8TOyf5l+Dg+pa6Hd/xbn3yoXb0928pAEzm82b7/DXvKbzmNyRlvaHGsc/lzqzpV
3YxWCFfo9331kDGGWpmWy2wGgzkb1KLck6zskw3K0qG5ASx8clDfeQUc1NQWZrlW
wqYCoBAfC0Or4o45ALGX9L77XDEOqzyfR91UdVQgaZQ4E4tMq2Myr87hVLpZZFiL
GcMEWF23Dj84mjEAescly7VbEm2A+DyGjJD4VIOUYZZyNMn4xd3MYUlSe84CTwuI
TfBOUiJ2YPcSd+x1iOSlpz+s2WAOwMUR+TLcE6qRrIX2Y4AeZ2QYKiYjO9SsO3Bj
VadX8lelAcsBSjSNZlGYShnUAVhTjne4bM0V9SXX0e/2WEzJNK6hShq8AZN6wa6X
9vhpgzm3h9u04o10pEk54CMkFPf5N+dhCT09HDK0Kxn4fqevDm6qMj2i+s0m7/4K
tBaUS3gH0i0PY/8w4GYVgZba+x2p0PBxZyNAqPVpR0QP5j63ROn+LEPbWV3C3ZJ/
dNCOyQb0aIuzGnhQYplmy0MdxQe9GXeR2Bq2bMEt60/gpb0AordRMS/HzVBCPFig
Kza021wVkqt7wCzQUQs/aYn0Q9l/46oYACuji2GyOc5T+bJVANtIRCFKouEbVumM
DJE95gxZ6HS4fe82gC8z0V4oHRNVIsfdr495l5HxBqXqG42N3fNiwq0Jzqqhu/GH
sr5MH/VEykjMCVS1TTpuYIKFK+N4qkBIlWHsM0ZRpRCMsTp38mEGkaMP7k/EoEcq
e50cJeRuyS5BOBBhqpPxCXCjZLCEfY1vB3/kx6w9h1+ZZOJp1Q99YFV4Y52UbhmX
QlwPc62v9chxMOaAoaCJgCMj8jrdUTiHB0Tqyh83Q9qgmqEoVMOdoz0CBe0jvbrV
7yxzF2eUmpMBtHPJ2hg5PfilN7k1z9kGxLFk58yJ51zFyuyeaM9g7sHEIAc18m8D
v6Tmr0o/X8Kbty4KSTZjyUYHN+/CUQQ/UEjfuMn87jz9xSFaAlJuzUdOzENrTDcP
1ktqcBLIiN0dHmoaDCOL2KE7+T15CNg/h3NMqxVIlC/mIii8gsKzlkHXxRYqqZ0E
oatwyrj+BLVoeC4Xu/ZMlWQ3GvQoXpO/bc25RpFcckEQbUGQXXZeSVyMQcPj5sXJ
dlKruoxs1ULTsKv+JJn9W7fdKh41FFYgUwpEZ1eLb+B8uBlF6LSH1adqdmmZbuvx
+WKftXayeoO7Qv6pNY08dXMkyX6ACtGf5478/ckgXFAd96n5mGDBKiV06J/GGbis
DsZinnGl2yIJwKyQUJd+9aiVjvLLfwdTuKF2ACXl7FcZRL5eA+rfF/nHdUPwAThL
I5Rz5Ic9eVZBbMNjZtSka4oKHZ0MAg+GTILyFGKfU43KUjbJlcEa2s0YPVrPRUFv
8FvvG1uJhIzWMblCjPH2zyMZ2l9uPkG5ByO8XTDEdQUWdan5xAKxVPuY2WrpYwsX
+x23yfpKoASrIJu6aBEGhevYTfaN359BdFkYjIYcQfeM5e9M6p8nVUUQoAjsz06F
jvO9P3ZQOquplhDWw5FcGCCJfkPr9+ZJFFhQ9S7NiOV7McW/H6zUqYgGAI5Z4Lsq
Qh96VyaC30bew50Fk0ZU51MlT9BVbwHYOR/9Wuv9JqY4MN5FajRm98akalPmgw3U
OwOTcR9lYZCmxei/9AIHAmgCaUFKsRRsCKZPV5xnzUp5r1SqUpg+zO5/MN48NE0b
pNlBVvIuOA2+qID8qeXLnsoNcXUv27UKWQvbH1enKRKRqFXD1rA9dfkmhaEItvgg
BKFzBXIlmetGC7bANRCvwxC4SEshDgFt91kbtj11tIwZbtGhJoa5EP6vhXVtw6hH
zXZjz7AU2th0v2ABzZDAwrYNr7z6RQOjvgbRoGzk5R66A77/5DQdPu/ROa2BrCiP
/u9m7UX9tI4h8BtBrVPyLV4JR/Dpsj7cqNRdf9Vg53vveoqBTUlaNeSR0wAwqlYg
/geqJy0QLfGCOV5vFrPdQvpaWJP2LPZUNXaz3haPliD5XXV+w3U2k9p9XVK2CArJ
krEJSpQTSQwP8XfIv5WFwni/DPXNPDU3sUd/63zDALZkhEojxKryWAmb8bV7smSk
SrNK6KZpEBYlXFMGLuujnsfedHbcqCRQCYRNrp0R2w649KOW4hGiITVjS1MWla/x
M7ysGHdK4voBLwd7nnLuus/Pe7w3LXJsYbYdOSsUTMVKzPbcZhluNlTQZvJop7vF
YmgB2cZNdz5tAxzAYomOPJhPO5qgZeWMMZkvkY7KkaDtZOuKY7hefPl7D+VSoLp5
g9N5dl3MrfZ8wfaPn05EgeqEbEpu8Ig/YIkUQKhV0iLVkOf7MPzmmQd5LE2Iyxbs
GzA23K3DaY2Ru0GRJdo897P+nizukj45L8yhs8ZPnv5XLOKO3KwlhmeBlWsy7fkZ
ZbucE4san09sB/WN/SHBy281jm+EGFK5aJ3gQHg4iqU8koAF+3URrChymajUJbtO
oXFUYkeeHrg2j6gpT38RCdmQgtw4VwwpFipILBdPRTB0vmb64hMkmPVCHkX/602N
0xNJDrQaRGz0FI2oyfCnTQ154FD8SK4Faof2XntlGzF14nCT/I53uVZViqM0EYGH
1NCzjJVgUElBdQ02cQiviQbxN+DkLVsioX2wMd5s3rChxNZDX0/kHOYAgSktMFU8
8UL3Majizfq7cHDRh/n7oxTYfrQmBCKxOkc0Tsu+aqKyKrZ278w4bZX5V3kpD2BS
YJgJYx0zB/+f078xSXeVuqskUEYeLMi70+F/6R0x9MG2xwmilaBt4+vHQczK3Eyo
LU0UT1s+vh1k6zMtkJPcFITaKkxr6Ow5TdhO2NPqP++qf7Chq/p05ndVyLh5xIre
uwMsEZ+GdUWGWWDxAwHgeiKBXdvKAxJxXu/25dCl1vL20sWWG340k5WKNvVhee+S
GojN99loqftw1Zluh/daxdIh4WL37r+cViwvWqK16tnqD1h5RbHCmB/0YGjOBDC5
E2P3j6eCgJT4VAOnSXyHBshAy8YZk45RFeExeaAF0b7Tw364mVdjY58ufVFwo0Gy
LoiFzYg9vvBf31co6ytqWuCghxhQpoIb4E6Q06+kbqC7v/w8FzdrUI+32GhdyFtO
Gc7Kow3Iol92WT1HmowuqcmJvnhTpyBBJMwKIfcdj29O0d1iniQzh0QF6ibzA8Ql
NngEPGAoK+l+fm4orrztm7QIxdBt41g+4/euGfw2Mj5A5XJ/qRSKmFNCh3zqYdan
NJB376OqD8Qrc1kiHcND3u+yYe6L+vAMq4otjZ3d4Fg4+T6LG4J2RDFBhYmKKsB7
yoqdKs3Q4iOFPH1Q0v+vM4AV6KTCXpKE7YXvn6LpV2YnhZJmWljoVQXc3Mx75jS8
5GSAvC6gIzznK9I0bA1vFPXb2JhDxjtGh5S/wbkgrC1AAyf/rUNpyopnO1f+B/25
gys/g/TorR4SZuQul97i1JQHkbedA6IeYQyKnQQTQM6TJimM+d9voVlV0CScpat9
vnVbu5u2dXzjosJxK4A2FqzngXZki23cCdMcS6dhvsEt72sONO/2trQG92s/7rD9
GHqGjmQ2o5SsO39qDteh3kmrPKBy7+ysnCnfEM1Al42jtkVsWKcrGejk6zuzS4ro
qJg6qcO+rVEAS3FbIj4lWyMpmNTu4ltz98YbFpQfHUsBXftqO8LkbHStn2k3UnnP
Q9hq1f8IaVAxrlRlz8nvpP+t7ILphebxwEtDR0ChWMOXC4UOsPtoVfgkHWJ7w1z+
pC6/Y+9Gf7xCx7IU1dOOpEVLFzU6vQwR1WHUs1gj2jiDOzY0fuKWHX1WdN0pxGxS
ThltbNER2pTsB5dm7wGdij443SQPqX3swPoXVD53TAu3uGZML4sMTgxA4Y+PUnGQ
openQiAwFORth9P5yAFcdsTm0aXNp9vo1mq6GZ3b59ShQk5hHfZSrpiD5g8THCJa
R9ToyDPCbSXp1wKP+C4eB7ndzDw7KouDIILQEKLe+HYjnIFQWQ47rv7Q6mnRm2fU
z2VCLi33Wbs4yneFquD7Dm/lon2hC4iLfhekSR9aybKlZwRZtDTuuEkA4MCcmdll
Z9GHRh2drdPd2BP7JQlw5ZGhST9+fXFXOJtpVyeLkAyoarhWS8F/Isswb2CIQTAw
RimNtTNuz7T5idCse+MIAzrhZ2JxJxidAEKkokuQYW+7McL/N7gqNkmUZl3zkrzE
nA2a+u2yOvS1ZuP0/3rQw63pBwnoXPxWzV5ehBBNJbRwQo0E7YCZ/ejpFyiuGT+o
mK44mlA5h+K4ySFP12d2u0RpU3lzmZ18D20KRzdGrfZbrWl4dAhMyonQH0Mjj+NX
QcRbxFlOBbCBAHrIoATmsrOOr041pr5FsJ0IxcjQ5sK5pJU7gpGeLxxmN1qIFO5g
IYH9cQY7AUzl/BKOaceEraCSyNN0/XVQilJg2hdPDRKiQphq2MG8LH0mpElXPSx3
hHl+8TmUCHtprrhBBb1HM9T4jxwKd2i2rc6O6V3O6tbMOzois8MZFLqu+IWIZCfZ
TTnhmjivyb7hT2q6bTqcTgQoE+F3Rj2YQD7o3YA3VXW5bXJMfnBjsiIMXFmuoUQS
jVT7Soax4E/4Ltm1esWuAmGRhNcJKOFMZWa/Z4hjmyEpwfZQPoqIuJLGLwp/conh
V0xTcMd+jYXSs9w3wGR4UBNKBYZWAxGbcHd0n9EV2j8J31NP0BEYdjN6eG3aeL56
aNny9d58PLfeJjygiebNgMsgiOYI0knIjcepi8Z+TaG76rJYrQ8+d2l75RYHRc5g
sEEZPFjBefH8S3w3yK4G/D+Mfi3ccwHqQUw9fJQkBuQ6/R86ZoQJ7RHaWOkDSH9u
8oBYB0ofJwDgjK3GbJyTPYfWwWTo2GpDlhDWg/9waU4u1ycERx2zb+pNUVbiLesV
Enc1pGAdKTWaEwrJzbowO4GyIRQH98XgdiEh1arhxra+0b7xGSSLI2Vj2mW6SPuG
fTsEhuIzx3LY3btrn8iafVWbMpmKKOuJqPoMI0I4eSpr/rTAi7JgEu5bVThWjAvk
UH6c4ClR0cNFqDaYv9wd3pdIVol6G95Oc9I+A726EF1WqYmR0202fWHKTcfIOyc7
sHrk+bm/aEbbuI1QrDobXXLOmH+8r1uJdk5b7/e+i84jDboAO4lMGYta5KEjTL3H
W4qPIMTpqsS530KuyBdfM3HkcyclIie3CqoN4XzUROw0+X3LulmOE44YBlsSTMkQ
Fx+pbhAQ2mO34lIIIR1YXdImSrEPXLqlp0DhN6popxQu6owJ0WHQG2Rb63m/LDrO
dNS9XcCcSBWH8Nb/2UaFXFL/QmgrsomrPJ2HL2eB1wy0Qq071JYi4WoJF7UsxRB6
44PcdCGHK2ueDPGfkiu1ub1XctpVZL0A3zxxMfeh8cxOeRz8lV2c49OIOSrbd+04
YrePOr3Zk5xAB2Z6VL/aDLhDA42dxh+A/0cVMtGwDV42zUQDl4NMSzLMgRvE/0d8
KVX+NrIGkaedvZvDqvEzxMNp9gDIlQikhCQJp7FL5kmpqENp0to7ItJWMzgnlbrz
8rvILCnIyD2DjxMaJHTfEBO0a9ZqzOGh5rO7NaDjw4TnSaBIXdlnj0Dw1WDYctAO
OQflFG8Lwnz0807uqBZtr3Hz09yadk+pz8yenfzoZox0nzTUqd/cxZwCY8icwStm
9WIVs08vaX0IvadI4qmR8Mf0eTVcO3s2Lm1Hl/i55I951Q2iFURU/aXcbRhpKtta
SsYF6HyrwozcVgBPNSTePO9TytdZtGhtqMbSIR026l5mheivWGUHT+9zhRa38GeA
OscRoN+kU0izNr2kh+ygfbcfbP4SHIHG6epiGdowjIxxNheQRWcDiihI2SCxRrAC
t3mOiflRzchX93Y1rEnuKvhWYLSkRzehKYFLlyiW4MHQp25mFpP70t+miCPjYkJ7
8ibfLLkYdlpFMpfmbj4AC4fgL6HTtaOOhTTRo5YjtzFEWp8fTJmRUlAfTbJGH0iu
nKmT8ojNLyUyNO7pgvPjC2Z2f4dG869B3UyCoeAnrewIFW3z37NIOFLXkpuzBfQ8
yI8veIRcSNn8GFYOgdP9z1/Yfl8hbpwT9ox7mjYoasAQC7jqgkd2U1/5w6G96OT8
eq4v4nXTsTzD50B7kBls3Y8EdnG7j3xcfG0IedENccvXofWEZkDPjx4+N5BemZS9
+RXUvZOPVqN0EGD2nRzRiWZVs7YJePCEViNEuQte5AAPKczcJgiL6/j6tH35c4BP
V+SpYHAr6U3ZSUWpeYoPN9WEJfUuks0ipoeippvADODBe83w0vHRkh7Xuy4VbWsQ
rqOasHUQulRU6/NXA/fpssdAc8ruw1bGCD/bfXSvLQMPmVJWD/MQn3OSPLM0SNG/
P8VmzbdkZ3vKg7kQsbOPaI5/Zi7BIzBcaNBnXGgS6mo47/nhDenkVpAOHAgk7wWH
c6f0mz3zF3i4uybD/lM6Gm2mLOzoFE0+hAQsXpM6Bp9D3dcIvQRZKhfq8Lh1WhSu
mL2NX5jIZCLPPu4jkbWAEQws3PMFt5erT/6RstdGsdAMKxnZZOHlTA9Eg5JD3Q6X
JBA5CW3NXEGAc6Is34tC4IpJkHM3seiUZSpHKBX6cJEbP61+VNUIBbo2GSayP4+R
P2zJ7LbEsPMqUHPGEOCzRa4KmQTUzz2JKbBakH3xUS5JN6rPV9N5nk0oD4nn0DzS
bC3JhsJOJ1GvbiRSm6CiN7lD8Due/rwMhdTT2LTUwizS9Y+8lbkHxGqxbi0vrN0T
QnzxURIH1Q327F+Moa0F4WHOFdQ9LQtJd7o0WmuyeOSoiYGuJGxbVZwnmYcFBgzW
63ZuXDl9LzG+LpMxAjVYvhIlIi1PybJSBdZ4KPEjTijYXR+T3VeMQGpFD5ulW4/h
hLpg4U+fBpYr5NtsG74n2U6LWR2tQjy2ra0Z1ab0rxj8tRYWzZY4rxmcTIpgqR7s
XTgD4bXYDWXVsSMclVnqbIA8PD0kqJBHG1FI2QvZcNLUHzIOLve3BUFKQSaf/hPy
+qMNtYqY2DxprwloVrWhl/630R9sKQHaw8Upyi8bccXMo+p0otFAEeyEVUS4vpQU
3/pMwVgkcfH30EtiBj8npZDu7DfVmjxY1iN/w9yD8wf1SBuB6TM7/6jvNa5DXCmD
dSmR1rGHXfrWBfNPWgsYXuToLro2hklt+eAr4Utmca3jZ8NMl3+uDo45ZUJpDiOc
BAjswkWoOAx21MrYxo/LyRPQLyd2apRRTFr0bh7GQQbwl0y8DRiwQdgoWEjstkrL
sY8REGMfxYp23hqMlEegUB6Dt0VMuutDPslPchH0LcVKOSXuVnEM4vTmPnu7/hJD
U0J/4ro1AH2RTWO3og5/7vodZhAKDsNDt+aKpoP0fluUI5W7NMzjHLRVWJk/kfuW
b0odmlZRzdMPDg3pxQgQ9ADHn6vHjf6Yt/zqtgRaIAAbPeJFbol8exPnMOQkQjG/
HEx8bikDurr3MdSj9hdruqe8X2kaQx0/wNn90+okG8tMMsro53la3YSk//4UIEFU
MY/J4aQmGzY6cFXdHV+2spoHbeiKVfnepHVXeIPjYMYdLtWFUGk2aqt5VgiKrBBn
wUSNcHw24rri88tUZ2Evp+LXcjDo7JnRlarELd95HJd2lJKGLzGLx1reQLFuLCKp
lRMYqQTDCYhcHnaIHq9w9jhGo7wzCYNIxyaTW9h7G1E5d38Zjrl3l/loqIzygJSq
40yza+Qoh/p0XS8fL/fJnFBOSdEWLNIDk/Htc4NiyJfmDqktfG75t++GmeKcAb0k
33cvxcSOck9qPbB+I3IjcGEA1B51pqxsZO3zDdb8LgKaFATQPqRm3YRg+Hhkif/2
mvz4FESmmbCeMk3ccC6g2GI3geMH6aCITsi9rbe0gtMQgKtaQgGslUatAMzZF6Uj
s/ccj8C4Z6MY81+payhvAPKLdvUc3pN/jaJU+11X33s+aupAmCpXecPM+Y8CJmAZ
hJtbuWNMCd+KwwH2LNRx9Eq6g5dlhv8dzDOmzZxxh3gAbJ8J6n4YOhwJxK11BxXP
JL/BgZIR6vkKUk6ueyHKtd/xWkklYrvb2/boisVajhnAKuQ1wSn0JkHO7y7G+Y4G
5/9cqI6SLtjMH3up43vYeXqXOyAph6RXkkM2pEP89TYaEk05Te+DWNrdA8CJjgeX
gJuURV7QOcuwQ+4Sztzo2M+TlXEhNhpQkSJJVqAsTDNDYWnxLU5hM1ZONIByAFWY
a3mIyIpkFi0+q9j0NgJMfbJSOcP3080VfYDt06BZbLKd48ht0/PNXxw5YBccPrmT
1TvPxA01ACcSP3/U5WxKmUuLD/Hw510cp4XU1vJjw4xVOLW8kz9dUDEvXzxnGVbM
cmAM1HrSXHQInydH62mXNfoYvenCfeUmI7EnKR3quRRGOCwR1/mh/WhNs7VCzq0+
DV0aOOhQcAM6UtlZ1zksod8x8razKZ4llFl7Fp4KCiLSAJoAvtC/K+iLFXTXx1Dx
9XRgUGrIpO0NqWnFcGLW5EH9B6z4tmgM7Byzu3YWa74ImzXXF86D6HoCAaEEFY+D
gs7PUzKt5s7yaTpzDvfUp7X3jYai9jSGSS420z/ByRIG+Eh7JpITpKVSNP1yekCK
Pjdr1AntHcR8+mwvSuLVUJaagsBwmFcIJhph38S7YRswgCeoRYpUFTFYf3EKje94
UHqlPrF/7zuz6J1bzVaD5AaNvn5E2FfcPcPvylD9FCP3I019pdGihzW6DxHtHr63
SsOmG7MVrTJPVI032cVEP+EN2HRfs/y0xYSE1no9q5qagCmJ2HLbHbmPPVeK3Kkm
yYuJ43UxhSczKa7nV0pjn0Qr0EE/xqtW6wphuQmIz6B3yCHaGvHfPbJT3P5lYRAJ
uH1cAxOIMJ1gsgvg6LjDcRbhEC5jXIOvfkfaL1hsrGb+cTCLTcS8WMYS7SXoOZOn
/wHRCPiTW5Q0mu2Na//uPXZo5yGnJV5Itj1qP27DTO2m3U10MRpmKOIrGRfyC6Wr
Vl5iPEZJzqa+tgzCXkpSL+Hqug2aj64r5fbpZzmb3Yzg3ZQAIhcXGi1jL0ec9SDn
+qskMRiHYowj9jhqHzB+23TevM9s+/BRNyfiSeJCn9WBIGcD6uyi30bw0yIkjvL4
hc06Cp0ss+nuVlzfnpeBfbuU4em1rgLqz6MHNKvEIz2pACJT1X9khgNsonuwsI+K
Wyo5bRxmuU2fSlutoM/Y22qoBy1fwI8U4XcxQClrrjIVpWPj4GB6O5AlFSX3lux1
Qg0vk052cxr9B7W4CjCTK+1q5WnmgNx0pAoBQQst0EccV6WCRQ5WGEbWntcGrwPd
bXklozt2FOGyTHmeZQGCbxpgvg4otq66BvfzQkfTpBhjMUicTzNzdFdKNM6jffnt
5IhoYSsf/Xj1jF7pgBRj2iHzOYjGWjYoOPTDC9iuyioybZwcJBCHIZ6NimYpkXtZ
GP9VJtNf6QswSaGrBPa5oDM83H/RoutIKbOCoMmt/R4A4ZLUhk9miz7YFwaDDfnK
6YKPkcTqBzQt84Y9hl/nWjoNAuPMmF1Z65ihvXY0ru3QWvbUonV3mi4IrI0FMJCQ
0bJpZP3qqoBOxCJsCgVsOK5ssKtfsEm5x5Bo1eBSm5gX7v0d+vgMDTAWAGX3b66G
1fb5+lFZs/OCGrM+pecrdBWkp3fn70wGmMM5jlpIDsZVyP2c8DCsdDLqCykuoq1Q
VtSRrQ4jcvKfjsUsVK8GqQ7lxpkSCug4R8McmcvUpQERCA/9pSJy/ZXpqrxWRha1
ojlKsL0buIBnX35OMJrF6AMxLDizMN1oUPIJVNenZnniMfcY/nbczJUO7jGFIOnq
lWshofs1c26TLSLQG2/PVT6gRW6U8jtr+mCZhXbzG/4r7WSO1hO4qlKNXVYd5LoU
b8rgTtIAI+2Y1pzuwo5zpI5PBgG8JvEIvQmlygE+t76CPZLmXztZcbYys9qK3SXH
DqEHPeiTawabcxY1AdDKGpgJyG8jNeGyERl9nWbs+jxptVVzxYmbwBvr6IVaPRu+
13QEtX+JU+E887+ERjYeEmhXmuuUBcssw/fvZJoKBbeBHZ260dH48kmTN2yl47Xu
xHYwqRKU/z4NzBBnEXRUaVMZR/YrGwF+mfk9I4anCUgqU888qTY/CO3EfI+SJP1E
bcTo+/oDzCa7dgX3oqJDH9Ha6xL3iUs7aSrB7P/QlqLh1UGE6VEKpphti5iJIIYf
O8zlYhxybE5C+OXammx8jC9F3/VFPOV3j9zhgJ/dgy4+YGU6vSmC/bQpnZB9d4F4
e/c8Ic7bAySpyKoWd5Io86DMHtAG2XpxlOgB7cY2pYerjzxGVDCOesBF4XGBA6cY
HOjHRRNRDMobPxqdh9znPUim6ZRrIkAivpKZmwdoU2ihl2Ee6ioP2deL2d2/f/+K
hl63dWMQIqUoLRKBTgVSXm6/i3B4ZCbqb/gsnymJyGh557CNt4ewxb42E0z75zY5
RihfYWtIMQdejYBlATh2SbZE/UmLjWvq0LzBGbJ8qwzNcj7FgWo+DP/7chnovpe7
D2PBK5DN++oqyLE10b5qekbehvMqfmIcR/YOMRLfaff+C6dZemzqJMAeN0Zup2ZW
Ox4TNskbDpruE1iIrsBTJwxW8KXSOiqJpeUyxvJOVGHz9SG9somMPlJ3lHieD0i3
IDVSIbDpt+B7+B+pNlXYCpFcemDJdwkSYJgeZKKteJSPq4cCUlDcJ1jMbtosoVsK
5Of0Q/+hI8+vL+ju+lC7G61581J1ZFnwa58mAkoAAVULoA3+8X3sUmTdkVjBv5fY
lBnqPHqRhypyeWhlvgCYByuTxQdcHeWZzq4lf0P+e5t166HX+sdeyw6o4mjLENmr
UH53IZF4B1bYKRE6goyAB+xK7HXg/SGabrxOwqh7NMuoXcZq6NgxKyAyVlhmVLue
cU6srnvx44NzKiVPmR/mxtRGKq50qJWuSWqGu3Q855rZjsBcGx3AYUxWgvQgKHO4
jl7FAWuvWctRQ3D8yiUIveBc6nLhpuEnortC8jFcGgZZ0Neotc4PtuxN6D4VwoaG
dS7VM6gj5iB0eK9AbKGz1xPgKJU7xrlWogf1MrKhNZLG2bpNEIv0j3TWBrNI+9Hd
3YwCiUVzzxLMeqyHBBge/ngpV8d7kiS1d2L0m5OPU5q3vNT412k+f9+4aGtxrhqe
I4LYhRfuxCZhHEBa+5JFyObsxl05+YCfzramKZBHft6CB/QovKRDThAAqdg7EDpc
XW6lSCTHfLu7C6QtnPQieMbEbf9Jbom+9SlHBwgQdMfF3OcttOvo0AsXjKKFh/tt
36NvOStzz0gqB/8OccRb7xNAZkckDQHYwQxSeybf5FHqgDDegrRbaX3YI/f2zG3T
UVPWzKSBPbZYHJLqMt+Tdqtw+U9APPNwL18fBUfBnbJQZkFz1VW78uXx5Q0/qoDf
jEVZAYdLBLzr8/N3Hdugs7yRFHv3tiTiGtHqllEZoQOGzAgkiYAu7iT/NxESKJeS
OLiHjkgjgyIQq+XcACbv743zNgsWQaygOnSDJzFOOWL/GB6FBsD3W0/HwGCo3glP
MjlvpuyXrxlERu72LHOBL1X2870g8DTTIamlQOGsCZmWvO3VuIyN5jHkGP14mKE7
xpU2sPAh9ZekTNw2U2om+S178x1yjCBayyDbFiiU/K64hqwwjltpA24Zdylf6dcQ
YoR72OoO7aD+uC/EY+pIEAbNyapbK0TyS5OL0CzS1ovWYVF7H6rXl0f/CLKtVRY/
XUzb3Is3iaSg7QLmacDSbVoB5S1BA7odAM00Bp1ZELn0cvfzYBV+wD9JT4LCPGHl
Jf+o64X8C10BFrRsQZeN9lazMHE7QZm4z3/OelsGdsFBEIWqyglZvu8fOnCGblYR
C7MQwO6+gLYp0j3i/s7089++ykWft7FrJ+IIcDnnIxcD0TuOnhDNVozG/WaaVM4D
feZAS4T1Z0NzjfTcnVXKklX/d0QWo0Ks+rAzDipkKzClHFz2jKO7PugXP1borMWB
q8INHTzK67bbmG4aQAJxVJPBY9Wln8lvxVIvWdS6P/eDbevacVYg8nnACoaLSxX/
zacRzFykDn9Bp4ad0fsLbeyg0Nsfb05Gop4/fB4jIVc4/AyDDFCdxccX+BwEVKcE
+dPcIr3Y1gE5KI8XJPM6y2Pj+WRdeAIXU4s0cBDvFKc/2tvh2uVIjgvg/NUrQh92
47v6TlBnFR57RcR/M/nYeu/omJsXO5WiTj3VexiKaEs37fZfjljkYmxgruW6hkAC
Irat+uPDa1GbY2YQSkKQsaE+0GI+o+eWRGhga9DfaUDmXQs30qyVSGrUQ6HJrScO
q2Ww8/757+r1bxBmp1qQkWrBb/eTSpyu2qJQ7TZ4B+Yk/gyv78e3FCNXeqzb+8CY
jlC/eQIhCjHnMu4Khy7mQP5cx6rbTtLRt8r5TemvCCOzu1m7BDuw8na+HPfrYT3Y
P7tqLHmWS71HjMAZQ3gH6mO0FWfuh/1M4M3m3dwxBVQCJB9rAXXKdLCMrKTMt9pM
yhldKU+S3ugR3+xyG1esXXkYmcVBMloJaQtmoNoeepDtI6cKwsTIBkLWS30cXauv
Hg6TF0giGoYMuBaoDh/lVc5sy/hAI2TyEkjNK5j6wMBE733Sy3oOAex/anGwFQxv
bLXf56770UBeyJjC48FmVw+GHZNc1vjCDVNsvZGIcYU6vaw2gziAQOdeM/Ta4aYG
3cJQAzmb6EPz/9CsPrMIL78vmGEOBoYhY9U9fsgB9Bg+QOFQma6znOZH9RDE/DrC
bqJRZqnaxPDDEVT/6jrJ6jcZP/St1zFFB2YkfmDZY2++e/LADXrIqASbs8OEO88K
qZR35HnT5qcheMvDX2VHV/qhSgi0RyHBs8q+eWWsyH0mQ1sztTYGaMADkDhp3w7P
O5dEhIfs3p5z3tPVTgPEwwaIu7/sJzP8/+KQlgDdC08iR6VGPxGcI/sfIClvmcnr
uYGkXcKYPgZgR8Rm56apPCfmHLMYMyR01+k8tCyZzQTglrVYpuD7kaeUgMYJI67T
WR8JHPT5AhVXBu8GooB2VSI9HLbT3wEXNTafKyx/iUpu1Ozo0dgoDhb8NjymjymX
y+I6OfYKgDoJivFILUWOSrZGdPFOFR+Sq0wxPCieTTWy3dr8Tcb57gKg/6QSySoL
gC/rrSjo7TCOKxT1CJZtI6+JexfEESo6bg/irtHIfPfkYta6TAdFZvy1AkCgVtg6
lUHWP+Q2qyVQLpEyFATM69uYZ76dLPqwVVkhgsM1tBmoUCd3ma/zDZQwqMlw6zDm
3d8XZwRetixMZqNWjKdxq0Tg6uah8sBhlgPKA4ozfi9y5mS7bxsfBchyjYsM5FR5
gYPW/IbJOAhEkd5asi79wWrUlaEC5u+KWzxLaCHhn+ztRDzJeXC4J2LUT/wEjY5k
+8JLvUXV8QW6weHFdz+O8G4xiA3WE69WfvayYmCODZZhtm0Rts/xvF1+dK9ehkPF
k9E5htCsaZm5S6ZMgUYLwbGs52ga46XE3DTmI/XJkN91FCCWIz7SMCBTXA90LeAH
I9iOrrHEQZi25hDLdTsYqgUPKEQxHhNkhjd2kOwJkz0oDCNo0POyMpHpfh2Vwo6J
ludVuE2v9aGqWGvu2+AcPI612Yx5nGBeyFNZCxT4r3xr9hh/4zf/03+GRpU5vVWW
gwhsb4epRJWFVk4ZmtEbvknUNnTkUyfTltzS2iqU/d/i/JwC373WOb+Xp5voykM4
2pUqf6uyEmalK49eFV8oMPJxQGcFhZpjlCxiPNa55XAAHEmCtqazU121Y5hcvdeq
Rq5GgHgO1u3OiPHIhICHoMh+FNVDCTqQPqkgxK4eH2o9oQHzS7t/TniNHaEAuyFh
BkZ0F7LwtXC0yg5Y+bpY13KgsPO8m/TxuYongOBtxySjotZjnubxQT+MoSK9ONJQ
EecQTE+DBZ5whMnZjE6UfqacZcWJnta41S8kKpTwAyebmpToj94PZiuteVk+3kk5
QXCaipD1uc0OVIiUZqDfaniWqyQhlu3F0cyCqWbnKtiReb2huMIFGbEYXcb7aMw6
8GpTobWdhGfIT8nGy7ffntw+HKGBQYFEu/97ayqTfV1M1FhahwczIB2BEKj6CdTQ
Aw3bymPxHftz9LY9HwapBLAxJsGpepCW/UVDbvBIGJDOC70EIn0kwXHIqvQGIFAF
m1rHVzLVWk0Nc6IKek8ZIqhBvze5bnxHLXx9XfuASGLqrcblo5oB3jhJW604f6uW
szHEQG8wI4V8iKB58q8SNbdjKg9HOpcODjyS5v53ir2q56SNn3xdDhQFc3TkqjrR
6miVoYeU1Da7puWo3ZX7lE2pGnpplX5emVN5DZYdlYuCSTYf1VrZQjGVNLOVmhpj
P464OonDVe0/73HECCEGj9bg3AFhJ+c58AN8JjuLQg0ree6g/l4PVyRrn+/CjXi4
HV3ShNvzGdHFsaTqrz7wPvAUONE544X5FvJe9U0DYl1ZegFdvDx8NjzrR0J4YPM/
/uCX35t88SaMPWUeOafNxOWYHI0xPmduDdpUuQ1GlDJX9r+ngVDwp9D+F41zRf6Y
WTYX/tUa6yY+P9qt6nr7hLfyU/UpiLQOgCsjC5y8ozOeQVy6jWqnTDb26mhE3ixJ
PNvELtCkDcRRYIoZU4Olgmb+HkTL85XX3zovsJUBU4XvbZsADTX+ndCVV01v/wst
+dWARuwxh59DGUjLy53fKJnTwzj0PVHQT4izMnwFBpW+buDSLXz/bD0W16fm3o3A
KZ1aXB4a9AXsN/UrkAqQ+pBSxXntHAZ+/XAEGzh+WSFDkiDNNQ7wPCqL9ZKLvekg
vid2daRx59WRuiIlHNzo/Dgd4p3Dz43SZYanRL8OG/G84+/j+s/vNdHdWdqRimSC
IaiGI3ehOJ9BTcScv/q69H+br4vBZM4AuI2xMjpVZnVitY8fu/BxjzZ6AXibrtAa
K26CZHF7yfZY0x0gbV08+zekNp8M48Ct3dSlWasQFLN1/RQ5/irSOeTwLC0mI2Ey
fGbyY1achbBXHQID7gCoYynYv20ZevGPLzMjvlIv5Lv8s1twGcGQRPXDpLD3FiUQ
/6oeXxIO2Mh/f+/BGZ2MhTa3a6z9JtuTVxSoAfkMzqEgyJemcSDjRoB597ei8CSH
9fST6E4SX2sZC1BC5sekrfg7foGgGDOJn/LlkeLZaWT1Dc8JXj3bVN3i63exU9/+
2eHpyotq0fq6yC/GqRmPT9KMIRn0W2Ljt49drArsWtyUZoXJIKywW9M3veUphzCg
jSNdRRJy6d/enge5oMtseCMtnzAllGZk4mjtYiKMaD5lsUCszEln1S/FjSIx01iG
EfV4IGBRty4NdQXjLd/SceArAi7B2+rGDdjBd5YbFSeX2nS9DmBFXBUyTc0QkOdS
jUky1He7qUw2fAanAN2V7Rul5C2cAEoyQ67J7ntQxuzQD5AkL0wHcH3QOBKreiSt
RClS/ol8kxO1nnM7WM3jzXSSmusLLKp5O/tgaLUzVMx6gevaJ2yPOVzKjh+I9eVY
fwmS067h82dFVZ8obt7dPjF9yIeE1T5DVlRj7juhfGbo4tHsHpDzaB36oexHVU2y
0n19q3FfHkKk7pn7JIthozr05keRBiWhDEAN6880CKaVhO2mSdHCTTp9YrMwOs8o
GMc/X6S5rpbXafN5lfbOgSnDYRhUkn7buU4zWkxwyuezPQnWarK6KksRz48hUwKt
9J7uF2luLX1Lk8B53tdllgA9g0EOsdXfer0VbgDz2fb1eQ5zWAMec/WQjqeQ8fzf
PhDRx4ONQDMNMw/z6UxF57cpDQH3AWfdQKHU6i+YMl+h7G1cY4eLS+TemUdpid1F
nI2rMKb4UIAiUxfjivlfGqc0UzrCpMjskE93g21Xpwdqc+x73rze91SdEO95dseD
aPnFhNSGpSSensD/YO3tRhhu771vNEIl6I0UG/BhHKMIjCJXxJWjUP+LrCQvt5NC
Hg0qF80pAPtgrsaIKfl03wFK3dvRTpEy94LZx2zBBxYvnr3GjN7DAsIlO6MKng1E
ZrRPavegjuRM1HDTTSpPAQ4yrSb7Ww+yByDlA+Gx/nk2zAji3oIGdFHrDKnf8qF5
WHcpOJ4AsFqnm7fIHjGUcjstnyw0+/4XVY8mplkoEph6LkAhK9kOW9McVu78WvM0
9Tg2TDVpAY4Z0fgY22Cjx/kM5WcFQ5Du09MittpiQXkCbPpuXYD9r3jVpgHYSbLT
rfxt9WVirjK/B1I/M2XGUBNcI8/4xYV4sfVEh2u/Z3oKBHw8pqN4YJNSBbBEkeAH
fjUlE+khxxCScQoskG4tN84ny6K0kNjUQO3nQsA+By7jg5Tyz8gL7YwRw7O617OQ
6QmWL/helN8hb51KgVnT0qmJpC+YmBg5uIR2JCjFGw+ET0bs1w7qV1HeLCFPEKsa
od4CUslkLcEyT6B8ZxLxqWEynpurTdq+iFTnGNLb2gz9LEUoirr8VqW1qjiLb8Jt
yruFW22i0HOFVV+LabvxRU9DJdtWWZyXkGi/RiUJ8bufrF49yQi0vh1K3b3J8+VX
DVUJTFYJ1O127/NS04LAjdrRgpFv50CrJfaLDEp7Vi+k0jGME+lFAVbmQWkx1KWS
9jGg8e6PddPQ+vxdiNDfNCbF//uq2Bhwzuk4x5EAtOThKSkjT+4C6qic1dozoxBG
vrwTGEFIEvxsrrbwgqwc18QjxYXB5llwZnGm5Hgi6+XeprNtfA7ZoDFkkrctNEFz
0CLuUp/P8im8QLvCQNnxP93f2w7n2TtF7wFP7jr8NZLslHF+H+Z57MtJqNTDSpKv
sWig8qbxnNIjnYHU+rE18LmwgTZDGmppG62ql9JsGOQttjDo1QtH3qm/L1IqN2N2
00QXPKFvhe0ld13VPXKrzpuNz9YwBf6o3vFYl5LTXl0Qp6decWYlX8Cl4QZtLA8J
IfzxVxVc7T7K4ejQyCepBAoQd1IAhQ4h1eO87oevPjz6f3RGNwLkz/uQXJZ6sKlW
dE4DiTqkW7T5EcdrlTC1ployLrp094nMSv4dqejWWxVwPHn9VYgk2bDWvtnEc6GF
DR9eL4Mmu4fNHiFNWMFS9fXw4tcrVLEHYOpLoWUwrIAHa3DnLXlx2THmaUhsuArF
gj3eVWgQhon6H2e+aktqaJdTrN4TZvymMGJ96mex7A7uNtNVRUIJb7ZQWCy4UJfi
U4eoim60x3R16vGkIkF/f9ZO5gms7ApfPHTyi/KNKrPBgoIDbxbLQaaQHwbx/zea
DBC9ZP4pJQILYX6gqP103YphvzIT7iPAwYB1mwjhPIotu+1BQzwXgar1Zd/cAO1E
1slVEhp0+mTtfhB0agg5bs3iGzwvdgVGqrEoWTE/K9mcDeqVtYi2rieXu9vWb+/Y
HnTVgJHtDf5hNAFjHdQJVl1M3kfx30cf32DzB05Ndn/hNBvbvQnKlN+4sJvKmEz6
X7XI+i6dlxjgZX17EW2mX6ZJ1/XCveWlvBmIPCURh1tNVv7XhdlfYMmf7+8M204r
DJFUcT6Hap9p/eGp76pEkFTMvD6tvZtzkovBGkonuafUwuerSlNRCZ/HQn9DRgKj
obaukVhQoG6Zo52k/Zl85exg6dYuuG9sm+jIwPcweVNA2PfNU5VTHEUEifvGry0t
LK0e+cw1RJNhhi4589U1OLDHW+bBRtCvpjdmKhezkC9oh5vA7TRHGHyqn5s30WGa
UDQjJGGCNrHO44pgaIHLi/IrHvIOVRwYCWU5i0Tun5LrVxHh+HBbDlIAYdp+SGhc
9k92o90AVmiZ2BHuU1S5Ypei8k+3+yjfcWEFal7JmZYUL5Dbj1B4mHqyXLhbZ9Em
5X+J63fSoRezm0AZ03FqtLKDhueIl6xTENRA2uOIaR6PTFrgGKRxM6TRH9qZ4PLh
8bK9seiva5okJmxXWjMDZwCKVYh7SUVNcPVrAxY6HSjDSxdIXEdPr9UmoHH62B8g
owGmEF5A3njdqd5sL09x7BcDrdZoDXBAOMUNqQTYON5rz4LOM2lJ8NcxsIgHmeAw
PKi9hwHVbFt1KRMmOnDUzQ6diRVr9hDqjiiibRFOiEeC4WuZDbnvaiAop4cTGoc+
b5lqbkc94Ok8wtnhPvlyzbJtjdKAbEC7zLA1SVwOvN5e4/ABmap5au6gejUmoIB1
7LhR+aL0AHGNIEe0JOqhrxxptJaqHFvhhSNLMXecLrx9Wpo7fbQDeWqWO/46tAM8
N2XFK0lC5/4oowiPewTnYIDayscv05POygzq38pWEhWlKv82hBmwUw/aIulX+ZxB
MyrduTywp0gCjMyt/IPtpD0gpuDPoTuvaMKg9TBb4sk8llwszRWzaLFJV70xp8VF
xuXl3FU6HZLWmY7yIGJWEEbjzPqlZWuV2sRRna6ghBGM87TBXFEbZf4U8Dnb7H82
St3d7JtQKsFPLoxA2RLX/6V1AJvMv5rcOUMqE9+2tqosno92IhU2OcfBx4BB91Bg
hUn2VemGwA1IrZIaf4Fk7PGueXhg0g1FAj7J7J1MtoJJ3OgcCSj0131zKmXfbZ5A
wDzUC0rc1Ba6EKeVJaqhsTTkVYjHxmoc+e2gIwAJ28vClBSirMsN3/DZ8j6KvdFJ
Orke67QzrYlCOcssawAzL3oULXUYL97ChSxTNOr/6QEGvhYaMvbWA/gZnvD6eAAe
qUpfaMFpaknksf68xyE2yfLgASZalM4IDcJ6DbBPzTT5+0G5rLWwEOV7TjiXgDwk
3GQaqKK3YSH5vr0RDCGGwAl3hWeZxNlhku0p05wBQmV57+TcLNmrr5qnbiUSh5n1
Q0AMDgzHMaHlp052YqrJ8tkmHnpqM7N0f7XBZRBKO+ltHHEMywoNlyWKmxAmmtm5
OG6GM+E2GfYAy8/pbVNJXw4p9a3bLKLR4Vp5VAw8YKKm8DT07443iXWHl4/rmUv4
DV94ExEaDx5FPqLqxOiwPagJYHkHfrk4mBpQ5eJD9upeBlIZC6RQGFtqMEaN6C1I
3pxiHrBNn8gQPjh4R9fk96lGWAC2knOBkYskp0SmryskVlouODhwern4tYTiN+L4
ZvYOUkQFbiLiIJf+a5r4KcdL1qHLH+mC0Jn4k10+Iz/MDoTohxP+P1gh4CpR6w0C
26mmQjsaQC57J3ShNkdhFTCSB8e1OZU0SdbmP5PfoyyNJGakL5LNRRdnzJYsj9Dy
urBDdd6IprDZIN5m5Yb8q3y3Q8fXWwbPCtSge+bEGYSClaKvSvoy4kOuDKGaj5Bz
hYtGz8EhHBka124g6dG8L/QJN5eaoJeVb17cY+ffkkkkMSm6PENhhKZzopcdJVIk
N55SfZn5zJnxCx5huNhzCJWo2JFh8RTsofut83MOcyJADkJvuB9S7SIIcXLGZqOg
fAFcT9TUZvPab4YNIYpqyPpbLYPkX08uZ/nWLibFAoDT1J2WzWlN2U0beNDLkrgt
Zl2TnjHcHRFehROwvQI9n8kHyf54jiV45zZ+weUnvkwESjq4CsGzajbIRWVmg/hp
9ViZRPFFsjz6XagqYqEx6FbTecVE7v22TLCXAZfQiRRB03oaeICR0joOHdtJdYfo
eWQtmFmhOBWRpRm8UMKuZIpQ+oy2WASBIFjatzpCpCuOSld1X2B/+pIhN1++ahQJ
YnE2JzcuKi/FyBeRI1Zd4a3J72QVyRCLux0kkPs5dWfTDz6mxI52hR7/yVyyHvCP
wZDvcHuJZbgMhJUGoue9ED6FeHD0cBWs+W32pxTV9p4QYLn9Kb6JKWLuAi9Fs02W
2/CPd2mutrOV8UjGjq8DVFDE7KkpVDX7LYnKPNRJMHUjqpXJPRcXI494koWksGdd
+prjVFgVNKyb/pDaLZXsd2kWJDIIdydsk8oa2X2FLCNPjniR/iEyYzdre/QqAWde
cR20IiV3wyzxDznWdxLWcRu15GVwP1goO9ThCkjbOUWepIkn6hqdhQU+laexkuQT
pAbF0KplHNxSlsUPt3Q8bBDE7opvQtF5V2TLMs6v+N6GQkqw1i+yqb7zsq2SNPcB
kohaNFx4eIfWTpaxmsM4djjLiTWH8BHCDQUaW38WY538H5j7nuy1hqDUmnDncrAS
RpGNUQ76kptk4pIzLW0gwWDqeaMpQJ6FdzQtUXg+5fFLWY2b7oM3GG0s+bg2Y4Fu
fyU5e5xVpl/IaiInT30FKvNSAsRWdyRTLCJpIXDs9bMGL5GDqgjnDXv8AlNuea0X
JBr+dxz97hm7f0dokkSyXx0yC3c0ixZOTuo+YUQcdzeBMKxk68EM4GUfUIa9daSP
uzYNfG6RVW/E3doewWqI4g+5+P3JAq+uD+TvNtcbLVe38xTyIiAicy9akULGY6Nr
MQPk7TsEDOYax6MVViGZ4kTbRtHihj+8qO7rqN9aYLD5KnnsdTOiFd6Uu3aCBjdg
31CPyQGuXrCpTU7TI7PwyZ2PI6TOwzdQflW+NsP+1pFheVbqKdL5ywFwv2oslMOp
fxHs2hggafw7EyEH6PStM6idqtwPrW1QqvtluqTG4ovZ3UqTssILHMFsbec66he4
gviSXK8YhM+sV1y9MnH9SS8mTfKVvXNOVyETnhLCZllNgvPnbCd9CKLyssJ/frPU
gAEIUKdWTWHA0UQPKzio1ag2WCnY+TJMD75PiQ3kzSISa5Xal8MI5ba9D+neAPow
UEDyFNgJcYuwFiNcj0LYPdIVRHXwqUjaKVqH+gfd9OCTJREPbWpKyF5DHz4GJYIr
bppURfX6vEUinhZcBeFOpbcF78anSaFAJpBKeO3c6wKSF2hSLMssxAhYu1ZOsCcg
Z3WozHl80e2UEFUphMGLRH8kAYprjOG4TKBkiqxa8GW4oIPVYqTAQZpBSTgrLNGy
B4oWa7vVcjjT0P2aChXV3n63jiyS3FIvpw1kbJTx22/P5a4TwxxnBHQ43bKIEuC3
MBqDoLJUIYSeGfffcDtRF9C859OqR4j5aT3922EK7TQcV6QwsryggBqP+Sgiuvb3
izGo1sZxmEKG7uKrPmcus4NNNvrVo+AyDPulof8QcU4lx5uIBVhUflxtfdWIRCf6
ufVvewEKut0m+VPnhnhGKyaxLNaqT8oq1pUQ94T/T/0knB7es2+4ggujic4jcsDC
DeDCMfQ5lDj/bIE16EqBXI/38Y1HSqSgDXxs6ADbIO0L/5v97uZBLZwDIBEhRDcG
7YuUlm4yBT+tow/tOKmoQzY/CSkrGtlsSdI+0mwob+fGFKzxwdUmPySpPft+8IRW
NpLdERAW7bBXH9TjsP34mEttGaRWbaFroDo3sXY7+3EZl19MBWC0xdtC0kZaR7qN
WnMk2D3m/4zNA/JWcpBLv2nkPYpYaAhfears6h+4zX4FDTUGb1D23ynpg+Srm9hX
i11JT6K+Smq5cPUaJFqu1/WbB83NQ1uS7tdAiWKpPvrO9/DGsLOvqBRV+mXFHMzs
cjV23D9KFuOmf2vhjbZZpn22u+SS41oCIwj3trHqZJ1wip3EAHnlS9UdBnksRumD
O2/0fS6a7e+b4OvcHtcKLoYoF5QPI+MUmQngkKJvygLTbF48YIq4ZDpflgoo3dC2
S/yiEiS8b3JB3lZ1eWvUn/keQBtvqsqfy7tPbgy/rR9x7XiB9Yt1k92ccjacbHFF
2RSj24BfnOTjlE8bkDArcueRw3rO7kiU9Z9eMDKDz7uJEohlkVgnjYft5+vChnfi
X17S73mPQIhF6az0xwxWNLn/XpMxq9ssyI6fCGvs9BBPyPa56RdhaYxaLW+uDA2X
X+dDniWRbTViYBlmOZ2+2Rgq1dwi7BjyJVJfdf0ZDoe+h9uP5IJ1nL/pUesiOP1a
dJuFV1s8P1k8QhDUJPgFMI4X6I9hEL5Sa7ngimkprnVa9vHaUlO6vPlptwnMzB9U
sI/FrBxv9sCDa9XmSvY/5HH3VJjQsBqbSYu74Qa4I+ZqCTvhE0xaiDBJhw7x+JO9
gWhKIXY5NDcQATjvx5V4stxiWYfuCjiGa9ROmTeTZI6HTwhnPQ1Zn097YG3xp1em
sdd62QvfpjIT0zqUIQpW2qc8xzd+73/ko2eTLUMGfFAZMZiPuGZxQEI7WBuX3TfB
E2pOz3DT1nvCLGP8/RU1dwYEOD48x/cR+R7uDWxYc74gdyLxqTnjiG+Dov0BevGY
YvSJw751Q3xIit4VLde/HTbSzG1vwB726xPpbscC0bTFOPd9jMiO0tAnyaiZa8Ni
WlTgMQipir+lSno3h4l6KWmXiI33f5xwVqgvEPFfgOizFxd01J8eYYtYmyCNhIn8
24YM5gjEJHGb72TIO4FcKJpuc3njBB7pOnsxTQg+G5kOzqPDxZrZ6Hriw4XNuQFA
Hji4zSrN4jqlzw4MqkO5KUQOaJyQvQEReO5NlfMxy3+NwrjHIXmynwwlZawxcRdp
72ObZ9rdurhTsb0IFOpq1ofalK5phxtUUWmV3hCtEEJJ8mKjLEgaWvYqsydP4up8
lNprKk/vF8VoOpQg9Evi8WsZqLrGo5pfrVEhy/MdZp0K3Ir4Ksdek+467vFnHILj
/A63p6lUuW+13sTicbnhxB1nF20n5RdmPE8jUndur14LRGKdrsgDE8LF9UqWdXz7
7TUCm6/ZG0/ZG5RQ8ZI/RO4NPGVfuy9APjZEJSIxcGrAjHNbL6K1XaT73ml2xp6F
zNxGYJp3Mwv7+3ttyHyzJjjFJQKGxKk+Jr2u6P//4VdHlqlus5wIucxCjH3hbw9y
OLHbMVieBy7S0IEN0y1w4pixpfkIkcrTDoXpKpcNJQR9k5aKhTUV51ki1yE/BSFU
1XHnKuLdfHpiRj0Pmjp+7xhc+lL1HboHVLQHy4L5fBqHgYQdSIOLXZeNklI6liEh
+obYmO+UqXPEl6v2Lils3KWHwKwVKGAs/Ndynh1iQc59cKstezDP9dbz8SDYXC5L
sPGbvm763oKXkEbeEMuTttcgII0SoY2hDB9DqxdxV+IY7PEtbjdG9sNlAsv3RNnX
30xuv7StJ7xeN50f1Epgso8K618ZAFWqRlKIjQBlllnVfVwELZvv2OnlN9nleiYy
qIfmMX+9tH3tbWJIY12m+1huxYbdz0TDBdOumRAnJBys7u0IQvVZe/SKddNb6L+/
oLvJ9GYQK/hY7swOYirJLXnl+zX8CBDpgM5aWgLhyZae72DWZRNNOUcxhyREwrB6
Jwjfb1BFLtKCmglPL7LT04qVWXwETledo6WPehkLFloIYmncnKRQblQXU0+GRTIV
oC0iAEltqFSHMu27e6C6BQZ2PvdZuePIxdvNiLW0FUfI6tgUZyWGvhJ2sd35iDPU
+pEEeAWHp8mbWs5pvfH2YgXck7dzjSI/l3A2tNfCdSbI8v4xKJv4eFQ2JrYJTUCk
Oac4TPSOn7RswASKli1HIbEwfKJ5MoRDGq0so1D3wVqBagshXfVvBlbz/WuPDRLy
ho/4aWwnJMlUCyIb+PtC2rfYCyVYCiHTHlWklpolBEPR6UGuzMNuKAwPALk6b/PU
kGO+FnCJFaYIO7y/qmL1i7GCHNnoyT9vW0T5x0bJyCcUJHZCuIx8VYlxEvY9Kv2V
4I0MIEymBqCAuROgcbHq2VsBkzT+F/OSeSH9Ba+Zu1uUS6HHvjMLvDjM+sJp9Z2h
JToEcnWHwkQW3gQ4974CFEkfU1afl6XQtjIzskH93p5kXyvXASuD8ojfYIfc515K
cybdmu8oD283Sh8/XoonyHSvvUnyFK6witL0ZswIpwDNNnPKnsYFSKb8FzlioMBT
y+O6RkR1EJ75BFhEDf5RsYflQUciJnF5owa0sKOC5/5ZBHjCPvEGEQBWj+06NxAl
cfEf6g2XHe+c6BPgsB4dtRjnS3sDzaC9fIUiqIKNwCjbm+Ulnbvb+FePCHE7rULg
DWEEYoPG0WQxTBa4n98cTjUqlguE6IC1Lw531nSEwryQ8mFloY1y+hUy3AZ/0zFH
6q4fVYl6Ui7TPFD6RrWRC4PvgmY6HuGmZz+vOwQqRfKXk0WzGpnzqLURTv/9Wk4F
33yJeYJtFGFcLKcLqzypxjzKtPfC3RBpsHc49lvSorxS79zORvfdliXEeD7Fzjef
itnh58CcjE0hz2NIAgsmUCm4yjsk7Ib9644O3E8KWlE4GRdKtbTy42w9WDRzB1NW
zf2MYp0UGuu35iZpllIrkogHvJ737sDa4NdN8KR2U5EFPS2XPX+LT2PKtilOax2q
wj11A0M8ZkyOPiX5eG21YWF1HaVs7yGGhTGWRLZq3lT2RaNiOr2aZkctaWJGOxBW
hzD4qGiXI/ZrAx3pD+rYh975jJADvg5aFFTE2Tk3kLLi4uLJ9lJaa3ZXhJZ+fe7J
VNZF6mmd4Ep1zQooarlRhuq7A6Q0qZ2QeD5Onk/sZ6w+BnWe+6WCFz/TM5AYb2Yi
ZKFU4NYdYffXb06zJrByZf8gg9JAjnv8AdMei1QfBDpoN8n4G2bwjJyiJZbudbXa
iPSJ8u1oYpTanI7muqJo1Vqgx4Wm8HabRiXV46gr+u/h7kQcpRzBYEz8F6Fv93pv
01AU4QlilhDoOPH/W86CTzOwyNpkPUljfp67KE0gY2HQWnJyuFYwtzeBbVCI/XZX
I29GhKoW0NEL4poxIrXNk5ksYZM6S7Ya315UZ4i8/8AvtoRF5TTVteWNb96JHHxm
t+yqYjgpVF/7l8c/hOvgyxXMXYiJQGu9PLRWKOF6iMVIprUcwbXC3mFJfPrzRazl
AeNA3lBhYeAHeHY9oJMYnCbpxCxh7R6WHnYLfGwhhMxgmmkJJmZl5BvmUKwjBoCI
D41GRGIwDkcPmYWjfMYm53ndJ4rRynb6vWU7pE4DJK4+MSIo75iBXxxmzHFbfOJ0
7OUblWh8Wia5ArrNOaib/sueqNN7MP/xGmHyfWI11g8CSloBiMF7udeRCUzwVpaY
EHpQgCGSaJOgFCDpRd9/cOV6qfXN+A5bQxTK9tM1FlurVamaDRo7uHicPd6i60zy
YM33WwhFYioS30wu93iIPy8MSdE/h7qdc5kUKMCMySagiMYm+XvlPImkSDULj7zG
Uw4QroLu23N92B4C/STbiqa5EGWMF9yPa6OKXRXV2uutAxDd3FCrRXuADk8CA27w
dfberYK8lerUO/W7UHlrSJrpNcQASc9rfbQ4iVLhfFe/jRJqkRWMXQC7+qKsNYiu
vIQpjfKzc6PiXLKw+/okk4vmIuJHddUSTSqfIIBtCu9qLNzUJAiWgdl8xCKhtZHr
ii+NuCJUam3NLW+U7ozVyxWbhhlKTujBurqf73OxgfnAOm0UYMpLzCGgg7rxymLE
6+GW/T53sFMFpup0CRMmMXNc9tTkQsg2clnZYaOoB/yWsC5tg8Yx0G0svkLOHfFV
0TtLB2Xr9cZLwSp9taDEg8OCGL73jYuIPOkuFZ/g588j6FA0/FkgZenp+cJOK3Wo
xOYm6OrBXZQSX2m/pIrbOEhzqtzRkMGMikR3JHFzJfIqP+qjMaoDXiUvf/TaGMzt
Pj/iEoOhq9m9dTfsIPjpNWfSgqgXp3NdGtdq9eer+NSjoVIw8RO3iwASbTFbNUC2
b+y97cBb+4dG6JCy/bigBu9Zo4vVREZsFv94/LyU+oNUZqKFC6QreZt7BnAdBPB6
PwqatQ544SKpJPBgSyXVLB7frJ2F6onbHUxyOHCM2xLMCEKa2K+/Kt/DqKiJI71s
S4xSZitPCp/NmdD6xmUhoseUAOa7WaGpRiptj9hUVZYwG6jJt9l4jxh9ZtmU5mki
5ocf7UHQnahmPCzuIhLFBL0GydWjc/Q3MuhjX35WK1kV1b04unEZx9kiTmnQt4Jr
XGkMCRLnwueaoxJvBWO4rDECjpSMPvArtYw3iEqUA2h8Sf0MMS8kiQNyNnL+4cNV
64exFgznXBu7S6KIAWTWavpiDE1sznUmDHH6+ZiRUNv1j68dwDaD0Q7040X49oVM
9Pvz4YeI+1jW2MfV2s8b8LgffMua3Ogob2vNhsdESgXgHafKgak06fsAaTHXHDzQ
/ALZy2r+tF1dLM3rEmXCKv1lvlD34UUa+Yz5t+Wr+XeKNyO4u2e3M4ZmYdsg5imW
HJKL2ansYx0Whpvaqq+rsgwx5hxr7VTlPxmDOrDEfaEpqugMhwpNce5l+lGjnZrn
CCty09VBVPdHmfm/qOVISO/E1Pz94mGaRJR3tiJ9/jTT8O/184COEItf9m78EgGV
mSODBG0HlJqfx0iLyOPBxAgClb1sAvWX42+/bKSoWFDiUrlJvYxw0QghP2IpO+oJ
CjqLDTwfWxurBKXJsreLAW+0rrzk73120RefQLKnQRTuEDHcwr2/EOYGNaiZG4bj
xYsuDTzikUUmhax+J8jCd4bUpxQuiOpfpjiHT7pxq6OzGGxfX/cb5rBfcFKXsAWJ
NljpoatzKDwpNXyF5HRMdV2E/2Y6WtNOAzMPGXp9G+4txGC8RTGUQ6oXPW7OgnrF
Ii/UnC3PWEj1LA+xH9gRmvayfxs2SsrAj/cndopN+srUXbDtAEyyX8LD0aQI96wA
pZBR2bpFn5LloKUoqRV72JSwWHHUenosHaXSyicdnXVMTJDU8Fxz+zSQT4qFvbXO
IVDwgnCyBqtz8zjy/ch7zhLRln8Fj1ZxD0B94U8aww4Qq4qZVojuusvVIZVTt+Xp
P71D4FtsOTmhZPrRT62q39A5+oXPVKm1WoOb3PWCiOoY2FZysxg8aeTd8jzx/eVP
p5s7PstepApi+c4iWmg+0XFWXgnJdI8Ra5Y3fPvzuuWXOTZ1Ah9ZoB2N6tCooGyO
kVhTxwAddTzAVrqqRyvrmxkzEby3qhlNBHV0c3ytLRyztviEiClVPOv0xz/2OAHa
ksDkA8yhalNWxjKJEZE6DV86Jxgqm+k2MYIYXP4Ti+KZf7DhSzXuHxLd7mni89uH
jREGqWARpfZnpMeISM7GMGOmgzeN53DRl1tG8ZpaAhS8MFIOyjw4ayDZOjQ2gKXp
jARdkA+mgnpHdXb103dEwoM4PFJkRweB1IXAT14rwZ30aM4HUgJCYDhZNbrtobAp
SoEyoQnJR2LNov3fkYIFn2grqih3JcbbQmTdwILRU3jZVe9o+7hA6pa/hn8MFl69
Neq2mYHQZUfusObIidPZhZuGlJJs/BuR3Qr0vJXVazUFKCR26DhIkZxrqDz9VGNC
LyVeG6P/GpCbu3jFnSOolgQQ4kkqCOBoVQ/ca6SwnDqmJ3Q141UaOb6FVsaBnyvd
NrPXvHrePmr8bhZZQfLpeXgyijFy7sE7/FrAIwGRynoo66ltpnRoKZxkRoK+D1cX
Bi4uc4d8v/lHXcer8TpaqFQcCvIeKp0bmIcME8WBiu2RGj9p94iAnwUdLG7DSWuJ
MRphdegs6MZuvX8CVSsfDRZ5WSADIU9LxLVc+aSUTB+NOL/B4beC+PazRcAtDzoa
GKNqn0nodcfrB/7EAOlsmgEO/UEOT1uHXyk+JmVbVXtu4gbIdzjcFtvsLmuW+4ri
OVpmduAMCUgl9IMB8Rt6PvaYGJ/V9HP5T2zVXcspBJ7uSFLyldzqhmdYsrFJJfdh
bnYlhCiktCB13/OGfUzVGC2AyGPs4tf6adgWHtbvzeblCm/zz6TG5NeXDFd2ZF2J
Yl8Ln2JnuUXjbrtfgJ3GQyEEhjEInDx/qW0yQyAyjmCiCCnBrBVO9VtDR/BBsCbW
jEy1CwforQ1Lg1A14Eza9vh7ABh3As8qjxvFATMADglPAhL+4FMghvyBD4Q7FHyF
euSTpUO1GITWpUMav4E3fYoAFJ2ChuTPc7bOIzO4fs+kYq1TUJl0ULrqA/Ktm+HF
wJ5HcdnDxPXYLOr7wNSk3wwKq8SvTgkmtZtW56Dy0LnQkP+g68XhfuL+BD5nEVg7
kg+f7h1EMOVWziZ/mLThuM7VWEiAvSrt5Sz8Y3MErrRfRzJrMJ4ceenJxdWf5KEX
LyEB1WUX0oPfDOZE4xAevBAj+DBaNE+1D7wVTbroNB1n+e2+TKWqeYc3bW6cpL+N
l3pWS9TNCDHaKTU+wvX/UjTtjfjXDGzr1D8DDQviwb7E7Gm6YEW3q+NdonyMsoE4
lrwp5uYrnIgdFRLFfWy9vXMNs4rP20jmrhcpO/UoAtkCWt4MMe+CjUbrbDb8Be45
PnzhdzOQRZ4OAIQPX3j3RKSrircHdH81eGmgci7OjUHVzD0NqsRXMH8GXzGU1DJe
pGfWxvCHUznnNjNK3BCuvpRUX/WNGmlUrkwbxJwLYxwdO6eY7ZCyRQGXvf7rbf7P
rZXYpkB3vX4kkoXuxemdqiTvzzWApfIjPe7Zu7pQ2vgf5LszXPgJmtrgr7pPSuww
k6uxk0uxHx6aYZOqdV9GTLxGG/Vu7uLWV/r8Dr6exqYHZg7YE3/GgNKJ3VKO69nP
KktpAtXct4K7wAqXjmfSre8lYS+Dzlvk7U4deQXjku6A6CmFoS4/DH506G4jtHmT
z7uahmEDtyhM9j7zCkjbC8o2lbQQ1+79GCnlSAY4J3zRvynUePFtKGZGrRkDtCno
KghEX4J5ba8xvfpol7l59RoNiIx63bAJCSvRuqCbolOxSO2TUX2fqU5wRCqYYqDK
VE+tmHk65TE5sz7Gj6fGOLOhzBYovbFeHW53FiQu3biXT/lPFkLuwgOhxgk+cMyN
Uwd+SJI3t7Uc3aKl2YZP8b42MbIF/9GBF/octf9uIwVTV94o78gXxGkOHu4CwjLt
NtJzrp6Sba6Q7LlaVN0O9FmHhs5Mv1nSMG9qJgm22ZkI6JnG63XcGJYcRb9KwwsC
dnGnXrWvxQK0Zj5kVyX1smtPP+yw7gBf72KA1uhra3+4yFvOd26CKI4oCSA52zl0
QvCmZuyTpmSRHCLYyXLH9lnmiC1gDjmVnSTM1bj95b5uz0+LOmJiUPgFP5XShjjX
fjYyr2Gfr4hLn99GmzI8oVCYfewjALBsMbTvCMmHjMt3pUTSyg+OWEta4xZlZdtW
2em+LT8NX6nKkdueX2qpltUH8p3cWTw3H28pG20OCH+jNpq7JLbB+RvJJcLgAkZQ
dtdqQ770sub7ZYXiRFnwg/gycIJuQfpYCjq/qmuQy3dD0XCmQvQ2/VRfcHy8ixUS
KsOJxNtLyNBfvTKByCYGv/K0mzJjrc6Y9kH/M1eAITEEgPVdkpsdsG9KkqhgmlcL
spyS1BF3H99eViqc2DMnQw/ZudM+8rMDTv80RyLfhaiguSHqmGDcpiSXrv6U+n5m
Sx917IL4zAI43SElSo855eYF+R9irXnTN5y+g8pVLVoje0j8aGhp/W4pErm5MFx2
HbixQjid132hzCY6towbhurfT0E2FHvcyOrNE4ZxM6op8C462Jl4jAaVzUEW9Cgx
F9H9DoFAEcRTc0zfudriAZk5s5IIJI64SuydBWkDndDEZma3G7oKEA4CNL/hamHT
vDTDoDhKZPPNDSa/Yeh+whH/Og1A580oeLIQ+fdL1umRGcOG/UPsKO/UT1Xm0SCZ
WJGhYU+RY+htVDmBr99vGRI2YCBz+n1ApkT3Ru2q/M8cJzxQPqhxYiEEFgPHUISl
hQpkDBVIac3+fpgaIzL/LFIyyna3/ubkEhQdL+V4ysyNKz6WknNTTfplxCDbAxiz
mDnSHEXxp5k6jL7/krHdByRvYzNXVS2Y7jmy9OoSmEONNWQNLBlW/VDZBpi0H+21
SrS9jNmRtJMCT1ZJpKsO4ti5BI/dv9lb7SGyLggadiWgaEO6d7HrFjjReUlnVkE2
hE+l4R5bu0R+Jy3prkU1oAyHVgCE4W4V+Y5sfRqJ78m3VfXrtp7gRzLtj8G21mpS
wO7FztaViHS2tXHgh1iobCr2BkYXDtKHocJgf4ViLDFrD5Qa6YElHjZ9B+uCBBO5
cHGT13yxOdrzext4jbQVqmZSBAgt2AtGb1pPNRtIPsQO5KYbT53RxFUA8B16DMYp
os6O13/7X9fgEYZlSX9xuiWVqsNu/hiY5YfI1boWE2l7c0KCmbFpli4cIwuOnXcP
/tcCpN0dArT+Iasysh9ur6DyZh3cC00kYQCU1V+DGjveTpKpsZqVMBb6Kh4gS601
29izGF/yryVWJKwj02T1xyAt4vRxZP3CicV6VEQu3520cegEMOJd/fMesmX/gCjR
5xCkZrFwq+6Yp6AePHHzF7/XKV0fNDvBS4a/b+8I3scTln//w+iqg+4XCuP6huuu
M73hNd/WATFW1Ij1av3nCa3NYeZgSAa+cJy2ZQg3WEw/230qbr4BkBihsfpWillm
wceXaKz1L2a/GXrGEwNe4vOa7Wo8Zp0CJUkCG5xzKjXKaebzseA/7wmEYcbTH3s9
0cKDv+XcqOmko1/RzcG9VDo2FnksEJVOtqPZKhCbW8ABgPnrVLaW80CeKqiW00P4
6ep2bdxEOR1XFdPKh3GL4u5/XtxUYtXxv570J8QggHO4Xks1zliKhl5f4ydB27/L
mACJAt3+FgduEmoCOTBFrH2hnjOO8CgmU+456/g8sE5pvctU3IBbwRicaEa9gaO3
wGMBX82GpQFsgzsAWfw9dLdEjb6vs+OGgI8yzinOMOSikxRFfgB5++3jDGHR3pNp
S3PNPfGGIpeNDZCgDhPAWGoFc/HuFU0HAq429Qdt/RdzBc9vTBqglwK5JElqy9q6
IBIAv4yiERqJl0Cyj9xqB8MivFaATgT33OHmllWnDgqqx4jGA6cdZZrVChU+8RaT
8dLOhflMa09aAwu47LKB9ATcDX7aUkzx2SMHbZmlFXZP0EgIoY6toOIeOTM4PsU8
NN5VI4K5uGPLUzxcIADJYVEY/U0GpJIJ/pMgmZgf2DgCe/UKVru1/wfd5sX9jsOz
RHDp8W1+fUo0fFDwCi9QduVjaiBM+vYfjzCMhd/YimFy+96L8R64mGGxMxBzxE+j
7jCW1sBKv+yUM4lED1sbYcxmWjFXO+9R1iPNVmfmPbF92ot94PxVNSHh18SBjBmb
n8kkdCobRc2+ebPNc1F+y9Ytd/nuxpc7n+/Hb2hCTNjFppi1r/rcZcgufHuvRMz4
k/2NcmdhchuJu1dgg/Z/LsVoM28kU644MWbWzdrI5xcAhKEMBn/iSgTD0Pn1vjOt
RBDL9RHWg251qC85l86VZLZgNj9XjmnfNKC8HACc0y66zlDg9/l4QPGFk8dOKsyR
2rco/yN3PZYhElI9okyg5KmczACWyWz27zvpc6C4iseUpOGH/9bGhahSoInRPtuY
NjcQ3Fbn83d2FfRAigY6H3D6/Kg0wGwU4eFh3w2kR7IrrbrOOavKnU3J0UKVBBRf
xT5Nn47WZ1thZ5YYTx9z+WmbPYSeMyTVuTEWsDvBxwn0jDfY5n0UQfaCk4CPD5dt
fVaUlLxuD+9fuGrit00X/G4bRBpCSB1w3grnRkoXk4r6FXt/emkpKf3MZ65x57TV
EMhkwBdLbq/imJ5unmTkhBsauTba9lV757kmHYP1lPYg5DbAtadBh81mkvhEr2w3
`protect end_protected