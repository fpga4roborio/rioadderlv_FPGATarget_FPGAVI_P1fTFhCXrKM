`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
ddtXksX2+yylW5zu6QL2Lhnb2d1sD00763mmSITNX595NcHTEkwn0zB1Dry37fOW
FufOhVzEJp80NC5qZ/+F0Vk7Ik02dIR0elf3clrjeJRK85K4e3Hoo4xn7YbFUIms
l/8VZSb14+JVGURjfswrIyCUotIzlzVYZ6gzoZwDXIi5gQIBf/gI+KxNXPaKV+PQ
Ufys/12rjO6aI/pPlqSm0hCvftmBcnezN2hk1UeXgOIuKZnogjOsf0iJVX2aOOWE
6pD/psybjbnsNB6kH5uFTA5frkzIzkzl5d9+YDm9OyC+k84E83I/7/j+rk4L2dah
QJOvksSIzN867/4Qt8qYTQ==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="MvBXkzurAa5VTw+1JJ70nePUfoQXBvZOku/SMmg4TwQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
oRtzZL4VJ4iwysPsC8SXYCzXS8Fw2gtZTOskLcDV+1B9Nzn1zTyNtlo6lNICRmmK
ZRVu2BmCc2G+fmzynYlNTnSa7C0Cuel6FYpxCBlOuk3OF2tzAmLAuDyOH3Z1Yjzk
a0aHuoCdIRKv7BrZCdALt03JeUmXKPdOmIlkVGFl8yw=
`protect rights_digest_method = "sha256"
`protect end_toolblock="Jn9CQpRhJt4rnzZPRk+dOpzAubz7omckX1MrFd4p81o="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 17072 )
`protect data_block
gD6l00tciPUa6pDNTk/+tzLxvdHE2s3DQL3/JqqujQBC/Ei+vcAB8wM3doqg5vTg
mdfn9XB1bLOis2CVSfu295W2DNwHfMSTc/8BhCDRnTlLIX0UCJs9Za0+LoM0rMrV
T7EjVWppbP+Em6PkVKCwlmIQ7JKaifJ+Y+kjw9HCGboYo5074hY+K/CBbfsBQY86
h7FrhVb0BFNFA4lVvsm6L7AA0j/naDd+crL+ugfrKagF8E6GZqJwGgV3juS0tWse
JM+vTi/QNwP83/YXl6tqEHGed/gDC2nonGv6+xkv9kDfHpnVeWj0tm7eIoELEE2Q
QVsj837uUZ22nWu/yZIDwMX1N5Y7AZb6o+99469WNMnBU0m2aTRojfxEMEXnULtk
ngV4MunhZIi40uGDkPOMsly8vnGIA+OshMVlqkRcesjBCfYeW0euoyi2v3j7QwkA
bB0rtcYdXOBDs5XtPES1tsyvTLfrezEO6FIDIv32aLv7ZGyfb9qIkIJ3V7eSn6js
iPyqL7Ozxj5d9978XfH2/FQgD/w9szAOAuQqAkelXNSaY0gVa7gZLKrsflmW75E1
mLXyKme/7/+luQeYmj9TwspHMOo2f07qAfc033+SA57afR9Kl7Q5pdXkojSJEZJ3
8JjySon4hI8CB0f5kKKkFuWJ1qsOMltNcR4jrJWij+C1qVTGLSoT78zlfrXyR5ci
D8LynlvPmzdLMdVAcpkYqdCH8pvDxrNtgFibx35yB76ONiyjM6ybK90xnetgmEUc
RJN2vjQ+bMHMlJIq+9nD0pRUIKwQ4jswTCSV0Mecx/v1FX+I1s1kupEVfN50PqOn
omNyysfZ9QhToW2wjrSZKQBvLMoyHfJz3iJ+FPEt5FNoLQwaiKeLznAsJ3u0NwCT
33h+r8846R8ZDYOxF/6eMkd77fmYhKCDTldCRq1Ls2SUojv/k4KwntFr9mkZ2PWR
VQKeYFvNlbdkgCaCgOt1XuuYsc7AP75BkeV7jdhy0G2XodOVGuOtsjvPbABSX2ln
nupzK3Z0QeTgoa/2MSgaGEWpVvXFzsNFNUzwVMhF5XCfZ5hmTegx6CcC2CZ9OyPl
ltzSJIqJKEvgPGPng28CtLVPbI8tGclhYopPr2Up5Joy2xmG8br38pxfpIikc+sC
ClYO+5aEpvXnNMbDiypVrrSFH5yGm3k6P55a3lkRvT3wB58w7p6ylqSiqQXyQtDL
+5Yu7ZSlG5VZhje1638uLA3HbtrIbO6GrHZxKKJAwCC7KRcJQGbCwiurC19tq6gm
oaqi2XhyHDaYWLkQI2tgDxiKBLaREQePBsWKIhIPyHLayTD872Uf5EkRKWgSmfmF
qaIBFVAh5oapZzq1zezfeemMFGYDEWatIaOb+xi+IIWokFjJ6lJ+Gq2DipKBFaNd
tROPPeZ4rNHfooxCQi0wDOM5aLnYP1Q1wRJ40m5Rxr0+FVbAprNmpXPOmI/h+gL1
1bV9U5/fAVHnPy9Ax8TwpjEF9H7vQDXDLRzuMNO6aERaqc2KxQchdj/p/wAQv2Gh
XtBJoWct3H7qSTDbuO/8dNJ6doVC6CIItrPc5Hr9B14XUkxZDyG+aqYcAWMRCKbt
FnlwTdQTySaZq6ZQnEx07kv1rRFV+biyJ1MS2PwaAg2+aTdSpqjVykS7F2bCy90+
f1cGjMNB7AnXtBhcpW6IqR2Z/h8Z28t20NzMHNrrzBadjGIvKEQQmFOq710n06XW
14JKGDRFoRhlxONWZ8Y7xWwOFwmk0hnm+1Tw5BDrjxQ6+mXMtsStcv9YbtogVaXL
r704t/3E1PaJEBtIx2PrTdHHSj9m7CzRmJbm+TgdrTKoCer9r/kBIIVxqMsrqMpf
H0aYfpgIIWbKvn75APNkXSaB2qwQpteJeB49LZWhlgXooQjuAp8tFg/I9dy0BYWB
27wvoxvoRKhAsYbXyHqaaDAQUPkAfDg+5IwOmP35HLju1dZwJ5D7Y2oo0yUcuJLg
Xz59hW1hBAboWgqECmuc4OskiWcfWsxj/OnXEjX9Zn19jZeaGjfeoyeesog7QD4M
kP7HLXKxtSqAVWc0W+1n4/KhshYdPAi9xpOXpy/1RsVUxqokLEUrFZsT3IoDKJGQ
1thKYE8Z+5IGZoM22SEQJ1ZQ56tqKD2m5gVy3fjCfBpY6ZRnu3a+k7oxABgDJ6fh
PPjDx5MvPe75HSgEiMnemXK/1v86RxkNtiiPDfh4yNjsvUjWzEx3ZziuMgjOcfM1
fIh5iO03Jby0JUv3tq+fA3nXpLuywTBvG411z4gzJwIJrAq6FXBVvHu/NMdKe8xC
7rRs+XBookWHr4zEGV+eEKonU4z7lo/brGeGfP2luODD2/6xqiGOY6JumPDR2iL7
zQNI3gkNH2102jugbsvZZUcBciDdno55+VegU9uqoru30QLsXK3XRZRJegjd1WlZ
TMIb639YQ5TyPcFr8oPSkXul2Qam0xbaFplI+QbuPyJLRbTYiFuN8E7vp8/f/94k
1/7rFq/HgRb+T2gUiSqNnzcg3V4Gy3mu1V6cssT36rnGa94gqA4OSyy4uABiPlDo
AnxYDf3rm1XWVYkdT4KL9mpWAg+v1UeZXthR1Lb75iyNbj4IzlKhkvrNm1mPE/DE
X1vES5KbuQcZuu2G6DW8PR8INFPQVS/ewhFkaUuy8Z2mvPXg68DVfvirXMVvp876
quiV7J0aehlzewxx9vl/PzbyaVCkmMv/FCFhJ3EVKGs9aDxKGlJutmoVZsdyQjhv
0N6YyFCw1rw+JfpH2hKPWy7om6VyoLP2ny8SHCH4RavE8YpBkWswPoGHZjEwtD7W
Xa2futwMppaLZXsN2krVU9tmt0zvhz5qDvAwIQUuGC3nDdNu7C0doxlIBpd5B+iy
eiNt4Y8X11j0VfN11cOZaH236AH6ptSBek4y6IZJWwE6EgJWab2l3DeErOBNALIl
6i6YZfKINun9NmYOPd77WlPsLZ2SRHlnMCKcG5pQXrftDCow5ppQRSzs/xbPeYkR
y746vuSxIL1qhDBruWACCOvQnnK9yG/VqRiM7IYrouRF5h+GOLMgZhV4n9+P4uav
G9OVe5N04Do8Cl4KFh0cfTg2viT3r5CUDjLfP4lQ9ZZda82zKz9nccBiJ7Y1yGDr
pD4DZxrzqNCgYmKs9HgWjifSk6grjJEavwZwZ+uAtGF/lTtgemoYJMB/dmtQbSEX
G/CgrGw1IUtWLezJqGMSO3LUGzzTmt8vR4NYBIcKWmJ7UnU78IfXPeaFiqoGDY3c
JwMuMK6oMzkO1+oRULRzn3uX5gxsAX+wPBSaGqga+cnZ9bmjLTuXN4KrwxB+nMmr
z9LtluIatRmha1/TodCOl45v+SfgxsK4KGmsEVutZoEMXPzSvHKEcVmiVhV9T5jf
xAByl7KR+eIBmUek69kDDmpSl1nBrRM414H1yYjdGvgQ9RwAsQD0QgNvbBBZ8PzT
rsnSigCVuqM7HVmdQpfG6wGRkeDgqCSYycgLFDjghFg+9atT/iLLLWUN/L5h/5XN
OrLZu9rqizERM8y8pxcVxeA/WBdZHjbE17bDeIQ6SWasTo4TG1Ls9cnmBaqeZNf0
Nb1TUlO8qxMgAK/YbZV8Wj6VYejm9Fm9GmZotq2fgR/dRc9EbowKF2BnI0bfmNw7
GXknVMtJytk40ppYIOxUQrdqUGxOPuaN6IgtaFnHyQUpakvWZiDyTdr79VZwtRMB
kqcHsq/cbozUESq/XNPBWNqOnKXUXhpFh25crxRk/NS9jjl1wdz+mzOoWZOYX4ae
N6DtaDUBjgMMWlP9X5IQQTZdwT+ctoVXJezM1cavpLvcs58mwv3d2UQr+8elOeGO
nn1NXDIWvZx3opYQSjR+3P5qsCQFvum6/lYBhIZNfFL78bFE4iBBiWtc2yfLHTiy
vnikXedGLMHntDWQsrE65dmANByNceobZ+HTAvu6g0Hou7gvQz1nVLjsKANr8Lb+
oz2to9h7V8RHhlewnW6Ur5aHLjGLIDMlBVAs2Of6TiVAGfKKQSFrf49PiWoLw9YG
FkSm+deQpi3xMF8LiXOKxPXa+EK8YBgkVLD3PYze9noefuW2TlgYO/rIIjcJD2aq
dHCfbKap5TOqxdiIOYs037BolHK5STplqB2pdLazQncCdWoV+qOZM7b8gpEjPFfZ
W61sNYTXjgY9h5WjOvpJ6JlkVYfk9YlqCKvbDPVi2fzq7stQy5+A+xMIKepZNP2m
DA5wArZ3nhbMXc9/ri+7ZWewO8FMxAfTfPb0u5MRoALNxhrIQ6HIEidLFFsEyRni
pA+Ko0DUDIjKZR4315vKdW1qG/mffZ0LXlIQjH6u6dMs+2wuGH6UHnlGcNEq0vBE
vuUq8JYuHp2S3mlwaXz/T4WMnyTrxwPFtuPMcenS9gNIrj0kHoxXZ2hVsSABEX01
LhHIdgJC4VWwQC6wgsOo7zloD3vuS9LGzuX8BQiEl81yruaYZu4BtcV0jpN/TaT0
+p0wg8SB8oTVbIE9FKrZ2zkdLLjlgv9Lp4jKvp8tGiV//XfWbke+opZAXLJkN62a
Lyn4263r07LnEE+Spv1oJhFRpCYlX1XQImWyEWthfm6jY88NLDturbvbcbvT+3Su
PVXZfafVtVTx0kFQFe1RSgYDIEwR7OeEAiYUi94rRXCRHHWCB1rozi0cFbRsGBZ8
taH+7YtFdlrQ8wUteSeMMoVHEr9Yj3bElwC6EMppw6tk2+LgvEMFl8lgLY5qR28Z
x4RjehA2iJk3/E5GpiZMvuKcC/s4wzLMfFvylWqNR1yXQvhQxqoE/yGuLs95QXvF
+UUyfG+4otjnaSbLzbrwc6NqfGGHaFtq1s5KEYoZMH7F11MoNBvTGJRcZGiZ3fWA
N9Prcr1lPpkuh4GIPfgupSR0jzOgo5kGXP/6NCs3uThr9RpMuh/bpamKE7JlFXze
Hgq+YsnOZjwBt02zf4B99+DWZ1GPOUcvfn1Sm97rgoGvcP7kZni6F2CRKywQynY9
XsYFQott/HS5fRca5joEoXNhQCODqaSzMtTupven8qd+byiiz1232XICqiemVcJT
nG1AOv8AVKxq7XLqf2NUIVyhUvaE1LP8ucBkBYO7fVGFIh8uV9aHxyfgTq6wNgai
P3eD4Zdwx3ExZ/QKgpNjvVN0YhV8JOdBfi7eEhZlnNLD/BkA+P3fXjhWW0y03ejI
2eaV5KrdFis9U/BRg1VxQo3YEhvwBnN0AQzVBtBQBbw8OVTuPhQQWrNC815Et8gz
QaG3Lxlr2tZstwKgw+wDD0o+tF8Ir/8ek6WlXltex7tJf7eNf6gx11cFEULeZ6t1
h2g0dF8mKNfcF9lUpR/zmZk/G5tFJhwxcsRjFoqjZsIrBAQrRg9aFRRN3km13Jl1
FTdKGnq4Ac4rTNPQFX+WDfuTtpOamvyBEj89RHGIKrpyCt10caq3wEQMRQ60yjHI
05JbX8bDDyopQTBWZGa3Noz9UjmhhdC2C99RcvVgkR8zx96jKLobGzGpaK4Z4M0c
W9Tff7tcHPD5LvZp5en7rDa4FrRs7SEpZYDIb4z4P3FCfSwTRQlKrULk94juAonA
vJZRjFXr+Znn0jmcYcCbw5Oug6EJFiwC+XR4OGDO0k3daVOHkj6bcA3Wxa+xRy84
jXsX7rUPCK0O048/YpdQ8iRkzdlqIdvjMrrgdH/Apbp6Lryqzk9u+qdmECoxYew8
+zBMuchtnM/z14Os1qV6jYPjX+0M3HdQu9PhaOSXw80PkMDwRqnujQ/Ja6XNbQGb
HFsj8dqWPpDUutQqCn6XXrtwLAmP0NWVD8/T0KG/wvC1iEQMRJmWFvw3tegHQ/0W
39QAcywbocuf+mLm3IOEhTKohxSFNLnWiA9rpLb40cnkpYHtbyca1gcpqxJe0PCA
IjrXBpvhHS9hvhQKsqEEtXF0O/5RPDXlfeth1gWDm7+dME38MrjDZpqY2OaIWudP
qDqlVQwEgegR5GQtJ1BaYkF5Gwv2j1Mv7VWB9E5CjkdzctKwtbkDaXeCcdyXf0np
Tb+TIbaHNgX2OyxQwZ6R7XRzjfmXg13vs2ccoEZGu20qJkUJQbQ3gLsZ3clEyl0C
6+TV5NZitxDoBoE8gHt8lXJjd5ckB/DoHC6WrrIOHiG8j84l2mRbBMFsU5abd6qa
6tucfF4iDu2+Lh5VfbI4cYZ965nptoQTRho9kBswrhkaKYX/fSN+lze2WvBT70gF
LI4fTJ3xuPYsVKqOkUZANT1JCE0sj8gcMVU8fsAn32Saia2zrj2lt4tf7njlHdjx
ktJ8PHqDH9DQScsklmslfofyzVs8C5sMQrZeY/P2rYeBNXUsro9w+IlNNN2CrqOQ
WyKzuUlRxQ/wpNoBUmpQz8Ndjylv7Uzx/2AQVMb/rvb/dPWcTZfzIlcV8CC7VKFt
U0T46ipCJu6ibehz52qIjWu3iZu+0isUOkomFrR2aoQllJWRO4cS8fxnkz4F5VP7
dLx6ce3hUa6cUySIU9meyW634cZghcpgnHHCY39ZKTON96iWPEWp2zoxvQJ37khg
cEzhWUt+EO5CabMJPfe+C1bRRvlUu0eZcN3bJORNZEOaSGyeLeo/8hdLjsmzgaII
MjnX5RhhmnWhCY0MdHtfGq27h7YNLw8wSKyHIxxa/i0P1wyf4IntLq2RalyP7DL9
gr3Mcwm6WmrCWG1MqHDBLzAv7mBiEas226NbrfwvdRrt+8auzvUlIN0PCI5Ne1j5
mLbNhX3KyqKg077UWZHMB5kG9Utucoo7j3Kuwr1ppOabaYamnOenqgXhFC0MhzJP
IN1MYl/QdPwhag8Mqd8/+k1p1NXXdxtuigN61DAtzCSZvW79AiatJw0qS2l04Yup
WQLhsdiydOc1fYDsUZsF5PpjbcvqcTI8irbh/JTpP8N+Q9n1s90ynkTl1lZz2zwD
iP8No7DOjop07TKFO4ETcIcBG6KsCg22xuH+G5t90oL7icgA0VwZXCTObMWI2pd5
gDXHopNzUuEon3i2geFg/G+2JY3H0SuHjVkUlGE1JlZjGspmqiRmKE+YBg2tAmBd
ydSTZHoRLwO4xm3HEsEO592Mwj3PioPuqqCFgnQt1FsR0qc7VYUWimVAGibfKszC
pJWaa2Da3APtO74bPFqHXzfOQ/e1aYXTFDib82eoXoWotGGTW7gbkfeiW0Lj9MtK
7s4SgcO+YWZI5VTO6ZIVbHlrk37PNbrOYFzGvBIU0u7uP/LaE/7nDeXarVyQQuv1
+6tC5guvsCEHGfZWuQyg+jl4GZLGw3ROKVjg/DNwADEp5moM7upD/uX+h3MDdld3
Zrx3BT4c577+OIJ1Z4XLXUnlrCj88nVVh0IyaFDUuH/yqPSGeDV2ws9dLRUHfiWX
c6bd8E+PSMqNi79hropAHJbQ0yfuA0vCIATJSZvole/5mvwzPP67PrVneJwURGO+
GYXtsXlcaCUWvYkxuZdUdoirNZu/n5iLKd4PzrQ16U67BJoMuhR3eJob8Og9v0XS
QXD5mPDulWQsWGsHNj6qwHk8hYVjb5PAhmpZam74e9IhD8bIueaDfODy55+0cyay
YFtnjFE+diTU4mKQicW57+CQWYsVXBY+NIfFXXfSEYVZO0vZDudZs7zMcWfhsBn8
L9aMhDeQsPROONT7WE133ISC1Nlccpd34nSLK0vrW27cEWb43/Ja811UuIHsmCUe
SsrqUMmwSPHK1E0MWyHcXkMSxsd0IFhU9doFl1xM5xL49eSOFyiAlYxcornjxb5f
uuSLxykH+isa+nLNANqTpwzFXNbayBhdO8JpP/ZIgB5RhiCuQdGs+1EoC5HD4nkw
0PXlZv9ELpWR5zzhh3ltiA/ShR8NBG7/YM+b6oCxivI1mK5BU+dHhpL6Liv/3nIc
qt3llVnNrj7MDTGjJXeGQ96uTfr/s92EF1AadLtd869Edwv8of43ZPY69UBBzJ6A
UHceFejRmH2vxSRIIGI83xhdsGZXpMWdkKgXx9t9Ri45ma1Tv+6GDPYakerO4Ac0
RejGKMEEkAgK3PU5IaC8dmp6z1kajRvTCiPhGV4+QBTJGXZFWENPIBtT3o00Pxml
6C5A6geJLXxVRBqRe4k0wXfbH+H+5TG8dYaSNBMywLXxTNalMeLCcbigryy/EIht
chh9buf/k9LcM3CcKaKhrtCo9a/mRf37OPWUNp3xhsPKjhyIB+fT8HN28kpATMVI
D1EcYEA8L4TSZmN68dECTJLQaS9nyMhnRWy9uICJsZF8Putgh9uBZ/CQqQccbtmh
iZiy0MFqHR2HslVSYsAiQT/n1zgCpcQDlmgnOXKCBL6mO3NW2/TmcRBdoSAKYron
/6iAdvzHkaim4HX3czJE2qhKqb2IjrqLa6chfsT5Qx+mJXo5l8Z2pEwKw/MM17yq
n9hluxmfddEfmSck6+ci7BSvLcnWJApS/p5So5AvjCKGPkYWlCfg0pvXtu1liUbR
aOL6fRss6vJ+Fws48kk6MBRYd25qgpP3PyZtsfYHljuUCbGjxJgDgk17/rTByhcY
nZmLsk/5ax0wsWjJOfptRi0YBX2aztVSn/GKuf3SeowLTnRufW6DNJCxBYOclPhE
/JZOEshFhBiO2BMoxUrGQHxa8rnSzlJQxYIdm0WW3JFLDwDbIBvkSSyq2Ok+2IPz
BS0MQ0aNxP9m0JQRu7dAW+zR3zQk+3QtNFTNi1tXxFJeFLcEE55b3MYa0q0cZ0D4
wpgqDA33JaQ3CUn2YC4wn6XtZJdkt8pRBaHq6dmXNVYrgedYlw/hMezGsb04OjM7
0PDy5a8aQ/70dGqyiqOhMAcsqWdonFxXTAvkToPBLZmpEoamtuMfu0PHbN1Y2FV9
6DyEakHYev9Zv0eyuj5caaT8xtefCyZe4J3ML/NSeCcuA64ETB0s9dUz6o8L2r9r
CIVqlcWdZPvPZ9i0DITMp/yNCpPRlKY1YwBTQDdwMlP/xsqwyKXnG8mFIHWiBLPu
6+jQv3sCix1O8GqqvC8Xdld7V6taHMrJXmJOScQFuoLOcPOxBq6qu+rzhuYzmk5Z
1FM6IMXiHX6rBwgzdZWoyq0u8pMTQHlkpeu5P2tSso5HCDXXivBjifPuHBZGJlpI
MU97Db3GyMFsKEsuPCr7e+VUla8ftVNoMxA4Tb1lVDikEYE0V2xCJg10T2J47vWQ
FHAf/pzm6LqKcaYUb3U2BaVEa9DsTA3eGnBY8MPORLbjToYBMNOwB86rY7S+UbU6
kLMSBuDyggGDNI3aj54e+LRed4UbPTL10lzWB3qihuJUbX0WfUTfmzbjdqKIYK5K
+3IsO1ig4IBvYTpMi2k7uFjHCMOXksxK3VLA8eqyWi55x/0+PmvCAt0XM6Gn2Unp
Z6LQ27a7yzESM980zQnTDoXgVWyJ5puuwOuFoVf3i688QghzZ39iHQxcrpuPpoxZ
pR3u/aI3jVepLow0VGcO1beliflVsouvWsGI8ueSxo+j1lfeTePyHisFhPUplZZj
CsMJkkgiNPEAxem8ogiQDKmAMkia1/Eh9kIOACogy/h5iwHq+Hf8hhHgpcJijmEl
3KYUA4lEDFhvVuF39hpAfP8IH0G7Kww1HN5aqNxRGajdV9Ckkz/vQt5xKB3Mz4r4
4FpMGy6HZWP9dkNOVT+AemOMXjLH2aAupPHQJyKzgaI1d5cKyLOIlfdWS04AiBOo
Ycr52QuRZjbVQxBoXebbdEy7DcjYR0Ddh4L5WR2za/ERfchu8K7OwFXUMKM5L4qi
UQ9QbgqauMxK3VYwY5F8CyIfGHQwBxzVGhs9efImSIfqoadJAL1ITmAqhPA9R02o
AFRAfEbnyifynUwq0Jcd4JzLtnQoWEHT3a2rXbOPOdWZnUzDRLM8CLV5dWjdHCpb
JlYIOW0c4AoUjLcE8rcr0EQa7jx0HRq8VTF9mDAlw2r1DHmSJZ8xQ7nqEVtOOm6Z
CzXKKEXYuf9kuc7KWFHHg7ro+kgRc1ZgLLLSisNXAYugScZEzgG7cX9rSiWPdF/2
BYooiu92m0mhvS+PUz/qxRudoEx8doDG4Q+O3cjnaiBMBW8W971Z+buo6p0tUGD3
VE6cMGo5oPMrwj64bNF0n248L7YchynOeV5/On+I2F33gSYewIYNpbGox/Nzu/55
LBAGKV1Bv655RKG6ITSp2EC0jGKNEicjxwjfIqaQBtOIpmYGG1A3mw0iQtyqHeRL
fyh+ivVEBw2sRxqS35kRJYyUyOnXJYcX8BQFMeL1sNxUlN/Nlnmt/3q2aL8gjR+P
nLKH0jsJ1USQPUCVDkg6wKzJJC9RHHEsJGummTZd2cUa+88GzaDjrSo4fwjqpGf4
4cAvNtMhRrn3BDpoiAA4MTgX7oFN6XiOXKE99hEA4vcKUXAUKL/nNET66TDBcwj1
EUpek+HpC6pfpzWqxkE+zTLZWkne1P9vDvE/J3J/mMRvOVw6fAzok6JKrJRGf2+V
TZ7w6Rt/rhIEEbzACo8peo3/tphmnEyFfzcdqIptCUGPIqQFObdS9Bx9KpahHYzb
AQ0VvjyKD9JTcR9+kSzT2pWPeskYhsDhJGN8/lt23+cqjX2EMpxuB7txCcmYLrCZ
iKcOIWMe98Q6Spc+E0N+5DGLPQzSmeMdyfCu1kK68A59e/aOIzuam1WHgmL5X1p6
5jDpa8DYbTVhGFa6csVK2fFznf20cTskiJIo/kUZNV4HjXXAXGsAYyD/y16WCv99
43U+TnvVp+1/p3BYcV0d0xItyEbXV14r5RfaUK9j/gjwJuWBRkuSKz9AXWms0t9P
0Zxvwy4H8/RSESqQjA/fyGvXyHd+qymOeEsziVkOrM/6jd8HKeFtkfb89pI0w9tT
G9GfmAqG/9OIdlXfgHuvUEtf5lUKS+My9Ca53nVMARiWTKcBbntjqeD86N1DauUV
v68qYCkn8vKA/KbbNLdRHejP34C7oM1G9XD0etxJEl+SyKM7iYfkrnbWRu2Zib7h
2/kZNQEJtZeHRNJb+CjVM7uXhSizEH3w3SgisE3AEGPT28tMuaFBwSbXurXMvUqv
vzAkVjbFRhEQM2fYv+ROl2r+Wn1/4BqdDjBZC2KGz75V2TqrFmAb1GlqkaEvdOJR
Dy/AuXzd8vP6jeQVAfkj1HLtOZ4XGQ4CvF18CzgU/axumu7McHQfsE2GRkb6ZnJX
+6w+Fckn6C3629S/KB19k4I+ToP06NXUgRN6/RSL8JaEHQlVyiZnbctl9XkqE8sJ
pn8iCypkO4naLHVY18wpOW+wMniyD4u+1DtOU+rzUDDH69Z6Zs8RqOp4lpyjTLcS
ApgubqbIZkd+3EqN7M/eqQQGzDOgbF2U1gUzuUlLb11lhlU176qDEyUWANMjy5Le
xjwy6Ne8UOrYjyVdtOR0pibszaSS4c1ME3x/6T0mrZZmntOLVqO3exxw6PtVQR0f
xUUxL/sxxSWCpXu+cgqcnrHV+xgLJvnYMnA9+PWe4YKt5hFJUoPmPNOdl7rBvAJR
t/BfKqxzSwDyDSY0z64/nmF6ZoFz60WcuBt1+nGYXAOSUhw7w8Uq218YhrgxM8iJ
KzmzNA5dHrexcZljgvITykV/rn9Nicpt5eQDQ5qfXAU8UwqRwXbg5PvH/53S+u1d
Km8tQoiRBSCceCLZrMAL9R3a2l08zcZ35Bv7+UZG/9CLu9FJrwfzct1+PxWQJBzm
g7U9HWC1lTVrR2fGOEcebipGbLM/bE49xI4tIuvEA2Ap4zbn8rKtc1mu+MAb36dA
KDR06E6BjGirYI+ISWuRAlBCH8Y+usWKHxdpb003CvRtrn2C7vWq4AluN7Qoayz3
4lXuW8BHTbwE/WAJJLiutNyVrrewkigtyyVwv49rW0HiMK1/0fGq9grJ8YBpdUE0
Pv6DmnIFCcBwL++14QOYzPqTXF0sVyNLlxIUvk5iWXNLXKTt3h+opglAJD1jJlTp
KkWv2OGYIejtTlwzieDU+fbsKMsGEzEiTV2+PdyDcxG7UehevLtxln5fRU67IHAf
ox6t9a9lXzIoIqSCnELvN1+YLuzwTiAChYLFi5MIOQ9f3aBjlDMYt4jcuovY5qD9
D2iCQmW43XPe+NsTK8YUDvFso+7Wr7BhdTfwER2xyXNKAeumAje6JJorfFzS30Y5
3DBXE7o0AEUQqmQa4/VfFfDb/yXYCkc1bff5NViMZUadDWqIkJlw648+0tc9Yadf
8Vo0V/DCOhSgP2ysnKN0OZoDZwuGFiwbEEj11kZXyy1VoGTzL+z9Gdl/ZKdUuvxn
7mKo/sZbQolDgTI77/hi8BlmOkdqOsO6iYzQHddb5gcFLIS/hncdDOR2kKnmJejD
tWOsX5PgR4TczUxzuxxS1FLDPymFYveQmXlyoElsylrDr7RzFbsyKtxmQ+N7NW1v
+0AXsCqrycN+CJ3ASV1sCJ4ZUssNzy3FGcoxxbUnvX4VIMmj+0CxmfEQHtIP4YN3
KgP7rjiWdFThK+uaa3+8mlvsUCdaUfNmdcu13mhfqJfu7CczHyGI97NWj3xPTX8B
5qWgpSWSO0pywUZ2mPdHw2+IIt927Bi6A8gMxz8en0hC1/XC0jRcX+KR9V7g5mnC
m212sBeErkUDt/ckbXUz/w1EgpdXfSQ/QvG4UZhc9wpX7uH1QDXb8NIX822lPijW
BfB1fNDLq45NJzELYamFD61VlPbd6J44Y4QKvK8r9bEdZt7yp2B+tjaP4DGBOjvG
lFAlckWJnvV5Uc08wJsnDxcNnV23ZAHtPeX/3FkV0eoie/KwWRnYMYOPj6Cy5xTN
n8Zcsn3Ejg+01BdKzDlfHqI3fcwil/cld+ZESaMGpSFMjH74EpB3sXtAE6ybkctM
b+FiFDvQwiM45mjVFtAuMPdZXevH80ccm2gzVU2nGRo3i1vMsOYzVbKwJO1vifm2
ZN2WFlwg0o3mj6PWHUlmPHtly8NhQTu5AJmMhQo0QEexz1JZfYfMwTdLqgB5G50U
Z6TI6acHlzx4Ng7j9AJe91/kyhSq/EJfRWVx8T3vjExxpJOfeA3x/sf6Y+0PxBKW
N5WnbqjODwR40LCQS+9Rk3OLdvSFbFTqDZILHnmCYj70aS252P25JoiJOsIJ+TBR
e0wWIxXNekylzOsWQEVPg0x8Qhe5Wc4cjV19k6DvNYC23IE+XhhNL9RBVblXoFxK
kUvjDQni1tTxj2aFnt11R2OSQO/wuBW0L9+S6+37X0mM7aOfd1Q1VstI19NvS5tR
wOadlIbw2aqYv5MaqNUkOWIiMPAAoPsNG8eowCTxRsma+vgkRgI+o3wL74DsmtB2
94RSNKSSOqDJycydnK8wYJ7RuJjG9EUCgXiUeF6gfwnsvTdKAPDr330MhOpAByhf
McRBIOwNmE2q8JZgTDeCzKjNEbgL6IwTA+VtJm5rvDgCUOI0brho+pUWjZ2fjRiz
howW/2Yqly/D25blFWYS+seo+hyP6DEwrDJ4oTrgkA1RwieSXGWYOodjQUbYH3o8
V31iwz+RscPPuygkSYbA7BdmkgUyVufw16zhGKAnJdPXXrcQhiiXKkTIGQdDRZIG
bCzRhw6Sw1UJPGAh0GK7QAtEhOt0Qe+QfbX+1DwidZGmSRsapVEFBIOso3hl463B
IiuFGOPip3OdfOQyX+rNOupLnu/qRmKNpaZQa7zMsG+Y/KgWHyYhyM9HX0sKGH+x
Xtcd8duZHw1S1yyLHe5LFV62LjrjIWofhUMlQ4g83dsMUlA1pnHwDy73KqNimZ0e
qHgplO/I42OPCUnLdoq+uNp4AAT8Qo9H6viWfjSEAD0w7XTsgqs4P+EG9HoAP6Jw
r0Ts+8eZMcc+vHy9dXk2wNm/MhRD0LAPF6EVURsZP1xrrmUnJSYOaUz++fRqF4j2
ZpWABZ0Lwu2J81C0O+DRqXiPhhbV8IkcM5C4crGB/gssb1qALjJu20kHYbCL9PYD
AWaG3/bPSO3vEeHMIDeZhKJwTurE7LFj8RREXxpsy6IRdgs0eojNRXwNefHe/YsC
/dobSjqjmD3o1XNznAu8mv/3oHmON8LszL92xKnY10hcivZ3aBvo+ydXWgir+2qW
VdcvnDPc3MjPko3DMyv1H9OpTDiCwU7GlhruNg7oKMMz+MfYr2nbLLycmISDz921
XKUbW8cSsi6+Ps2Rjlhg0Q3yxgrJS7nhweFrbuVDOj+DIP+yO0V8aKGFFeVcNBHd
TmHWEs9gWrWqNwekz21OHqSx7KnVSMeSznp78/ZHHzSjfhTSgBO10IQkdpHJaoHV
xNNoNvEcPggblS1H+P3Z9onrXfsyaWD0Bu5VONZD6kw9U187L6TDUUrS0sSwwDwz
LYHh9M8oUOjGAIgEO/E/nDUY4mOU2xcltvi1xWjFRS+SO1WiVJ0NPIsmKSA0SWKw
It8iNaWwxYQyPJ/PGjJye+YBMg/WwIzZYwQTkLqck3RbY+PRjsR9srK4bSSq6bRt
SBEU7pWmhQ4WE2UyNRRrmr+ianWIHwpSPrCAE7Mrm0mE4MGNCX5QLO7focPOcaqf
71uOAZ7HGMHQKyUmCYABTMiLJzvzr1diBvuOSbsZidfdv57+RahApY7CMJjOlLBW
sySLZz9dGMA5HZYrh0fdYxIfVogyV6DA477U/EyK1QYqT8ym4blhYH1wmSUKmkcB
/2Emm7lpz0VnHHapxLQjU/JOQSmPw78YR3I5DICa19qbHFFEhA3cCVEIlGKsiek3
3inBoesZafYESo6CmZ79z7jkWKLtEMiae+rOptBXqfCTQvWMH5wqV401MwHNV9kj
3G+nJ9NbK1VL66Th9t8DJf0IhLpzPE23YDXaf0hEsDwN2lgiUsmAA7lMq0NeK8iR
yqSfH6TYwDMochA6CGaDzl5l3ZGYiGZA3PG3AjwQSOymIXR+XEd2f6t1l+Lw0Hpc
UrRCkR0aKtpE3pR9B61ko7+BV0k+pqTfqgIj8Vz7YkrqwwuxsWEc/nAJsbjrL0rH
pk/AYtpPnaNNFw3TEL0aZJSQkX7Pmr1uL+vkNHchP36QtD7rtV6T9ZQCphYL5ccD
aoWFFb2SSAvwwlIsNW3lGEYiY+9Peu5PPlClRGEqjtVF4MrWCyon7wsCIjIhOkam
18otQ5dje3ReVH/GFhw89LmgkV/KMFq7uecEulubdiq+HC0FPpwOyDjriNyA5dIi
Qs6la6pCLqR6emHcVujikQBhTEVKMiQNevhHKRUfW4CbLAZTZC/G1naW3+XEFKBO
qSsLnuD6jGAi81lO5ztvRrU8lNLRy5UjqxG4UcDV3Vme48uWASTLNl9G476h088M
Vws7rMV682ywYBx5uWsOGyDco68fkxwnwc1gzwqQIyuMBL5FtOHlqs12DpwxQGba
qbN5trhh9WAgZja9r3kEYulXo1WxWb9qT1LWFjM0qEir9MMOwCllAPrDCVYt5qWg
zAFpFioTYhitB7GAK71mHXQffO+XBDPmaarh24mznbYWTCYC4rNjrOG7fMDo81FL
7PB/CCKG1M3DD+8WRZuP41cW3V/5V3CjQVj5Zuyq0dlAU65cktMKMDiQleOoVJ5C
Se1l6Sm3EfkM75d2XgIM5umaDGLWt1mN7YWgQbR7tt8EakiV+gtilJLEJoaG28qc
VW6Nnv7Y/hcdoggh1qjRVWTOOarC2UDLAMWE+bkbDecSeVXGVNywNfyN2hX38a3f
uiUNV/Jv8EwuMFj70SGHp9HXMtBB5Z8Z3VzhsVoUz+ZYI8Lwigy2YjDLwGDp3EXw
VLRahOrP/AXU0ZTWw8fuN2FolTwnpQLEimALQWMLlNQvvRrhDY0hgjWuGizgown7
CxbOgIdXVB+5mRjQzDmo8myEADzfxOqLBoaRCkcwZGB34GTCCLJ7n6tUgLTMz6sb
9JVGO4tNpD2Qb1kVpMpvBg0gJfI0kcVbjtcuSjxIyBwV9IJpXyIB03n0E1dti4Zu
tVR6b+HEn2zD+dbdO+LHngCN+2LFySXD+d4ozqfkRdaGi5QKy0CiOnq0weTfZWG3
LL3N1mFxbtX9/Zo9WSucn6WP4pT/qkLAG57bTViBe52NTC40po2wCsT3QPqUUzt4
YvdzHmlV6FXa47HeyK9xW4lmYaeSjamPeyBhl4TEaCLgBNVqV30AGXUCRU2P0moc
f9uCWuXYqe+kaaP+qlLRyUSygiU3hdli/jXDE/u/U+28WFIHn8sh2aQdPQbu8dHt
tojkDsGM4DNUuWTP0Ejlcmd1hvldhCE0+velVc9T8aoOlHBX4cwbxnP+bvgOw9w1
AzuQG9OKmFx5qiQpsKas/SflPDfDCEYuSS9LPYdegph4M5Pu1gHOC3nmQZYd9XH5
6UEU1mZMQFZOO9HhULQHZO3n0D97vK9PoeFCUwZ7NUXWzDdRiscbkfQHhp50imAW
4cJ1/FiJOxvSulrevauUQEsMNPISlQJpIN4hbKMIvJMcDa30N7iVn89uvV5gnBoX
zU+9xANgIGANkHbCJ2h3HV9KFwQo68sYHn+08ETTugVCFjIqTggtHkB0Rytc+W6b
PXbdOJl9uqRK926aRAQcfBML7W0/VHxo8nOdyeJ8mtsAYSA8L4Onc7RoEI8qWOp1
DSQ85WMm1U4Kt9ZIzHiJtG6TWg75ELXeFdmClQq9eVYUEdVmeKkIh2UWqew+3qpF
nKq9EJdKnk0DHNl6wPu+vAqJbuOe4QUNETZ7v1gOU1V1s60Sbxnj/m4i1H+d2+Vx
dGpCqPDzM+At+EZFZ3bb5qHvp6K5TRW3C/8uYFVJi1Asvxi+EP3dKGy31zzOpIvW
RGCPQAnuWFUbyWyOpdQINr2nID1qwiwj8w4mQlohlgnQu3gre69rcYI/chcTiqZw
O/MPlmseV9nsW0Fgz/ux8VwWhsObZ7esxNm31DIk+rTIMxBHyts6SwZ3yLvCx6Qf
kKDJBh0zn5rKy+SEXDRP1JV6uOxOZ1BJ6KTHQWqpI3Tq6FKhRtmHcdoCKT1B7zAQ
56/XwBJz1cDIgmiD2S9Bow53eqIm+dfz5KymEKpVJzaEqr3O/Xl0ZtlhDpV2HRgW
EbjTuzC93Gq2R3hQgcqj9xYN+z2jITlusx5C0mEKonzK2rgfw7dOGj7iS5re/wp5
WN1VnPNP4T31x4uJ0pbk38wx4YQYLUloK3et+kfWJh3Geg709YvQLZovd5wkPwKd
7YNt/glFLSGViG65SqOlSenK+G3j93+y9VtJWpXxIgqD+KbnbRPtq3uI6mUMjZKh
tl+3OT4P3Y6acKtnlsMqIXgL3xVyt+guvFRYQoz441oTqUePyj9ZLa0yxFORwku5
5aGKejfvpyxOVjNxydgPUXV1yB6qYGJGoHj9h79MBvRxfQh1zF2W0aDhLGx//6ak
jPTpeDswLwy6oyoTOnwLSwuWtpD9d2sFdC20XnPOeAoNDZC2PqxU9Qx2jXq2nVLT
23ej/YVVx1z4XL4gr2Bql+A8fLd9PfZbT7OEEhZM832Anvon/dUa35cy2MsWURf6
hfVVjOWyW6BAZmFUnJPzz1SagbG6nRutQ3xlkMh8R7nhOU5Y6toVRG+L6eZTWftZ
n1WNBBZ/V4tPZ+0+oeVCPSJ6JMtVTp4kwxkgdd7XoLMenyhDulSVTbXMGINt0+El
2FpcJiP13wDN9TQlrY5cawlsdt34jZAZruIckbi5r57QHnYoVldKeyF67vp3kj/X
hscg8xUFiIOgO5kBAnQxFykWXvDctd0jsog2s9347obagZzGbCMPp5YiNy+6d/iq
JD3F8BDwL7G7NPza1HOuoyRMIIU3znWqQE5b1h+ohpqvotLaSOK2enwd3h4yAMkX
GD78QjA2gsroJH0MbAhIzrnsuTAui0MF5Gp2LTXcxpyo6ipWlKFTyYPfv6UEFZ/I
/plr6A1GhfpFohObZrgIA/d38Bh+ImMPNvYd8Fd+jcmjYUOBpeTUH8evIwkhzu6D
GukyuaG/jdQA/PXe4AIJuqTMK506y1jMULP7L4ZJwhq+EjATMZvohLx8am7v7mEw
XOGUruI+E8yS6qYG4lZE3LtwLrdVtLXJFhrO55qs4eF7dfq4+gM8CuxmY49cm7c+
1h0MEhfTNtspJDTsAmmOT23jk2PN/8pTOkDi0N3SPXmgrAONGcYV3r6rcaTqkpDR
MUcH+dPVyKXyEx94jCKhPLQ5bPQgtnNvuZxQR0BLN/+LTz9/0M/cDOXyv+7EiQxc
VWUP/1xdXC7xUEY0LZswwQb/81rBBw3PwWydOX+hglvNvqAhEeVzfzuMBhBVwH5D
jzmjLVu9wZ+5cmycey20D6rTlUjgAq0v+fUZnmuw9D+ksdg7tWeU0tq+J2gtg9z7
9+tNqcQulw8ktyzcNYreH0yOBinoILM/zBh6FKTdS5YgmVi92+ooW8m6CP7qBi3M
zwBJaO1ieVe5Q7HatsQ2wxSmQcYvcYWsNwzORVO3v7XQOWxC3v7aIm4iIDOHZxu5
0IsLFGqv1iU401FNKZjSMHJYBvys5f/gkDcGceZAqfbu1PrBfH9tCCjNbTTKBYPL
J5FQCydouU3ClC3GW1xVPEKzWE/nc2h6hToDrAUvEkZc8s0SgLrois9rjpYkIMbo
coPYkdMKtEZDFpEQtJi5PpD3YnSchJDBL2nMZ8P/TqI/rOJNc+yI3QdTrsyLu7BF
/Rlals9AVbdWPQ76+f/1TrWl57ihN+pz+qr8ikamPw8Rck26f9WSsoNEPNCoOZJX
p8DcCFoUf7YyUOqh8nd/hKVLA/zr9m8SWdNr9O5K9eVZQjf99cZBAYDxTODUd+th
TWf0wvUth6oW/Mtz7qwE53ETcDwiBOPFTB1DR54cZd5RF7opBd2RDzGrv7/x0tUu
icpOvwl3u5f5U+dBfN05VVth3HUgg5rdtr8U8MZqguZ182czgQn6BbnwJRWOCWm+
FwZcTRXTAP1UQCe3gEcEV++qHBC+D+aXNezKzcjtr0f2pozNW8OMLVo3meHauGaw
8OAZxf+bnlHHgvGsFEpEvVMM56elb40XTCbQFpX7mMAv9Q7SXfktd1l0Yk7zlLkj
OF1RovYBRr8wyUVdrsNBPJV/4UvoGYS+aS5yUI7gQ3gy8ROYMQu2rCG+7M5V3R9n
X1oOOP5N7Qix6V2YEBw21e+QgWEzrnZBOoWqPW/os1HsG7FdlELNe+9pOaTKQ5Bu
jQDxiIVyaewHqfuNzlr0bxDwdqb/AWDQ/wy1nTQMXblpM3CyJGai6fNbCqs4mm2M
aT431Tzrx0PRwVxfI/JwPOToSo9im0bhPZajYfjp/ME0ICNv+EjYRP0PWiItAwCJ
FW2nNhJU30O9hmNYYABXMVWBfG4KUopvshYj+0ew9za0W3oUyMfpHsuV8N09LJI5
zKEKwCKL0MSCOyiXm+j391j7jnCgvzPHGKs7lUCYyPvYK5iN+dR+mN9zA30vI3BF
PHuEequYEKySzUSPylSZYLwgXyZ3GSk/M1V8e3CTcuw5l4c2xcfIKoplw+XujqsU
jbTZ10Cdl1fppXeAxZgdOPeaKIXF7UKgcOj1heF67AXfL4f+PDRI/THKsalsXVaO
C7UiWkPdGS47sj7CtooAgjPneCFCNHBOdSgsf6HFRJ5f1o8Vs+KeY6YoRfwbgZOJ
wCDxsXfAYtzK5N+q8IQJzlYkQTNrC/PAUYZ1jmdM4twgvL71yZsSrQdhiwCsENGa
3GjpFtxktfzQusDuPJLNqZZEwnNrxDVuyI216FEjDmyQ395WqE7Z7MD4vEhgfjdv
7IJgYWMFROZeTN1p0Be7EMlkgcI73Tvg2iCmM+duzn/hZzKIZsrpFLzui9IiFYnJ
sECvoPmt/dE9z9YmeAX4Tjbxa4Vc7utA7NfVHwnRwCB3ZN8M16Op+evydtvxh8pH
YMnmEA2FX6W7BKGvshZWzioNBwOwrY1PzRDWbG91GK34fMay8Rmvr5uR9KaPO9fT
Jfl8F7DuCq5/38wHVtc8Dqxg3C/NehFMZMzoOOI0VCte8LRSSR93U6FRRErpaRuu
h3kg+SLtkoLUy47GIU7w3mKwXZgX8H51ffJe8s0nxGabnjsTvN1UMsif5aIVsbG+
mVWg6wsZ6EeieLGWjJf74vxGxOY1cSJAiL3yhSTcFwMmNbSVSiyOLxtOW6SCztAK
kozwLevVkku75ZDLp8bHax/gPO3IPuoK4qOwPxSsz8VX5RbeRJbnqS4Y1wY+j+UE
XVPk891xZFT/V9nFxgFyq1NjSh/1Uw0+GHUNDp4k6moP6lH2hlxwwFWS1vNUSy3R
WmFbloyU7qLCVAvSQbLbLlOCbm2NTfdgvVkm1CNhe/xaddIaA8K7AzBI+GNtVbMW
1cyNJG7pc/VXXXSbiWHAVvz+xfBfzZYXKBRE/qfIC/StoLEtdlpwOfQrqOr75nqY
GuDyv36y4H90ItIBZY6D+OpLnxWiLAppZKhiHcJjLnIF/NNPCbLZBGrZheRe1eVk
PPIeDhLa0EtXMsLTCBM7Gk2OEvUQxMW2ooMt0FxAbw31V0WO+Iw/416DNzrzf5NX
jKjxYUXeiEyCZD8BSFbLL058shzN4qifh0Ld1eo+S8sob/5Oe7TtSWbSq3TCw9ng
4VGqLPEDs6hYHFfptO6jF6svXB1X8EhGJFDzOO+Y7BBGbAiKNoesb9bFVXs59B5z
D/P+6FPWkkoCu60BaQwGOCZXCDr1RXll9CA6QanNOvwtde8Ow3A06/ZpiDGTrDUT
N/uxRxdMVZ9lGxYt1QKxnt6Xi8E9fxF4icBGe5Z1LcqSV6kN8jMqSWOiti/ucHlA
3i5SQRyS7lImkntZ0lCrQVmBOO6vZxbm/+085gSWUhDeuQQ5h9PDv4lQ18zsesjN
zmcmxTjup62abxAtZQV6NlAzI8iG1hnChHQdQmCbqyEMu8k8u4Wtm6z/XjBocwqZ
+cNghwuue8+X8Pu7Y3uPwjrjRz60f1X/eUQDbmA8fD0O3/NMjed7AcjNP3kUAPrI
E8KJrQtatTzwi6kZ1yNlXiCdYO4vH0O/qCQP0uCyHLsk73GZ6AhkHeFPVZob+ZNh
ljI5T7f5/KqGGXribBRkEhCEI3OpJ163Wfi1DT6tkG4tXPtx0WNgRu/Kyla6FnCp
6BP/ONrWEaier8rkxbq1ESvyBv24xsjaMCP+QJTKTPpbKNQtFj06RIEXkimD5wMT
yPpWQnGhsdrzLG/ZijHTUIBQCC1u276u+tzVMip2qVLJlrLkPVZVg+VANTJMVvuO
pt8ef/ZBdJXDOPz2gXRivNlfb+jcoJfbqpOZIDfd3+OJ04Btw/M2u5nmOy5gpSfl
JncaduVBc8UJ2A2FB2+8R80iQqjcK8LMXMEMMnx8pHLDwtaUT4XRokyvI5j5LPkX
Z1iuNtX/7+wRzpf+J6XB8BRzqvdQoaot5VDaCtWZ/kwQNcA6v/gsvPP+URRAixXZ
I/89BJM06YaS5pB6Ip1rYz9AnG74aP5YevdVDC9SVH5BwbLxxY/u17LzhrSsViOC
Y9RGKQe4tN07y/qK/CW7UyBKkqsUAt3LlXR5xuEEUzDe0f73l+o+iZYfdmZSKh2f
hicaeZgKT3fGhoedV9oFyaoAls4Nc+v7C/0uE2eSGz8qiC8UDzrvT/1TF/ArIrcr
xRISj258gHH7HmTYHvVyEiZEYcBMgGjbwnedUMj/jevgYwsAB6Xos1m+hljzVmfA
vSLkZLJkblY2qTRTebNhMWnt3OaR/yhTmm3n6EnMOh/o4kv/8TlmNJhbHkoYLE6C
9fBEhHQBfB45aOEUQk5wej7zxRkARWQUMR1XKyM3Gqlh/ZJh838EputpejQYemcg
aPtu4Bxu9JviI2MACKny+qPZ9N0LSfvsHGUElFOZRk2S8x/+vp7DoZrYbcovc/ly
VjZfMasSBPeAvidKjIXsKaBxgTL6wMs5q0350nV8CZ04IVimVrkhf5PFvWrDOkYF
gGc8ZUfELe83RYwy8tlD0zTsqRsBwHGFLbMwInrH1GFzXMn8IzuZo6tsv1jcrgi0
5GBak5QXXzfJrRUMpT3h1XzCkmdIyx3b/cka0dhGdjPKtToRCmqiOVBkdG8L/dbI
1coKt3yi1JTfa5RAEfliS/P3GrYzAJU0Duwl5LY0WwDGZqtpaIRBGEhSmESKMCWM
xCPOiZdvjbF760u8I/VaokG7+eMaazBehaRtXVHEubLo2wmf2SXM+VmEhPZusOwx
AQ6BEeCLmMdO3qFj4M4/PchT4B2maqf0L+8WYMSVNhyL3iABthEj+PQaZXdyK42Q
oVnAKnVko6a7PLTdAI5/IRaNIYcZC1ANY0ijq40qheNfutLkcoL8P+5qQobdWw6o
4aXY7CAYodLlm+cVEkDu8RG0eDiBe/kFvKRD8xClj8Ulz8iYHm/EJUWg7rgWDSkH
g5aXofGzRdzF8vlZBrXpmJ6Ljuh4tXVyIKwZDojyldLgKBQR+2kAfhttW24JMNhH
OSNxaZHBgL0REsEsChTCAWpzPETTar7eeEQUUS+jw74bQ3fEMmU7orEPPMg8wXuT
Tegkm/QMdkn2QhurJ5/INSw5bFzPr3QhjtQ1dxwaoIg766W8dYgN/Vn5eM9gx8sL
sZK7yWEuXlBeQ1EPX/1WJ0ZxzG/X+ZIP0CahqQQM77jpkSraV0e9l0C/IvMNS8RD
XuUJuU+ICyTe+Wkv9bFZFkAr8Jy3f6npuVFILeiVM4t5qscVisksypPUNxCDLzXp
XJYEmeaQft+OEUtBghT5tkHSKo+yOFPCJ7bXl1vsRCpMF/ifuW/K1+WHsw2cl0mt
A5Yh30jaGiJDOLFMIiGDMz28y3Ev+HOXfzJtRopEyFuAx92M1SJXt+KA0T3wTSY0
HAqYAHcPm1uKDMpFqqFPm9a04OOtSQJbIwYQpTqSwSk=
`protect end_protected