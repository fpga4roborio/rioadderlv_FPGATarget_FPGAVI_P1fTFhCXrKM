`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
ddtXksX2+yylW5zu6QL2Lhnb2d1sD00763mmSITNX595NcHTEkwn0zB1Dry37fOW
FufOhVzEJp80NC5qZ/+F0Vk7Ik02dIR0elf3clrjeJRK85K4e3Hoo4xn7YbFUIms
l/8VZSb14+JVGURjfswrIyCUotIzlzVYZ6gzoZwDXIi5gQIBf/gI+KxNXPaKV+PQ
Ufys/12rjO6aI/pPlqSm0hCvftmBcnezN2hk1UeXgOIuKZnogjOsf0iJVX2aOOWE
6pD/psybjbnsNB6kH5uFTA5frkzIzkzl5d9+YDm9OyC+k84E83I/7/j+rk4L2dah
QJOvksSIzN867/4Qt8qYTQ==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="MvBXkzurAa5VTw+1JJ70nePUfoQXBvZOku/SMmg4TwQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
oRtzZL4VJ4iwysPsC8SXYCzXS8Fw2gtZTOskLcDV+1B9Nzn1zTyNtlo6lNICRmmK
ZRVu2BmCc2G+fmzynYlNTnSa7C0Cuel6FYpxCBlOuk3OF2tzAmLAuDyOH3Z1Yjzk
a0aHuoCdIRKv7BrZCdALt03JeUmXKPdOmIlkVGFl8yw=
`protect rights_digest_method = "sha256"
`protect end_toolblock="Jn9CQpRhJt4rnzZPRk+dOpzAubz7omckX1MrFd4p81o="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 13424 )
`protect data_block
gD6l00tciPUa6pDNTk/+t0OO0nC/UTtBwLB41d4inuAUA3i/ALrNyoJVcBnAmEQW
ptbcNp5fxEUJjnOxnedyZEuEBxWRieZFQnkRdF269oNo8RsKA4NfIvwHPa8mN3P7
/Fa2D8tTrIdr7BRBGlfbxMZs8qAPJlfknIxAMI9rAGt6uM7HnsGO5vSM4QiMvepQ
H6cg1SLfgn62KFrELhuOLU1n3Q2YHiXj72eJUFnAGjem00RSpk7mKl0mEOUTl/lu
kpygAMrykc9pvwYNkHPHoNN/YNmrQpv6uYfAsw6yv4TCABxj4q4SrUkEBADsuuuD
NiYdODOlzN828WUF0wKqv/S8BAxMsHfzz/TbvEJub58YVCFbrOTALReadve0Cts4
qXRKCH6jInkpsZPn0GMvf+ChQdoK13kMAtwm+Ct480RtK3c7MPuBb3uar/cXmcdM
PGOoPeVxiH3DQbFzwAysBHaYqPxgwCIv86odQpjFpHK7PCjkdv2VIPvXBBSt4A7N
sZtpx39cxRvelUkNWL1s7b8W949oLSeb+hv/V1Xq/FdbwErt3eqvwPPs8RUJQxAX
4nyC1OGv+JnyzkvSa+lWI4U8jQ55RRs4UZotp2YD1G9YMci7jQBnPEt3nN8oLUqS
8SUi2LbSQqOxBRp40jLm/DZK235plsRMsR+vgjP0n5ghgVJBDkOCTf6R6IiyUDJ0
NGPiAMv95K5+hUxcXZiqWRa3F/UDbNqyx1xVo6OB/XNL7yCX0dvOlgXitvU0cT7H
2q9ATajQmKT76/HDqjDSSDEDCRACG/gSHJ1865nv70x/1iG5NLs66jmaFnlLMo/r
dhrsq3C5SrBXO/ypHA9Q8xSKDjZaaR/dzX0ldD4DAX12GT4NBpuYn6Gy8lozSxVb
X2ylUD6Z3q6CSuqNhYDLB+C1+U/z7F1ovfekFSHqIM6Y5B1Jj5GlImpgxFWe3cRG
RQAQ8Dcr+yFcj72IXPvUaNW6QcIaH3krmRrE8d8o2F6dPGNbkE0CmCZ+G7rmcOzb
GY2VIdZbGOKCGRP3K915aTtELsKR4Hs0hivaZ3hNTcxlUBIUvPqfdKJCXtgHfrGm
0xNXrrSmFQ2wDoP93cy0HHFZbmpBsKcquRh9NwSb2w5HOUgf94SwW3vKTlrmeDe2
ydS3SY7stMLt+hlOtDj/od63a1STT7xhS8NE+fwLSpz5F301c4DX+i4W6ILG/U/8
RPvg+ZZMVHGi5g+T4RN8i1L0V8SGVpX4IS4GTVCSn9GrUujJPA5MCxkpA+FqspDW
mAGqEg7RqztvTfAjlDYwuAawOmMH544CTpPXmNOZiuQGl9IP9RFjzuzslSnXA8cD
5UctRUvk+JVp1PteRGc087E0HAkScFsn3/fBPsOTBJcykfDc3UNEh4HpCIi2o09N
n1CnlOkallrJO0DnkdroM2rJIIArJf7/2f6EHgBNNeE3lOEbaBJHO4krMp168qQw
Q4z0uS0CSypMHSs7ybM6GD9ouDFE0p4Dtu/b1P7EFJB16RTJNSJEL2Rym13VwE6w
KRHW7/sG2Dzd+h+g4tdq+s2X5MWQ0NagoQVJEAMvghILDl+bBHmGQKDprUj3hWRZ
CxrVOBVcTmJIFpcZ1Z0ZG6YkcbrwA04PF5YskUgaYP/p1YZJ2T53nMmjDhHhMyyf
wKULvrYQzKn8MxcNhFtHLpbZrotexLstNmGLhSr6CZSlBfSthoBfTNAnuN6XQSH3
JfidmKi09EnD62EJqB3/vepETXMHMNQKwde5lkPeHPuZxykEXv/MggvMbE/znxgL
ikF4pwLlgmuBUYt6duG84VP4O0wcLlA8n5y+I4qyizGieFq0ZaSfeMryAC5nPWlV
J6HzfAOqslZyu8zv9AHTRrsSdU5fsQYF58BlDwlwp7+lc7hbWMBQWGiHHPLDz38Y
P/PeC/g/Yl+JspA4xpb4hwbFhzoKXmdj/bCKbTUlfBRWXChyqz1gWnsw4gijvQmQ
ZHTtfTrITaKl5gJVBA5MS/xu/LiwzdOE7zAhAkhUhOrZwYA1FDpDLtnMGLG5HRXk
Cyr7KeROO+EDh51uZfTgnTtuBhGraJjsBRk6w01is+MqppaeSWtCWMboZLOppF+b
6LZczaNlzStzOrfxxm9UWuCavqYtTraUIkeq4UCYQHTz1+fB29Bz5jZaxkl7Sp16
eq7bStLMTykiJYymEFW7wwzICSvHTz02Jnde9WqXgFP4VGppwqk3k5lACeiICQvo
eru0ZBdHHdlrRTtllW0SJoPeyi+pBxR2Rp5yjCc3pO6Ylc25FWlK+vu/YSPvbfwJ
wFf9MwHpiMYAsZjijzCZXze1njQkaEOuxMeFy5lFlM/HnAaseZddhZsvsxevy81B
D8CI1Ng7mWgCIEOn98jW74EnArEyH0fwztp1Q6UrJhBLtt59Jus1ucn4j+UFfTwM
Jq9I1vqY0wucADEMN0x8wypzOlWUgFRzZrIPpa6H0LIXlX/5tYtygFieHhKOM8KX
pvOxs9X5v6AYOI9ysCBh6Y9oqDKQ/P7rsSpQ2KXArjn5t7ZlrondWjvVBwtUHLdk
j4TzlG3U9eJO7iGcn9WK7po+3Fv/h5rrPZh5ISfQ3oxQytu05nYYmMcJOZ73OD4Z
nX/hQDRiQ3QREeh/GEAbWjJOlidcY3o4IJmRXTynyLzn1UZjuVxTuh4lifZ7iAyN
VlyqiNlqmtnry1k/szXn1xyn/GROwH6X7QmDPZ5oa8VW6GYW75tMBap1N/kfVbPC
cq8+irsxJzThT1yQC5i/Ox3mseVT6YDfmNTKp6Q6YrY//rxCCJygEpL8PULAjl9N
eEL23agsqd1C+wU+OrvsNAsAtXGHbDM2gw/Nji/sGZgbkpnq4AzdzdasUfwlrhHE
kqBLhvZZnMVekZDsSyBtz6zzGF2nqd7njtTjw6XWO6lfdEhxKKObSgwnce1dMiiJ
T/Vg5auQovFxn9k8B7AqCWE+t99+Addkk10TlxjgyaCm/Jk9UVJg6IDkgEbhx2xd
SdDHENTGpQrnA1tYFm549gvjojssAZg1VeZL4+7IxYwHcx80nkjQnSb01klWVapH
IPFAa4bP1/1e6zqWGnquBRj3JCZcZzCpfqzKnLyj5ZM593mUwg7EPXPDWECZg6L2
0GSqE27V7Us1w0GL1y/IBWLRiCJ3lUa5lUpR2hCdUl+MqkV/oy+1aHMCKO3UkE8a
Lccg4h0ObKhTZh4JmrL/zWIzH+euXLo4XI+CjmxW7bMKHRYFbsuHku/DtiZ03R2/
nQP5IxEDM3/0gx/5LHcR8OYLw2rRObE6O2H0cumhRhT2bMH8usWbuWXRxH6/SXRD
CFdrMKgfOoqDN+7yBFDgjFZy9Tw5ommZK09qBh+Z4saZI2Yvhe0WIPPhnWpCqBMt
dGozd2lYbCFFnzs946OcmoW9Ae8TAQWkmdHbquA2apH8WsHYcDdz+HxQ2P76YQ0E
ReX1w8MsO7DGgj5hxN2hTfn7S62N+tLIwxzVe/TYVoJq5ggp/SF/LEM9zCTDq33I
YlxFDZMr1lZq4fwIQqEIg98Qzwzc0GmurepQCO9gmaOIa8LrhJUz+4nI89clAFQr
WWFo4r5c7iW/FoTYe3NWGO2Ynzo6DHBDYErLK3QWhNGQ6PmZtNxZXpzlfXqEEpsp
9F+tp00/8gxKKdO6dOkqomoHM/oC0lq79C1XPvI5xoo1vgy8lh3T2dqSQfLYT5Y3
QDAAkzxXVX/cfRME5qbSiVqaYTdlPP5celIqkZt4MklAmEDmrln4KVowPMmYdM2W
7WWeD1ERv2kK45PviaSRKNZnMdDVv9ZQZSVrpwrGYPM4vfaphIKZD6rVR6ciWeF7
vL7WvvG3HVpGQNpuqbkJM5lCXYllgX+guw3wMJpKzh8xAzs/edgdbS7Yydgu39HU
RcAHqJ+oP5xoEVQsWk5pnj+HD290OH8oScL7TXETebWg2nIi7oaTh0zzYukPsh7q
iQhEit4c9al11dl6iqAR3ZCWjd7KNb7efoeNdZvkvAN5fBhPt+Hd25RSl4k56xSv
1LSmBOmSk9ZQs9iEFtSOKPSbU7vTV1zd1/tCCcfebTF2hvWmyZO18qOdJ9nNaJTt
daajB7HXSKYp/X/rWf31iaGQnsOKjGgq34mPZ6lvf6ZZ7uST4NLIZxULaAH8xVsM
CwMZosvNlPk1/k6yBstyQxdXjB/sbXXRLNBCpRAI00Vvq+yMCZHxAvMudeiG85T1
Ey6Q2Q/LJ8EqhFJIaiSYFmZDEnl0ltfu45Gxp4YMkvnw4MLqpvUbI7yeI2hUtZj/
UETaKkonEGvl1iLLo+H2QwZH1u9r8gSkaULDcAcBy6DHZBAHmZrLf/CBjihHgN8A
WMN+vEq69Nc0VavCXs86dGuca/DpUI+SywMNd9J6rPgJ37oV2BW04fkf0/NQP0ye
nUAzRInR9QSXERG0nOjFZ429lgIfwssumRIZZIr9MUEs+98gXWXKeLozuN1aTf4o
HVWti04+/wIEnhPrh46GvE5LopL9rBZemXADa0aFKMLy3h+ZKpBKvoHn6XzJOXmU
pc27FgsXYd5x/KoXLlE43cxUgj7YM2z5OvfIW0u15Fqu6m61RgG49T5wvl4E76YE
aPPXsLYKET298ziaN7FA1ZdARAeXNSudKCnVEUlrbM9o20bO+v9XqDW6o7xGF0zN
0A75rvGqEqnvkU+xPt1TuSQmCWsMSxQmosGbos8HXyUK+y7EijpdvMwZu777iwBC
Qb0m28x6SRNrNP6HBuWs/f8uYxetUyZPDQzAP9l6uQJvql4bgVr3nzQonYtvC+dW
LCgWaQj8W4rzqDANEwMzujpLqRrakt2uWjYUSzbtSBLo7rlgn5LGck2Sv+vfXGYB
ffhYmN9ZVKNoBsRbmRUz+ATz+/+sq7mllG2uJLT0G4cny+ha3PX2moG/nUhX0D26
lA3UHxOjFJmKVjYXh8xfLk6bXUf6BGjy9Cg3qifvzzKqqII6p5IwchRwIhZ1H8Ll
HUjXKJU9LQkkseIN3FuD1EGirNcqgK1EeUqtTlJ/e7uFXaIZ5KnNlXctNJaHH1S0
CL7chj0xXJxSq+0h61q0VSiSkQrxzLZ7lFZ+AJ7VvZDvMAOwhhUGIZHcNHZHFmws
rVnYO/+E27iZQr5oNUB5KWiPkE7zcpXUjwk5K1Cb0HuxOJMNo+9KKl6t0hWdZMLf
s3/ef0rgTK6psejcID/4mESUZfnvdcb+vvDoMhQKC5fE420YKt3FrFPvAGwpQ3cE
tr9Guz+rkqH7GuHkU3/X26sb3Dc2s0R8spEB+YNDPkDp7ykIPu+WsyVXL+wzyR9s
pIDd9OigTE/fYkb4gnI/44a0zNHFCHcHZ7Ih5rgxPHU1U/79bCoWdCoJeeS/J82v
zUZ4Q/faFk5YPqv5EYEMCPpN0NZx8tUpH2bm+rxe2DYs8teIyzU/iLl3nchVn73M
zsLwpVmcuWh6IECwNsfdEzDzA0PpSL9gc2KFk34SN/lalmbqdazOBHHyJVv/l6fI
YveNz6PLKOlHj3ESg3mJz/8WEB1/fcHoUKkA7/fISuHGJUjKIesQQVmcDdgkAoQz
rjZ/RH8yPfSo4gjj2y3uvNDgDHLiEP7wRAtyRF/zfqcvHQlJAMtOKOC5le+0tNhW
zWRjgkAX/HgAsrbE1dqzcYKb8oCVY+oXV6B/RgKPNMrBoXx4RhRy3Oj0kLBIiluV
xNwGIsFwLl0k29PxuuMjRXta6OzPz95zVjcPH6K+P3c58iVQZ4PKvtq6/PX5gvBt
2ZA2nw3k1WNt4UBgDkY9KAjvNM4vxpiEJUvmN23CdO8ywNSig6wJDYxh9VdRy5Ds
1sjpWWXRckVm+P4qNSN5BFXshkysJlCqhG2UuCZY9lDXDOssg0YDg/LrDHAgkY1V
pgWMnpilLFlCfkz1xfEzJ6Il7yIWMYCNzo/ERXHKX/Gm360Qvnte+EQGHbk183UJ
WyZnGpLTB3g62PIBtHfPIbVwGDxM3yrLgSHh0yCf35AK9q98hBGGLwXwY1d5smib
ACY6VxoSBu7c/2Vl5rsG+wmY/o+8zMn/bnE07A2RF47T+d3Qq81x5h+zJb0DL+a8
8/hDmgD9jQY7oSxk8/hNYoEWqTYJihQWJqKBMwkhiEm6RNSjN2GE3RsKWn1qADUL
cJGa6LGnqPBh2ofqHdtHpfLFQjiOlWqK4j/DYz608hrjrBhhhhavDvn49lpy1QZC
T0zvsKM6YFkrz6/TpjApzZDmhL5wzUUUMmQqgKCCgQmpDvTyLEJ0PXRVdjqRlEJo
s3xiO/ja4TgAL/VaDO5OCcIjhfo8/bwcFxeVWLyoI+H7bjlavP0RWpkCjTO8Yy+r
vaTAIkrHlHHEZaEao7QiujTIQG6GJ8ZKSkG5QHbbCq31kQuxxxMfSm6NQVAP8r1w
2jv0rkQVaTtHDUFhwnKPosPa21D6iJY9jGguHSPdxrknKu3FNJvqLh6HEXceAsIX
xRMWvSYmsIE/W9uEv4A1sNgEUIxh12FhYe+c/HLXSqK60nnr+3+mnFhzYstryGbR
trB58QcJr6vtDxDs4FqjPn5s/XawHRNBmmyRwiwAH3NWTLHt73hLEhAwafH+sSoM
z63+Z6Ziw4WrcVXdSC0MGyPNeJYj+JRWaS5DGbVyRxLxHggtecq3ngp/qpGNg6rC
pHSjIwuNLKaLcyiYDXXe3wD/e+Hr0CyZfDpsUuu6MQ76eJthQJtBx8Us7csYcv9d
KiIdCu5a5zOwe01lXBScm9ARzYuNU2ByED+qICOPoGpQ812LoaEdOrN6i5MpCUUY
r/yW8RPLnDVkqhijyWsfopC/SpW3yMpkflonVKj330045d8pyULSy9WqaO064see
ZCwOc5JvjQTBnK/bqbmMXx+iKjRO8q1G7KZO53GthyKJ5l1f6l9n4MuYD8ULAH9N
DRbO6fb0j8ecfBS5YxIxNceWhDcsqU1RITDHze3A2ZbpfNQ0LEW6QxMOd87elHMA
dTd4nHqamgWb56Pqz5Xxk6+ASZjrKV3JimOX2RQL17/fZtrZhPjupZuubSJiLMg9
0Ep+QAOj0SlV9sL7RleG91r5rHHHmJ09CaPTwa4kC2HeHtMxsGgJ+JRYp6hdIjpH
MoQ0Wm0r8Hbx0sKHntfhqMBxJxnrxLXQTzcbj8vlOjfi+ISEIELpJFQg472e9yUl
vzL21iSh2ndgXWI1YtstHfOlZKAqgG8PUvhU68UYDUvht9YUwb8g5nscbpnGc76T
5qZNuYlDtlunAGaXsWUTT3lPY20zifLQcSXJg0UJAD3a4VGCRATZgog8m5QoHPML
4ORGxZOzzvk5mhcyNv8MvQ911IpORZEG7Ol5DGPTTyzudA7ruc/98qPGWYOMUit+
Pst/y68QdLkdXOZQOykpMsJPLj7D2aLJatp8llHMWXivoS4CFGG+RYK+wQj3qrHR
PrX5LSs+oCfRBEg2RQu/m6IutXbOu/9fnF+dcwAX6BOmVC9ufHhfbzOSmC/9E/vG
z+Mfm3MhsI8C+jsut9NhsvTUUQsqhodfBDNV7MpEP9E2UjKuFs6a/v23HwV6Grvi
8XLEtU23oojUVQpnMAcKSnRz8Tc4CcQQPoYDNkL1NnFHB+JdzyMoRGTQ6ZIQe5qj
+urRSk2teAAr19NQe3lUlJUyU9Wj4bqcABh3oXUkzeNyIC+WUxbDS2xftg9dzC86
vI4ESJdn0Eh5t+ceCpPNLA1Ywtfo6xbchWUkQlwCQ58CAMYkfCLAEQPBux0bsZrS
Up3XGSLdhsnsqN1niUJ6JAlvZQiFgzYTaoWGg6WF+dK0jM0aRrCys0LTSMvS+Jr0
9aYdgoOkVjFWnGk5GTrcbfznxSdd1J8InUuf0rlgj3TVCNUHF11km3h6gJ48XWkR
QfkCB0Mxkl2pLn/rnoikuo565KTAvnm5rqYGHHFZGeFg1hmyupRnG3cMEjTnbazl
9jfTw/Eb4ft4ltMLzRbyDfFAn8evFmzUIDFO7RrjPjKZ7lRcf30lt4mIaNLm0sx3
fWoXGKXYltyQC64ocpJp5sLLEom+4oXOvc8Il3K2OlFM9V6Vx3+cfskyM9VSn9nS
TwG4x1kRjMLVmaP4HZl35K6E4pHntzYAby38hWrZj6VvysanUnNTnlpS0m/8EAlV
aOg/p8W6vDzDyTfjkeRzI1ya6vnot19+okJyIVO5IM8E1XrR/7WTIEZovDhViK/W
6yZOhT+LA53JnBemMlFtOefyEdsHxpyztstO+FglQ45nWGPjLMg3D+3DTKwNnIYc
7Jnc8/CKr3rOpCjeTeQGzlfyZNl6bgSngewayHJx6LclSOEkYm7TTYNcQzg0pqCZ
JJlC5rUEDOAZT/sf4mBk/DBsiPp5XOFbSYiKHUt7Z3GANmAcMDmpd8kC/iTQmdP3
SX75dmmWalAnHiT5GF+17nnOVJ7TLwcxg8OnK4RgfgllPuxxU8WtLIbUiRH6epzp
J9B8EHvRh+nyZzePe8sxPZyG9hvHQ5YQ0sU1ARs9r3JyzoPodFOAq5CKezXMn5Y/
l3/IRUknXu08wedaGiJ7DGls83w7XN7hSYXfn5YEHCaO6duAs2nj4HYRClNMSSxx
c6HnJ+dCtTCobsfmtGoOCXL3wXunQ2VUC7+3J3mskdSWlJg8ej/JCPV2ekq5Lq65
jEX2oOb1Bc4PsE6QsOdYi3mSSmsr1sSY2vHRZcQcyAaR79NUH84It6VRbIeEz6SO
tEDRxvl+IdOqg+PpgDoCB84ZJLsMfhKn5rVfWUTR20CKW86JvbfP8y18nkr01eOA
AoauPLn+j7mnh5s3aR128WMuHEtLHLm73cWEFxWs/bc3j4RilJt7l8sV5jsst+5V
x09UUlDZVGenCA2HdmpSSj1JyGs32y6DC0cFD/BtL6w4nnPW8ojJ8NvMCgay021t
d0uVeK05iT12KijmZlmERUnEKXw3xg/NfOvY/igxJnszY0Cy6kMCqIpB3rOSD0Iv
hbIbogq9xLDpFcac5sPXwd94EeVfvEsY0RIhmyvfxTRt7qBotH2FYbQkgUNpE3rS
phYfBKA5f6vHeY36mo2Nliv3j2zaZwfJwye1FbmttVSTzz+INERRV+v88MZOAjWQ
ae5NfZqxqOGZV4CAyG67RrYVC5Lrw4aDkyownjLzo2aLmLrPV+Wp3fwiNYO5dWyI
22LbWrXhWiXnvCYRejuKZeZ/ZGN3Ra+97GJRH5uIUvWvehtcpLt54f8c9RnRHHA+
Skqv3uprgB3Q8vZtlpRxGGzoO5SQ07smGbN8ID/fFLtA3Dz8KaQWptlIUUA2UFNe
O/UC0YH3FwfaklPDDmdA/2RmdyooZg979Q0j5zA5moDHOwtVZcARwZy5QstVcTPw
kvFu2dpjcyHdl9U/XeEyOoy17Nh8dgypC+ysupcwVvMcJWhc+eLsUCjq/caGKSOL
eTPIeXap2n4x++7hOUGLC2DFTfrejhIdHF8sgb61CaKBtWLLlzmnj7aOrjSzatTq
bOX3Z0urgokXBtspmaXDoS6tM03b2OI8bkI+RRnyZKtfYZwyvWyNYFRpoNTehDnX
DQQ0r0pyBEUEroZ7dU9DLl/0ABA2GBu2kddlZa4+F/90dH79buLi/di2leUW/Lou
uVxtTHM+pnKN08m2fBQdH9U8S0A99K04ylQt4n/6NmZ7sHAEU7MXuScTu81TLppv
7fE8d4/1TPGzBe1V+U0lNv1vG7mNGuSJgSpCMAficlP3InZWmzmn3Gfto/g5BxvA
jgWUhLhemxbxfH1lX9gF8gx4lvVPfMTjQn9QHS19ziaL/9imyKGDZ/ePKC71nM4o
Cvk6ICb1xnE1yl1XNFaZtrHkMWct7h/b9NB9bN1lIsvFdizse3T0MQpf594FOdI5
0pA1M8swYblM7aiKI6V11rqpcnDzO6DaddYsgVvvueEL6mXBPfSX/XLS0xb2Wgru
RqhgdKfucXeS1V8caVAjpgxXLghPuFFrC6biyIX5kwVicxKKHxv9cUcDgRRiBk1z
CMlOwXizdgRPVnJJWGaLm4PSrYtdZS5VbF5uVYibHl0RSfbIQxlPH7k23DorK9z5
xM40fto+ovLLCO8us4dSiPX5AtLGafMLC37/N719CuVD9nB+F/vShT9f7uBem4mf
xp2mpzEb5HI7cfJy6E8rJK+bH6pHvD5TrHc866iSxg8jr243sMNIniXjsMBemwlj
rqTvRtGTwOiS/SxzvIVPKwf3zuboKQh6NYlFpyvfTT5/TjMgOTXmpwtB6eOnO0c8
fMQ8bn1YPO5KU6g+8Z1mtO+brQj55wrvYQK9iZflA6cP2tZvmJQaoEVv5dFBv69l
aOCPX6wHMat+0iNqimhjUSqxLtzaturNz0k0FRDH2os/b+18bef8ltZbQWWesL4I
KzfB9oWk7gGpRNthdcKNdgcAaPh057/ygSJlgV2u1EdC53DaUW6VUDxe+LOGTgeK
Rv4LowIO4SIYq7Xvsm9MdcY07uhCKQIwRw5Wde49X+MjUKPheIRvCn2p1qn8VwSn
r1WvOAM3InIblA2fynl1178ATt9uAVlUJZIX38nRoW2tX9xO/Gxy74QWFG+bH7tG
8mz0wr9gPB6D+6E52C+4yWDHBkafnNiUSaAX93Q11m6rdOIWjuNfMDsdAw9aOKLf
jQAL6e7qG5ef4L0Gs+MLc0cdeRTWOG3+XLfmp9aalTPOwnqcGhuTGVBXugJuukkc
4w56ooMT8/COBysucDCivHITKY7Q/vohyILZQejMowCcasD2QeFh85VsUy9A2vCK
uHMAwztHuKJMk2DcSOYI/QyAN26aNSKCjYvOpSg9pm/p2iyHxdxFtMrh3pYVg2+Y
TQGUsU2RcG7T8he1StagL0wzduadZX4W1EWi16I+FPlU31MEF2ADpH17K9kh+6K/
skZ9XVL3TFEWd4FiUcNuMhm3Kq2XV6CcMUO0gwMQas4q96ljoHWX3ub3XyKKEkGf
6gO5nJZ8+Yr9mnGv9DDoEIfKF4XvYv90nWfIu5h/xSI8WTUE2qGjJsY5Rq6FkqdW
OSEzOmeFvhKJSh4IYm/VLwDM4XZjNoxmDGFYWMBoTDjYOmaM+JL2oSYNPVfs3WNO
8Q/vUn+CPSN5WX5OQyquoEShsRnPR9ZP6RPJS64OnV//0q3o41g6vhcQ5Opm2pyL
KEDXtSZ2cMmSuYWrOPrOB8D/BeUVWACi/hLfILL2BVjKprUrDgWdbYat6aPILwkO
UO45m384cdaTTPp0CYCm6DjVwqIiiz1fs0DB67bYwGw8rNX+yk6DWCTN4qGAEwUn
W+ztFcXIwryDed+NzwQsAzQdA2jNEItNyGyQdopzztwgS2GPtYsrgGIEpnqmuZOY
mY0L50/eeCB7BaN5kvG9xApqn0i0144D7ygfg+3x2FQal1euSPRg7vNznc4zAsBf
NI+XNMfjVOqV8ysYLAIOMF5XWAyytVaOcuOdLk7/NjdowSWj0AxaJqJUBXz/u60+
0+k0Zx+d90A5RyKI3pWRLWEGH0iDXuLmm8bRQIBr2iDPndQRxoxvpmbUpbM1RRLM
jthu07aMBWrwK0fLj0VVTxhdznK7l93rY/JSPa9mRbgSXDo6F740HbyTNV4LFQZt
ymVaOrYiolyRBHwZf71SPBiQYOizKHpKhpz+YVYJvpG63z3xlANI3lOUciDNYD/Q
pV9V5GOsbME4kmHe7wd8joeaMfWRQI8ADjjgK9g5ZjnO4yrFl26NqbcrYAO642RE
6L6EUXO9/oHrnuzyb9C/qm9btGay7lcQRYhDyxJAeXQEilU6bs6fAqWQ2DS98Dnt
Sw7dxG2EbQEF5Qz3b7hVeiCeaIV5zn38m2CG1Xhmb4zfQJq/HIHy+rCydv2Y2XYp
CUc4OeYJjf1vxDaGokjAR4cO1AZvGEFhz6zwF/a/4dicRWQUfQlYme9JqhCKwdch
1aU/kN2AROOVklqZs6xuLy3VHV1mYgGo3DW7h1g8N8DPckSesS8A6KwItzFcp6sR
KRnw4mf6bQaPmZfv55KA8+GzcusPkjDNzjbDimrN8ecBPB8Tm+viV7/ei14Ls7lR
ivOQuySamOpk/fdJjlpkQR1i8o6RSpU/zzK5MAMeen5K0Cxv7puVdK6Zj1YFCJ4C
c5QeS2XuvxQUg2/rLTs7dhRO4pS4aWi9uZV50elytuGqNTfD0rqmOXM2eZmi1gCv
dNEfojxYCHz3nYkWP16PfoeVAeDs7U+qcpA+NhXzhIFW9JQ4+wTTlIsRSE0YrJ7y
+houT+FxuNrGB1Jnoe3DAWrV60E4n43yDbetAHeNly2AhYYrur6AHBHxGQHnAgW4
F8yYFsOS9ChwEiSrfxUl0MicCiv5ULHkph0Ntnq1PK8pOeD2PYNO50ppYeNLcurE
FXo0RQfL36PcYeA9BopiufAnUxJtnP6PmragJiYQlG8zqjxj9nuBAIuognzINybF
Ufl5JiWViO3pjbOwd7BI3ACyd1Tva6byorXNcZ6/Ls7IuAV/P8sGuhQbHZ+GlMxA
2obxMoDgX/EP447xGTmK1n+TC0AH/u/8bGWaB4Lk7uBKr5Rew2ygTUVafvEUKEMy
BgR93oafZQTdLBKcv1Emskg8sTVVoEDMpjdoE4QBWEY+CKUzdek58ShSBRYHmFPN
NQu3mtI6KXzVj1c4rjdf1iEA62o/KQSSCUs8mjjYkiBA0xGf5QFfj0xWt2xBEo2g
byQi5mNCUMiZLpiyWKu+NQ60KG3AmHf80UaSGBZwFpDzL84/vn3cUowdSg2GsIIq
Zi4pmygJlqJTJy3L/43H8HnD49qgKUw8mrox+eEDiwfUP5yJNv61gyBmbCykUroN
UNQ9r68MYvaXsuASpAB/wiP9BJXeakKxsRXKedSpc5PGInHu/jmMo37S5r+aLUI3
RTXxD5Xq1kiu60LnxvduWIKEGVpSFkTFZm/D7odGcYPZXUIMduMq4QscD1LKDWfp
nr2k1XJatv2jrc0g8M+L/uGshS0SBPCiE1Cwh8+8oGtqJhIcRSUnF+2EP56tj5ip
zrvawJHQolbOdB0YExm7vWIBiYbI4INsztq5aR3hOdr8Xmzcv2XCYb9WyaI/EL2O
2GsfWvPfb5Dn8Q38H4jNNOA7x6itIeukeDTVNuXz2AocyI/U51j3mifnvCr+p9VJ
KE98Y5DUfe9KbwgXSDolql2Jq5PZoGfiFNB+Awu92AuwLBh3+EXl9QzSBJFrxqpM
jtYyVHVc0BQwerLCpTZTKhZIZWllu2rnVqY+gy+Nq19HNE0dlt0OUzBsJeHJlaK+
vywMdnDPgDTOCabLUJYmoo+ezaDMB46K4TfUtCDml29E+C+Rb/1GqZvKKGU5z2hn
Q9WRTp7pX2QAS73Ad5g5NWRXTMAWMibtqzf1O9UYXcvHsM0QS9pgt29kR0Jan77z
KdUor8Zy4MPRGqAd8EcfE7zHWXkCjWRPiXgy1onpeMhjllDyCWxYdhjL0+kUXSKy
fuwnpUSe25VqvX3uvCpU//BJQ1NHh+RCShWclae7D6jvSJGQ7WohNm37y+DA9BB7
OgfFaQV8cm/fOjMUq60RJ82tzxXvKMLrgj87oQEsidwesXliwPIjnHM44n0qdTFH
OK0epgWW/On4f28GWBHt0D+Su6dhLCFUHgn22S46rQ7A3iDR0NyvA+4bhWUL+VGl
rTb7iJ9is0hNbYke63MJ9Y2gWLOVxzvkZDPjWkY3rdLUDj2vH5vCSvlE4UCTkyOy
VCNt9JkKY9mVwalibKnASmmT0dZJd6T7QkgxjFQFr0YfnQRb2w4ba3b/7IlnFjoI
HoJA8uAqflYWIEkv5T5z/h0XcZkJEhTNn4XbBs07R9JA5cu/e+rO0oIt2mwh0/zv
MatZ9ndsgi0qjFz7fw/r19tvKG7lGNArU0PmRMpuNYUU4wZ858e8G16bu6f8rmaW
b/+qRXhyC6SrIGVLD+Z0/zAgcxEd0fZzAu7r8cKwFgCxBHrPmRAAJnvdTtEO7pXk
pwfie6XIIdDbOhO89ePPCqJjtHEoFaK+8lL+Cw2i7bm/FdjJkLw1EN/+Hvnet+B9
L9Y4SUPIESZj6mFEtw87DMq2oBeVCe9NwBovsTS3e5DlxIb3VLSIK4G+f+au/BMe
OWpxMkM0EZiiy0ttQ2Yu1KpPRJLHtwGkcF2ic5wSPOuduUX5TmByJXmCDmY/hKnC
ymtxTufTXCtypkiQqeBmxuqxGMFS4cT/eNr3QiDhrRjIDqdzfYUM3u2l3MYx/kmV
GTDBV+dWzFdfuVPauPQYA3qR8RltVBL0/DcgJ6kN/E1PQZqJLXOvOcgmFJeXV0Kc
MpNvE1qbzrN43gsTy0AUTtt3rM+hwo3p8QFUh8qPTD3YJVQ3LNEbvSVCcpvIKx9C
+6kpC/Zpm0wH7xSC/s1O9l6ZddAWj/Je1fXO7hgdbbtc03v62yM8bgAo+FuhG0EH
aUXucyS1d/f5vGTWkiYkqi/St7NAaj9wRTXEifdZkzTvHvMnEZuZ2YH7z7zGJMKJ
ssvsGcl+nXGQpzkusdkvTPo8b911Mq1Qea/5AScfsLCaoaklPRB8iQMqRgs9DvYJ
aTf2Z7MS/2EQnuno1q6NjB9G3XEvaDca6miUA5+kbEitVNDxb/XkXQINQBuvlRMM
0y7B9H3XYH32Mi9WKqVUmtGAWjCw6zS0o8tQsWz0tYRxCJzp/gis52MiLMEd1Erv
vnbTLP7RVFYV6sEsj7bCw/DHtTUNUrd2py8T0ZwoDh3o0AdX+WMJCRC0olLNsVbH
S3esh9+K4u/EWaVz45nsbTzoSwtp6KPbvOQjdkybFGtLL/pkwVQBPG9hZrF7bxvm
cZ0NvQsGlvXUF7LFGg+zNCnDdCaCToJKX/36o5UuaFE6Bui8k6WV5BjSAufXdyH3
rgG5yssggMuzfltUPjVaWN5r2Cuupe575zPPJG4Wa4rGV1fhk7bHc4yi0jlYjWfz
Z/RptGUTgRLRf5GVxo5XQCGY+VkslZxuVEr8DmyzXc45vsZ3Y1s4bZtz9KfjZ+tm
y8oEqWy+P8wFSmxAQQ8BsdS7GWq45VY41xKseyyk5RjyNhQGY1nP0JRWMKsCb7Kq
epZmKy/DqgJY6qFTZntZ0CAI0NZD+5LJKcWVXvizr+C+GuNVWd4IuJVKwitpY4Jf
IOcyAthsqgN5YSamxUjCPz7Gb+G1OYF6k6oBvTLNZFuCTexLY4Oz79r5sdZ1O3jo
dJs36LwT+76GJXJ0RHzK6qtxul/DGCNK8tOrdJQr7Vl68VrlB6F3ANnXXEVcTNZN
eW2OaaIEbK0Up3oamSrmJHZjZeoO286dU/78f076gnHi+WpwMJAEY9HvDpuUhAN9
fEcQxdIcEo/HsvYkyYKHrq3sbwo9fqVq86CqaPSIbCgYerfpZDedOMWlMcJ7Ewh9
fW39vxXh0LsRJnztJJumFIm6RFJ8RD/DZZHJOZpGpdG7ol+yMz4eF+cnhBEbAMaK
1pRi0HCuZHx+563Y/4+L0JAoW33UC9pc6rN5ntzHrH3NFcESRBDHuvuD17aCryso
G5ZFkeHBKLijLmE0+xqA3TW3d9JxAfzLVW5stk1GP9aDLpyNWuNCJSW/rSlY4HAq
sEMY93rvDV83ub9DFz68VsREK6fBkhLog7g7oWCRsOp2MTshhV7KPR07BuFwT1Xb
9I8neDt8Hmvj9i0c1wgT19V8xtseGoSx7tkvlnlcEY21/kDOnsJHDlI8yz9c4ThT
P3QMLPQqlZlXZxmdY0TiDIQX6s+jd4KICvRSsGoh83b73ZicDeMRt1gJ1GlRKDtS
zlulDPqhY93RsR6AUSPXCN5fcQRye+/7fpb1KRySHHUJuJ4q3jPS+ez2Q2AuhYZa
yHQ7E5E9px1fH+vrOlradt88jfsSu64G8R5SztRjxzdGHSUl+4Oay5e3nj4Czgoh
NJXzzcp45Wk52NLQKzNJiXgpH/K66YmFY/rtk+KAyjPR9sTvUykDE90P60EtEMb/
tW4seIsiGjehquxxd454BEBCnGfE+nUYp75kbUq7HaGS9FMwpfFcaPd3aQtcwkhi
k0Dhu0lWN6d1zIX6eoEK2XsBDM7O8q4Epqc8pL0ALQVgXunHyKhMfCKa5JSQHNMC
mWunqYELTlO/t7Gm6tYcwbltLalByK+E62QVLqZNz8PrX81CIGgZogfskWnIxWdh
S72XvH7sypCK6Uyt1Bm3fnv6Jh6OW2Dcy/KhX8NC8DIbMLdyyjwKQUwlrs5Xxue2
vlUyGGda8+KF2rNvi40sPDdjcyHyVhkSYEDB7ngpF/AdqkXySffrSPvoNmoagXKY
MD3qQuCz+dxGK6p3xTcU/LCtNBhBKmdc6/8B4NVP6FMK2qSNt+PVEXKS73+yX4QF
xbDBfz7L16FZx2XbeK85RsoGiwDf5R+WvLId1WbcKra5PIw4yn+5tiJ7azcdF5SH
7QiIAf3E+2i1q1AGH3RG2dDR2qbBWc2aZvsmrUznisCWqde/3N5C+FqYI08dTHig
3ntD5ts1dZARxZj/gqVXuCtBX1l+KQVdCxxzrvl3q3gBm8lIIkreGiC1ABaSBloK
n8Y4HbjqGFPS48ogZRJw9fmkaJcksvq+SNQqMaFu3oohfznntKmwPo1kCsw9Ac6n
mP+ekZ746kH7R6vJ1wUWDIL1BMfF8zTeThMPrkmyBxTFnZrwExeqP3grqOvQgYJj
W+0Dw8g1gUR0Dp6b5wyMduqpKcHGPqrLh53N3lRoKUnGR5lW/Sx0ypPZcmLH06uU
tmzcpb7DeTH7RTSnvNpHIJa5n2zwWfZvX1HmSKrBMRi0ZH2tnhQK8Z+euICK38yC
9Eq5mCUAfF8h/83IOHKbyYz1BhGWzTucBVhpUMOcxiFqFgWRyXFUiFECJDh9Pc+j
ffAjE2Nh0TnOTdEdAouVghx7NFGG4DRBcNXcTaiJDLJ/ZMG0FhZvdFSAzFsqAtOO
eV431qphaTGxQw2aOZcMyMYcFNTE/EDlSd5FBrqOkwZ+PVDKWYnbP3iHL9IzAmx3
rx9b6A7zfygmy+cz+1/b3RJi2KQK+0NXAoS9XO2jNFFuGJIKhiQoiYdaauz/MLbT
a3CPFXYb6dXgZagdadiWxPCVCeTFRkUi2BjDIWIztHD355husit1v0R9za5Q/TY7
QhTVsr2krDq9AMrryky+Hjq9zhhW6wCR7iTYEFx5KsfGYqycag63w2sbStNeCQZI
LYvWAxicY9zuwyHydKg5AEzxhNIVxGW/PDckMeWSpbio1vMKZ8/w/oFMjdqmOyl9
rUVZFr9AX4OIWC+nPRGtNgpfSQihwmUSsTdUSoPDn9Tt4FIyhpokkK6+mYxnm0mz
ezI7974vs88V9PkJC2TR0czVLr8K4e7K2AtoPxyj6dqM/Ljie/IhQQucgpKtMmYP
LLyqFBK9Nv/A2RlZ697TRO4GrDa6f7LekUKhU2Qhc1XjiboIAwyxtPdT5X8PGkAA
h2YnH32YJEphdSX/KjIaKR5MUZGROy8tzAcCRaJy8agFVs0yUf41vzfKb4erq5Iq
ZwEd6LZBBcOAAhBMme2sJoFZlP3meyXQ+mz+JB6r81d8m+KfzhlkQh+VPjRctP2/
8q88YOvdFBia+aHmktNGQFYC6IpUTeetZANkO7uTOL6lC847ubK9A27V7oqmiLRs
/aj+PXqqS1mIpkfvpN4acXonk+rcuzeF7S/msJlD8xrw5VAiXNYSoOB7/W3/01Cw
TNfUvPmJEqCMBGm+2QBdnRTsnN+968X0wS0WR/ysZ/je8dNqPL6UNat8IfMzo6IR
LezjZHhVflsTkphTjCEAbEous3xEoC6DuyBj2GaqLfzq2UadsTdB7uqwlCaF7Ysh
dW2XHpEwQklNl2soQivMfaPXzrGAojlq3tzLnohxXXAPWZ3ajvkm1CKw4OX9phLX
kOf3ecb1H7bsa8meVxICY/KUg4+/SsZD7nq0P/DAi8c=
`protect end_protected