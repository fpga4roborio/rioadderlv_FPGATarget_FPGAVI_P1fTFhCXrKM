`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
ddtXksX2+yylW5zu6QL2Lhnb2d1sD00763mmSITNX595NcHTEkwn0zB1Dry37fOW
FufOhVzEJp80NC5qZ/+F0Vk7Ik02dIR0elf3clrjeJRK85K4e3Hoo4xn7YbFUIms
l/8VZSb14+JVGURjfswrIyCUotIzlzVYZ6gzoZwDXIi5gQIBf/gI+KxNXPaKV+PQ
Ufys/12rjO6aI/pPlqSm0hCvftmBcnezN2hk1UeXgOIuKZnogjOsf0iJVX2aOOWE
6pD/psybjbnsNB6kH5uFTA5frkzIzkzl5d9+YDm9OyC+k84E83I/7/j+rk4L2dah
QJOvksSIzN867/4Qt8qYTQ==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="MvBXkzurAa5VTw+1JJ70nePUfoQXBvZOku/SMmg4TwQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
oRtzZL4VJ4iwysPsC8SXYCzXS8Fw2gtZTOskLcDV+1B9Nzn1zTyNtlo6lNICRmmK
ZRVu2BmCc2G+fmzynYlNTnSa7C0Cuel6FYpxCBlOuk3OF2tzAmLAuDyOH3Z1Yjzk
a0aHuoCdIRKv7BrZCdALt03JeUmXKPdOmIlkVGFl8yw=
`protect rights_digest_method = "sha256"
`protect end_toolblock="Jn9CQpRhJt4rnzZPRk+dOpzAubz7omckX1MrFd4p81o="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 12608 )
`protect data_block
gD6l00tciPUa6pDNTk/+tzLxvdHE2s3DQL3/JqqujQBC/Ei+vcAB8wM3doqg5vTg
mdfn9XB1bLOis2CVSfu295W2DNwHfMSTc/8BhCDRnTlLIX0UCJs9Za0+LoM0rMrV
T7EjVWppbP+Em6PkVKCwlmIQ7JKaifJ+Y+kjw9HCGboYo5074hY+K/CBbfsBQY86
h7FrhVb0BFNFA4lVvsm6L3xaIu0d662ZT0qZuL3hYMPrxcE0DAmAvQLxDYIkcFo3
9hw8a24aOj3bsixQuchUBMbPLU4grlfB0qpeIGbotQRF/+y5NdL+rLHW0dVPIR53
ExzrXCSg9UPlasSImtA8DkYfxQ/9SoTfeEOS50+uHIImBBckPxupT2o6vnwZbAyU
yFRGhF6XzASji2sDowRoqipoR95hPv+Z+T1GCcyFuQ/n8+NlyaT2YElLYzZgpAtr
hr3VU32hpiKRUU2XDiXP/rlLnFlBsoIAr96D5I8V1VdyGbt7sCOhyEFysmp55nLy
AkuNmSFYA4agwdFWI5xWfJ2YlCznFjtgOLbWCUy2gEJ10g8gnb11oFw2SuD8weRI
5A07rzKHMdIByP3xxdgPeSaZrcNHBPZ4P6b8tf1Awr/bkm7Z7zdCJXwAS7oWeERF
H9lDsrC4Jp5VyhHEQ7BeVP2RNVHMHblYtBVL96S8OfZWQa6tH7xEx4sDs4R2UL/f
03tRf8CfEESAlRMsWwvOwZyrteNPNocUGE0sHmZzeU2f7hJwu98w4p6OzqC892dF
Ezz8fEaogq3upZvCq19rH6fwXr+4oF3cnyXx9N57eXSfLzy2SoeWWuuysgtlORg0
HRJdUrvSOsWm0VPgnwoFHjD55rZL+Huw5cjOTNd0c5zg7+YOTZuO5Kt1ZzFl/ryH
/kIgAAFiPD21kM/ARDvL4Q1NfQ/VAdLPFd7VABTC3ZxCPC9/R4DYf3tgEpQjMV7n
95cUWwo69Z5oeUuypkldHylQgdPQ8efInX1MPGb+w4w0Qd11PRgzea4pFuFDXVWN
Tk1XUhUg9Q1TVB8e0UWgZi5Ob7uh9u2dApN+nxomFTb3X21gJ8B6UDWNTKZ1juBN
OenAvT79EhsSdZ3LiHIr8n0A/ZUhtA8Sy2PFdPGXxKRVagvVKE/1Q4Ei8CIRBfnw
0p1EnSs36d4RcEeTkuEIS7qLWaLEd0VOiaZZxmB48IqTT5hWDWvIF5taevabTKyC
k516/XWKgOgHEC5cPNl8zkOB+peWBipK0aYBCI1yQqD1HsZL/fJMVjIgecS+5Iyd
/K3kHEpDeiaL8HB4DcfM0AFAN3HOHNfRLXd4/Xi494otx0HSukiO4+3Yknma1iOI
lgXSN6kaMggNZ3nkqc3T00im45hUpvh+gBmo5WA6SwB4aSY+Ct9JRhwLgh4l6uD8
1mAzO+m4FFgNXHlXVWbPOqGmlta1RTg4fkeBmN0aMQNKFX6uHFpes0hudiSwha2B
Yemejf91MEjTsAD5+y1KYuh4ClHWMSKOgQYhzHILJbZOwvsT+ijiH87HtIgJM/gT
GzWsoYQ66iiHv4z+ZeKfdNmbvFS6BLjnyFaiOrI6jyOJWwlfNgqlo61aYrxMb4ce
V4jDw6bMtb9kzDVtsfb7zu6VYIqQG7FgN5daJfrrGTPK5BAI6JDoT4S/793Qpb7B
Z8sTmzGcZEelm6IZH8vzfbo4VlxuPSofoNoEKCw07G9KkatOhAzCCTPrYOwmGX8m
WPIXUppbW93a9q0eY6lcVOGJ70v+XzKJRSCd1H6lKEtdeoL1zi1IYRov1E2S5kZK
jgFYa/QZjlZlHJVHQcv8OgSNGd2eOV10E5gO4neSqcVQCs/H5ZMCypy9vSjkUr/w
ty6x7QaiCEto3O1IEDZK05uVJ6V1ub/HsvSoiDKrJqZl7BkcVJxU8OZjqUmX4pFP
9svB3CpORNW+HOqcj1Ttc/68ZBRlKEB8MRvPm9gcoo/uBHwZHubPFVs5HdWrHiJa
DcU5k4ZskCu0af0ypG4OHJ4HFXbJIteABw9FhX1fq/TqGGtHKP4Ja9H6VzVRm2Nd
wDrDM/6KutIla8wKVCYxGnzL25CR8hML28uaHJF+YcNmzmw1pJp1vMcv7n78C0jD
lFLr8wtyEFUDj6OXPgKbjr7XtmKbZlioX6x9MXTTmk4S76u+WAsudGAyFE2wVfL7
fcUaj0e5KbiCiLiVvEhYdoG9DCLW8sy429G5PUe/tXEsI06ALOdJ9gXSSm8DehCV
mJh5bmeJM99beDiegqK4bQO45itkyE750wqmcoq3IGbL7zzznI43dYuxPr0IU878
4ONQZ3F1UcPcpnGFb03BfVxXsHQ3QTe52H7YgnFOJSuDJNp67tHrMNfr0ZiS1x7N
fGSyGhHy+ItfaE2KspGJs6rtUEo2E7YPZIKZ/Hc4CQl6XsoL0xWyT+7c2xG2UQ2E
NeV3KjD64+ISZmkc3is/OGYPFdBhne49Rrrg0fIE8U8m6SS2Xli/2RRrRoFz4HUk
P0ByXWa7fBzKLWZ2tNxfE52vJdRw/gMj8lmqAzLA5whtNgOVto/ZLQp5EhUgH/L8
81bPfp02YMs8hsYSalsuPbHQkfNKR0tfHNn2cWF+n64gCGC7miOIy3H8i35XfDie
xmKL2Ih8Xap2n+RxYLjGXSCB7ftjXyUFFF7fVbv59XHiKFWRKfS63oa9WiM0nOvl
Kjt7M0hUWvVaKWiDYM07yx1aADNIM6i/Ia9Bg36nPhJeWHpvv2iIbj7YZTD4ERKj
cEVewuToNnckNUTGdow+1LK7ty7jso5EdQnMhZpIuOgO3TzBREFtHHHzgIs5YPOI
iGQAoDgaGR9ENc6Co8K9/86OE60WgisfJgSHK/noF5YmVbuquHIqalrHcRo/nxck
1wej+PvYnFhORE9o0b0EwYAOAimZ4owdOugRnDv8Ti3Q2eFOfLpWsOO7L50t2SwE
ci++BABGILN9igs42XVEtbp5zgBsvYFbwhXHcf9ZeYcuH+UYmJxqn/6KC/s5m+uW
CzxmUuZ0iNjeJDvxae4WRIylR3cXAKQ3AYX1zKqyKI3lXAT8BElTxE706ST+6kwT
VL+PDzqAEEoZjzBmcXzw7BsbpHW9Sb+4rauye0RDSIhu2NGjnqRdOl/Z26l2wdJW
ysAVr3lMWcz4+wdpdY2YH/e5QnU93r/irn170N7pIvAs2GZsN5JW21z3T3BhlznB
MAvCgniX15uolgDUzjHjg6hkJTM7TC/YxsOnbm8pI5FnNYRj5llbnM+SPdnCggBN
QPiDaGVrp9LqDvbZ/wA1cAXD7C6mrqTKw7DjyYAPLeBq3eB18XnEbSHwHnUOOiYu
maAE7+24ooqnAZqBfkU6L7YzfpM2rY7ecQXrCCE7AJXYdRr3ng2omrvdA5QY2D7p
yJ0Ww6rr9RFhOwiy8iOkPKneHNOO10WHnHjPDlrGQ9lmQBIEjHrcp5mOcMUePkRr
hjByUBsj+yYZXGOI4DExetCNZSW0KyufU9A45CSew+P4M7PlglX096gc226crnQC
QkQ6B96CAGDXWwNLgYdCLbo7XVBldHuqdbdELm8B8vpaBn2Rt8dB39MBQ7hy2Bjc
0Y0r/IToSyN9K+SFErfw5hmK5W4wOEnmRZjHnVRdfCO4Z7wwND/o+l0c6pcOsv6i
8e+xygDkepb3/DnVXJMqIMYtvBkQSDcEEoHBy9Kn8rsgMU2aG94xQ7j5iFDL7BsO
RzjjFA9y5TyQkECTCU1l1bHDhi23SGhINHiDq0Ju5lOJKDxIpwjOqtWowXLFgDlS
lqeDiKWcOjNDc+pxw8ttBk2uE9kbJIyBmzX7rtwBC2YAwfi36fDUgUwvSQhQwZnG
pIRJFrrUQt6hJKpCbuNYr6VaI4uaOnT3AoiRtRiIpbxgmKWIOHHsVMYCuV0hNLH+
TWhwh/5QZac/xgwgq9Ja4KZaTcLAO+4eEs6QSRaof7/Sg+WfZesVDNAlyftyW+d8
nGPgeFSQPEZeFiJgFFV5UX0CXvNwj+01U3GsKC3IOzqprM4ELcLiaLaq2qwSX7RP
tjWFz97SicpLdZCuXFTT0NgbZ3UhmmYwApC3noDbdF72qf4jFtq3Cl8aB3q4hDnd
fi6ZJAozJXqFcsPz1RMsGGTj0VlpXU3e+hQkxl2Sg4nvRy7/kNNxsYZuv65lLkOO
vbXxw7DFb8oLqeO1J6/hnXwpU/KKK/NVihdx8l1RZCpm5r/vXKJXEAB3i3dnhm4Q
Lei2P/R1KF2X5/U9rc9qu8fZPbNE7VIgtcKw0U84zI5lgaAHYtDkvaY14HKzdSgB
tZxCSG3auhZbevECPGOS8nSFaFJDPEMuWFLihqbq/HM5B7re4jLeHrRdDSq2AQTD
i8goHebzCzXK29ntbwBsFQ3l5B5J4IyExX5E3IWFnQZ0xYCnT/JKJ5pxihswmHCm
wHEDyY/3E3BAJM4kH+har6p1+NQGOKS1CursOkI5ZIHQLeFtQoWKxgBD1C8ma7TM
A6Pjk/UlsJEmJeVPYbi4QWDhliTkU6Fe5VhHI5feNwjQkuRLybOA7rA6pl5dZNjP
+gi/odD5j9ld3+wP3nybxGDR/69yVoebOM558m/kcm5gS/N5VvGUfgA29XQxJNC1
ALJdijyMGG7dMDA3/vkOuxAEZG9Nl+k+YCIIK+ZZNgUMcUCgkcVjkk2fZ3U9iwy5
nwW6QG+l4e9pMuUNGqgKCUXclpeDS75eVVEgusXRMYA9hybSzalEd/3IHo0C5CQF
1TTbT03h/oi1IGl9JwyMJWbKOEEo+Cdis/bPtQiRaFD07QEcLhuEpSA0cIYG/pgs
txKURgl26Acbo3ru/V04ox8b66p0RtNYD2XT1BzlyurgwqYK05iEm6edncl3ltNq
kXPH3v2FHjqaOkSD7xSdzZ/e+meoE8nZN/+7Ozt7AHUtpzzWgpFdhwIOtTj0Irjr
LCY4ANCzBBdDIeITTqtFsKG7kYv7H62qyFXZJycPEDVdWo00XFrAy64uTIjjb9es
tjB4Q74QN5FxxMw4SZM13gpP950g9GoRcsoOlJmAzR1kQEL5XbBK4pu4nRgzk/YU
LJtbQxUDoVJrQXZLGbqQI+yrGRFCCZvbz1xZ5kvf/MlzHzgefez3UMss3ijR4uP6
ebrmksIkPRubJ9sisVY1u11YCic7ndafrdG6e+Way4VL8MLe0FHusXcD67WLDoPG
nzSUlVyOvKTD+7TcGHKJfCGmoVtALauA5kjeKyefIqPbqQp/qhBvO675Y3fTrv8F
Jtaej1/ybAbqv+3QyCfaEDuOwDBcMJbUMTb1eTb3d2F+zmH7nGOXSX59FxDgUQG1
8RYtLgVBQkdfKphTxQZ6Rvkg5KG2TBGgRdsY88UZuNTa3svhjOczxTfHIRMpnums
KasZg+SgpiSEnKe7fjYdNYglS+HP84g3wcj5VcHoHMygZA/C4FqoFs0JNrbaIJkK
ygOXAw2D1y5Lvm7bnA0sU6+t6+jGlZrMF0KAnURHL2AyNFQxbuHXxwZvqe9+3OYd
guhnqt0PNArVLixT/YSow6F0qWz4ziRecnvIGv20EX0Qoy7ztJCz5WDjrqo0g5Le
aJtGLC9l1PgOgn+FTCzZbfal6CyyP9QtVALWR7fMteAAY/b4YGWxPqgWQakK9ArX
J1BIIpDXk9IWxIC7eEzRyjeOqcgLN9CBv6I6CZZ1GBRXMwLYFxb/huzs23H55T96
Xlj4x9+0LU/L99hZOIOqJQvFCa3Nl//M9RWBpNFz0JTWd7pGTUFUJOszrVmqCp90
EhwMY0vG61Fuld7jXJIHlFboFAttwbPm1HRAHA2cT5i4DQS3m40PDj2/k8ux93Cr
IDEm7oRumdc1r4C1BMzpXx8mCWaxuXoJ9Yvw7iWfL+HekSDmg6ENbX8VMjMbekM4
oS+PaSmGb+foa7DKYsPWf5bocsjeDqbwCrPdRtcaEE/ioXOl/zAMfmLsuJ514OIg
appiUz6SNQ1HsZabrwu4g19Vslfy0zhJgvQ+78kjGd+pBL4V6bKFHKKJuMu9skZJ
r3l46DwHCDi5Cs14ufZwrH2ry5KW6hC1Hp0MVpLbgHEq+TLPLuWniycZ55XxeMFj
OWrKGw6cOIvFgS9MyWQ3TuBVuha4W9dP+hteiZLI9lCSI9pront/aiBIo9X3SFko
AppbCAickIGEcC2axVeiTMk4fBp/1p4HpyTE4nkcWH8xPw3K0/hYxOC7hJ0NrIzp
oX05aOJj0XEMKRHTgdtCfIU4KBurJIOqS59wt1VYvl18ttUkKLkW5W3c642Y+SR0
A+vvWnxqi2YuuS1ErLld8rWKIugqsfoKmCXzUrVyWPVsmaDdn5UfCAkKLqpCOH83
ogs7hw6d9vGm4mTM8G+mbUtEq24ogStQN+cnWqEUSjlY+Onz2wGP+kDzIRT3NX6J
O0tmILljR611Rz+QFfcdVoH2R+/9CkwwZm+UVgIiwXi4igOfzpT4uOW8bAWJFCnw
eaSzfEQgQgGubxYjhuJRGoOwn+T6vlxchry8URWedk/HNJuCztMzBKDIH8+hpiHM
1BQcBWAZ+WKr3TWkuc/4SkFX2JyOMIYFZoj23yciVkY6n0OrvTKY3GqQuhmEEDsy
K3QWav7l1I3NvBO+lJJdk8UhflfoTMGIkXW8y2tCaZ6H75Fm2VUr6wf9fuAMRdqK
46FQfHpc4TDY0tD0pfhN7GUtK6iboAkcRhkTolN8x1UgIDvz1gmqLBCGcaAvGoEj
W+QiLA8GmKg0vj+vmE7tl+u1XuycSQImAaqCs1vbIcClNOZW/X0SsX/G+B2KwQnV
nlLOVc95kN+fY3mxRCxytcOmbBH9/i9AvMHVAKP2drZiCSBh66LQ2C33K6aj3YCf
BNCQhhr0T8+vcfZAwhrRZEeBiu9R+dvoUkgWPHM8j9nxexARHWbXwXTHg2ZZFhL5
zBmner3pQnVG/+CSMCHkVJtFd4oKyeLudE89MAfACrk0AmX6yvO7x9T9KzpRvuGX
WPzaa0oGjEFFE4xYoseiIUVnSdckY9bi1QA+gPMcQxsdVDVWgHTDFzhFIJRnR0h1
0ggIHiD+HGmaFC5HrcHSD/k35Jmr0LHFywnprzK4hLE/xWsxPU6pjIuCujwKTbX7
lPxT1hIhsmxbIFl+NiSc9x4G9FjjcRnoE45dF4xe7Y4rFtuDI6wmxRykOtpkTOg5
DZF6G1KjSeu+JrRW41S7MNXO8BHSdkFQnjKv4Iq/Q71w7zMNq3187yPDO3XyvmYT
ClksonrYh+/B8JpjQJ993OWPh9/t8Zts6+eoVyUVQxprrzKVPm4UlcdIvYxuhTjA
29gINP66WV8jjLYSUWxR0LQFheNmAPdnXhSMUoyBkdZQTjp6ZNvUIYQBfcG7zorW
fzz0ZgYiJU4eLY/QgkzPYI8kXgTOndmeihy90q4xKMvR7N+EGCxmsi5RpKSkMm/s
bAXzAR2OSX5ZaCqVPvK/SMeOKyMijLk9OZqS+9Di+AX7jAZvD/NIPv0iwtnKNgvz
Bq5kQ0TyxQ3ODyGLPQZJ0nWNoqDpV++DnQCqCTSG6wsdVC0m5Ig/i0LfoqVDbaec
Lfdj60s+h0mgQKCV4afDtaAN/lDU7DxAao1k0F4LdKCIWtvWPdLC24gj+xLVZZqi
SxqgPQ2owYYtjk53xrIThaPLFt1ofnNPocdevEuWfCJEWBnPSd0p3OKrBSfjVfwR
/IZK9v8SA2RZQe4IKaafxBO26xpoG1vTXaCnnwQfDJNzEp+NHSvnTGU0pDlizq7V
WLKCiexmZA3MuGHWGK2Mggxys+OPjyxbwdc3iCed1Tsh9M0/wPnfeKy4ehRkSS8L
p/wq/yeCj0rrBd7C7OBRD87IzSkVTdXPaYwnC9rYLz9gN914GEq6L8C9ovZvwePe
r5FLrCDB27dXy2iB+ugFslh3N9y/dxDSUoSBwv/BcR+VNZXLekrHSMKeiM7ePDMc
6HXULNRasdIH/Uo1aNCP1F4kmcj4w5sItigVyfHHNk4PDvoBxj0nfI0eLtytnh8r
ckNLOrfs2WxAuDOklAVv9uE6j9T8bCymce7gxo4Q/UhCF2azTVdW22qwKbLQlPMW
x1TzkoaKl5Ug798fbYvEzB/HBnG/gddX2IdJ7ITmbymyUSntCyxMQRXywYVhFoFl
nCAambdvkjGQOEudDdhKxUT1gr9vJKL7HOhDSsjxvkoeU0pkaEIe6vCfF2fFznii
Ef6EGe506T4+ij7uCs7JPLgYSkqmV9MgSA56gfOby/TnO5klNfSdtjZDYkulTawE
FrQNM00T93m1dA1xBgBhfz9QAIhE0LeOE9wk1JLXEK+2fqZO55c+SKS3eMJFOqR1
6MBXbb4r7fEbF3k0HuFAMYqOXbdQLxYg0dWW/nVq+vXM/ADC8Br93XN8NGyaATSR
aJ98G4Dk0OWWfwjmOzVoe+oVShPxeJSLwqT3utO6EE5s8xrnYZz/uaNxMdgAsOq/
05R9wORtORG/m2c2Bo8d/rTiYPN6Hgp8ozcrTsbrURFN1HDpSUiyy7R6TYjyIl4z
EJgZEFlf9OGipHWLPXJ2URaZUzqkSF1shoguqTdSKVJGus3de+Yeb2+rc14klQS7
ToJpDLSQNz/NM/NlWERiRqE/7a4amL9t0TyvQqHs9w4m9LjjfI0DQOulB1MgmCgs
ju345JbSFTLrBXkaycwNeM5qYhaMx8jo0Dzs8FR+/h0sVAK1oAOZDmNE2NgK2CtX
59TVvg/822LLdkcD1BT3aQPDVCBTJh4h5cAeHy1hu9YqHwG2AGAys6CTbODx1xrQ
bGp5JbIvisWvQI21IskGNzXOWjAxyzyBRlTgQuX6Rf1jBkoiy96tu1875fcfp4mo
uswOpv+HBP5RNPMbLxMzYfMtBbdLofquNh/ZI/UrCViVUNRVXPklleWNXwhxzg+O
4pIfI1bT6jSJcH8Tkt5j4jdUWnUrMOiX61qElEqHTiMrvT3eLQO8WJjeef4PlP0N
nf1Nk8NngYcRfqEXCRekxIZWEPhzRmfy8SKEwtMWjumqGjljnplYlqA7LBYWUEgK
Bz8S/XdyuiVIWvcct796K/Z0LReT1cI0HRGYjHH572EiSvRGh0h2Ys8sztuE1Jwt
jQK14C+OdeRC30JHwChXn5XnlUc81xKTU6E5JTiMmrFu6NahQJ12tQfiVUf2ikrl
3oxBJy8hua0gGUgo7g/00vndJH7xiFsQNONDUP6FeM6WJXQ4EO5PdD8/xPgbmbQ5
bIhTcJ7PPPh1Sz1ayjj2IMk7R+yDQa7W8/CKubtgiChXBsPkSQ0yfiJyynK6BmL1
dDwHB1PdvZtCETcIq6vy4k2qnN/IjS6fxztjyhWrYZQCDcshOhO+/7K72o5VbpyL
1cy/FKxqvkQU5c6rToLZxxgLUIYSKyXwgrodQAfTR6imGpEUh/vJVzf8kK+89mEn
WhMCM7m8nxfHVBryRn5FQaKc445HDnQW+bEk/dxb2ruRt4PD7Ozhhe5M7mbp5CL1
KAHbwEYIRBmPnJykpzcByl7aO2hjdLUNLY7HGSHBuKUM7ylKRlRGUIEnPZXSSlat
Mt1hntP0cxFuzehnOzwFm+SnFCceGkbUipcAHhX/PCHc7+J1ZUXP0nRrByqjJfp9
11r6NLarSHBu5HpERuyYvp7ufUuJoDsWQiyETtzfvK+MvC9Te2vHPBQBQaIN4I5i
Gjo9oaII5xvzIrB1UEDLsOK5Pe3/BF+rIxzzQA0cKdieqzJveSnBEU+QTX/YLD4r
N8haslLX45ibNcCp/ooOHjjbDSGJeBeb71QsGGRZa6miW11b8keK8y0b1kaGNOZp
OZnhTuwHz0l4iFVOMEanRaaG1JMokWzF2dfz2yFfjANNolbLDGB1U+Ujw3nCS8Ec
dBYLkS9drwRyUKVIi9qgLNiATcT8BM8FtaFLznbV0HE5T85hmV3mjrt0Gdroq3BT
nbCUuOCfxrauNdcMSM0nYBNmpI6chV+8xAQvwxWZwa//ZlN5mE/uyVNKu19goh+k
8f3cOgQE73f/mzFp32oBcNf3Tyl2zXRLXDtsBsOIp9QHvBaCdIhR8jZojt2Eh6er
O2mAnidysCOX6l9L8oSNP1Wmys/QDrhmk+gIqr4HRDOhmmuxkc6kh3GD5P+Ai8Ft
gEbqDkrWCvoxFDdzOtBLmn/GH71BIzwJ9rA2OeHAuTyq1k0RCV7PfNvfKlawc0+h
HN9jvpQmGitG7fBoyox5Bwi3NdB12s9UX+Wh+3mFM+0M8Q150wBRk5svBQteshe+
b9lwXPRL1jQjsNi8Z7oZjV7kXBu0zryEBq2qFM8jj/6PdOiPowhqM5zbdi6GQ9GE
0zsQMCouNu5aAtQJbslhcIYdTYyiyFQS5qLOqRnv8xNkH9ixbiV/B2ERuonMkpRx
D9qGgDNO6sbcvER7ix5JjNf8QiF9WPZbL6wLpnLxc2CTyTdti/tIl9S4pIjClZkn
PGYOLVbGINwS5AceuzlcaVNFX/eneT7Q+4PdMqrZx3xM/kaQG/kWa/jK4Ue+J76H
4J9BpaIOzi13nJBIROBiTI+ws9eQOHV+u29wfFwSO9cNLaW5ZiH+CvufhOZCnL11
IVlRpX599kboFr5YMdRd0dTcj7e5a6Md5T2txSbcbfF8ylDKnqQ/SqLck2+6OIt6
3r5HakLtL4CyTW8GHKNnRyeGZvZg0m0g7FrXQIOTZ7QKhTj9zTMHqwQcpW4wAkM0
CTf00LOjlRYL/RK72cDb/SA3bV9mnDIj+b/lFrBUk+grQXZa1ZXkTEkbN+treLV3
mHxu6AazsyQ7ZseSXXVUjJq05mRYtVlMl1GQ+3fC8riEVqFSBuKeES1qlD4KH6by
s0KCZ21cBoRD62793FkP8e8iZv2XwAKtAWzUIt2aw1+1C+DMfIkT7mOMg8YiTqu+
9jFFrpuYOxAfyfCmFIanN+1cmox2rG5biK+MNKv93P1G+xe4+xYHRkgzidUZmGnJ
+WCz4BCwuxIDwrpZY2JGLbN64fxwusIa2m0e0OF/6OoSVreU8LUGpobzrLiF4FF/
x5NcaFSDs8qD0SjigNr/tY0Bq+pbC01dSQOzRYYqk66TOOHZXDoHNj9AqyZ9y2bF
lM97Nil2lQIZpnosg1klsXK2fRFZb+cAjaHRz6MlmMA0KKWNRxVjdmDqh2Uo93Wb
dF0hrIOJLRXTI4rM6TXOe8ywAggX8B2bUQy1nC7JcJI7DlvrsU9VA2TvljgT6IJV
1JIKrfotg2A8cgSwdowhToNSqTfTT1BUX1MxyfByk06OujXIzsHgrL6AJXuCIP2o
0xqUKO0UAPIJ3MgRvOO+ij0INEomKvY8168vBjMXM+LZm6hFrZ0tl9PBDkQLBFET
wn2n9nwEwbU2H8XmHoP7ck5tzsnWq+PT+I475ldkduGV0ArUSXo86JT9romIY9B4
xp11nWlng9qW5MDnJexRSFFeZl/dQDDjHG3Vc8k+QM/vowGNYq1IE6YuibTJc5YS
ZzxDrKKDeD5m/+4KsJqeMlK8awYu548vTmWYigSDgtiGAqYnrj3ae4YGzKCGGpfF
mR4vRuc3yK1JKiuVceP6G20HDzsTAxXF+RW9Zf7I9LEcxixypDYg6D5B9SCuiGb6
G6zBFGhah8NI+MqXaj7ONpPmtSBBEZ3S3xiS4yO7Ir3E+bEpl9KTHPtgXpVGl6xM
zO56NUCeG9FrOOrmyftNr/oy5xRpUHt93qBnsbF2d338XgfWvlG2TOKv6w0cU4zd
RTCkNl5sVbXH4cpUP/BiOabUW2b7gdCzotTsxOxAJjQzdnL1UmKcEHHD3J5F6Wy8
nyd91xfYwrt2SFTaEWrLPu7YJYEnTBS43EE/0Tju7jhA1RlLgve6loZX5zGoWyAL
Mu5Nt0/ODUxyr6/dAVeYVSR9BVuqdIW3mqAZ3aY1teIYz2MKADls2aVJxrCR33RT
cZGu9/7ITNV6xLgs7pdn+11YuFKITeS+lG1Mr1HxPJT1z0TKJlhWouFiQu0bWU6E
mO/gjaBW4KG/DGm7FtKZe7+/EsVUpjezsmLkBf5E2p4vn+6WR8hp4j+hVcfL1hGO
QRCHpNTNRrCqOjBmuBNULHoZWWqYm5/nxantRt7ysPLGCLSrIZajEatLRYLqO2IW
/KdGMSZsM2Bi1Mqj2nV7kTNwCzxSkIFpf1DKQ2KEg7FJN1wRJS+trqFaD0sWE2ZB
+tSh9kKMd+LIFvTrXtH4U+yn1kdR+10Ouk+cRSvp6mC9anFn3kWite/4XqW7e7MJ
lIem211eV3k95iPQIYOx5RJ0y6K5UnaCpS/yHSmlw2F6TBYZIMeKnm91ew+3AzGA
nve10WqX7KaeFWIMkkz3ZKlD+z3R6ygq7Y8854ruhuxkVZmv6YxO2hNdyvoHY3u5
WJaWgEmXETUE0eQ3l84XzfKMND8V5SvknZofdqtzonl64O/TgbxRGTKR6iwA4bAW
u+fC9TETNa2UfoNiHF0gQp6n6ELOzQCJ4fbZ3jAgH3pFfooBbMBmd7GZQGpTrpXW
pzRsHmYXs4ljIGX73gD6gkgSijtiesoU9LvJFRkJpjomVZphmmGocoAzFa42na9d
r/5pbF6mnzvYWmnWaMkpHYMVOkyOtBqQDjc5113WI0SbVDnDVQ7wSJ7+0N/90+Kh
4R5bK9B0AqJ0GKYMa/e03GAgQhz7FizsLO4myiuc72SZkkyTf/jaJNr5Veu4MFUG
+HyMv01YiYveS0dOs0c9+J/GGI5bDinnsx+aKXbMvMT2mn/z0enHG/WW78WYpexX
htHCDVM4VETx3VCbJy2ltp7S4Nl8D4xOi8Uhj1nXBux1V6XYQcx5vrNEeuQ1yUKT
6RgJbgAZI6dRNMO0cpv/fmz79q2XkxeDOkEeV8ziYf1/xsjf52MGwzckDtdQpmYR
5fPHM4LT/L1PfUq2aH9PIjpdYVuEUfh5YpMoRJmY2M8ubcHtWnM36V3OlGoDWAce
Puon2lJuMInoJRQqHtTVVcP/VWFNy8V/K/qC7LXrH5qXrHex2OuGkQ9OfS+rp2oa
jSDF62ijmFWf1oLPM5UFqgK4YkJjksr4lXNkKuSE7TNI5eXIH/0spaIxGCtJ6rJi
BwVSt8xbmpWq0W9YhNYJ0hXimtxoOEsI1R+H6bS+HPYxe1EZD++xkvev/mR91Fvz
noBfCdZCqsnZ0+klEo45twRAY+WqmbA/HkGoVhPEmJ6AH+OntYwl6ZCoTmTXexAi
bFEclRwZUomAO0GeVfoVFl7rFIs68/5jsWAtXOFq2QyEOuPoepmCLi/0MG9u7ouY
KS0ibeBTQYHyRwO/zokTibkMbC9pitaYEoGqjEzuQtSV21BnLOtmphQuWEW9WJBI
WkdO84SdOg2BjvsIhFao2N32omGLXLdEhnCo0axskR3gxbGYe4wKoR8XH2As5fK3
xaWsiFsCUZiN4HpEmiSaV38UKzkLQmiy5EZ1VU5EANO8m0C6e1ULOISfZ/ropkFH
e+BP57bJgDhKsZ4FrTJIcdZggxnYQa/1U4xHk/3NQYsSax8jOKRWxkDZLcRRoM5F
UeTokRWqFn0kuWru5nqUdNz4bMxuG5OzEWdx4vCGxlnyBt3Mb38CKnTT1HCB7gxA
3iZHBfLHTcBUaky4VEr5kfPTd33MplYq/BFMBw78q4uxrTxSqNQA1lshZR9KMImn
k8sFHemWv+AqsoKXTv0+5LsnEtdGEnwYJMukInUPSlq667A3hYGyQaN6GoZQ44fi
/qmFpmCcdLD6naXzLcn187bJ6oQwzhHnDQWar28EJGqyqMThtoAXVI2hnGTyzsWe
SBLTSmDbYev9sZuHzmcyArU0wiqlCMNTED/i3PVZi+LCnQrUmKcydPCT6QZh562h
/d2jFNiMOlWF6fCg4tCseRF9PYUJ45xYrkxOH1TzeMmB713vbezbVD6XF58AZmzB
00b2p++15XeBjkX3YekgvA4IUkSa65nkvAWtA4Wy72zG/3LZsgB6ZG0iirSyx00r
Q/yraXqC4HcknOxGOia5jA7H8jgiEjDPR1AdKWWta7E7o1Bx8Wpo+ehHdL+XpCt/
B6K2L24kSd0aMAflkAuS/dUz6/PvUC8ch+ylO3qmMW5gtFsrSn7n2SLW1oKGarqm
YYRSsVTuXX6aUGO+eGdWPyLgfrB7Idm1m6VBozB1Ed0eZc51hinpps7oAPYWN6DW
ksQj02jQpjbsy4lx5+8OgKJX3KI8YIBvnxq1pLqDBg3bFOhStmlJjJ3Enq2UMIUH
+cbJmLkZZBoVe1ZN6yD/yyeXiyrzO7hcxuUYYHI0nBw60NdglvGu5DOPFZJw/tg+
AUFbz955LHM+u10cEkg54z5BdU1bog+TPL5Ly8hKqTk/591U6kuFvuBVT6lgSegD
ZO4iSlUW5F5W/mvuzHnOBCC64g8iTBRPMXCRXYNcvgob1UbpYo7QMIodKwqlJmrH
vtWWT8lkQZ+bfJdAxWzDpFiqUGFYZyX3lsm7+C5EucZnzqtcbf3QWVUN6wHt6vl3
5loC4kGxOIn1rL15viuNPS49KnjkAwIjfuVBKt23kohve/lrmjEJtz06GNd+rsq6
HnPpM8n4cogQSyWWsTMXiR0GLCLl9ODiYQbeQftn92ognN4lZZt/GvgU3q4PTsst
MKeQmHEUgY9tss0Kjuqc+Rou53o2Dzp3EB7qKN5IYDAFoXrOq4JzpFi2ZQap+5HA
lIPFkVmfcPVNZt+c9LEE5B7ahj2TcCfmXU4ma3jpIf2gtAdCamlehq5KtwmeFM3b
neZ34kfKkDMzZnzhYO9h4E0qxcm+R7IwFTn6gQNO2qrLXMj7CRLu9MB6KYh1kow1
Q2p52RI6KvlSX3MSIy1yml5/iWgdbcOp10sh1CllAyGtQtgVFgXWFuUHyiU65Mxj
PoWzbnjQ582P6/R6sQJffEH/D4PWE9EhVA2U80aio/cgDRi6Ntr452uy7R2oTfOw
MGNCDzqlRp90adaN5kJaA9P5ItKCdRbuPD69X6Fvzhq+E4DzW4hpOv+a5Xaw8NSK
vO+VN0+DsB5zVh4dI5E6EAy5rrtKdgeB4AahzhBhGINHLrDFIluq8JkUT5Fr2mRK
9J+u0v46QDVBqRvpaqKnl2AJOBC7vDdiU2/9CB6xl7graafNy0tWi6tumMl+nsjL
CyzyS6Wsdj/r8FpGLFGxdfS6sdXuKrN2IM8l+15Wlmbj+SEEXkXnkO/zrhlttKbP
19Mm8xttqGnLHqfztpiyLicLJ+T33uaFdTzm6m3Bzc9LvTZok536KT4UU1OLFhYl
j5Wn0VmuQclzm/W3BPdBvcd9WuGKuMN8Yi7yn3pLVvadOo+vXtVSGO7qmpI5nBm/
U6KkWmbbLlu8Fa8fCsNzX4FvYYLwdkatYIQ9VGEJ204abWDnxCv6lD386xD/6s6/
Tl31CyLTJEyQYPRIMB94J5FZZdP0H+0t5SrFbQFQy7rtYx2MpaQCmhwsIXcY+kkV
5zUHw8mxpf5WILXSvij6cqWqCwMuLMeZer9/0Sw85mrugyhrN8Pbm5AFYDkLOy8b
WlkPUQDoGTPZzhRgo6f0dnHzm/fO4WCtceQdJhJg0AgVPyzEznxOVVhP7hOguX/s
PADlGMzCot838EGlDKLMa5LS+HWzd9kJmvftvR9Quby2KWcIsu8ayLehzwis5UXf
wQfn1NoxIY010fRXLGZW53hzjfMTL3UQFDkXwKtxU0nAwWuZMoZ97+sgc0nBSwBq
5EyZ9MCLHvHFgeVqtun9UQPIv4Yi8dS7QVUnjLuaZ+/N1zbwuHBQm8cPATGOyUy4
WEIK2CbGDJpuVDHxoW1O2p3U/jjdIrVq0Dzn7OGFhfIT7F7ZWqnLsek2LEtk4E+y
0oc+CfHVPCfJkalBp7qN5hlX9Cmsi1hSkEXvop4DgezJ9TKXIUB9HFSpfNm3VEFM
uruXz80rq8Yxr+9mdl5yj1mhTBGIj8g1HemmwWS5pkvuh6b+hWed4HrM+k5shS2A
P0BLQrlXcgybo+gWA+/5OhW81NgcoQ8xcs2Ns/e+xOWWtPmDtn1bfh7yyiqA/+r7
uH7ezXNP/5Ug72GzsEoxjM9l2U9Kbk2/DjLVROqwnUm2X+S2ObQbSj7MANNboduM
xOTqnbT+qYDg1bgv/lIG1zMe3UgU6/w1tajGSJJ8yQ1gRzx+nE4rDETVUvibPv9m
FanOwvbQwXnVk9y1BGzVQGxvQcQHPusfIGbAIuM1jQHwkpVK/M6Gms2EeUm9hOxp
1/kXXjFF/rsTN/NINgsbQvBSmUhFKMBBmU1zHZg01JXu48QFUv803MM4DBcmYR/L
LgnqS+9DjLG/fzhD3HchMEHy8THX2AY16uGvML4pFYmGdeTo5PIFEORovp819OUq
4G0JkZagr2iKulpr7oD3UcOfo4NHH4aUxzLyd1V0CtpQoC7DntUk0+FmlbwoC9ly
HKJnMHQfVaC1XVvxuU9ozcfeO5i/4GEEZrkQTVzY8+rj4KZnIvfJavpQgqkwjI90
XQvAw4TYg/fUIydhUT3y5YuhktKDieFRkyw+2uJadjtbvxdn16cHaww8Oi8URWE9
iq2Jdxxz1wMNntsjJl1NS34vPfIHR/GDeJ6xxq47pcxwUmoqh4u2q9KtihV0h/eO
c8stnujA12aouJcqGrVqgZnwVx3Jny1kIKluPkg5q89+ycV2uUpSRRFwuayIHRnf
Y/EnLWq8HOLKVlh+jkLABEWCVmVA4mfOhvfhWmy+iAKJon9TVAn6nfxYsD590Sqa
Vomfb/Eft+a2QybbvT1GfU7kI+TJKmIOifEfb64uHPhMo6Ae3B5vTSdTYQZNROlK
zlWCSInfJK3hTc3MtYffrH/bB5p6ggPn/ZOB6rprQPs=
`protect end_protected