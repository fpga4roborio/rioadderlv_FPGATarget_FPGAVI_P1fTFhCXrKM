`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
ddtXksX2+yylW5zu6QL2Lhnb2d1sD00763mmSITNX595NcHTEkwn0zB1Dry37fOW
FufOhVzEJp80NC5qZ/+F0Vk7Ik02dIR0elf3clrjeJRK85K4e3Hoo4xn7YbFUIms
l/8VZSb14+JVGURjfswrIyCUotIzlzVYZ6gzoZwDXIi5gQIBf/gI+KxNXPaKV+PQ
Ufys/12rjO6aI/pPlqSm0hCvftmBcnezN2hk1UeXgOIuKZnogjOsf0iJVX2aOOWE
6pD/psybjbnsNB6kH5uFTA5frkzIzkzl5d9+YDm9OyC+k84E83I/7/j+rk4L2dah
QJOvksSIzN867/4Qt8qYTQ==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="MvBXkzurAa5VTw+1JJ70nePUfoQXBvZOku/SMmg4TwQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
oRtzZL4VJ4iwysPsC8SXYCzXS8Fw2gtZTOskLcDV+1B9Nzn1zTyNtlo6lNICRmmK
ZRVu2BmCc2G+fmzynYlNTnSa7C0Cuel6FYpxCBlOuk3OF2tzAmLAuDyOH3Z1Yjzk
a0aHuoCdIRKv7BrZCdALt03JeUmXKPdOmIlkVGFl8yw=
`protect rights_digest_method = "sha256"
`protect end_toolblock="Jn9CQpRhJt4rnzZPRk+dOpzAubz7omckX1MrFd4p81o="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 35248 )
`protect data_block
gD6l00tciPUa6pDNTk/+t0OO0nC/UTtBwLB41d4inuAUA3i/ALrNyoJVcBnAmEQW
ptbcNp5fxEUJjnOxnedyZEuEBxWRieZFQnkRdF269oMCx0sx4MevpZ18u5nPztXE
E0Sz2bS8m3CppTnYrfl8T90UQ/yvfGGZ3AfoEHsFODOWECH4IID26DjTF3ySqVGS
tQfA0BWxokGWLjX/qt5IscHBkTLoRVKAkErXxWgCxVlI41HNsAO9CantFlQBoyOA
B5ifWgFJpWQITyKr9TeUazSQ6ejc593lDCKzuhd8NfAZUkLWjkC0XJzW+eXato+U
cs25w7rlNGuup1U6Ghs+83XJB6TxTGe5vUcGdwZMYzNFouejYeY0CklFIK2wORAQ
4GjoxlPjLa5upWBbOLu7QUM9slyeec6nqOVNJzeADepWMB9oRUa3VBAcKnxIYra0
JZmR2rAFOXv6SivHKUW+cAJ0F4aKWf2j8ofShLRj36aoPbEKdVwlxy2GWmVat5vX
IibTNiZpHyeQSkaSDSzHlzYh4ySKLm968q4YwcqIYhPL/xf3jUCdsaYxuOmpWpr5
J6dOQ0AMvt6/zucNIgh9rG7/xJm5c60mWnyWxiiIVJLYSagOOJWeP8W404caOetQ
VtD45ht+JbrO7/i575WPzKH8kHK9HaJ2aZWq5r7NiToQZNxVdAH5aOlPi6uI5aLP
x77q1O2JzTZmW4SY68+/PO4lpgvjFiMDa5D75rBiEtIPVvq9C/0u//992KkWD8gU
B6DT32X6sApYlXfAqMqs7zMV4wzvbTCNjZMEhMgz044wx70ANYutneZafbQXZ50F
fcVuAo1ee/i2ep3Fz6SA2liSjNW4KYgydSYuP735AQfMD+/NOx1f8vnvOSxIB5tT
/TSSybidKkUBtEaOEFXzWv+DT2uUF/IzF9/3YR+mEF1IKuHf0OLW2qfraK4Cy8Gi
t5GUq6h2XAWdcpx9/gqdcf3D42B9yYiBXYAsk9D/7AlVctpTptTcnzCU90XH6TxM
BZsyNZbBrLVSbdeINl4u+qTcUNNjGtjh9qR0j3LwqGBu4pPv9hCjBK86DQs5UxwE
Ib2GwjPSk83sVEtw1fjcNkvmGJYA8hLK48RVsXWaS4ACj7wM3yiPeUjgmjV/E25Y
Pv2TF1zdwqpouqifsFz8vA5lRaa1WH7H3qs1v3dZ0MC66jZGzYQ/q/ADZCuh1NDo
GBk+AyUAEpHfMqu+vAzIAWySNn4X96SRJObJ6lrN5xUpAgYP/PQF1KEcS6gTHaKf
s/y5X4592Cd+fsQZtlfgx6WYto3oPgas/fTZw3ZTVsjto1dX7SnbUwmYc1f79H+/
hq7FKKEWQfXj0P+wf/PDTa7o6jUjWE+gvhezuxX1SVNC0C7LeZuIyaMyCC7FlzAn
8R1FwOMNtKi+GF+q+CjJTS3Ew4iF0AtKvwBxwOK6dCaSvqxNupZ1h/HSqSfdsJRV
yB1qOq9dWMfrDG0PMIAcNHmoZfcky99Hir61UibgjKXhtiSDE822IlMPggX+YFsX
ISSLtXuovWd99c6JW+/TvjcW8L4PTRUTuIPWISUlJmz97CY6UuCwdLsoGV7zXR3w
/qKEOUg9e1XBhhVD1ZjACuN8bEj/M1P9kQfPKbKMsnQ1Sben+2r3e5g7Ei7JmThJ
epOLjum4wUalbdboZJC0KpZ6UiOAwylNkjdMsQaHMXAUA/W8lGJdYSnQjZz3kqki
1JCF0LSzinO3I9pktP3uo2fV+jWZLjQRAAo3HKQeP8gHcQDOgFYnDz28+n+KajY2
jtbXS3EcMx1C6Dpf7f3/xaCN3qjuMbxFCOrnMc/TkdZBep+3FAp2j2PvgKNjF8+j
lXS2IUOHmSqI4NnJ2bxiii5NGvE79oua69wUSBbPQmjTLs8MuEqkfWCgwAKAss4m
eefF9y11OTOP4kNJ4QgNllkUvKFApshopKCYdGBYHtWwDxP4U6aqkWXz/LJS1TZl
HRrYJrLlhtfyPT9vgLxkLTjW6uXkQqEtHXIFkHw6nRwVUqJDar0T2k/uoWy7bRbu
dVM/MswhB53xOoLIANDA0Fol1byPbp1jXL77Waw/az5mr8g6hN/hJMdSA0MFWRWf
Iubfi1McEnH9a0mUpc03luPrVkpSEqOzi3gU73rR5lFUY8q5GZjgbj5xVq6hSZYq
8673mRyDv64n4tKHrApADODBWhSAGiDQUb34nplXjh+MEK5B2e91rGFLhdJueIEW
O21krM+2Eyg7MguBdY/Bvr6wu0GKz6gySPQSrj/o7ItFaFwb3McN2o6pZV1mP73F
/8lrG497+Rhhcal97g2kBil3Ay/ruGF/sQEbI8yS0v2MZtDQHV1r59Ci/rZGfQjC
YyBBqU2Qnzd33oK7nAfuSmSWNT4XTn62MCYzt5YYBS0RRtjq88asjhLbSpP2ET5I
pzFtq1QfurI/xaniz5rrM6zkStbqQLbe3OY+cMo5YekGsaQijGMp+m4pL9lMt9dy
2tnYct6J5vM94LdybDTXt6Fxq9MRiWd8/UPTNyMLfbZkll4MjZ181PcbEzXmplgo
/84KeFRMVJPq0LJ/8vUDzoeHQT3oa8B7+awOEfF9a/fnJ8+uZ1r7MKbDOqL6j1kC
vefcR4CehcC59nlEmmJgLDXlwVTDYeMbiUNbxqJ8sQ55YMCsCEPPo9qu33Q74ssD
X0k+KoaR62gLBfnasTXl83614lyQqJmhu1l8KHukh+dl7COg+UxjqHm6YvWgJdfH
0JYDiMPoW0tliQ+rKDhY4wyrKZ4hwnRsJfI33YyXVi63TiGYBW5NKPZBq45rsH9n
ooxHXmUw/hgjLH4cOswgpVZvqWuc3VMr+SUHI0elYHZtfDIZKkgEeBpZk8hM3stz
6tn5HIl6ePRJSG7SjWeWTRJMrQ2NbrlAEGi8kcD/ZWyziZ6ye7oLnkAnRsxd/src
1LcOQEMleAaFA5utICJF82ejxWF6mXRaLLvJ1d8sRuDQnZFkw7+dztbI0uXgyg2C
9grD7O6wcOmsQW+WHoPFqajtj64T4LipbEvmLsTlCIwgsxVd8uEBKl+1ccdF4x1l
HYA0Ito8Wrd6L85n1S3/5+x9wnIDylvAMy4w2je52g4ABjqel/CGsY3HrqVqsx0u
1s+gmPinbj54M8CNRTVocNf3BcM0zaZb7CQVlhWpoaNczv3uq7b+cR21wSu1OIAq
L5vHLf6rKC2wKXbLPR3szj3JhF89SqDHuarIAzr9+YA40sQ9yqOWrwy64dypLT33
/fOaxYPOWDKAcIamoFvw8Xyua55pOMU3pQwyb8cCpOp7T6CtJO4bOwMlYG4hbGNl
ifakpzVzo/ZSOHYWWOm2kDGoN7ejjPPJUlzb0Knu8PW7pQELf0/TIcFe6IXmy9FD
Qtq8XtGCnH+SK6Hx5OmpM4n00pyDb7J3j0+r2uB1ziPIZU3LLsccAeyUhfekwtR/
8aZaXPQytSzYRv8rVsUTklMPUOG9ps13G7CB1H/F7uazF1rFi7NA8/iRS+DTpR05
LCylM/8gJ28MKIc2md9oAcLm16HhYn2xn9MqMcmZEVeJQED0qB3k34zXH2O7BBW6
K8W/rhc6S6c4F7Zo261Wtsl0BjlKDMHngKBZOVcSEPCBU2SIuViefxuXB9D/Jrmx
2KwX7+ZMj0HYIMxZFw80GOspjg3uSoM418QSBXanu3h5ezZ9+Ux8rKythpFgN/cm
q8JYl7y8iDnLYBW5voT9z/MurFLQI1hygpU8U8jLqn4l6COZcQrg4dgn2i4LEfay
F+C+qczWvlRQdUqHmyUcts4qyCzFIRfQTVerQ3dcsyM53u1TV0y79ttE5vtCG8QH
trNwYs6hWN8WtFbxGh5A21kU5K6qD7UyLbGgL1Vb2Ck8auWS/WZbAajIDHNFDcIS
L6kLHJ/mhmIJL5Ut/O/cqBIU6hrD418MMqcsNBFIGVnaE4TAETD8+BXx2kxvWxMQ
wsdywNEJqewByg9/fmxUv/i1+JqQV2QzgQlBwbzQW0r0g3KWT8y0y8cdWxuz0gHA
t/VZPhBsKeuM1DrvJcYIHbLddeV6Lhw4M1a5sIKrL3XbjcT6KLgd3aTKoBUq+UZ4
rOlZoinI+kHFDEtq0eCsFLE30+mL+jIBQE/bCtuim11NOQsNw57M1L8nnSm4ermA
MhoH4f04Me5LxJhTUO6V0OPkey0linLq4V5eBPLu1bQQpfPL0thhJQk/g/ofaLAC
7U3f2x9qYulrOv5c3tbq+xEMhkfyIdHVOFF5KNjK4xhmQhzJhWquQbDEKOGlf4zr
J6Lae+aDwaOwdnos6RHBOdIwrNqbDl6DIgaU3HdsPUTNnCnwLKyJFA+8r2Xp6Lma
FMByaDrjf074Q/PudcQ4c1jQxcNE7/YpQMQ2KtBTUllOV7PH3Y0wLbvgqD/w1U6a
NasYy6QeoMkIdxpbpi5f1g2oMsHk1ynSyS/mwJRmYjDhCtc10YbYmckqRzLdmfuR
/YwaKThILUinNkkKcGQJkckJxsn5MmFJ6nhwxUHMEVed1da+knbqSnMMoI/YmBu4
4KX3MzsrmnL4Lh8dKAdOjN76LFutWvZh5J3C9ZOmAFGbglMhd6hFLde5Bj9VLp5e
5Apt1+V0rYNl1D4x2yy/+vTj5/VqjmWQbQZDQ4TaxEf+qs9RGCnm8HedbUspmkqx
u3cRt87mC+A9bGv2UgeM2IQtP3XMvzokIm7xqCf1l2EEyuD8sh6Xit4jiQ5Av4qw
WUVLWcrIGDx6zmw4v/yGtuEsEV6YWwb4aigRA4+jorNg23gpU3cAUOyezUlJh06f
BG6N3lzoQtbL+a4zVvwcyoioAOoL7bOQ7VqfX5YGkGU5ZV0lW8jamwnrkg2rBkCp
Q0RE6LujDNpvzL85bIDiM6SNUCml5l9gSST+uUwPdiw5Sm7snIldmftZ4a06rLgh
mbFtlHSLcr13xJFPI9pMNqftZGKIxR4LfASaD7RYEZjau6KVGX3xoMLIDn8SH56L
6xew7ppCMfnKorMYz4tK3wFf9UwkF9TX9F7CKHFwl60RjyBcS2RZpiE6jajq8XVd
KmhzUTkpSSAhQ/M1I9tKD/WLQXM2DJ5QWehE97VHP8kdePVc71Ub+MfbfknkDDsF
hSRDsfqiiZo5i7YZHu36XvWALTwraS9GoMFPp3/ID8abboDjhnJ8k5UuyELMxEmO
fU80c1qStjuJsimT7/ALhIpaAMzg2fdCvibptSYBRyI3lRuL8eZXzTLJC+LmFW0c
wzODI51ftG8m9dmNPb+O5ttofmefvu6tkXhxjyE2cjX0CqadGA5oyto7EtKOosT7
kRml7Ecy6hJzvD69TVg8QJAZiRA6Yni8GTQGJuIqpxiuXN6KcFiMXCu6X2WbqGOa
9e1mkPsGObw2QEdMjyFr2Tp61ghyM0GkuqBFZemJ4SPwBgvxwgCaRisnyt2nPfRC
6Zh2U5DN/4xpZ36DasbcjcprqNiLEDLV+oc2vRZOcyctMtsyUq3Ip9NfmEzah9bU
7DzH2d41VhDkOiHK0tf+gCATiijDf+RnlVi6lEx6a55VgIWpijoYUYh22UIgAgN/
G1Jt2VzUb+8ULUKh/Hd5G1OF5mo2C6K4WwxZgQ7ryTCn60nPi9BOBnjPjshx1Ix2
8lsKSd2hfmdHuAFOl4Y238YbZ7Nx3JjZISYY2ezWEmLoHMX+7dwU+HONP8f8TsRX
re86JGsCh+FV/XrrJ4dCVtFUzNy2ZX4LBEwgl7Ym1qJMEijNIXB/3NTpD1blTGBI
a4LENSS6IUk5/c29agrj8eAXjvIkyf7IK8WX0hjwBB100O36UuCxwBMr3rbb+92V
11tyMHX8pheO1z7bWnapEfcmVkvVEQ8c+LkieUJiVSoRFtdXPalZLjMgY43R+mpX
6IfW9aLRMfNXf9jBLVN4ydNEzMnI/BnCEJIV+84cMFksuP2tnMhZKDXLczIqoNxq
Fz3cG0dV24UWpyy8EKQW2iWnIYy67uu75yne2py7FvO1XDoC0JRI0cEb97HR37aL
qtNJ3IKcqLAi+ggGUUFCd5j3vwxUpmgpipGuSE4fNSybhRipLu1nobDm/vaZCgX0
/GyC4bD3bMMMfH8aCcOHcuc5H9QR5sUmIat7olrQdISjTHNUIOKxeMhOZR2x3NaL
Af02A7G1O7DDFydQVxpEL1kU5QqQLXAb9UgwNO8VnD8Bb/1MxEDm/TWiCcQl+MzH
LE5IQtFYgKQkvK8EajgMfTt6gpK79Pjq0QIITqkADWd4r1cijzTbFQRIsqw3scaW
29MBc/M4VJXYr45xlLQSUIzL43l8Fv+W4b2ui6ZN+GsCk6dWWV47MqRCvgYaRafo
e8KELV3HSy2CiQFfq3vKJTZlecy8C1Jd/YaP2MPWho7I4Plqg0+ABQ0VfTkqE3a4
kEiULaGStPYfEWqM3XfiyjWz/2DBHSwE33JjmgukVnJI1545yZy6syR98deOb+LV
tFG4e/RjKnB0qGekHcbqZNQApuNqhXyYJufNowfjVpjC0z/kATu6ZtPNxbH6L1NM
9AFvIs8K4ByfGpAkpMqUyvUYRoKn0MlT8HdG6tOYALunUDobpzud/fr5+dsp5aRc
Il4ri86zLhFn8XH++6lUT4DeLyH4ERTnf6aUxIOfoBl5cxuiKHfrPYqglh8qIXK1
HWPcjJw1FpGP9UFebdZL1ARNE1cFck37gaDJ4ZFMhTHbhNQhNaf4W7Ga+xc20Yz4
EQv/vcGxu6H71OPkF6U435pnEq725dwN0qhMouWvvkS3HPzakNCzYjXN8dbKzFHw
ffg8jZ+A7owcv1BAQpwQv5AkWabYqIZFHqsbZLn/zHYtSqtTyzcSZc7saPtf2783
+XuDOHVEUIoXKnIVOdfgZ9d0OPVQHR1Baj2x4PAv72I+G7lk0OopipZ2aScCsQkM
1e+cB5+5GlwBCk3aAon3eTwKc0RcgChGrIlRZZitIJkljziIGEt0BxsIDQlhMYv5
M0PsW8xu94PRtIeLHlKIjhopfefkSz6cYvq3Am+Ap8fDLyccYfYhA9DhQBBO7zKT
P2Grb4H+rb74vf7ri4Xw7/oZjy6NL3kJqTlrxouVzV4AUEp56yOHJnfzpsoOMKGU
rgtAqAJdGsYhk4FHehLvoTvVh57b9/r0HYnrcJQ/f2Tb3UpXiDdjWe6Bdc33EAug
5Hq+EHAVRV/T+YoyVVrTYdCkDaBfXFV8RGz3sICsY83XcO7elel1wP6SYh4chrjR
qPH0nDoAVyuhAq6MAMWV3y9LyLrL0iSwzkzabJKaZS7mhSiwt+oTM/g8aHQN8flq
u9EdKBoEIV8JgE62rRlUlaHFcQsmJce4Fqzj+c9waWV5RjfuBwvXUFfx9ykNaK5F
ZMpdvvpCvVDAjogh5tCd2HuGHC8JXU53aK5+38JWEce4i9CM7YZFkHizUsksITuL
gPtDpROv7NcW+KPeyXdHjstdEmQLahZwMZ5KsAr2iRE/aVxx5SpyLfwIOOE86Adg
vYc9zy5LRw1tXoAbPR8DNiYuD77iMdHFV3KhSWgZnN5kpNlLlD4SO/P7Y397pZM8
FwOHFB0B9uJICDZJka0sV6M0i1NqgXYGk5cUP2Nq7S3qXP8stHWieo3JOsV1EyfE
WsU8sRx/0cONjGbojevStaRSQXrWP1J0kUE7spHMp5sbOrQ9Dwmj80m8Y5+sUjiV
2KZDyOt7SBNow/HhAUxEKp6kz7nxl3jIwnnqfRcAcgNsJpGc2XB+BvtR62oNkHYz
/PFj8njbhQyQq0W/j5/IwN5Xnm0hGxTLktvZNmV3SRC4WMMuQqG80Ie3V8LoUXL0
91Q/YH3xSOgKvhFSbL3Epvjzt8kNvyxg6ncH4kHXOE7LTSxeSdLHQz4ua16rdEe+
yBYxb13qwJuSNTdG0OUAqKAe2Aq3k0d1q9ztuSlZAOP5MawvQwoLh4+SSpjdzvLz
gwD23wGFjz2Q2rxDMD7/Eka01dxZOFwbYjldREN0WYECluRgaaCdzIfky3IKjB5c
c4Tv6euALwWBPIFFTNLnv56bmuh7BBceOuTtNeSMA4M91OYldZgyxl40I0mM9Elg
P5CACmjLL5jQnvHZhDsTeCNCTUHP52jxusW1T4jXMjY9d64tE7MFrix+GegdDkYR
tO1vW/mM8xOD4TRDOulwEOsJDR4tl8Z32qAwp93IXilcYMtgSi9t4/+cKZeHWeDJ
oAlESirgVUwU97QbzaKPuQ51OUlJZqe/jmyDIH5KO49jHrrKrUVD9R3j55glw12p
zPsAc8qk/OQ/Cd1t5bbpemPuaTv6b409/1e+qDTpFsA9PEG3CzUQ4l7PDAasYSjQ
dvDgEZM4K3Qf2Y7nR2/CedScbqR0dO+zRkW5g3yo7TDNeEyuzVFCQL8ranvOUxPh
9AgcmOo2gf+HX8Simj58Uk4JplhEN+tS3acKEbjtz9CHSyIRE25+Kpvx/4YYPfoi
+kaNGiRF60cqg8g1g6twoJXXmQdC7K27yMJwqo82U5skhVv4gMZSZzVYWwD8oKOm
oFEaxno32mIGuTIpDNqUGPePAz5JdiVwXqdgdjqFNs+K9xmqcgbZMWUNMSFINsDC
/IY89bMXu+4oJfeKcQm/btzNtpae5Q9+H52tgOBibswsJPdrWawSjTLc1tNE0Cfi
IRSyZ/u2jbrjUWz8w5EBcEoaIjQ+3ayVyGup/NIrHAhQEiHf5DLFYyQ0e4FgYXo7
kuvRplzET9jshmuyf7chchWWDipqteB41ayweRTTs6C9QLgzpSDvRSOlI65wtNPC
tzVmUEptShfbpCerhE0JP4zzSV0iTHf3SDsImhGpLoWjr1Jj3PJrAL0l7VFlquxO
YzAAEQVV9d3lBv/MBDGz8CvtBdcXUE28LjXYuq58cKKiWGKuP1/WZaHQf+o00ZDO
j5w2CzwAPHEuw8zZJ1rNCtc/FLJ76/l7LF021K6nwfyMeaedsANw1ve3y8UeMbph
WnOdcIOVYbcksQfUfxXq24uOJ0sZDPPtieTaXXR7U8rnlKGkb6DIzqAZFsNzENkD
vlRKn4xWHmzjIOLip4oRNQu94J3bGjefk+MEaQVJbcqkpHud1NdIS4+CAI6a4dFV
UUale2vp1o6JAtk9DCIrs/i8eNxeGbHISKAHPD4ibgjfkWMaCeYKh4B6gKVWksS9
75ZH0FXIegCglFzwF3Oe1gMdY/3nqH4Xh/sOZYx9WA42norHeBd2c02m/MR8VQiS
lLkW9NrxoaxaSbQ20/+B+UuZFD3tahQmxPtc5tnjqyGkSGxrYZmEZOk+TIB6qtID
LK2rW95WjBgAzpN7Ap5ZJNAE3A0kCp/AxdLD3hRfX2c4DGgSJOVEonjyE61W6ObQ
fuOGJThFtVFFiXLLjvlxQ+wHRgxPf6AI6swBaSue3DUaINfhn1H9lFz/lvQexBLD
oGx7XSWILraCpn4nmUdC/Pck+tTsthtHfvn1ajQGLshrhbRX3nlpKnnaNl116Kd8
sqfGQa3l/mc1H3S1DZGUPc/Dc16LpUMdNK9nJu6SToZAoXq3ogUEioJhXT1vChJB
ku+Ls7okhaKJwaL0NB/6ab1LVDPgSpL8r76dau2lye2WIxOVGNYE1m+C/1zLKyN8
kmYxi1cwskdLOO36WlMr819gRLoWD/IAGKgxceO9NpZs0KuP/DdedxUorMFVUg8p
rwaMkDfNgVItVV8eV8cA0u30sHyqn/SVc7YwjBE/noPaTR17jF6ttzzltvopuw+i
o5zShGCTUZXQ5wK2ntaWdzbrs671mgfkyaOQrxQOZmkd3aB/EMNaHE7kReKtarG/
Fe1rjrqA6vxLeMhZDxGB838JOUNVzu7X1ImyK/1mEW2M4GyStt1ezjmyO/OswmFw
AoIEgk1iWOAbkAP1TnMKdYHRFp5sy4N+1dtm3tSMQcoraHZwEHZpFFixFrzEKr1D
0lWwVXy7PQOJ247rAQYzjKaSq7zWmcNSRRtsUB2sVP5pFVtBw0Fi+h0vRke1drgI
HDapUSpMLUxUtMLeJHSlFF95ciIY2XYD1QsuWyjwmXXdd5gQKyHxixA+oo9wGqr6
j5LmGTmWZZAP6qMsa13QBQRz+i6cJxhtPdYaZcSGPB52VGd4SdhmFtRlb9oQLIsK
gC2Xr8cAMScqNsZWXAM7X94YoO6XR+Z4wIQngwsR9tnOSUb0TAm7fsQrHzBtsHGk
RNa45xnUljGbRNxClgvUsok184eOFLIhs7igRpciF1XvO8wXzCQla501xeNcCza6
+7MqpLxgv69dGuDRFsbtJZpl06twsa6rZG8qMxms5fUy+aEc616pKyc8WceAMOEQ
iEZvBEtMNnamo2gnzTnYDL+N0sc/d9cLhvgA2TaI0t3VoMaVYDJYCldd8C3BnJzC
2aMkV7gmB+ft2Yy+av1vuO5dj/wm8whoY/ecSbtvcA8dSAEITlfCM8VLhu2q1KGY
xnTOnKo1L2kOCflj8fd9enng94JdpVoE2OfWPIvjjn1QmTfLLLbWomeaOzwCizJb
3sPGh8XMzt8lbtS5ST8Q2G6WSGkTUxgkzqXE6aM6WWRPICaB+rIs+z/GyOd458Do
8nudHbD2RjMZaV6kdYqaJmr6C1F37vBCMciBl3TTZA2JVOKqg11H/rr2jZwB34N9
wUaFLAs9GCUTYYGLbTSvDeHQ1xT0GhXnQbmYbkozAAS9/rJivE3K6SKXgkqy2wG+
DKcOET4ZGpACZR5MQHZ5oxUiHHZF03EAJUhGe+54g1s7NoH2UTTJQNOvjq/OP+8Z
tmNVuUWJ+m8ueaEKWzyoOmikisgrBzyR3QiEhyOFsDKE0dFA59N4Lp5NeiSdiLei
5WEuob5n9Bs+dPAJEKzX6GuoTEuFVbmABHBDL59+5+rQ8nXVgR5nhbnoRrCs4Het
FeAVkL5aq4X+SUfPwN9QXbYRBadQzHiTwIdQr0yjnTUuBkxQuPLFvicoFB9Trb9h
evBG4JJHaBZvarw9FN2nLqmzVjYDiseEQbohmaIqmHwmn/Pt1JKRXw/CsCLzm+kY
MF4E8UtzHDcbHG4r7+kM9g3VX6HnOndk/NSBHBezNxVVssna6qNs1/6MdD+OZm4T
0bhS4TBdrw1UPCMvzjZSH4+FhL9iU3kwftHeU9yOeRO0uBNHIdXQ6WS+rk+c9Wn+
+jyKSR82PbzkOixmaM94vxLXdquBzodsF7O4kKv3eTCVBBa9JFFD5vUt1G2+5+f6
ak3a043g3QJLiQRtlTz3FsP9AL1X9RK5c6tna+TVbXKpIYIGjlOtLouJ3MBIUksv
kazHflW2OI56p7/FMOX8qsiql/DinTP6kRAgHoU0qKs6Rivdxt0Rla3vt9pkjhqE
CG2MKTe3YUzS6o8w08is3iXCGaTWpfdGzQ/MEZ6ywaqcXojK+Kt5l1o0DPTykbFx
RlLXie4litjXuj/tC/Y7hJ1F3Z6lsKKGOPeXKBb3lXM9Eg53Dvupuw3r5fUGpTY4
am7A6LO2sPGwoaPeu9fIw3P6X2w0ViEXMwkNZw+faQ9Dic3m6PM192jPa7trTJFG
IsHWGWGyw8USa36Wjffm2uM7WLkRJ+rkDcNBTQVuxgaQzYEMFrDFRF9RjSAehJSu
Cx94a1dxsKv38i+HdK5YNSg2in+oerSV3l176OHa+hyK/rqA8HnsD7MGStKBoBjn
eDBoq9ed6OR8PtPDhZungUglNtgWPSItUYG0nfq+DY0TbGUYPpWVlHYB1GZVdTXr
+bRtb+6ANb0D7uxOrLfEmHUFF9ca6hnTVlJjmWDLc43Kucco21pY4AWc8bQD3fsz
6o4iynMEBkuerZPOeaESKT4/M/PIK1GzOKZNVUJChis2b5KZSP0C5X/rrjxQkOVC
BzYl3A1zlLvWH3wyaaUsJsgVZ0qE6s0Bm1xYCjQYa/eRZRs0jcSxByHYp3SXNkI9
0Vmq8GijRwUM075ntfynp3UEkoKsEArx/h5LmMqniyhNI0WExb6fKE3MlOEqXcwi
G239Zr3SG5AG9pq3d+4TcwWmRhR5Sw9/nFJyxHPTzTiBQpXa3tEqJzKJT435t5RM
zBirteufZ88+273MqXM8StHbCEhV4OYsYOIa8RU9XCzs6iFXoS8QwsGZwQHM6rps
8EOcdAaYeP0qKz1dTYlMJuS91u4MnVWvID9W6cGPmxBeXNttlU3qK03fOZED23is
KbzF/b0kG0WKqDz4PxqIozg+aT4LCJRn5ukqk5364ooJ+Dyj0OVuWH0qsBioqyha
VHoPdqqo6JljFU9KZq+Eux2IkuY22SovNPru69tnU7s+yIwupa2Ws/JXZRywwMVQ
9vovv642gt24ULEZPmVhOtjKxelgDbO0UFr0Eu6jFXjVA4uiOX+/WKxsZ8YhQtUG
pBkKS5IQr0sbzkyFhuYRngR/1APJjJt8cn5xslpna/fDPwbpgI0pAO1jngvbrrg1
26QWUITPzdI6iKlcD104G1uXc9VL0oYuzII64H1TH1JLycy16lgi9zCqH3e7z1Nz
jd+PlfYAI6nw6p87Xx9XUv+8gPsTLG1QsMdyV8ykZhbd94IlpZiagAFFecZd5GP7
aZoHRRw6gPb1pHfzOy81Z9PmoyF+9vMM4fJdenrdZUy6HVQDrrTszxGSsO6BGLC1
tNbh65dLuCxdVcKvQcNQAzYF/rdcoys3H3P5SFzbg5fFIfBlwx0CEUKescsy6cU1
sQtT6Cd2al5ZR/kdwl2mAYN683ZuUaY4ULe/51h7CYAlkSOF8+BGpPZuWsGQ67iw
iWfMpdZgUsn0FFwNnHzwFPdhVbFIg6ifCDPSiiThHzg5xsEXL9a7NoskZeJKR6We
55N6ycCuUByRDoqBGTt6lCOCy1YNJkBNq/7so6mnrKoukIyc2nAGNcF+C9JiPCwR
3E01rQQX4Fvw409YJpMd5xgkMdjkMeIN3ZYNtKaRBpv0X+HVWjpv2o+OjJNg82iT
9GNYmUr074QH+i5sYz16Z/hacGQOSQF+/Ayx3kSl1HFKMGbzObc2m2RLONZHvGWW
Gw6spM1hUwxSBsGytzkZLOwDw6kgdrg0VsAmeVTdpLLPnPE/p1twrSGjQvBXfaWG
iKZBM/A93YDNYXkEC4S7rp8Tuy6JtQpCLTmIMSB7fMTHygQpl+2m3d9/izocweRC
SzcalzXiZxQtX8lCfXaZB/jnH7StDDdMNbnjW2m884xLL7KBZ8dunk00/5w4PpyJ
Sf6HoC+bz8fXPDlN7wgHkhN/5xfdRYuBKK5ozuA9e6jT3wrrKF3A1qZX7eUWx/og
YG+8b7Uvk8Us7meB2hr9waG5k/zn8e6EqfX2Q/y5QorYr3Yt728ObyIGo+IH/bXV
COgD/esQ1RweR3LVO6C6lT8G7apoKsbvytituGGGTxCeHcupNf9NTTCKuIoNZTDv
32N5a40gD+4DVd2POfDaiRdpSHlLLyM8aW9vY0uB3C90ACx19eYBOQQ9gtipHAoG
mhAERfLrR5hvQeimTmgoQ+6U8KFpFilooas/ya9XrdUtbYK60OXJ/z9QFBf9Dana
Xv4/9mLPxkmrEvfXpNUX6DD7Wf4R+RJW9khkopV6op2E4Xx5vxHSnJ6ySflhJiSG
tlYpExhnmLtaPYEEQACM1HJ5tJFlZzrhICsM3PG4B7zM15NWW8TbK0B6zPwfWcm2
abXu9j/2niFsO8Or0tITPdAZ0MXGw5TLopd6KH6h6yNUtMuzK2zEa8HBPB0ksUIo
OmsahqDPeV+4KfYZ+QOIcYT+MPLrGBDqY0ZI4FV6/yxokdsjxGIAE/LsFqHhCxsl
r0pLU9VS0Pz/fImPuU8MEB0ahvIoAOe4iLQCdKIhtNzfq6MwWi2qjxQE7HlWwo9y
M0AAsvqZYanneunmV9Kpux731rzzURkZEJ2VOylHyjN2ETtPUCMBsXsTmmgnAG56
kgxYIPW9BHZXCgdbFaadittZOa0GS1/KEccRb1/lRFXn/xcRL8vY9JvzI6SyxmXN
yC3uMZ3fk2ZxWvBro5/Pa89gbILHOEsCcMafPTOrtleCf9gqu6mJE50Dg78kl2Qm
juJ+KU++yc1cLjCNfrBJmYZWviZ0mfyH301rBMAxJzNCT3F/wzskPjOQ/xTCjQf+
41zq8uYEPuHLK8sSmLvLssFUX8MPAFy+uJnf1IVLOa+uB+HbJQzPyYAVjO0k1EP+
te5zzWuBuqY/1EJUQEq25X4p5fUf7v++IpWpSuUA+UEvwpC/3J0ShdlPJYFzUGz3
UHmle8WHounbGHEFe1gNLfj31w8oxJv/WtCzP3j0fTLMK4iVjY6nL8T5RHwyJagi
yVNIhTSyqdxPbgDQq0DBy/6lNN3YBmCCbuPqmlq1X+iSfE/X8N9/WUzhaCevgQvZ
LCPahVK3ooGG359E1brmnp13YBMyy4eOCgZqXtFdbXLZ2BgjPjcqHi1OG1YkRDxp
qdw5QA1sQcVAEzTkVIllG3wFw2dAs20L2dxdaFYzAr0zSY3krxCVCy6t+lELZks7
fmoZU+cFsj3lGdgv7jL45DihbJenCtGRZsexhV1dMGJrZ9fOXXMLNZDGqP7tDSNY
hSrrl6Dz0n8WM1I1ma5Qs6k7u00YipWXwkat754dVxNELmwhFHpAf49DBwiNaaC0
l4zpEgq3bjfSvG8LNyJzKxj4oA7Jn1V8xNTIKw2kaLcpGCfrUshIT33JyL70tsR5
/cFpqBacTYgRqfXEOZ/X7giw1lQChzSTWXmYj/vW5OPL+Ss8a85sNC17L/uyRYpv
Q3dbNCRkHDsY7shvMS3lV0z4l9tXLFC56E8tEOahtL8oEjal7IweO1UiK42JzITa
tFQ8F5KKJNM5aMWGtolkskFK5I6hQtfw/6hUuE8qII46IYo7KkU3mYvyI7jwiFiG
1E18raHhGDwAjElPIyGGerMiVF1nYG+NippfMyvrm85745CG1lpFjbpvT0OVUCp0
C6l8KJDcYhdShbrfAnVRDKM7a8xDwh8zQJZ4L9/9l3C6TIpwVbOogZCTqW4rm9Hb
HgXcL1lJOH6dGIHU7ABQptKqStylFYNbKdfuzp5esOiVum9ETaYmvq4jaLSw64uW
hZiXlClZcpEQ8+38FwbdSDDl3s+MKvN6q/0Zm8vWn1TGduwKMGwjoV51V2AxGVEB
GCBiLZJqnXBgOSM2zGKuzvdiixAcdfLA/zfZtx+YXozGENTKqNyD+4ot3q4iTU5M
AYljfFM7ENEhzsofoPzC/2Wliad7lr/r1nbzxOtd2uB2ev7Hbq6WPpbNbDnYedxs
d93Kbjfqd6n/iL1U0CwRqZ3opOoT0MP+szS0GPQB04fplhiD0DpJmEXrBIH3V4b3
ZPzL0apScGBGoJe49MLtmf4K3pZy64uSWvJsJA1YYDFwzXAJxXY1KgBx9QPQaNA1
nxfD/oMDbqqrVAZOJa1jf/am4PQiVrl4EMzcVc8O/GFDrBiTVJ/9qXZ/mSo+DkFV
gg3XGGWAd1Cl+kcmPBbOun1G6tnP66FL4ey4btcOuGclbO/Y+TLRwPCuNA4IEpDS
GZRx39Q1U2u1wr0owfgRF/IrnGPdYuY7UN/VhUjrhZ7eKZzZx4V01LpbFX48ww08
arNQ6WQoZIHCJpEZXp/Shf1u3mMhOELc/qXbBBTnaLqr5huSccVK+YFEcy0tv5jC
odTfFm3PeGwIbmvymu2clNy+cCzM+DDwVZsw8oGKkLkaMwO2mvYQW5yMRPEXfqZU
7D9NfCxl/lEpFyOaYNKVynLBPiLCHMlGc04N2tC1IVt8r0og1lBDewkt0cI4ihIu
OBPFiS7Mz5z9fvAoV2K8ocjX2Lu5Ww7JRfDI51jBGeuYDUEmNg+nFnAHuawf4zfy
J2xEsO0OfvDBRmLRdqx3DX11+Ny9IiqlFPXOnM3xttp9Ud+IlwPw6Sz6VPzOkzye
OLh1fyUJngNoinRyjl2/2RCpqqTqC5/MI9SSwt9yXKtnH32k4tED1gCkM5pbaiFM
8Uzf1OBUp9zsMDvYBCtxmx+AraFdi15ytSKNb3enuiipTF90nc48IPCLb0Pw0Kud
HybtRIkiqUauQzS+C+R6S5MAdt1n9xrvKNU1U/IDuwyu4os4OWaRoG9Rnj7PdEIk
hK4B0MxTkgV4G2+GfYybDI1imO2vH7JSknk62NPHdUYYtvaueUFICJ7G0Kv+PEZQ
J7doArSpWT25Vyq+Je9Y9RHoQnVXUn2vW9TScgeZ/HtMxOJj7S/jNu1VzuNv0RXk
CJWYybA2RAJJxBl6e3YEqFcdt4xqpe12R9dh/H4GSLHBZnHFcz/xUWRBCB+ZO17t
n3HSYW1z18UMfStFXK94As1mXe4pyDnceYCJtE3+xqQZyj2Skc4T2eJjSDjq/s0Y
zoU8SsdK/MEqcHOf+bAmnmcL3Ij5mKmoUMWLiQWxjuxn4G81LS1IjdW/X2My+vh1
NqMd+8hZNNCoWxI+dmCrGnMzkiyOszmlm9tWhnO6n2XKe038Yx1KebXgjGff07KK
dNJphb60wseuuTS/jPzvHFKeQxT6RC7vwsS+TyIO7sn22JfGMwAi8T4vgDto+mKV
oydDnzC0KZxlLCauX4ymP8vl9sBhsJyd3qwX9sFs7tEOngUaO1n6uTjfha7SJQP0
AE9pyFCkrvVoeUDP/di44VZfOU9QuMQ80/sk7mqvefIS4QDkqzbj5z9bdhe3LvhL
EvELIz+IVaD6UP96DqGF/vByN7N1kCr4DvEckYO05W3L8w696mG2BuBoEUsGOSB4
22yd16Zc+WLEY6V1+TIvtzG+qRvaUAh4NjOyb1WF/FOT9WMm+iNSop1AkBHIlEMK
EmfmPc3ddGh9a6hoUp0/deKnSafTkq2CuEBJ91QW/BXoxQ+93rBhQk+yHJGof0H8
xuFSFmgUJvTNF4+dB7jr2nXObskCv6CRXySd58ZrPH2pA8jTAJo8SeF47rAYpgAM
41zns2vA8KrQcIES5S6H+3sKYVCpORBY1nbx5Lsj+NM2jos/Sp0IHyTzf8SVyqlK
F/NH2+v2JiWwCjGVIkiQcER7Ky2Yjs9Uzcu6x4+LP4djIMTTppoll/hYCLTW01gx
6HyIDWbbZBGjIi7E8AraBgfbKQ9gn3v6Ob8jUGEYoCcI3cXF8ODu7Byn+oiClMny
7Hc3iv6FVlAj13kfg6NNNKFzl6bAJHlPXWY5fN86h2UBL+nmzY6Cnx2UMYlh4hMh
X9VbJv7Khy5zhfs5Q5b0pi+5FlvEvouuKD5D26EfQWdLC0dxQ3fD8eWGTxUml1Ij
vPb3S61ry+FeulBGFUb0opWccZM4+t/dlWip8V+Y0rb8660ZS+ZtFJQLclT/4RnC
8E9l17DqeuA7K0DB4QqXubFdHolu4DkikOzXYoPp4WCfVvavY/GAi14Kj/eObZql
2JANaS+PYTyiZnR0hYX//IzH0TH/p+imTUaL1vNXZ5ZLXDRG3kbDgtQYRtt8Mcf1
C/YtTt8iIT4FYag6sC+mquIDEmCwp0wbPJJxDne55/4cTrYZYWyJDKtQCGHhtm0i
1SGmu1FilCRyP7dYvY+sWFtGI9Qo29FsJgrpXgbsEeeODJNc5zhfsz3aPZGVJnbc
ofB3zfxhC/lzzn+FIhN580/AunVaPMnNI5RvsyTfdqLTstYZUP1ad1hf6PleCQVx
MzsGBg946e0vx81q/KnobGyS/JkWSxk83nIiEmI72AcO5QWVRjALrAfDF2sVl0Fj
Mw2cckAeVUXbhx8uw11+JeRe8j7YsjQCEHDHmWBItwdfNXIM989mmZbWI3s+adBx
kXyHfQoZwQ4l57CSpqqy9xoBLOtn2gegIrF5mat0+FU1dFNyA8MJQVP4Cg4z7jkq
QEuj/Mfw6Qf0Gmf3PvKvRrybxvYyv+dkbpEPBec6nfj65vhF+PkQGKn9kTA9dk2J
xhb3GZScD5O7AHgdDvNZAgIQUYpvM3h3ftHNOwOA9aBJVG6nQB0Baa6WLAZn4LHY
gN/6sj+GZTzGMrVaY1A89KS8+z4mfu/sxH8KsMY8afRoCrZPAefRrntKs05gXASg
Mq/oJriLZLqvXS2Rik7+T5tGrxUc2pCureG76/pDQAA313xCiOiTgInEmI1fH3GP
fVgSmvB5BEgMCboJijL5h7ph/Lg3AwnRbK/jli0zpmbMAjxvis8Kh8PXVH/g+ZO6
w/1dEYHg4MJ7BKBd/KVZP2Zl+gk0AhTLmVGWS/dp7FwuSgewSzgoa/jeegek1jiH
ETpE22FNt/IXuzjm8zVesMm5dkoyc0NnxuTDUjlY7RXZ5rdckHam7xomVoqntJuX
QlCGtWnwVnlZ8BpyS0s7gntvxjaUvx/ckNEge0scCipGvQYuGIN5V27NVJ8mmxRI
+gBCEkJtaUiQETlJKqOMeUlkpP5Noj+Ns1bmqbmjJg0EF1L36v4oxJtksTNV8Ks0
oJWEFI6+9u7sE8GE6GwaMQpXBvxOfq+ti9qGORGRObw4D8+dmEo2KUfLg+jMNdma
kxSquF4blXwZ1pHXcBOMaLOHCQqMv7B2ub98xj9typsLYOmz7x0InSDilhXLda3Y
wbwLSwpi6bjzlT/Werym+ptlYn+inUJQBqb9Rq4O4g5SRW/AfKaWgy+kXFhsa+ch
SAKrjx7OwuBh+Mc9X+QrDcXmdVh+WAcp5Fy4eS2qTPTjY6BDlis0O2/KkPTfBGov
QsOUMYScjJ1rlhQrjQ1kRJClQTjaXhy2I37wabY+pQEvGH4pNSrjiCGwpVRYwhes
HFfm7z+luc4Nq3miAk//Bhy8bx5P44nsRAAIarOCAetSDR+0jFKZLQTYqU5nffnt
Ogvs3sjqNvVkxdKZ5rzXfDofa7ZBAlzTK0oVPQFj3NIcOYOX8bfPVPFC2Dxzd0DG
cyLRgXoOztBDgztyXWdAkXVpMNHrqhipotYQHHemmJjHiMNLglbrTo/aNhjNhCNh
LP+pdVJ6LA+cbiXdM1isVtFJ7Ek+4vNBPBPPdJt6nDX8+uxhZK/tCg+nfyaudQ73
yR3vOGfT30mDdDqBgPLiNUDGe5UVYsa0+T1bO0zmaXxLzH1HPJdxDSTvw4GCNAIV
Dfxv7P8j/lCk3u7FFhP+Bpzx9S4JfK2ejYMB2ZllTga9eZc3c44FRTqriW92zPTQ
bABAncZ+KsWCBNUCvb80tp4/+XDEByrR/rjHqyaxY589TSUFu3THdIMAd/q8dA/+
yqdGaqTK7qk7Qx6haFsJ9DyGTKrkcf/Q7lJT04C5BoBPdMU18PAUM/E0EnE4SwUF
cc2Ugf253wtVJE1FSwGFVsW6yqw5jhS/+nSGPe1MAFzFa2pV+ZHwIdLaFnZtlPej
sNpgMZUlF/IbdgB88tJ+Bcqx4bLtlVdwEWrtFzjWGa6Chg8aT2RiPV9PMa/W/jf8
DnE7TRh5SYoi4/LAVZItsRhQGIbeT1BPpXhYNYxN0u5or3O63g1Jq7HxYJ6xo4ZI
33TFXamqmhKEYi29h9BTJ5hTSig/JGsqYuXUGbsryBAfVGOrV7T+nW9+bxwqgcIF
XyVE0hMyyPgHCY63TLp/kKN9GRZN9UTpY46tBmkNzjWHvQVX2od25fNpe0MWYlI7
VnJ64GmwGooU90Rx0S1ym6P6JTe3nSsuzNQL6eMwBbutT+ysk0bgFJnz74loTfYT
GTTQ9hrdPJ9KEs7JLRZROGfZTAmIA0M5JintHNO52KDoCIPM1cppFZQ4EzNS7Qj7
Js6vN7hsaDgxMVAbuBL6Ya6Me8Ua6tiHHB7w+JKhcSIQ/7TeboWuRx1lTSK2y73b
qNkH6dyFuHizKpeCsZ4tLgyU6EeKl7nLDVnLG/HQo7Oj0QauK1Y7IkKlHRRbM2Bj
w7B1nfgrpForcEstsn3PGI8b/yK1HFzdRaNvxFMGoiLq4NoMv5Qhl1w08Wlr1qnN
OzSt1/B71jeaLw51jEgYyF/t/8btjO1MmJJXIlM2HXmJIFSh6at1ZkpA7YIcBxaa
ff1B9jy6EuNz3pA4fpf44MSwluC+07zvr8r/YIjxATCI0BSnUqML3ZumD/CgvQNX
rEyDJENeVAKW2ojrX/z9DWbi+rSrO5JTbqtpgzWanzqh6Vl6a74bL9FXhxbe8GfS
AxtTqxSgTfsTq1qhD516Bej+1Or7nPDim6hbQasDb2uQu54TE2IzPW8JhLHe+WC1
Ibyrde1JSvEI6LObHpJqFEjqHlRWWjXKryKNALnU5MGvOy4RAOTCm2DtVHxdfZsZ
ZFOfbuSLGh8o4qnbhIwkUSI5ZxAgU1zJnHyCeCuQnIpUqaV0mDWV4PbmkBsN3S0v
8emEUK3E0TznVxu+b35k0u5m2qyqHI+58P0Z7zyiknIoUObEEDc0vkQaWb7v5oc/
iBITroIMT0jmRUAABf/VHOL9YUe+1p2tWqZmufcJmWHvrVeCac1/tCPYn5ZekWQl
qoSgzaOMaQnUS6y8mKirwcFsdGLBC8GvHNOZHUVlDAreHBQYf/mog6M7/EPSTDve
xE43sQ9Fqq948rrlTB7HtCiMomrNkd1zhv692oymzLw+wsATDn8PYP49kO0wFAf+
9P9doTw/crx+rQS5VQrM08qzOrT8r8RxXGvennM8kDRGJA9RybuvgRaAI5ySLZIb
Vcrst75JGr+adBqfiz3ug9vsVzrATiILlmGG77K80z5EGaD8wixp/nEfNu8vbvl4
VR045QlnBzjFesfFVG0r9zWvh0KXjCzeEZiUNcCosqZv0J9n+Eox6SBL5nTdApxg
XPQk0VAXechtnNQmnqMuC4J3g+BWxYAIl/K0CHYAfopYn2jKj6F4QvBQAiqhsGcY
gcUaSfE1iZTCyVQW/7w68fzBn56T9PoGbVMfNsWZh3gUjXApPB3NdBtx69DD8Ize
sFaF3UUBfypezB+EvcATwtdzdkviJdZwDXjPbA0yGm4FRHSJ73x8JzSs5LHrWDvt
Xf+7cY26sNVXXIHn0dvFcb4Oh4oAU1tsgmwwO8ysIrcmHfo7mQ1Qqkh0lRKBgVxx
cQZP219WlioH8g2sJbuIKabP1yuQGSMJiwPbhZ3BU4rExLQaeB9kVwaioB4Yc8ls
XGkLwUs7psUtaB8WZr2Rg3B0RCd4Vo6bcVz2xnjQ0b2eSKPByF6No1Cm4pZ6MoaQ
CBzfiKDTsHEVCZE1USx9WJv/PfXdLPvGfeNHzOdnYbmhlKJWTF4WowJ8Lt2N6IuC
qG2VIxI6yGubExys4iHtq2PRtAqm87FERePUeealanqqbrNQjKaLnMHapNkaQAvL
qto0uYJzPNLbpVb8yPbDWr0LT71nzzUpnDdGr51fjs9UPbTrgkEr9mTmd6jTrp3H
IuC9z+MTwwO0pXAUVVolgc7c48xnEcSN0+NW0OQ8cjVrWUkL1W6gxGBuT6wBd4vE
ECmGYdeqN16+cB6zSyes8PuFnFbXLwS0tiuVDBtXSzKzg2Vx0lJQ7TNSSmVjxqzt
UUPFiBecUFoGAFkfGy3LVk4iF0MOTXvTNhJsV9ZPqUGrp/RCRanLNQLD7LwgnwDu
XMeDt5uJtVmdz+i4Z2827M+fcCRJBYC+rKiQBBIGW+vISQXLWxXGJ9reD8OZ88Li
LTjQ3PlMvHMOvb7jRAe+51WchcKHoBmSLxffZKtx1XP2pKamhQZBXRT8YVsS2iUm
tLCXadWylm1UUqcSuNyu9SQjOZBXFCIbM8Lzzt5DLTfliv/5Pqo0yAPvhju630rC
+uSWejuy5V02KW2H0DO5PwJfNL5w4DMEeBA9qqWvZVisTaT5bF0Hh7zIC6z4FXWE
k825zRua4HOm/mfXKGVSFqXLTJ1WT6/AS3TSk0B5pvZrhgbLDuobK2UnyKn9Cz/g
jkcphIypFtEK/J3VwmKbUPfiSIEvNBWQd2xEXq38DPeYGtOZx3WPNPuY9TvOTKXh
Oe0PH3vnFyZ5UgyEnVTIOZ9mMc4K/uiOUS/gp4XMeQe6cMTcz+XR/PBfaOYAz/Gf
ZBOnCAhyv4GaGV/JMnye6Ddps8IWSbWYL5Zga9TOAd4lL+EJqDkgBVDJlmQWID4l
qZ/61Ct1IN3YZvLET+50wSAU5YERrdisCWeiDuq3CjtQUfNoFj7Eq+OLlfS91pri
E5idRgIPxNQouEN+kdJ6OGJSRtyGV9FqHuwJnHSNadaa6KTS63fYx0OVPf8qR4D8
LXgPQTRTTfVKfswyFKXKev+CT6ecxPQjjbGuVktatqCUK+w0lZUuhZTkqnW7zuvB
OcyMBKYw3HnyJHN4+cwlzE03hsPHuxhvSX5/rRHi9wuHtmX+Vis93Kmatx6Uli/J
mBxneKwmjxy1vY1h09GHbaPGSKRtIt2g0y4WfHHvCvXR/BurHR2YqjGRmuJL2RxP
bkmK5Sx1ISL5/fYMR946MIpFtBvkZ1Gqcn2QE3hdyczj7FZmX+nlj9AbPxnYW1Cb
ac/UampuBVb0f6U/jv8lS7gvM3JHS0SfEsRPYzRuMpVibPqjeQyOTyBDLa9SWENN
QWeOz2PHFKj9yow2LEeoxP3QF0XLor5AUhuoTFzLp/fdITy11YA8DRKLuEIoN6e/
BKQ5XYeyUE+z5tZ/mikTVFNQkFklD/Tgqui5TTu3Zxif6sUehhI5E8iYObNwkas5
qPvFSfYB6b3OrCYU1ZyVus2baAV4vi7ns9jFo7Sx4sXxc6WxY1U4TPUbdSHJKR01
THzWMsDYYzEKPSXK2chv3H4oM78kbHmM57KVZnUdtTWPiXQ54Y5FFVhrzW4ECb3k
QyCp+NAzMMoIMIoPo+JQ2WhtMU0YYJW1QYd/YX+5A6SNnA0ZjnrbYyinZ9juFW7U
rMCspo/+Cnw15UpM2oj6TzD0S1W7JgbDOqzSLyDizEde6WEC996PDhbqyjXnzOHW
jW0UgdnS7On6G9vmQvCyyXpORvaIJuNglbx0jx3p7+Pmrd7oIon9E5rRm4W8rOq7
BJ/HmadcKs27OGnwRb+bDDUR6624nCzsfJ1dGgw3NOCiSU8cw6f10HUS4RG63sET
z9koKMX+oxlbmIgGW+Utnw+hjqzSmNJS0I7Z5OuiJI4whUO5ydYfWWXO9+ENCuq1
N694Kp2K5P8kcJnePYMuNkoyRcIXIGbNJ/hV8a1gEmeKCWqxAyBu5Tz4a0J0ADxf
MzS/wG33PVZNEJEgAbPom7uvBNaCN5E0UwdWR1eH2n3FfcDDZq+LpMR2PXYvKoN5
coA84Sbknmh5nKRz4QnDDwg0y04Uc0Qo2Q9AEXVMh3a+AfBhRklY4vKXle32n+Zq
TBRGpcdg17yibz519qYOLa1Katyv0Tf5znNNFpNAY0+EVgmaiEq7b2S0s8b+A1Nm
V9O65ycCq5LUK5ojycnjVfB/d/Yg4EcCRDChEVckaE5CR46aPYOjET0XjHn8K6Cf
sFOP8I8uoiecOCtZh8CJcDP75mRE9Kgtz4cdO0JZO+WneU3F/oK4ToNa5e0ZuOSa
H2ZEmihg2rFA8lbgskTHXkJTKpoQgIhX51PpBY3nBuMrpiPv//pQNYP4dZJzuuzS
8yqYZBlB01hXKqP0QM8PB/Ud5R7l1RZ3T1pJPZx5LGOKtYnbKa2zRhhj+Sik4CvZ
dI2hLFjsi5yywq7bMERBWtukfyuAR+4ex5iWOaTrjJM2aWRUP3aAKMb5oxYbG/4y
ymQchL6Te4or56gvSrCTZB8oVWquwu1Lwd3t68eXeHI6W8zzesEW9aXSx1g0g/8N
N4veGIELBDYUBDVz+JP1Ckjs3Pi86Zz/dM7zjq6NWdVRm3Gj0lc22FQp7YaSeljk
HapsK1xUIPIVJMU9+4gjwkq386vOO6nhotUA60EUt7FRCy2RGF0wbW3DZFhBeidI
FZKll6b6uYBr2U7n+NqEgSY2XqMSg+DkZAWVKY6za+T348mF3YVCK7/BQltGfPub
/vX49Kuagm2cmSZToW0FqYlH9pXC9GdIv5IAy4UarfCGprD0Wa8RXZmY+nYwFWwI
6C7OP9lSq2+UQ4gECf2XDHs7mJ2q1Tk+kioRF9q+eYZ3H5pBPTZjNs0KxtBQQfDW
KFJL4fvpkuQfTe3r0WLtaG5cxAhfjL0IqSOdI4lgpu1yGAfVu1FxXdxcZbR/tsBM
wcSKv49dUuziDOaWdyn6i5ZuE0CG5PmP1a/DjMNFnh0l5H67ZMu9XDEbHH0PzQmA
osTf72Gk/kNy5YZtB6koXDa/ohxDEqHT8H0rkZ9IPVm+stcLxjjNHl3bzmZyKk7Z
zVrNkR1lvC+jnwCfOVd5Er76gn9S+yQCkOMhDg7NEkMuAG2NidTu2GC2WE6yArhb
HgAKIchgHSp+I45lnkGB5aBR2zQfq6ilWQkn5MZcKA9v2gD1mUXQ2Xn2Z4VVTeyz
9cY+CT6Ie29HpKxztX86WXYB/BGZgl0J1R5U5p2dF9DovqAoxqhLFiwQtXafJwPV
VJSAyZIGmx1Jb4KKnpep+VttgKPt5+QvrOBW/9Um8NE5pIJHUhn6se2wL/V1uKYN
iE3f5N+EwKgxcpGmNw0emAQxBrKm/5U9sNeS2BFLnl6M4XaZMw755hqG6GSKK4na
lY0ADpm24tg8N8ZcoqtZEw9t87Vl/UU/P86urWoGu2qsP85bSqrvlW9SRzoqlg3O
i5eOJPfrZ4N1+Qh6TEpKXbhnj9tOij+GOY60huHcwXOYQ/AeG3W11Te28h7L8Ued
m9Uw7IDZfDq+xKwvu4B9CkQ2U4sDMSPCcehDG/LCLcpF1WR7tpfA3lUt0oLJTu37
X4aZy6cG3jAUOSorWNrrYIYFQ0J9W7+iKFGyrHWCjWkKRXBX1D/4ICH8tKLIAGmB
K3BYlWxkuc1UoWlzfvZi7MO16s/TuKpS4KCSVYtgKq6g/OM6ideMw2hMPVxsb2cD
Xnkl5wODM9QI502EJq1VyokgflzQiE0gipn4jcadWXpDQGv/xL+doGLOVPjNAk0O
oJBYx6UpN08VuldZ0Hcmg9cNInvKmmMzfS124h8kmiPBg1gj3hCMByCvr0+AkpvG
bd7SyI6NLUVK9vkAWRFeYep5Ui8Xn2fqkKvkJtOPhVzk34DyDypM0GkNxPXyZ01N
986SM+949m4e+rz3qSYeMW0XtoPvz3FEnWZlDNAivAp0t7r+ExTp6lzJCzWtidzy
+9nqMx6AlxKYujD9W2nQMNXJuYbfBusZUnKJl76kp7JOqdCUuGGOGF0UKGoopF3W
K2jD90uzzkgvpL9dvST8LxoUwPQNLtBhfIBP6HufBfbZLy8vjNsCRYp64TaHlZl3
BVX1N0cNx3ldBVoZLTQL/pTk62eU6oCAUQYdHJJ9lNBxt9sGYq7acXmZCsCprlYF
0/1ee7yUwxEgNMcUZVx670g9JV/9ZPRdhJ9SragO2zAQ3J5Dk5lObuEwWsKqfIGM
oux7ECuiVbhqxzLkgmNbFkYiEPi/natoyBzFgMb0hc5BFeUc/umiiPY108xQzClK
AGenePcdELfiKZcfEdun9dOQqdfrLn1iW2yMPPAEV2z2ebUHwUmu5tAQblDSICvw
s45Lh0q81sb5/YwKYnStFRsNOBp/MGVd9A6tec/flVcYpztwAevu3V09eH/WLeMo
w6fkBc52HsPogeKujek7Ui2H1yGl6DSuaBoGZCWwxuJOpOvKoXlVfLSii1GACCRH
ca09Le0qzYFMUtBQ+WhKcjDOMNk6fw7U0ZIAtkdZC2ebdHbDU5Ny484IKCto4aAc
jkwy+Ujc0aBaNJsuNiZgOwDu3IhWAZKKr8W51JBlR5XXpbEjIvR5mq2I2SUdwGoR
gzBgegu5L3keI+t5oGHDqVYdk10noLPGyCmXY92VZBgEa+XPnTxt3wlnvezZAGg4
tOOrB3xj4ysl5OsxZm/1RmsOgDqHnjDlfWNqf07I5V5a2B5AY99KzB1mMRyINl/a
olfZd7msB+f2zpUCE6JSOeXZ/NXioLOdVOM5VqezYiR09wMMndCQKliSuvey1JZX
PMKMNZCUHqz9GziQwX38eqYthPl3WEauvTsSYGLP7E+FKXFy5zAzOWV5G/Kb30Aq
gYhOE7hygbGboLhfzkmM5c4ks2uW76MRYGd5oF+8kUr65PUugtlWqpioTK67gsqT
JlZioQ/AQATPYfQeui6v8lnrn7vRkmqeSfSIFVFyCcZk3cW8jiuGwlQSXCY2LW+d
7DfS5dGtEY9U8DrXuOVeY++gDKB5oQAKV/i5DcBVyJw1bDnW3CjFHCArmpOOVIDA
L4eMqr7+3Cfi/rEoJ8mcYvI3ET+prgaNOuzZLcV0neNYkAT1Wl3LtzKlFJKZ5voA
ovEapiCLX8p3opV5LYrXTXByj5kGnoUULj42ywLSwzL8Dlk9qiWCJZ4CPyLl4/+W
0eBYz0odysYA8EPfHT/Ny4GlyBk9oVjOHw3s2S2FZMXzlzvxkt2DMCKSkLPoGJgy
7MD21V7cmqTBRW29JvJ0uuwVZKW6+oK/iD3TkpCMmrGuKoNIOVfSnyAytLlvPJMX
K/tJsCZCPj3EWQbvjN1hiDuAwKLT369Y4doT1KZq02oF8tGEEcQ3jtW5YRshTMqL
Hv1a+GkNQXPyJygvncyDcnaqGcMZoUOKQuit7n/jiAvW2eNE42aGXMV/uMJOB4Py
JFUfi1uotX4J6ZE8N/UUtebU3xZYpZdmKRnWqH69sJtrR7W8izpxUpSq9JbvnY9y
MdFe9C4d+2hesDAFDpvG3RHr3wdc3ZDC0LOCyVsZJ3XwGEZZ5fWl7K05EcNtLj6U
PVWecktubhc3havxAhkqrw9j2uVUH+EdmX5RsPl6LlvXqN0PW7YHhIZsD/bGw50K
W633RQyKLznt8yWY6zckkUy++N0KKhTFDhwTpTvytyszYqnitrz+V1NcUt4AxYvZ
3OpZoS0NbrDH6LB05pzUY+ag1vsJjkH5jXV6OT6rQY8XdxIcGKokY+77FFG+1U4s
kHElHFOZTJEb5ZEovQKh6E01ZRyGjfKNtOXLD4Cm1V4Npxi9tFzRQCUxOwfqpOT4
MWjs9lvLjF/A+cD3+LnuL8tqPqVIpeHoiaurAuXl5eTVBPQS6BI2vWw1qDrO1d7W
tbqAg3G541BkcMwDcH9ZyOafJp7HP0SJlkkjnJVGH5dJUiwB+4a5tTKwTXISA3bi
xOdmnNYZ5qMG+vaam6oYSmjn9H8cyNs0BDODp5B797HLoNbbRAyJB1V8ijfSerj3
U7ING24qerQFF6q020qnBkt33N4DKXOdpRbiTwZ25jdfIM3rOiBkMRk84F4G1eKg
lkvyNJe79WtpYpWIYyFTKdF+mhoIWeOf+GrQkczL1b7ESFbYaDUnYZgQjfeTPXUO
m1qAbklfU7ag86H1Fxd3+mkr/O1PquozT+u1ooaKmbuMLJoK0Cf4kU5n6ZQba1I1
pZtUiZmdDLqM8TJ3uFnAbAY1R5OkGeW63qSNmxvXwYI2k7rDhgcxEwVKp8in2RuV
pnC9AQcaA4925oqCqdF/JWV/LHaYoGwkHE9NkN2lBji7tP7874641qsuLKSYHJ3N
dSJQdyMh3Bq7ihwS8AavOkcnb4MzJc6e6dscDOXAxqV0tbnYbnlRCMmAKIagxVuT
3516ch7qMLoWqRE0/xyUb85ymdDlwB9CrqoZujvUov4JD3ObyfbGFNdE2XzxBdUP
J2rpcdd0iRuKTDSinuJy2XOq/IOxOnVsz3SkOIua/P2u0lK3MStnw/izjADZp0Lg
XBXWVfbCNeiiQvFTci12luvCcyU+WAZQTJVyD/hYp/G+7vSJ9s+0IKL3cWGBPWHe
iN3Eao5T7naiWjQ+03BOuGUNX+19+Jr6B7aLbfBDNfxiwdQ7H/nvIBr+wk33H/+4
X+bNPRb+D5fGCwOqW0voKKkrpGFfp3RCgiRZfIq1WmbbLF8NntmtvTq0pUss7yzE
GUbNqQmgPLjuUWlJgg0chDWNpq4UOCNg26fkBLqSBdW100DpCSfge7kOsIFYY7CD
keR8TwfrrC4pHOrnQTf9Wj92hpNu5xldHBdI5yk0epCO9H+0ZEzQ4Qsu7WlsLZrY
Cri+uXa6njYjC/aOv7wHgazU4BWXL3E00wIXk9BaZvv2PVyHw1zX3VCl3RbCuXRU
+TcH2tW5yoF+5ahf4vCoEuYd/4AfW7CylrsKs9fp2JxnHuO79RdAKMhO7ea474jp
oA4lCX4s0OyEvdnQGsDt1ZcG8jJviN7QcaLXYGlQRLeRYVTjvgkAr8/IUTEHEVhh
z51eWHsptlEh35xeGGe19r+Pva9Jh5MH5FM27PUrrZgvERWUFDULunbJk6EuxJZP
J9+VzPzIO4oE0XblBzNQMgJChVzUEbCQCr9SYinggBJGdNwCQYXNcYs7FHsSL7IT
vF1wLJKzhgFjzci+u6lkFKXRclZZQMMAHd4C6Ewz0kbLG31tl9NJFPpPo5dgBMLR
lEhH6V26ArR3tol7a/Xjp3QZEUq4fqCnS6jlmKgGwNOeeqcD1myHQBOPPB9N4GLQ
y4Y64+I5E07QqiNs8Kf+VCJUqmwiGM1WO6xAKbiqMPTokLtAm7Q+Oqz47R4YpvOM
R7utLG9JvHtkxrcW+oHVcjY5XzpQTEr4m/v7uSU4M3PrWipqvLlLT4/XyQH2cHm/
Fa7kxfQ7bBlqwOIFMFFFEkBqsooykMyU0QpnjeNQ/mwQujB7Yd0tRbpxzjMEfLcM
tdfoAb523ZCL6guk1Hv1Xmq4otezrFd9BsgbvugYdwtPv+5pf4Ai3ZKwNswkyrzr
G6LIyGwFmdJCjhnI9aiSHGiPnViKe1BL113ri0qGBr+CUxV/hrLUbYFI/L8G50yg
rfLE8eolkpFFgBXTyUgwkpTSnvplFKEZ7gBqk2T0sn9AD2/og9+H1/tX2YiEWlh+
JAdie2E7tPU2yPHfwrBOzf6Oecb4vamF4Ct3CIByu1G5Bdw8bLyQe7jITqW3RcLG
ZBHHyJkE468VerNWF2rOJXwJU35CFXn4hksv/jmNTj5HsoEWncn28hPboanx1mxY
wOln2xECmaWW48a/HL+f9zcPoR/AU+xIW4R7XAd3cb1Id9TsKkcPAWD4/R5a2cRP
1HcNIvRusZ2fFcm3+bUi7lyhuS1TNYx07a3GlR2YCJEh0xByPLN45urqJ8vX2bDU
2N/5cgzFxxPjyNSJI+q0id+Qv+VZhoHuDHAyzud6QfR1w0P3jllG7e25UDx/FXyg
sS4A7Utb/v1meHWjTs70Ezs/v6Sa0ur3AWw7pC4SN4lqjX5ECSZB9d7FAuPz3Pw1
D3K1HA3K949WAsE3PgQiInLnH2S2jODfuex3Vs+GizP/jOS2aaRZXNjjrvplToXQ
COyaNemtl36wLdCMkHL3/Xwaqht3Br1etY09S3ErwzlB0lPGid1NEqC9IH4SxrE1
YzqR/SWAqj+4SX2aq6mzUjW0MZhH7/59qgSk1xqAKZ1oY0uYwTwl3zw2edgDSPWU
sjy30pkSjrDF/xlJyV/TeBawC265IB2H5nx6Kt6gIG0H6u8UEVJv6XoyZHsTwDYH
kZXRO17+1TlarbH4CFtcWg/oDSTXHCGgLzNqdJIHnlQKFuoBWbPUeAW632mfshn1
EQOCWjyivjOJK4zjpLs1cvxqiTlxlDziLAZiJh6icOgdEEEzdf9MVVwFkMeF70BP
qlXyGm5LfMPWiWobQ85HjaWCtAJJirDIRb83u5XAnmx3C7bku3cHOtwUk1A0S20G
hd8gK5ZpRLds3xMHQ/eH1p/Lfh8dY2ek0DH0n/Hcso46zgzfQruqN33A7WIREufX
+GcdasK0vUwUbOZe3O5lU3hhgEioFSwgjioKvwkSLQfjUrvySvVKR0qu2zkDxMEX
vDS+hUwGEalO8Z4CO/BUvWrkSeZb0mK023W+C0+MR4S+Q6d2Tw6ya7qi+2TqLF0N
asYUSlnecLDAZWLHY3rrIslaopJd9+Xi2mgB/DP/RSb7LR7kFtfmVKRck1qaPMIu
9Mwcgd5RPHm81+nI+2KgW/XWh+VjIVRpf8fDFXcj10YCwhQIVGmTzY1GQOoSLBxG
iuobTfFu/QJTAPMk2SmND1+VFdzgTbun0EvNPq/rQ3auQHPgHTc/hsx16fwxcoKv
IhRI7VP6O0/Az3C23oFibHir7e+gH93oxlZb66fl0gVRLOED6QPe4R9YfTrPVJWu
nNOhK6jyHYEfRD59nf/iSDUCOuUZFYdpxAFxlHymRwFj4cHm65GEadxpi9CWYWPq
akeP7CKd3TiIXhRMNjN/GaXk3Bg0PXv3f7f6xbX/kY3VSno0C7eZNnLP597yAJal
8hEUcy31hHRkhpYlKOijxmnNyzY2yklE6BIZRIyzCEI3t47xipeEwORwkzIGGsP6
dIKLYWQpe4wWs6S11SuBPqssBs1yrO9EBuerDitWa5lZW0geplEkSlllEuwRgE9G
n54UE8oogal+y3MERZilfaAiUH6O0w1yE2GErOdD7FxVWudEGWaQPxEqExdYq9+7
Wps1rwGFNK0gwViZkSs06PxH0/xOCdVMHHR2RJxoVc317Rl2lTftu7B2XfxN2v1T
LjsifVsjUl5/5mgxMRxLNsR4bfSX6i8J2j3xqkvldo6dQE+z1NSN7UluYnMocjpz
fGowwl2jRnwlXUtxzVLH28JepuU1R1AJpvISnSdqBZbdbE2TZk6QcRghr+Q4YWTu
FoBKX4j4TKWRROygEUKeInGkMiSzW780KljYgnNhLraLbxld7WMZ1vafnmihxHdx
unkLrIQvSPEn6AFLgQDDbK2E3afE/kWInOK3VdLSzOvzmXqE+QtKrT5bFtnI97KL
G1tOIakKSvjyLW0YmRDCayD8G0gfuJ66Sp3E9AZeKCihasKNwRGAfmoIV4V6DQdH
NmhyqB2KraX+HXILMig5PEzeKsf1oAAqoz9ks9rpzNGZiWLwOnMcC/vojaqVcJj0
I3D65hcCrvQo3VlIJoPCnEip8c24oEpzyXRFtLFSVesoiGr2QSFb93hAYG7nwStS
R21/fUBwFTed8ixHPOehqiCvwXuwlrRZfPashVEgfFAt1PQuw09UipXhcFyxXImv
5s5lT0gNKMui6ANJjnHHAlfk4e+Kk3r6vHKNnMu8brntASR7Jb5+OVuBJapQdJ3e
SQkBt9cyfKLajG6CThNDMMN5J5bidYXpWE28KHgnXgI9CwFtLCNSD5oSmFKWPF9s
3hkv8MmmE6molYVtUyGwvzcD96hCw7RqfVcfYNuI72e1UozmC7YuX/0Du2I4Tvo+
ez0hDKibc3erik5LanWWT4agLk/oRt85+P0cbS4hCg60XFQ2Gsj3O+/xPSHAvZNI
4sifcWEv9WM38InZeaeHoezHS0jb/PJKMtKSlgLyLAt2DYiiTLwq+YEYM4D60dtx
UBeZe69sW9/532sejkhc7cCCZlhkz0rQgyswSmRYnJZ4+jFiDKYN4CgaadU6TLsz
KBIYk6CttC2/LtJb5C6rQIavce5mY1NyHtJkbIqYqkSlj5q2BPqw9cZmIhMoCe2d
Z0iWx0hdZo+IWfYG//rcyOT9ZJvL+QPj8cSWgsorhkWmhaXsayTMjOqwUMggmHYM
r/KlqBqjFNoO40UH3MNPa9gK0OuYn4sPrntzlguW86ZCZ8RQx1CwrnSl7BnoO9Tk
yy3CfhsBy2mgcUMPcBStm16dt/gmr8Z82INl1KwN0GKK2iDXyl1VNmMquCe7akUW
zJwiZ9GFW3nke+pbfcVswBncDLkrohxn0UPQTUFpZa5uNuozmTERKobAbUmMDAy7
JS5xiu4o8Wl41ivrnpJsw4BDNMdJ1b+QsH61bNDqU3bfUTVYcxx32SDZd92EUaJ9
F285O18+G3T0I06WYbVHWQuJaWP4lTOyo47O4AsBdfTmxwSjlv56KxBbbcvHZNPu
D+jMvlL5jPD6FnYiNyOweXSUSWjR1rP6gfiLYXmr2mpheIGctQjVn+LW0F3kvz6R
HouxyTP2kSvB8PzlXZklcr6Kz05wdVTe5+fPIBpvGdlsJP/AJRR4ClK1emjuCntI
UCvCYCv6dyQW10fD3CJPvUvD/wOY9mwgO0K3EQAtUtOH9jpu8NSFGECLm16Jum9b
HFO66aKeMJia399lLVeGPmLzIc7OfEHgKmurtz89tRrD4QJRntaY5iu3Q7khfctU
JIE44A+yPzZtbs5QgBzQynt67KOip9hvybm1QgLqGmf5dOPkcYVjHDE42Cpguhle
qAgzXbzlLcy8ddyKBYN8G3+9uCL8c4ZKsds9+IZqfelwC9diAj0bidEg1wvHB3cx
4ipLErqohRuNQ+DyH9RlFezrCiu7VchnPuSauTSIQg7Xp28VX10XEU5JUgh5vcDB
BhRCKeZXQYUWrrqUHbvRw/am+9LO18UblXt6/MD2EmMVkrbHk7r8aN2tD+yhY23X
tslJxzTBgIrd0zk/+zkd/5Ams2M6tk0w/VQi+56W58qgGad0+fIQMi/EzzVGTTRA
Yb50aOzXh+xUWaFcOXmE9M6vWfj/+IiMzQHWbrc68gWYUBLJGQAfruZYpR0echEA
Q6uCQChN6panTqmhoupt2sGIqwABqlL81d8vM17orQKI9nFqK/q8GJJshDPLMglf
ZSvBAJr0o6Y2dD8lLPfPpsJDPYym91J7+69h4fMcM2kTPsu+/zQ/Yv8wac8x9kKq
l5HQGm0IvYv4f1le6B+W5tGavbvVaNhrtTRAA9+icom2i4iomZna6zG+cCxtQn7J
QGOGV0Ws1C3ujMIcuqBIpsHMs8kxflv9VWNp40/PjJhrxXLlQHzKX/+7HkVRaRdF
+nUgj3OWktY8qrq1mLnlxBtlbObO3NfKk2chFbSCcZ02IwSuuLEbbwkn0QmmZQtE
kcm6Du1POd3KSAwwJsZ9vO4Y3new8C4mOVEAeNa7g1/zLUzd4o1HuLUWQY3AS6QQ
/JmltEdcwHMb5y7OtZXpACSpHXGR9pRpcmfA5gv3Dj98o/KQ1l0FCEt6wAWkFNuK
ZrrJCDddchoz1aAtYWYHqrNmj2GDrbgo8v39nxrZFUBHGQZLFjBBofwxvu9+TinZ
iFNWyx1yM90z4dQ1R9wVoR0HITL1rX8WAibdjCBO6rnxJbyJuL2alER9wpavkA8d
BH6rPBhmTegIX2uCL68kaA16ry2ia3ibNTLK2h+19Hop+LBpsPAcsorwyQpvstjv
ZAdcHI+kOpXeo6ieraVm3JEHmRk7G3Tcfzv3pk7JwjIx9w8kkkiZ16bAx+KFl+TW
Ecbx33NQ2qyiIc7I8ACdq3KY1hKKXigKycCXTDRnkq3CWp8m3V5knkE0dLHn1N5f
IIIzXM1vbm9C6tkIb7EYsGImtJO8ourdr9/9ayZRVyHTRstdLyAg70NwQP+Z4TYB
W7v+CBEke/6vSoLgCV9aQe/prIqfFgcKWe469cqN9CrP2n93En91YTLwHDrZqDEg
FVHZ40exlOogL408XPwSMH3HA2wTOj39+M68vuwtWPLqEkiUN9Z3srN/yikX/8b7
+AUT5jM8OF8LF1w888/Qcr3qyKLg7du+2EqEkFOsyVtWhEDxHD+VkA2GgNx82XVh
UIQ62ZHe2jl1wjQ1XNgDXQEj+qKWpSv/CNVxhhuU0BUgpT81RIYgqr0E7c586P7w
4EInFNEI9odAfEURCDj4u706q/aU8Rvs8ntK0dziQUltzFGbU7xgyL+ECLQ9RcVr
8SxsWhGTUwJYq+ShxNBPQcMNHHZrQGG3dkZqKxgDAh7Hj+g1JBG2/uXFKst1s0dq
H4rA29FW1O6A++Ra8DG5G0X/F2hmfiyY+KkKobS5xeneu3ECdvy8QR2/yEnW4amO
88cFeVvnwh+Kg6ZFd+lgpuCoPAC8XbVr5hCKDlZzSUNRZV1iIe2/pJCGOGPOF2M2
H/KMkBWAYbyzt9BYE2wwVHBUfkYRRjRT48iFnpj4i6B+lV3LbY5mruG2wBSXSiVz
Z9Zj0v8hEnQLbml7AeL264QRWZeKsu1CAMTm3tnsndToIa2I0+DTzHhm1LuYBUa/
T41zMLynXKIHmpBohTvy/qF7Y39ucPFcGOU+x8dkpEd1MtVgk/gqLeafcY1JXz+7
mddH8YN12DMl6cCJGfKikgiIG14YkhoKL66PO+AVplMUZALbeq9QSoXv+gqASJzj
roIbc2/oBoMlrEIaHKh+tXgxB1biR3wBQH0Hlfz2Hag0rc9+LSy1AEP4ATuC3Asz
x1yuKhPiPgtXdv/32kVYsZnbyLTqoqMI4GOq/O7iMQnv6Eum0vJmaMtUHaGl6/vR
Q40ypOtn9oyIFREGH6QCRyF4vLjdi1dRqKUiC0iPPeCSsuHeIzOKb1ezWO2bxRwg
4X3xSbFLesFtSG9CrXssiR/opf1vUxZngWpZ1vTBdqas372zdDZK6/nmD62bCiIq
1IqRCp2M+tHTHlwwuqMSc4xwN4GLwqLdiEf/7s9lFvOLInwipkFnXT9i0jH3YaC7
pVXRi3W625Qv3ADy+mQKzdDJaF7ToQlH5a7B+D2EU6yKMwKx0FJA++LhZLJJ11VT
uubdl37OYEIAjfhmnqFJHfZNI7ZZIKrD3iDeSxyszSRcV+1QthYpaFd2hEH/6esn
IN2iKVc8iwgoSyYJjPTD90Fr6UA2AJkY2dcq2Ok8rqnDYK8Ad7v+BhRtz7gAQZFl
UKXfZOBUY8dx6YyHgpU4JZbNCT9yXHRXCqDNWsT9sLhAscITHaGOl+JXtQ1fa7bG
gq5SzaQX9+eB6eVw9MQS9YGN8uA1rj8GVVaj2pJDzMR04EHrsxLTjGxl1aUA+P0n
TFavnBdHN73hAHO/3GaRsEHYHst44iVL92cWm8WJx2HH+VOudEXDN/sdGuyYpofS
1tUyeXpuSoH9pd/B0X9JdQiYRNvCtMZ/V9heCqffav7EIqVMQgnpCFCnwYeDa0us
QthLSNgTCQnuekXxtVjjOqWTTg2Zkz+QY48qdDYLMq3AubrZJrseBD+5g6lzLKI8
QxCEkfjPS5IRrsBBP16RIt0wfpz8vWohBj8f8rExbcZ8uV+W9DlzrCQYOIiR0LmI
2s9udEFvI+V7uwj4i6HYT6fu5mDYd6+aP15AL+Vw5w8of7D7ycMJZgt6D8biRHmX
fzPrEUpqujvPCKxFgd1YMc0ksQoyYvXdLGEcgg6E8QDkG75DZrwFHa61om6Fx5nk
vPdzpNyp3i9mwrTufEEwmUupilEIR+KppQ+ypWsrj/5rnZo0DmLLSar7I5KA1mQE
2Mu7DcoGD3R64ONBtkKKS7sE+UkZc8uKt4X4mO/eXFegkjhCGMtINt36tSXN9QVd
bGGL9qGM2x/Ys6XekBghP5pOK8MwtBB/Gs+r/CaJxGQeLrKI3llLIOhKTPqb4hjR
BqQQNAZnXoFVTddL5bp1CxwN6MmBTGcECEApwwo1CnceQsu+QppAG33PPKODzE+C
Zct0aKXiWpN3B5KZWjmIa4j3AhK+0FlzRIJcUucHxhhAfcNp8AVvARsNPVjIzuB6
Lo8r7EDfnthubb2WRR3YJ5QzB+XwLMssqVow9pvf977mxIzbooycTIiyC8Pws9vY
XiOt7uPtX5MP+uwsOnHA1TUcuZDxohJvL910kr/vorwlSCnrpEILM+pma1TvN6ZV
tYYxa+epuqPNU7+tw9m7ov1l8pG1C+otwxaOIA1sLAeXr0tz125Y5ZqS1pLVD8wd
qgZqcOgUMei8S8F8eGmncHU+oiUAYpUdC20pLOvPG7eKWFjaXMGs+8L/j4qoEuH0
2laFUbatV4E3ODeLZNsxKGV82nQ6HwPmGQVVvrKBARtWjulGjXt1u+imz3F/nLCF
MjnM3/MmQ1rji5K0KJ+bsJjdqFOyGseantwDZVm5Yb600cFhj/gcRCImVIy6RgA5
/vosywB5Uu/Dy+HxXwz87b1Oo5PfbB54I6UADDW4ifL4mCCKUF9wWLzrxzyoEZs1
EQgLhKjgIKmTc+vWlQW7wNrTKQtBe15DCyFaz/xi5h/GzMlw95se8QkCuZPhmvyt
QNpZoU8VyElLzcPtQTH7zKFYOIK0egmt8sWhFvZmS2mPPXuC4QOrVXR1ZiasN1Oh
OE/Vi8iL18RN7A1cNJIB7QlL2R8eTLItInrNo+xSsyog6uUjzKMuyXVBQ4L/8k5O
RVhrn0hEGSIhGP5TW39y/NVHwjyMRojZ35AyFQINEoBFvZAH+61ThUGx1YmYX0rI
9i1hHpqmkBiICxpuYZNn46VEaDrnxuq68jHNRVRVoUjrvGYvReJGi1jkf5LJ9RW3
6ofC31FG/3zMBS7FTuvNFcJ6kqhETEHr77TEBQKHfqY9HIDzBIC7+civBYrrH98U
12OFtWgnYwMRG5Fi877BToGg/PahWBj1A2/rl28k0NWejmNAjv5fCPABtfgyN/WU
UcrpOAKWFjMkyndlUHxL1HIvtALI/NZG7z1+5yYvlZ/30I0QWcUUYVkJY65f5VfT
gXMGatE3kAa2N/sizMoXtYgHxSMn22w+Wjfjofxm1eOhqsBanPpCoYbl8i8P3pxo
YGy92sj/ilJ/lNDkqFIbH4YFjkEjqYEWgv4DV8yx3QoX1aozVr5O2sckiJa1l0Mc
GnXmeH937wDbux0Yp0e8zzXbEu04fLTf7c2TO0ocwSzK8fgfQ+u0Iz5yNdok9mpM
BSHg+3xOSP4rgmjpI7eKgt1LoAU3l56roIlmnsDjg3zcHFUU3btseYDHLMpPsu4f
/nHCJm6nBoShZm9ncRlx4+zi68qccdAJyDM6ePE6rEdPgjB08OzNtMLNaxOL3PgC
HJbPWM44HLaYPivYT3F5lZlT3CcdxlyUlq4cbuk6K4CymwLH+/vnu3UUvz4AHWYc
SXCJiNCAY+wforoYyM7wAMf7sLaQ29mlp8DT06d8XeBMJpPnWGSongb5HOYj6QuT
VG4rVZUSkp2qL/QwkZ1FRiifa4B22zfgBPS9VfuCekNzOFk7n+pdm9o9mD85ejbB
tELgPM8zz1PwvyqJm4xHDJHrHpunJW/HWWwmheegg34wtcQqsRg9E3AuR5pDQQQT
LdzAlgwd6ekZbu4dsMCe0DOR4Gqw7iN3J6lH/PCTBDC8GcFsPwtOQ8W9MlP/4lbd
qBTt3KXCrfDfQCwRIt2Nnvwn12FY1OAjuhMqEtTWVUe5H9uDFJ+DJJkaEs9oYTPk
cuzt1v+CYMo5p3HsDuDpU2mAUInYoxfejMdryMdxJCMiW3/3brfjpNMMOMxM/pKS
CAnaY9HZTvwSzNJf6FutvZ5MjknRSLC0guqfQ90+0B1l1vWLHFMf5nsNhK7ju+IF
npMfhcyDSTXqeqtFSoS9FU92JxWFCDYIzWp4NQB4ZIbcWn7lqsw0zvl9wyovPpgL
QkAzmZU3rhVBJQaQnsW95dksSbkDbnjXh+qE4dQ2FfqyPnXSfJx/MinGZdCJP69S
v3OpJlybiaVIlcrPAi7+GQI4GrsFBSgZdc0KApOKQueyP6Ug3YR80iFOrRLnXNbR
oARsWkrsRPpMpnXNEtPK0bEiuVD2tUcTq78NHlYmY+cFM6RMZlHUpo/HbPYQHJVk
8jGfEchjRNL9aDsOB+hFhFnBfUZCGjRXmw86/85sBMArWkIyAtB19Q1zJkU5QI8e
RRE+QhdKFLe4saVzwSp/J7y59t3YEZrHGaDzDeCmU1CNLNNGb8eME+ydWwlx5y1F
bM1GKEyrFwmcPL+RhuKBRGJ4r6HaFPRRN/F81j0/2kXAL5NzNBfFiwXPi4KrsqAC
hvJhz/8s6KiLt/6UKTWkc/jN95bBwz/LBjhnYT91qMeUtKXUZ7fBLI5iDJ0Pjrsp
s6mQJvyzABqrbhSh6UIMWndqTVunTIY4fIzv66F1iGeG3GPlxjRd8Vij7C0SuNdZ
rsFfed02yIRe5EpL6btDwbjignJ4kibvb2vs7Rhs9xyBGGtYwTy2qwgTjrlm2oxw
FgD8EH6/CmkHKvNlnL5en0rtiiS/EUjR9MJOlErxvSQRJh8WBRFe044ZYDMG8nrx
d20DPuLsdTHeiFGH9mCQB674uRxjdgJCa+Y7wsc+9DHgisZT1lN2R2nlZzjtxu/J
5jCyjHJLageea4kBLHLveZPwZ198lhKoRHV48fXTrNfynDvd5CzOxpHolrgC+dnn
FpCoqw4p0evaqGj/O1mZocOlIkvoCUu5pXbeZ7bQcl+LmrNYphWmyVYxUudIcKF0
sXPQopAkOVKD3uOX+/Edu/SFz6XgUXfiF1pcmz6nb01gqKPOXlvgRq8QP6ia864+
8zKHD9LwY+8rBEQ9cEo7ZrTwbheTdWSeFbv2oysp2SPdlkO/yf8xgARgyVWs8+3V
89lZi//z7YrmC6powjfydAg7afY9Y4kMZQsAs8nlACSvUvJBWoaCNAnZeIGPjKt+
735fgY3Rx3YPI4+p8r6P2kN45qAzK/30fY1DK4RxlFNBUfqwAGBMMXFFMRzsLlXp
xa8f8BM7KW29JGr/JS+n23By4gk3IWFGFqH03re2jVXdhvQrNaQU4tMkimJHC1AS
EA5C6HKHIahvQ3cTPTY/iAcbTb1zQQrHPjQ9rlS0f+bVmFDibV8VgfxNjT0GPgCM
qcXYmLx3HUd5hly2m8qpeybreiAk7lyq7mAxKMIA71s2sDn6zR6koeBGgKpBI2C+
34v5cPgYVPfyey4Qq0hohqU7fcku/VG0wge+snR0I+Mv/OgxZ8F9ELA126ydYLK8
ozIuD+0i1WRB42+efKApteujQGTn6kjllxSpkD5ubWeswHWDc3fw2tLFrH6yrfTM
mjQXQwC0z9a3hq1O4em1GvFlFMFKmxZ5oBCp+QNN5RcXVH2XZ5gkD+sUHTvzOsF6
sFfaasXppXvJtK4c4XbXFYQemP7MGw4xlzzb1thM/7YPrhVCv+M8u7E1fwbQ2j4H
7h0vTl0gsucdHFzQ7YB1OivIbPIv11sF7CAsvLGrJ120Q5dIDcy8ylA+UKBgfSsX
O3PSZomYW1/HKPjs7TORFf07e5ma6/aVP9jaAB4tbYCI0JUvqez9evoIvsLP42bK
Iz7Hnx/ruOVizYCUm5U3yWDdMDMjd85vyjOwy1Efqz17VkzZ1P3+gK85xK+q87/V
C1i6FLOWQA3VEyEt8S8I0cgvVxnxtsFcypRarx/RI0nUF1ww+37V5f4Y/F/yGDzP
hU+xDa3wEi1z71BB3x6Ed18m/vMNr1swGKQGkVuocTdoYz+30FWNleF7q1ld6seW
YBTH9A5iz9oG8igX39Zo9O0sQ0DKHZ51UR4ZhiFxs02o9fRPBjrwI0yErMZLdchI
n8Swy1F2Qn7A0Qg7OENn7S5B16h4Zjwo19eAWZTaAZ2mExUWkl8Pw7K0kUU2+AHg
aaVV1zi/SrA0R7YH4TZkdvQLQCOVc1hUMs9UfhP296cKuPVo8L6WGXsvSb7or0SF
+FDQhJ5/1pQZBzIwUOyLaWRUPV+2OgkQ3zMb3IUaaZNEBJHqrVeKyShiB0y0G/G2
fz31i5tZJVOjdNbf9cBHGWQAn6vHNtHftd5/4ROgN0QKQcfZvebPluQF0uU2R5aq
Hbm2xE+kSSRu3xkjfJ6+wqlXdaSRNC5H6rUhyjKAAvaGP2ZxDlgT/cJY/ixRj7VA
A92jvCLJYOFB/JGnvRtUWhzjuI71erd9E4bOggl4FC8WKbjT0AreL4QgRKwubO/M
Jr/PsKZ1cw5/KymmJB3c7He9/pUA7xD0rIZERNMDR1I6v8ZTmYWalWNzuJJPxzc8
ZUqI41gtWzCFnVQfADAd5STyrZEt2Wr0lfQLr+YziQd9fH6QRpLAV944+wrdc86p
ObDvOFI08wD2YyACSjeu7OW0MfbJhYcViJHG4d+KTY+dTa3o71rDXVefP+c8zvWd
7LNISu/k/PewQO518ABta/BVdfHpue3bVENmoRQVfITAjVgWVM5tQAOuiptinGZC
YA7ltZSROaHvXNH1iXpcA2RjYnQ6thBMhngUlphXGXEVcMj3llUfe5NBlC9Xqs8k
oeSYq9bp/HKD17g9bohI1ZZbCTClgRqs+YiYRZx2ssCmJVDnMMPkDWu2E7ZPZiPz
mB0aHExCAzjDsH32OXEm/8f3+KGDZF+6vzE8Lq4BbUu1A9JA6Odt0Xi9KlCquTg7
I0n7dvXF4cbyYy6BI9ONy+cGILUaVy1+JCh94TBJLfWPR9GiP6w/NyqOzh+Y3z82
teEeot8CwKMlmqVznc39UWNVrY8FlJAadqvaqK7saao3alGJ2PBIZRArElzgxE9h
GOvtqmSV5MLkRwQBGrCy43RIqonKjCfiEyyASXHn8y638EH+TVgvRa7abRTPLFq3
8tZaa42XHPxCTTU6RiykG7XBj+Hk3ODl1cP5nNPO2qrxTQLh56uufz8hIE/nBMLc
1bFlrH6YS3wzTp/dDOwRualru3D7MyIC3dEspaTqNVyGsNiAg9ofqM2uMehX0Qoh
bPS9Nyx/Xi0j9xOB6xqMVHAKTI5R31jxicHwbT6ttxTEvxwxO3lK7nPaHT6YIeqT
4jNB3/3VO2R+t/jA7S+zxzpjkF9Jsfp913EAD33gmpvNCiv6Vf/bFwdjUIhgc8Y0
lHNuLJ546Dt9ONDZ7fJlHV99/6135M7XnoazWmA7zoSm20S/q6Wj3aq2MtUgiE5N
FJ25TCjDQt+74PhUNdfxfcJkhDr44kxcFV13G4AMOxLk4vOaX9jXf+IQ10OMS7v9
ksN10SPRcg3soJy1xGaxYId/7tqGPBHyulO4aJACfWVI97QCfH0DVwSkpP9BZCru
ztdgXJJQLSh2kD5NZ6PbA7J+7hvWbQDF0mbVpjmbzp/6gQt9R+du9DKO4aezs54s
pD5qbu+SYVTkHm39i5xmQF0gr6zOdx2KVKRZurr0E0QMyXweVeQDEzamngefrTYs
CyA6pZBaPoZgbwzIQSLT1boFe1NxlPMbygJM6LHy1QHMKfHLWrjsurwnLL11xiaj
MgG64XXhiAraBSJSORuJef17WXFpePhC5vw6OnQdYnEVDofKM3LF19lmHzIpXy9h
k0M0QZbnoqGdsaOCEYRLuIQaTNCgcPAxFNyNwlqhEnqiJSmSOFsWI9MnrUfUPvIi
7Icj6EmTz7Z0LP+vjJpDybK+O5FndjL1S7yS7aJJ6gnFyJXkbfQlxepFBn6Gixba
4y1W7VGFUf6usPAtN6dBXd3kfQmGqTA7Uxb/5wdUJFwAsjzcAcJ8xOY8iehmEXiu
sVvbQGltOuK0q3il2k52+lpdTqdEzaQSFvlsndHzB1xdsPMH5PBQB4ozPNZMhjCy
ONCtPfMAtvXXf4wpJ302ifi+3+MrypTeHEQMNsf+v5a0HpJIsvHgNXoeRU3ERrnf
MozDwZlUDGD+OtXYS1DAQg6r1lHKob0prYbGxuqmWmh+NucEc8RGO2aF0YGnS+aj
a012LqvIB8rwoHD82J4t8Fpc0Fa0dkrVLJG/nOJP9CO81+arUrX5+F8fRiYYzX6e
IoWPt9H52d8ik397HxN+PS7jf4wvWE1MRrOZTHLCTEd4h9FJo2NQir+FkJClRsEG
l/Ua4z5/IkMNgP33SLu3rjfBs3Y933Xap37b9X1kM7aZqiZ0HZ7yikVpLDJrJ6f3
InF16Bx+u3SWc8Ie5TZaqamEuIa5mAGVUWB/v69Dto7+CzeiLgzAGE5nTPlBUZGl
2USJPuakha55K9NKr7qbMC07iJzIwNDbbiMh+Aeq+Mj43fIcwpEi9grD1nVI/43D
4CoKq3RCFUzCd/Z/2iVLOmXRP/iQL6Q8VpWCAUxcZRIYf2eITTlpPJaSszxDWpAV
0/J5ojro8wmDtIBbu1sQljSyETTlGhRGShnDcGvt+RlkFWenW+EV8VrMqvw6ufsA
dvp87bdk0ppwEsD9UosLiMPsLhrBYLwUlAV5FMn66Q/vEtojCHKmspqH7HPx6SP/
rrfwVfj1p0xw9uLoa+3U1QWBF96dpYVRah0mihXHQiaDWcWJpgtyo2kac+OE/TeT
NTKjIIivAajK8ovoTfO9d64Oy8dPDLLcaDmtYruoo6V4TWY83tmo4a0qZcaYNr+5
zRMckUnDBqi9J/3J5LO36EUWjD2b2+8MFNi4GmOhTlV77H+fefGC8WDrIu2Jb6y6
xz0G9tTHe/N+gvLBzWCmJmznTSJmtF7zPTkUJ7fAyWr/24+oj4gdT2vrUCPtSavp
3eY89RL+CWmppgf1glBiSB3j4dQ6r3aTNiLXxssrxHtPR0C/xvxYPSll2ORT3s6Y
9DV5jjYCqmAAS7cmtlp4K2Q7jQwYlqDSRJ2d1fzDE4mE4vavyyIC5jlcI3J0HsOw
STiyv/Ye9OBP5cpi8BbKEdB+oatOL6VUoyPPwsFqfLlvyX0zLiffE4E2flETDKPU
oQf/nTOtfOxooSCSjYGmvVHEwm8gMvTiavWoYRlSkr9NBVxaHaVn8ky//4WSrYqY
jekmy7awma0FlAjCnXKqrRqtgHoVs08K2FFchUTjpvc0ftJlYT4ncuV/BNPUfQwt
INDhrmApGF0sKBv7CMwtjdxZf+fNqvhh8dEEecxXHsHccZTIsH0WXzrYFY/cybNv
Y8/2mWsCroCIeLUxPr0CgVpqMo3FRqVRBTguCDKYL9yzjEw3e1/nWnEDmFiO2geb
UPgCkjCw1hgL+7tRkA+0xdQXFd/tecmBYoRM4OSgMm/UnfEpHJH21fgT4izFOlQ/
9jEyC+z2mKFAfAYgxvRlLvcK9nucfyDNGob3oq7F9zYZa5hnMAuW6N5xADghwflr
LdH/QgPjUi27BDe8102pRg+RtzPxPZ0TYDDjhzD3Q/1IuEeY+OGMWtXBN2qQwk/o
KHMm9eaVSldk11rlg0U0ss7oGNLxBG5Zp0SkH5CDzpYIImq+anV3JaEkDViXV1d8
3GP0PVbfnmtyaU8y1LbN61TAReMQYai6wppolNko5upSkFy5igHvtXCIn+XfA8xa
cXXouyXz1KsFbxaO9ZqXUb4PFXXnVGgRcMMNmw1pP4pG2Md6u7AZ+j2S/ed5NDKB
CQVdQdKl4niqg3D2SJRtERcNo7/xzSscJSKMbwas1kzvD5RJ40RtEMIxadhA2Emg
/EEXzQJ9UHL4ma1zZ6bvxmDvOrERyYUPUmfXV0s954za40fmgzLbLr7xJeqSB8vf
Ivd5xVBE2Mkl2OPJi6Mwla1g6Rp13/8dtMqW9BqmXcVNlzC3IQmvd6jztZOk06rP
y3jSulb6qM6hMwRfK9mNRnrk3/K/UNCtg7x4LKDCIv0Dr7i4nb2zsysYuuZURvHS
juf0CythKVfgOscy1+dHPPcgOcLa7qpC+2gKib1RB2ZxwdTd/ECN0JZwQmaR0Hnp
w+PFuofr7Uh/9C6Mu/omaIGyJ5/pXFocNynAXOSgDItwFv5Z3OgE7/KTy4/F0k7v
cOYroIo9u4FEgRxa1ez+pbQKuUDqO3FN06JWDc45P4hBdpnM8NOBvuDtXLoerfii
62EWBjKJjFkPW5uCIE2P7jxvx0JNLx1ylFyKr7Z0WkSZyNmbZ365kdQhN8G2Ioq2
wYI6EQ3svICLsBIL3S0FyNQs8eBxV0Of/3pu+a5foNOFRfYoY8dL8IYR7T/jDRIJ
nV4pYrf3B/wK4kUPbgFvJ+my2E3/GuuzORi08JY1++Jyo5+UtmZSW/8MjwxGjK2B
qk3+PkD/pDxR7oFaNzP206NoYcH0ipsIFbWyD+AwXM91JEeCWdzgHLreI3ifIboH
8XPj6yvQ2LiSKyPuFrrQedWNmxyDiVX+sMbOUjNaEKhdo5rkdz1VmoeZkmSv5Z7F
ehmx9Hfl1RTnSxUcu39Z+G3Qpo+2pHGzNqURi8AhEMibJIdRGVFLILeNAp5VADgG
fAYkU5ihbJ5NGpFkOx+B426zy09JDaXDjV1uw0ib1C9HVJPHJQ7+wMvTwTV+ysLQ
n6UQHgknmFxDtpJPK///skp//oUyh0AZcHg5RKVdf4COzv5bVOcALYSD507cMnN/
DOo+uUnhjW5f7xWr02siM8kGbM9TxYv9CUuWcETVh6kTd7zTbyLUb6mxXf5vJJDC
HUekBZsJ/xO2LsFJQ/peGwdn/O5MVkFa2dLvyvulitmLjXCEeNCykdCNnbj35vhP
ya9qSx4MwxjF2lu3gweuTEKrWJcBvwMOgUQp2KZeHjlJ42ECB1pyD2ckJID8uDEq
e6FENY9YiumtKFOKLJbe7i+cea7H6VYksf2Qp2UoZOFI6WXoXtzNvXPeS2EDn7uV
15wGxlPclihgGNoQm3FpkUzLu9OThI3L9I1pgMm0xtsoPJPCfCcO9dPqZMLKWSGD
LWQsIsFsZKxrK1T2SmTRPNH+jWkQ/2XPGGaUblzxJiLJ404TeKNfBhMG0u+MVabB
BilrWtJu9D2XAqvQvbxusUTD3/sw5Nq/FAkwZAaKFZuPFfBVP7GcNhGt2mvQn/Ww
aRO0XLJ09P5b1hX+l7PNHC7JBr2dzNf+t3sSfyyYlMVlmEeaAEnCcvai5a/BQUE5
GkTi9zUBTTrd3FgW2rbvlmmqzsirza7SVnUqnLHIucQwwyKriHU6n6h7P7pj9INK
QTBZWgZVXrzo13rpMqXLAGtPflNm3+G+VxAw2r9bwon20Qmo+SqoexFlqZWj7xbz
OI9jYX05KcVxysZNaxttQ2mhX/uDrDWxyJiRQxvtOzDIxVopeopeG026/EGK/4RN
yGUEmmrda5lbHr/2DrooF8BZnACBFJsfhP4HeDKr8XRl+tGuwhNZ8Iuax3Xkm3Bo
p/jEA/Xti9cVIc0Aq1oaN9AKXS13VV5t0Yeq3nGUh7cmJRPmTM7dsPTk7Xj2tBZ5
IjXKTgPkWprcDk8JbaOW6UYiD/E3XDnOlm7d3rMWD2u3FRADVWm26/VCLx5wiMyQ
JhZLmmt0StcWAo6YpaaHgMD/DvjSLmtxkTWDPmG/Cqa8l3i2gNHc7BjwoAWlHBed
qY/8wltOeTgDJhLoQLyfJtgKk6FYnZ+VTpzziwqTSysMyRs/XixRNXH6+EgmzeRe
8+cuo6RmloSVr6C+vFZ2gaalI2JUNx0VCrptB99AamWbcJ+Q6P18xLN+SjDAmL4+
tQMpEn8ilJois3DPJiB77SLnsDLh/yYLfrckiV2q1Vn2TJdpVAC5QnryoM84DH9M
vRJxZNIY0ZcFttgELxwEk+Q0uNFGST/Fqrz3MkXtksbbNrxENhuTeBFO7K3ve4UY
ojSXcLlZCzdOZfEhkvA3SW4nC/zcxZUqRl1ibwxQH3kTdL14YuzW/oFzt6dYn3Wi
yaOlDy7B9IaIbzsV2OWzf5b7dfMQbOMOK6jUdL/FlGIgJQdXOnReTohzs/f2mxfb
HOyjgbBZfixCY2n8iSvuMBPLRztoK5Cc4fkpvEZ8mG70lw1JXg8oid3k/PJFRDC0
i2JsDBGqawlf3sj/0SR81+eW1sEZRKHn3ejVs8RrxdsFRBX1dlbM+D7DMx0sCuyP
kyIXp0xkhEpFb5gOsxHT78sg0J7+Qdxgv1R3zb8+/mTDBgtDXoICYGgbAY2VtBoY
x0zuyJ9YVDu/j1O6jh63hgEzPfYNf6pXDhHYEwk6zsWu7PG7PI/Wu88RTK/Ezi2H
qQNMDi2G9XdWjz+7/t2IgvOf3oAWy6W72aV61gj9ePHtgNiVgzLQsgfFeInD/1Ie
Om0+LwbAuqMLf0jqGM+i07PrajDG7wtlioXJYDEvGj/7EW/3BVEF7YkUtXa2N8GD
wAWYzt/a6mIiZJu/nM5tBsURGBxmiMh+ct1aLqY7iOAc+Uuk9CmAMfSla7PBnDJj
Wcnfeb0ndpT5bEJMNAIKkia8zDHQfRxJqvnpfHYzzgTy3DvDDYyCl4zZvDHzmRVf
88Pw0k5FsZiHSoywM5OGJgId2CX65wkYJmEb0A6EdQUOP409Td4RPRLtUqlWKB+q
YLAghChD6rh828viF9OXwCgWkedj2S7nIDPAJm6+dWEeEESUXsl1E0fP7c4S18Sv
tSN4BvCWDYd1R150iRN/2dnDxud5pEiVuutIVX2TDzvLlAtslCQH3VORdEuNjYSj
vADuAR3v2MK0e80N9UFZOUHxVmyr7FK2taO9OSyaGplrVDVKKw/3Kk5hRLwhJC1O
aadBeWD7Qqy54sva9w4weRS+YAbI/lOUtDm374Psm9U8EdoAOgNOreH+1bXhQmXQ
UGkBJdGyuIpO6hjpQWP/CH3kk8gXbZ0rY8F/nJ8+z2MmQFIBVblGPvsEjK4zs7s9
4JGgXM+6+8its/ir2XlFdZD1CfWSiBtytygZ4ypTN8Al5eb3A6AVzB7//ykrEx7a
1Fl0XrwJbIMEDEqWCeB4J3AJq1qVJdChubcjJlJCSQcmi0nyxxnn7CA7tNEdVi7Q
B2GYGdr0KH5jaCY2Yg0EE3SJWm8bukXDIjnbq64Zs6UtTR8ZRH8W1s3fKM5Sz91j
OE5MIT/G05y8Z7oB9Gn2IwJJ42Kv08A2pj8qvN5M1R70rJPmAiaqWLFZqrkwSS3f
0HVOD+RKv5kxKywcAPKJWiS5TOhLCeUHD8Z073my3o/MHGc7SLMeB4LsFIgfdIzD
nMTChu3xeljWAapASb+hR8HLFwZiEE/+8HnXr0tx0rjrO2xEuG6/3nTwhHx0JsRU
aBbrqWnOR0TlwuyN1wNWHs1dQeaN92+/9NWkcneXZljReKW3Dt/unJ5q8FJ3xU9a
Dgdw/lA/Ar9EzEckUZQ/3gxXDD9SBuX3XF+WJ9FIGShaq7wk3umzEUjtArNjtwv6
RZY1rjnz+xiGaxEwFMJ3SAlEIetkZrepHt7OBmIKA3tdzdG2c7aG1SiTLkVmse47
MpLyHp0yyntyexPiiAmOQkg8y8ELWQDiJhkZvtTp2S3FBuWzf4say+5ndhLO5ydK
Vkb54GmPiSNRrZxMSFhhzbkx8X3XlXqEPV0zmMP61+eF/92uaYB2Oe9Oxk1cTig/
/7ZFAW/6S1y7qGy+7bjGPrf1plOB/lfKJH/8ecmeROgnXq/Wal9ig+BqCLxLIYTm
lIpfz903duAm98Z4nTqumHHWmacaPLyngf40exhD+SECAerpC8hX56SlEtb+2NIl
lBZTx6uNtTLn/qOtx1KVYAKg6JQW7Hif7s7ALw5itSt5LEGrnxdbF5m5qEXAUV6C
B47rmGV/WcsTCqxJVfImcBw4Ajg5JdzmxfuSbUFySnfCh/7vyHj4GuVDX5LY+D4Z
7iV9lDadctoJivqgUWSCIQ==
`protect end_protected