`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
ddtXksX2+yylW5zu6QL2Lhnb2d1sD00763mmSITNX595NcHTEkwn0zB1Dry37fOW
FufOhVzEJp80NC5qZ/+F0Vk7Ik02dIR0elf3clrjeJRK85K4e3Hoo4xn7YbFUIms
l/8VZSb14+JVGURjfswrIyCUotIzlzVYZ6gzoZwDXIi5gQIBf/gI+KxNXPaKV+PQ
Ufys/12rjO6aI/pPlqSm0hCvftmBcnezN2hk1UeXgOIuKZnogjOsf0iJVX2aOOWE
6pD/psybjbnsNB6kH5uFTA5frkzIzkzl5d9+YDm9OyC+k84E83I/7/j+rk4L2dah
QJOvksSIzN867/4Qt8qYTQ==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="MvBXkzurAa5VTw+1JJ70nePUfoQXBvZOku/SMmg4TwQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
oRtzZL4VJ4iwysPsC8SXYCzXS8Fw2gtZTOskLcDV+1B9Nzn1zTyNtlo6lNICRmmK
ZRVu2BmCc2G+fmzynYlNTnSa7C0Cuel6FYpxCBlOuk3OF2tzAmLAuDyOH3Z1Yjzk
a0aHuoCdIRKv7BrZCdALt03JeUmXKPdOmIlkVGFl8yw=
`protect rights_digest_method = "sha256"
`protect end_toolblock="Jn9CQpRhJt4rnzZPRk+dOpzAubz7omckX1MrFd4p81o="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 14112 )
`protect data_block
gD6l00tciPUa6pDNTk/+t0OO0nC/UTtBwLB41d4inuAUA3i/ALrNyoJVcBnAmEQW
ptbcNp5fxEUJjnOxnedyZEuEBxWRieZFQnkRdF269oOPlFUIuoMSjYPKHVkK4Twb
zdRyiy6iypSRisWdVCYjWQHDAyLX5PAaXDh6Gw52a5t2D9eXQIdMbvHks1A5h8x7
RwWPsT9tOktkv3sJyX14BZpgUJxDqcUOUVvX3dRNj8ob/dX9nTAfuQiPJ+fcea0e
7jk9If9Gw7D4AzfX2zHU5naqs6XcuYSzUe/huZaaj9bivaXBri/vQf03enCJARik
W53phvJJu6uAdYc9nxKjOePjpuTQX93WYgaVdEuHqmYf0ZA97FTrZtrAs9KkjMTX
AKVj1KTvQNB56tHD2UR6llM6XWeTW4SvRHi/oY9m1+92gUX48yuGnbuXVEiqKmmX
Xv/SwibNa60+HNULGYH4H4Tz+2dRi8SG0sBkJyv/dP/+TRxMcjUimBpGZETWfeJn
1MKPaNwDEEb+aJXRnA447BdguOxfoTnK1M6VAog97TkdEnlcdH1eR5JamO8Ji2Fc
1iQbuOJLOiANXxrvIC7efER/tAe9OGhmUbzv2iiGzFoSRH2jyMoU/e0uYurZUDgq
u2W257BTJQ/RXBHNpUVE3Iewof99gu7vgG6WDZVo5o8onl3QgV8RuUt4h90JnlgS
fujAR2HdcHv7UoPKjDo+0JbFmD7e0Pm4JEwMAgspXIWY4c9RKVw8VZVz4YIKXUsC
TZAjSahSCza+yW96LxonMCGf42PwLR3k3EKD5dJMt2u4tM1tSp/BLBMjFGj4b+YP
tQtDqCzN/ZKvHkkSYaDH1ApbU0EzkAfcXH9rv6kP0P+OtgQNLr7p0wHzSRO8QZVH
A21BuUkqDnMuo+OqaDfCjicILa6WcYGtBk6TouQIviyNhRSAS52Sf6dMu1T75lXt
esHwSbNevlOCJo6lpyK4kpbNlhWTg0qxsaLj2uYxTeQDpo6mRQO80BMeEtKHC9lj
xw1HT0FmLUl/N0ngsziSHoHV3vJoTGzjvL9uQ598NjuHDH2MfsLjWQo322KPoa0w
NjycBsdkWIQrIZxBDCL0Q/AXRSQfRnD830TWjDJj0BVE4a6g4PCCfvjArQZoP0JZ
MmTG4zXwCW90mezUhuY9Qv+pU2DZEJiyygLJDk28MSdSBkw9Joh87JYmfBn+RtVb
2jGnjf7cv2nlaijNfuU+t2iUGXcp0DQhGGEScpEdzW0rfHYBZAlgyrf0ovzVIrcI
A1lOh3z5XMiTkVGrE1Qya23cWC5Ni5s4aYjhcO3RKVfqan2W4dwO/Wymmumca6k2
tdJ6VBDUXK8AP/UFR8k/AEoLOS7JW1WCsil1evN3sb6/CoFCJ8oLgwy+JBLlcwzf
2Dajs9aCqRuad+yFWHXDjbGuEkbmIP5IJCjXnmEFgpDgJAgXkWs0P5spFmyvm1ec
cZPmw/UHP/+Osd5No56KL6BUYOdQGnd8WGphMwXY2QEuOGi9RNAUkZnxpFf7T8ot
umAzKF/3FcNnm5n6mAGNKeT+4pBr188C8hoIEaAC5H665OwkXTzLvSutS8I9Ed/I
9iC3+QmDGFmxgsk5pIvaT7jrt9EkLTUe9GKji5aCGsHfYyyA5pYkRYED46eqImIa
Zo37v5vSCEHSqPQxZRBkrItvXv4TBdJojRT3BeZtsuEvn1KUroHMnXh8yl4eIgBv
Vwt9T4l93emvTIbBN8wlikqDASEJd4mZ0ZRfGiz2dT43QAgpHQYt2JQFghilxun/
U65MlcQGfFkb7CNp4dpjzKkUTBVHh7wTwqKZjJFoNAI72DCoVmm4fuhapXrq5Ntf
OKImi6OSXPCkaN6siJyo9iFJYZ8mT8Dfc1vf4Zt+cLfQzZSpql+3xf/VMvelAL7g
8hCOMP/EHKpAmz/o/6XKTxKeXP0++LnBTyRv+PISnPE5tpa5oYokTU1CBArbDCyM
jYuGBaZmKCW9CWA5yOaj6PTKJGDa6PfSZ/hTZQ2vc+LU+y+YjeGRE35T/a5fQhcZ
3+VpnZmZOsfIrViAZbjHLMQair7TmBwe1u7rZ1imcAG/eO8d04+QkiH+f53FBxZu
Gz3nPLgUb40SmFfm4mRGcNYxK5JMhLmSp968mYp5zknyMKjYkvYFJ7CcZymxGnrK
9uMCrIR+HrFtVOX34M8e3xbLOGDqAaJTXIxCL+JZeegFBeCHACPha87ZbOrfun3O
TdwqA++gCL3AAZKF4+hLKGXaQeb5RHw7ETGGIVTR9bhMegyA4LUgeUiPZ/qMPFEN
WlMG3+BtNy0cER25E+rwp+i6SoWM8+4IbD7UVxynxFdhQItJ8yr0btcB4Gu4KE7Z
4mMmxmMS3BxPBM8ey87Wjiz+1M12oc6MzY0Sj0IquNDV9E+5FIn26otEtuSvDp4b
nc0mECSzsHfaDzDsUHguIbuO9T6qgNx3CLXrwypR6gh9Y1N/e0u/HMrGv1/EMLkf
pDGrVX5QzMYS6k+kuYunNAvQcKSWyKOl05vmaTuN52kRucziDg0iERtrySbcKc0B
Tfj3mSyPvjkvfFZ0NrY3SLNqi6PVvCpkVkuqaZ2955JR4sL7tqjbyp6KpwitYRuL
VAPOZub8SeFKMIGERPV6/f7CrdAZf6/cU/8Psy/PtG7ZNLAMHwP4dFG4Usk3kSnZ
xa9fZMCHTPBU+lTrOKxMnKvI/3rO5gQZBkP7M8D3mI5w8AG8Ie6N4OE4VwAsB4It
YfQx7hig0i93rFMNT9PxH1n/mpjJE5w8d0wXIjiYm492wzCOumYcRUP1a8a/t2LX
x537Z/DtwC2Y+Y9rRDm0VZEhHZbrt7QdpuHILE59JJxTfcIPrZfOtf84q+MZlrCc
umlZarN+FSCEr7+Ufg/EhdqFSI0qj06UUbpbGbOv3LLGjzYZI7ZL/IhoWDc+0CIi
PLyRsHt7F2IlOPGM3nlNEADRd1EjeQ1uQUpDp8WcXxx3DinKvG2iGgk/BHxgYiYD
w0JUzLK+GoCiGaexVuSwfSqMgu5zonpR/FtXKSqW9EW4qo0b7Oa8h4Yj1jRfEV5A
/i0aroNnQoCjvw2kWbgQWA8eBOyAQAdCe8wX8ywA1HM0q3OIOCC/Wqcwvps8sU0J
8qn/1kePFTOQ2RiP44WStFlO5OBVkHMMmoNzVx+hc26tIJrVt0aZKAS6WOtC8bcu
1lhVnARCYp7cMMnRkm7CE6hEswJ0+cBUTWuAnGDpN0AO5+t4+om0yrcGYfVm8JSc
ZWCScTip7hBvqfLW1YaEnJKPR6APe9wynmY53YA4B+bi2PkA4XsMxI1nYiWxojH6
g8Oy3BLV7iCI/ALu6NEMmY2nRO7Kyx2C9TZof5nD2yrhMa7za7ODmevdAiJpFUlx
m+UyOtR4p+Gs2qekgudRJt7A8uZsvS/9nw+1VjDIfHcI5dVD85sGlxU8Nrb3OCGA
Ao9yFvfKp6aBnbzbm6TlNHrggu6DqN7VojjzR2sIpL+4bTSYavjnQ80W60ySd4ep
wqxD1SBJxwcHjZbPpESSBxvPZk3IXsYCrl8ohtC3XPGGdjrcDTH4SQp1AtVxGUYG
Mdmd72lbsy/eEYeXoJH8JL7YEdWKzFdE3GIAsOPnRGPsAtBujzgTFGcT7TndP2xf
5cZfljRxracJv80cKYtrnWwRROIG1GExEfwS7shOBMmuhrnOZqtYgUVfXElkSShC
Eruagilqtu1GHv4f4eZY6VI22zaI00R/cwij/vwDu67iNAsKImktfq/BbgWzWuU7
bmd+cHMe2StScRYiwdAnaPz/oI8CAAqVnxrwHazrmh0DdTTXoa69OWJjxgu9AUlS
vzqjQWlgBbwGsX7yRcgiVaawp1+BCDICOnjPTa7GpTS0J9tSz8X1JmcZ5JWJRkHS
mYZRC1gSeYutN/RInSBAesLBXhBWWqDlqX3fuwjg2+9TAIg1ldS8cwxfDrJGho7h
2L8YlLpjMtdtGoNq8G+advcj22rpRz9iJzowt3iNMbFtz3u8kSHKCuDBefDGz2Iz
Xwbc0FKQHCE6lPhVdDAwaOEiYb17Xaw9+7E3+dcor+k27/4BwJgtPv7bnMx9eOLq
V21kVeikBdKs0IYYZyNQZmhuddqHcF85LTo1n14oleiOihA+4DYFBrq3+4V7G2xA
+KP1zW6MrNVWX2+9Ww4/NqjA9uvHw37vnaaT58g+Paj6S42RN7FZkYEoDP/eDC/6
8ZNx0983gsHF1D6sbW4pz2wN3WlIQjDp3I6Gkwgmnubj8Y7VuOwPGxAGElnEIeOR
+CImXAS8zVodOouUXobEIJR37hwycxtcVrTZJG9lZVGNbI3IizujyCWTbqndqnBf
GtOKbj0WhaL9J2rWhdOqRyJWWBFeiRE6GEk5GnAHZ0DIoAFZ55Fw6UEdfYikhWDz
qA3uydBWJC6c2AoqKG6hfGTyNlMhE/4NpswhbKBlfL1oVGenFaGymZ8tuUQh0/LD
z4gzRadXunN0sOzL66pPQr1yuS6Z8ZvqaCFve8Tm3A3SFjlOtbS2UCwEC+ncp3M0
5SwHn0rCgViQvusyO/7qbgIGE0ibc3YvmqKOaAwEjAyXncWoV54BfG0kIG02s49d
yRcAVeIjCJx/b1LtbLDDwdK2kl9XXfOLcVs0LN+oFO59TYQCKf79rzunphzd8mHu
ZeeenxqnCDB/Rtt/VWW1sRe6ddQ+IBGOxWgz9CRaj/3pmzt4aLy9em7wynWhtDBG
HqZa0HGp5ibltW2nXP4yRawejOeafEVpdpAXbriS7UsVwHfyccGDIBkenz6AkWyB
/YeqZ2bltNV4thrmQ6LNrvze2b5WenQ5pCmKpRe5PzftwSVJD6GNthF2SSKRjz1F
REU/kYvBNnrUWn8B/vD2Y1UDjkq+t08950f2ZTU/pgj5q+sKlf0KVVncio48rvb8
EAyRyC17VRt5XdX3dl/Us73TzgAyiyoUsHxI1rCU9svcBSR/ZdIrcWtap9kpgBE6
9YsxgN/4c4DMAVR3Ranvs+G2GN3v1Nf9gziRnWQF4+W/y26YEITV3XMaFyvKt82h
1VZ/Yw141qwpd74el1tE2PBXUGn+AIZp0kCUAuzFWFFbqK4FLTZzfc444u5hqwId
bCLTRkBfDhDlrdSy761cHOBj6BqXkkv1uKn1ombG24K1fdoRd1viGZe9X5Dq53kR
eSuhiQo20/SnjordjogUt/xAnmFaHvXTv0yrdRmYy+KXVY8hruHDtBR++NjeK0z6
1pHCzowONQfngoauLOcUk+NaAiMLVnW7uDdpDm8cpvZR9wKTgg37Sp8EGI8Ehf5e
7qjzOCooKEjPNkApWgjoh6zTmJyl8xkV8PaU9bqqtbqsEP3TM+LKk/v93cCr8qrp
H2SJ9M7zqBfUdHJ40xtCAXItEx6QggOxKSjWmqD6iqCZeFT2jmu7p4Rfw6ni1J5m
oqUUA3wOK4gY1MYAvN70C5vDMM2pNP3j+V1ER2ONkzhd2EFu/lbG28fFSEuLpdUB
f9eZ8Vu5ceNagLJfuEARXrOBSp9r63gT5SUkts2mR8S/v9YvntqG36MuWmXfx0T+
W6cZOKZ9gXuBUqUejSx3T4VUOy1n6sFu1pAloYf36pzBZOPJiI3mYMWfhxvHH3Xr
1LMQm08BjIRRIHgrApl7ydKJPrgJMYEJAS9IL6+FVpWQD3MsSiYvYjXEF8dA13un
yPNPiJRrirZfXHL563rSB4B4shl2/1WCuXRKb7C4FKeTc8sFgZAsWkd1n3VZK7OR
7C20AvBL30+DNNvGQPTKt4Tx4MKOAaJzZr3IjB+2RPGVQnmHjjZZcUHXI8qD0gX/
3YEgfN40t+F/EfF2E3pfbF5yi3pVfQBouIfpydqAXHOGeYv/HNzqEFxjHXzoxEZr
WJtD/Qtizuha1JORdg3SV7CKmMuVThr6g+K4dINCySWpZCzRqqUih5ETStTjjIOI
B2o/zwW6PkK8xRvLUR5VNpNKZf3S9NfVsuBUlVZfHqpIk6vAbrRruS4lSqWaC2tU
ZMK10QTY/P607i37rqQF9gEoCUJXKjQg5Itp1xspjLoTw+k9L7ccyqqhRJZCcAKO
kc6TMosM0q5opeDt+bfbLp2nur8/iI8MeYdcknLyfzYlWwQi589pwuuUZDYeNFhq
whxoWnSsdhD4p/3OFSaPzasqnSxpmkO8x//qcELYoNufwS1FfWtOxh9NFQWYYcsu
SSdgrF2Pjy9opbpkmQlv02jO1s7Lf5s99Ro1hCmI7k/Pc2zAgJT3s/p1WGK4Ifjl
6b4v6VpjZhD9RZQvWhLDljBDjwH6oWDI2wMI8zPz1RSavRVYVpagYdrWDqzyNd/S
CU+3miAUQ4atLFbla8RRDTUtE/ifrEBf5aN+WsK7pC0sxfVGrGcUDvX6jlujESQ/
C24UCTBbZ8v1XlQDJOukj9tJVMlSBNDtCg0JmnGFmLQ4TDjj/SDxdz2kYOqbecB9
iD2o97ReipTRwl6OAPkZhFMOJyV4aCnU2Ifgf9s8RXJ5mqhNeDNx+zYQMONP/gKQ
BYTsH0kZl+36aEGQl5VcDJj+mhKfNXtQ0v8xhnXcFOvLCpkys2zhdVQG+EwmKFY/
aze12fqFQOoW9pAKIyXiukunKMbRSRmLDesJT6XnH5/IS7TKMwUyMzjq/3wSYEA7
e9WP/mZQWnEP4MidfG/n4NPDTgFsoh2rchkwd+HXU1zpqsK2soiblrOli0TvSZOW
RE56J8BcLRMrNZHm5+vw87Er4R/qD9Y9hjGNkKIrVM2ojk1wuwwyj+Hn/Q3Ij+kf
JFEL+VkjniDTAWC0EiwGLTVxlA4d7dc9Ilypwlmq+vuNzVMS/ol7q3802RgLlkMx
hXrZfnej9jcfqpQnnuk+7puR9iLmgKz+bspSTjypJJszQjclB08rZUpDYMjYYWoz
9OfwL3aqNPZQz9qMiqoqRpYYU7uYff/hKM57B43V5WsA3XHkBpFg/gaKXxKkRnoM
I3krng0SE3fo8QZUANgtDN38U+E94yjlN6ctmcIoXfHrh2MLfR5SGjYxDvZFlubj
HX6VMwrmnGTv2VuuIkck/ulfgAIEpgl0GG6YsGIU2K70MM4XgmoqONufgpERcsfx
Q2GfxhjRo0uOnlXRoPPAzO3z4n5I9Mc1/paKitHZ71oeR4zbRikIaMKvesfCFnf7
aVopj+4LF+3OhGKBzUDH4ppmD13/iPmKrZpTen9gDgMav9ifA8U91HjQRaNFlpUW
YW4O+qY7yzl0l7HvUuZtZ8CJzPKrA8R5cgnqFnRl/XBEqjzRRFQ9vCmmdfMco7tU
88kEqSoR+MNTrWYfXAxNAifYBXG8plSoggrKMDm6QOa2nGYHH12fsJircbP1KskO
nNWM1ETfCTnXosd5v2fk/cLLdn2mSn7NVTmVIKD0s+W5KXyiNBAgvCB5z2R9p7nb
vuj+f51SYhwIVreUVFGZaV4kLp3aBusOs/rh9Q+bLujcfM+Xfog9rHuSsVgGNfRv
Iabwo78M4xVKd/ok5FB5vCTpQMh7xXbaJ/cmpTi2v8K4RmY2Z5n3GZEI6mwHTNzl
4rFjRwNI+Io9pC/i7sldtkq5h09vWfcv1w/b3TwjEab8aidlKqPGLYzKM6xPkx05
DxG0cdKrB9KIRSrOIUsYCAcM2w++Ch50cpxtuyYsXCR0879Ze+FwCGiBS4G3pob/
WepOxdVfr63mWnJFg9Ygle+rfS7Wa4b68D5+SFK7scrIi5JqhS5Uk6zosPO24YX2
J0koc1BI3VoGTSPkAW0mwFUqvXLGVx5lUCi7eKGotDq23pVoRAf55MHPI5zD8DpW
uEqVUnEHSolKc3iyHx29yu3DF8fIwplwPPoPduCYvdcIV628vdRZ68PssSC0IX0T
Ayg+ZypcEUACHnhVYV1nuyVXz9Iiq6Y3Gcx2bMlJgvjH5xQBWmoJipydwB6UYY8P
u/I0jUHzKT8mMn3cIeCWD9+eMZRmE6yG73dpSNDHZF0dhakdvFlZ38WH9XSsGaIN
fLkJMgf7mVgLYzTioRm2yea2fpHnoXntFQ1VaiY4uRWQFAWrNx1DBEAfBbzmYjjY
Bxh/fNQOnmJB61kRfN55af7dzLZXdbthyg4mrd6hRVNiNL+qD7yvhYWHAXWiuBc6
3LbwaPX0Yn8vgYG3IPeVkAdYRz2oO5T4rJ18qVnPb3GHpu6sIxn/VgTjYfOsGq6F
J4sjDBa6N+XhlpnlhAbxI5YXCDy47Vp1EBnuOgR10qiHq1NWb2kY3wzleDr2REJp
8BkkGyxQqNUh6u3IJhXZ07z+hHQnkoX6j258EbMmsE8zvrYBQEIFq5Lp9RhIGf/N
NlXrRv+JqiWQXXSVQbxLumfXU9AkR85W5kNX1Evu2Xdk5IuT02VPxsPnTvrEkhj2
YqBRY15TYBO/9e4zACfr1toHQxQJTOKskjIShcd8m9FC8AxS3aBNtQhbYIXS+b1K
Yv3oZZ+3vN6Au+m4VkXvpb+DB63qRLcoSx1GesIZGEIFREOsopaqckeHGofbxUUg
/BwX4sh40rPD/9/Eb3IOK2LQrPu0QN6n0kjRhFouWwBQRzkzx+MPruJuUHIo0HiR
cADfiWBSqKXitGVPcSidTLxhMI/F8xN6ghwR5DWDEICCMrNwtK8sQJU5yiYTlu7O
r3ocInCnebXt5WW1iV+qWxewhwLziILIJG2RLsrXfwsO2G46rJMks2+KtFwvWwVk
nEWFO2Zyy05Bp8EIawQrL9L77VA2GFtF4lbZMAkZke2LSCveSo7JiVUrH15C0fA7
BoMv14FEaHza24+3Dk4TCWRpGUrS1sqt+XteDIoCACTxgAy8wt0jf8++KqL/4aZc
+h1O7W7oGi367IYngySLMiIRdIngHjlmqXQk2tf2wLllCRbGlB940/cG/z0vVXnW
ppovH+02TRHlcryyBZOfWxKvPQcub2jWcW1YIUWrvs56WVFgXjnSQF+UUS7pHdWn
n3Fi0+NUOP2mN70Ny1PubRSIAs7IdCAgEoZEyEBN3TL78edkaK01r54qXh96dfjb
3tPphHSKIVig+K0ja62N6ZeKgouo2Sjx6QNUI8uQiqBS5wrMe9y5vy2zCeZMSYoz
atO05nxnYAYxEC8XvSjxT6gdk39EdGO2iCgCgh0GqqWE9fV2mbMz1tLeKA/UPBVI
3SzSxbPPCw0flSXVGVulIaWg+2Spzm2tzfkGFOsGlXY4HWWpOnygzaXPd1rXUTpm
xMP9W2Cma80nZc4/m+tfMRyia00yyFPwn6ZxxzswArZImLcnUyfJfqon7gjxVNvp
FgII0k6Y0lSaPOZ9IlggR5dVKtAM/vE8apT0v9mCYRZpV0bz/r6way4Nq9AknnGX
iruzHhVUANv8/elpcw03rvjWFfIaxlSdRMZvEGd6vfoIHxxDjRgcfIwXZlJn8ad7
hSMrUdYRwV4mac/AxC14YGHjcJVxdwDgvUd1m4NyVVLdeNaGhRI6hlFNUeJ6t8ku
+kyXO3fIiaDctvuUciSJFB9VgSlRMs1EpBBxrRqP4hVR7m/8uGHDMUc756/H/yCZ
xMZUvBn9K7LH3RpUEG0eLcbHu9RHKUjZUYxEj9Yyq2+yzextHPrfVE39o4KL5LTz
jDc+95AyssIaoTbPrf3BgnjXf0sWlO+7VPYrcbGF+AtXTT6zBBcQf6vGI+LWPobP
chqrEoRMMu3Ty7MJSioDO9VLzXlgRI0u8Equz+DbW5GEqvi3w3GVR5Q4f4OHItYs
ecmm5ExfLcOD/MC1qFaDLliI9Y1Yx43dZlzh0/PRLsyxLRgl1867jsmOjy+FK+6m
AR74TzZVzxVeKHf/OLSY5SZybINXKgCocY42sdd140BcFMASuBIbuWvaz4F5a28x
PDXrCaJY39mUQenLh2VD6iEtbp7QqW5p47I7+pP2NlXgvDT+/NrDbmZF/sBMakNH
0/9Gfppax3heikMyVPnDmGJFMpg4F5MIWbYJ2nx7zKU4Lno3H+3mMvmSzBpFa+54
HNgWmFmKyw8HonvmdZIOB2PqBuUrcFXV0bfeZeheJX8fqQ1W7GqF23Pd6KLPiN4O
tNZwjB42S/pWn20Rhjz+By8GBIRVib0rzQMVyPkXVGgqujMOltMfNfIJmbrMDbdF
CmQXl6jtQe8p4ShNHQ0BO9xOT2h4JCzw/0ZfMJlKaL/wdcybA9j3+E87J8ulQ1Ef
90GwBPgduIPvHxlt1rGx2rsrGt2HavUAJjmf9bN1f8rsPE30+j/hpKEP22YY7T8q
bE3LG401PrGYHy3GgdGjgxhT5zh115+mOnh8Mg25yPLsvDICsa0rpJyWj3ODgLOc
h8lbcSlKHPRJrDQk1VFL+2ekxV9jaeDs0itFLG07FWy/dF8D7vDubcXHffXlsxlO
0VgtLA0uT7Jrw9ajucgxdcv16T67oHVJGAFgqn15jreQc9VTqo4APfk8BYbdD+wM
TihPRuHXm42dnYxNA+FeDHsAiXzFS6wYIskkK4HgJ6Nwxabk63GBDrNSAg/WSbCX
qmGgKjPAAGj3LwvwB135bXTIPNmQC3/2MAMJ6Ixdo+RQx8mGmPXBGO9kwOSdhPhq
nOAlxqJVmcJluCrxRcw4xlnYDr5xq+zhaE8tfJF051OLfkASpQllsLppngqFDTqq
ViK5nW80VpBBtC9TZtrBP3mpx1i+IWRE9JztnSrkTLWzsp2L1bkGp18zlmhXp0Wc
l9MXNiYX+g7Bn9BKcSBShXBzQsCfc5vLLE5T98oMdsS4y7Uf5WjJfXXeJKW2eqdo
Opfrt0ZJgh68filJ03L0f3OtChPGxiLS16LqeGskJ1rT/QL9t4wmAqXkECweqTAl
R7RMO/yiRY6NMhZCikaJmV18c+uspYMUdugSE4iWv7mFvKITjVSw2p73+z3C3S04
TVH06edg5PaoPVM3VY+FyLLvpMIzcMwW8pBq++w+go4bz9g4a1ITp557IEPUhdQ3
OlRfXAu6DtQ7Sl9iB3CH7joXuLaj/WWRqP/Opiue5S7wF9HO4qzPRYge4jIbplmc
9LQ2m3PHXlzdn9suW+qaUcPkdPV0y+BZM26BukyBPgvGprCCskDtMiSJFjM0b1t0
NTlqSLMhLzxSb8yIE+nkwhAEUfgls/9vLKsymCj1QPGTg+vuY+FqjHxJ0we5ZKOJ
TLssbG+Wkg8p2/jq6/Mllf+C1Vi3OdbCy4C8sk4YLEXtj6Zu6TEsASl2gmM96/Pk
gcPVMvzk8HTCQjmhqAioMmHV/U+NOTtXqDRYKhJChSWtQa0jfNtaWr9erIXE+qO7
9eztbpKoXclvY8kE8ILvxBupQLY+R+lMOHHdK9y0ff1UjYCFtEGXNCT+eiRT/KqU
L42hnV1R+EQy66/EVz8rwugXGgpKeD4HjXWCJl10eyXoct0e6JGZBxjtNIxYeEnJ
hYpBQ4kRDuqrmmiRjzS44JzGANWfwtE6d4NDWI9efkHt8DxILsBXdwSHu16/PY4K
am69dTeHaaQB1fGjhnsSHAsOznPMseJcgqPrrEG17vC3PEY4FSGBajmHo960G6u0
LygXDIahH7jCOQ4Y6FUZ0e5ccyfFDmMDnKfF8dWzkT8ihmGR2JlTYW3vFc53Olxr
y+mdXtgwC1mKPxfL9fZCvg+mbskmFwEQK0neL04ycHOqB+D4ftXpoQDLDHqdSfxr
B4QGIccTEWc4CynlhxSL9UG6FpYsP8TkN/yGHroKuxoiVHxtkSD6MS1ND2H4Hlk5
1eeobMHt4oiRtyAzU7re3OwftrKbI9S0gkloKq+lhahjmSWlWXfp7w4RlvFqviL+
16uhyJsEKvRHeMJr7JU7XqG9fQSV6l9Qzrfw4lVPAIFyo+zDs9hzEae2dfyozR93
D/5el8+j/yttT7w0X/UctceRJLa7JkuaCJITaZWTc5O4hlQ/5ebdlFBgk5dU+LE1
koj2YlR/yf3P4VJQ7EfFsxXGLk6/Kxc+0ACPVA6hD2M2x+KonMNlKgPHooqdQrdt
oDhODTs4P6XWt4vF+2Ntjg1Qbx0HY3Wi8KKr/YtHJBdMnlBuX4P22sn6gkyZSnsW
Pz/DQ9ozTSzsdG6529PoLklzy62N6uMi/3hZtefYBzgh/CQMECn7L3CRB1eGGDHW
G9qjBNfw7OaIMCii91oZVns0vFGVJiCUIjQLyUEyKCwNrZXglEgo+/4GyI4T8lpw
D9iANAPY1k+jF98QI4Ah9fICu5tNPhI8ec7zhZN1hsx0/u3sIZsi3I0Or4gZz94x
BsBGGnfR1YufwySL8e0rrGcp9XESSNFjAhAy0MlT0bwiOwxzZy3LWyIZz4dQsfki
M6EEGG6hk/+e+oZO91bMMVTnnJFJSOBB1jaPI1U/0UgNWAOM0XiIr0YcMSQ4fMce
qOQgQ2+/w3Xw1T3OfEqCLwW9tucagxAGDY0KWNU/5eIiO4oY7bLf2TO2ScmoZ+RQ
IWfYk3sdEovgH3rp853MUGf/snluTOUJ4wYYPye9PRupzXhM6IW+DjFcQj9AjXow
TCEq3vjx+qjm3kr6vPE9v24iNrpCHYw8F8bwuh4opA0Tss17JNkL+e3T8KJhtxYI
1/aOLa9KiampQgNuxLr+l9rFnZ7AM0drawdUHEjUxJTCEuNIOAwU3a2RWh39ipFw
1sLeWgbeZZWpEoZ1RYHDWbx3ipBQDgCc8mWZKp+dSlFr4wpeLA845wOHB6OglXN5
ktZMiwLz4qkUjziD5PlA1wGYMlQONh0SpQbq9Vn6GqltiiYRAAtuyZY4F7z35/yB
HNF0Tug4RG7ySLJ4mHETR54V3xgBMXYMk+kRCkkewFWA8i2n9LN4XhQpVzPsjHg4
SslGbCKuPtVXS7OHqUeMTngnHPy6V9BM3xNHeQRMgLQHMFb+wulNC8JKpyYhzo+n
fpWD9CTxoossSvpUw8+JD93Gn8vbFXUhZHRUT0ROqGzWlxWH2LYw1Qx+l4oPtvGb
e2VYoHu4ojum0KGFkfVzGIy51MH4zCVOLpBmhIsgbKSOYc1LmZvvNpJSG5JG9fIc
Ibx+uEveTaBuo0eUcC2+tP1WffB985b5S3064bxOhdXlePu3HcYBl0uw42ZBZris
gvMjw9bx3MbXSv8ttFEKx0SvHqRpU+uKVMjgFCeFKaHEMBZUKoNvOTG9u1gz829j
y4rOM8pgQHj1OKFjgudlR6y3aZvePDFK+qqtZyECjp+rWp6v+XjotqrXfxX9NSAQ
PMuYqkxCtOzqYa4qEgc3PQwIy5FEXMsZ98vSU66EOXdJ9eOoD/hDKs+XOFh3y0SP
uLT6oby6YyAZtS0RmcXTaTwpCmnEZCDbOfQBm/+isZr9i74dwFKewT7ODzNJVOwm
691CqIhtdfuEZZ42SnJGp1W4JTateY7zF1M7bo1ZDAgpImUg7LhBH4YoK7CuQd4a
yevzTRdA99JLfrKvsCS7ZQeYxY7iuJg7Ef85i/JlMhOQH3Z2Y901xFhCuJs+nRDn
/27OpQJh6Pfw5z/6U30m3muHCvXhiLjxlLq7X+vPil8mDhxLXM9O8umR5Y5DaWwF
oKA8NzpzYXEcdkYdewt6QIwtz3RK9oOFZHIBGu38bMNnlJoPPDPiiaRyZ5nYx5Qz
pJvMMBCokFVzBp5WXwARdRos1c0eAJ5SeN/qJ7V5hQOESd16jQVzJGpZ4V2RMlnf
eb2eQEp0WqTJ1e17St6pUKQ75ZSAMFdt6/1g0l+KXhVjMU0W2bTI8qMWnWFnB1oz
KTZvjq7meWGLaekFHVVfVfqRx5++0azI9PM1/0ejF9Z1F6sq4oruaDDNZUJXGLXh
oM5pfjwy8ayF6B+4JNnZL5uoAOiqs5wgBhOMCqwgABnzrUrmrBbWQHPFFv/6nv2D
aqP/tEj+AEC+dKwepGzBKtZIHSDRDxckoxqYAhWbuDyTX8ClBdx3ME4gn4DUAp4j
ZkGF4TYE6fW2mohy3paGG2RpS9VUO7vYnyHgQQov8EQSSPd6XODseyVp5pjl/aWG
qz2dnBNpw5AFQsKFk4uKiRHM4D4JS+I4M39ZPfb+SJvM37Vn+qrOVw9QKvCn36Vn
9mGWsy9HGJZK9YYYKdLBlHSYGhG4q8kkuMRlwpNlBHCnOCvL5PhpGffnt5SFjQm2
PSv9rnOBmpOe4KDr+bn6rPGFFkyZMtfxxkoSW4Dv/vWm0IixKalw4IArcCpJzZXJ
7sB75pFRx/AVe3Rkh6Nh/62DLfKRChDpo+XSC6OqZPOKP5+TWaeYQCmttm/F6vTL
04abqbF/xTcuNGh/+QEKU2xGv5jw4gLdiOqDM5ONK6mvOQgjcQSk5hW8K6WOeIhH
FaefciNyLZipS6rb2zaJnHGXZcKBMk9MW/g0Ambf1k00SPvu1Ch7j+KmrZ9Ln/yy
Gz4hujux5IRMn2TvcrAHQ1OpTfaRIHepY5cy5AbYw/ps6i9hziWCoydIWP2ROSG1
WTy8Bb7Le2XhKhUu+UbVrjKveOknpbs+sx2BPOJ660yDfs0j0a6Z5BPNAf38/7Ln
nCIew+TWh+01jrrKBSgiNPU6TfExO5PQhojY1mzRatvLxezR29emILWp/ahrHn3D
Pq862GHSSxp1MjnrfjJeoRBI4HWKUwHBDNoo2FG5LAQjl1KVUpdSIxbElcPlmpSB
6svjBNyy29+FQerbKS6+r9GciwyRvTg4B7WTNNoijoXpL+nvKnqZJ/W5SHEu/V9H
0Mmab7H+3880OT/sdTxvxZYZpL1oUnI6LDg133PqOE/O6hQB0I+8jiGl1xMfUvnl
t7SkHbzk/ZRk8tPHxbW8vu/auB4ehL4OB6whAiJ7zONqteV2Wip5vYwrj04sVK7M
Ei/GDCLJNvGhF1P/Zk4TZGGQYfem1ZHd9KVPqd7fMR0BPHaEmyPdvl6lfZaMrnwi
GZrW/VUYzg8Kdn85sIPTD7U8lSRYck8ZjwEXamzgimGwdU4cNjs3qMDyIOEq6UuA
78jYaveRgLcnRrMR2XqTkKFWFZeodkqnGRau0QFgCCETWZL3Ln0jNBYL++iKfENx
UintKaTT60xD5gBGK/i/7hYWtutbY0HToBlodUB/nq91DMmmPD8xNavTQTBd7+xt
opAOlbBeHuJlmJpFM5Gc0BnttuJqbWCOuzk7IDSbM7zj83ZcjbTs2E6w4/GwH44y
j7ZoapQMcIPhgTugGHFYKdeDmU0qvijxap4wQgYkXNoyVB0WeQG/8EsL6bTqb2Tx
cKo/+fELh1SkjCVUJytplN+Y6CqARdMPBDERfeOFEKiwKCWId1HJuydYwDo8N//r
JFypyvWHXicXvRWCBlD8YCSkxx8UP7AscSLPbVHcw00hcooZkY/AqcMGZkDQWceq
hdNsb+LRF588Cf0GTAo23T7luwZiX6Uo3h7gjxY08eTLk/OK5vuWyam8eU9sBY/3
cH/dsL61VY4AnARGxEqTjEcR7MPkZtLrhQ35PjIoXeN0mhg5lV7dYlIK1RS0Jvib
14gPcel/Hn9sOcSEUzCrr8Y6WpoGrVtZB1wre1GPpJLVIJUeAUrRtvUtXpfjMQSC
0+0lpTeWe/TXIPkI/6Gu4REQK6SBB+O0unJMANZq8UvZ/EkEQzUAIXUT+ccSSBx6
sfgV0xD5ykBXs8FTU1tpoNYQ53lTkIBzEdq34CRhbpUGVouY1FGHJoRkyaOuiW7N
QbjrB2NG1BDiEZM2VbmhzxixRHwQC3O2SmbOHWEQmjtdLrFm2Gdz04yxw6IBqhzU
QQwDc8PS6oA4FSoNi5w998CRifn1kUlQXmu7BXwOEPdZPa0CaiB8O/LGK3ON/fy8
GgVaEjVl+zLLfqkNCTbp7pspEJ/xh3xZmgf5iNZsNHENtMvPnktuodaJIk08nyk/
hTI+oHmb9wU5gI/d383kQJ62pXNJvhmVFe5S/23wThphz9fEhWczHInkxbBMDtc+
trZ16sYkI6R/9tRfOKcTTfJh4Vjpdw3fL+/f3S9imhqLaRnYSWc3FG8mRykTH0eD
OaR7Texbi4MXA+Yygp46EObRAfP9qxOleHrXd3FWRQAJa6GYLCd/nWR/G12GaDNp
JxRKRGUyDt5Cn7UTXYJ6S23ozvLqwMWCRBbaEyZtpfyB/vSD7mHsIlD4kBDhZhqn
gTsYQh17otwZT3KVOrNAipgmjoqkEZ2ka7ilYHJEerR8kNdwxgm/bxOfaf+w5Fkq
cKcduA1R3SKvxraZcMNkBbhRyybuTDdHeFjxBbl0lgJtLaqOtYWfd56pj8mWNBLt
5lHTCEq/2BLXux0XfOkKMhGWPYXMHsIhWQ5btae0mnha3yudylMrR/Helvk01uyU
R/E/rQZBEKsgl6ofMP995s12FIJTUYqz4bSpxS+Y6CS/9NuU17chZZ0XlbkxnldW
iHTkpO9aXkP2LyEsqJYaOgM5xjGLmvCd/KAo93LA8UC73vHtTaOWBWL2eNa59QW6
lKSJrAgn8VGGhObSP//l8qiBZWOvvgxTk/bg4tS11hv8WpydGkE/ul0pYyS+2y/C
R5TMZGl+dF6jCy3SIjoqAoBBBkkm9A8/4F7HfS0Vjw1XU4xfW5eC/9vIFfGuEJbW
SiBpcrfEAWSSOAX6lwGOdIPH5AlU3qi6YkOp7pzALleL1mnrW55S4qlnITz7sYkq
XSz9W60u4Vb0tz722F7eURQWwJgNndazJKIV4GH4TeMqInf5XNBUK8y4n1CifTGm
mEfjQo4UBW+a7Iys5sR7zj5mYCDCB+X5RTTsyyGBjwTCLeeR/piyrGu4+zULos34
0F2Rp/a+VsfAoC83yooX2WT4t3gvB7g3MXGQSX3rW4LWjJF7BwADmjAWGtu8fWeL
mjwZw9oiGxpJ6Ng8AA2rJkM8b2ASiNxQwi9BcyaqHyCSxY4+pOyqYuacmRowSgS3
z14uWucJbXZDQhdXdMF23/DQQfuegTq/OrQfVuPJ+tcfra/NdOb6XDDcQXh3JTRt
LbC9njt8hRB8+H5Ev55ZrCXxUVRgL4A67VpU5dRy6BbO8VXUbzbU4ZvMt/1dSWUS
LQxS/HyHePskmGYFvYT5Wl8HEIy2DV2iVlEQyOtrMXSubZNvKOCrLI+6ZIKTQ6Tx
fyJWgZSiFv9CpR5zG/51/1SV/tWFDK6hhckaFFI+6uYHlMxtcReHf5ACi6umtWVH
qu9Q2VxZv6WfSJj9UIWdWBeINvYs2r7szjEh0h8V1ahmyvenHMQhdpetVQ8AWMER
94LVFAJpm59dHd0Yn5Gy/D3XcnvD5h25Axpj5n6W23WR8JnKpfNGG99w9EZRRfiK
Da3+a41nBLPNbQvszviyVdSb+0XTqEHOqT6U4VQZ5ZDLjYlXd+vY0sat1ziUMnok
MKlqyc1vTUGpfbSgHMczEFsa9TUEk9502gcUT8AaSbBRrfgWoo0HL0U09D8wLxWh
nTWeCxArXS68ocsuBJ88c0croKtmpPXP55hCKK77SLsURaC/0FX9AAQHoBp0Tm47
bZv0jtc9pheCdv3BoIhEh6LbdX8NRl8n3QRLQL1vo8BnaUMCMHbqeNVdh9HdfFHV
L/L34FdEQHqxOMAktkA3seAhceV85CP8VpCi8ICZ+KkH6xW56kbNwzY5ufD+4cvX
9wY/fzrkrUxAt6TegBvirMO9CEzVwcAQzPpNFMnHjxfO8QY+EOqNJqeOU3VxFnDR
kD1OKU0PMWJRWvkyeSjRngVCsGqtRxiHhkwHCPkRaPLy4y98cHsywzBtGMOjyEsw
CXnPTszXFdXbQMrtF3dSrjjc2bHkr5x4obDVh6dK8iCG87upTEkkzIaxTw7XZopk
VJF92r3QXDD7dHzZdzoUc5moCupQjyCJfBLQgvW9fRJBLCr04ZJx79S66KhSzVQJ
8S7RWMTDN9oWF0/WdPHJa6qgIEm9t+xZTLUY1M5zK9lsrxfKJAa6t/fC6A8tIshj
sPasG1FTypfFcbccZcyAqmfgIn8TJgshhuVpWLdNl+Me4j4KnrebNrRwgaO6Z0Ho
1PxoeveEiPM2i5naD2j4h78M/zAiHKzULxinclJgaIyhhv3JUlEQQ3lzaGZ4qKi0
tZvNZDbErQg787AYv7zHLMZEkJTLl8/2p5jcLH/duokVn6k4zee0P7aY3tVY9HAs
FcHi98Kd8dLecOmo1IFeYpUc9MTjZ1+ubDT1bw/KsS4FREeSvyad1Udd7Ol0YcT5
hT2LpiQowUIaPDu2sHZdjH91NpqXn0+8w817D+bsKNXrmLsfb1DbuHfcy7xepKAN
rZ2Q/Dpl+dO+QmFdloLQh+X4Fdwwt6Cd7hbbnNW0dI13jU5BFRfx7aDWxrdTsVJZ
sFxZsINmDL9lXvAfx9Byr7lDym7uliBgp+tCCYiGB6EU+s0X4RW9zkVMgYDT++nK
Sim776exJmxFcl/juLFtAIK6282gav+HX+nsrQxlMEpIBVZ1K9HEjGxjkKwkRAXY
rBNaZQGEwMhuZqOb1MygDnCohVS0UXQUgr9GtHVxMHHOz9iVyO9/Fp1rAOtENtTO
elCqATO0xpJmG+kFxEo3hS8de8qE3+u68NVdtXx30jtQ6pcjpBtUk0S3DW4SM94i
qS5wcJMUpCCHkN/Uit4iCsc82v+7pJEr41yuIpQ8VJ+jDb8k+x3QAyKPkIZ+uLDS
gxarKw18Hp1tuHs0q9KT8ngCWdKkmn2K4UckgdcoSjK5UBt3eJymoorZgICzmmHZ
79533IKuJTuxnTvtoS8EQ6FhvGjWFRTV313Bo1o6oDQGhrJHsVNqG408bMHalG5L
J/z9eJxsoBS2WZ45PN5rmk10mYAHWDjJD1eeZfNfT7lZpHholhpmF7MVrUJIZqBb
MKV0EmYxJkmjWzwNq4mDslxHHfYxrvo2Kv9vRQ5Vt/SEOlO2+C0WFlbmchW10ADq
`protect end_protected