`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
ddtXksX2+yylW5zu6QL2Lhnb2d1sD00763mmSITNX595NcHTEkwn0zB1Dry37fOW
FufOhVzEJp80NC5qZ/+F0Vk7Ik02dIR0elf3clrjeJRK85K4e3Hoo4xn7YbFUIms
l/8VZSb14+JVGURjfswrIyCUotIzlzVYZ6gzoZwDXIi5gQIBf/gI+KxNXPaKV+PQ
Ufys/12rjO6aI/pPlqSm0hCvftmBcnezN2hk1UeXgOIuKZnogjOsf0iJVX2aOOWE
6pD/psybjbnsNB6kH5uFTA5frkzIzkzl5d9+YDm9OyC+k84E83I/7/j+rk4L2dah
QJOvksSIzN867/4Qt8qYTQ==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="MvBXkzurAa5VTw+1JJ70nePUfoQXBvZOku/SMmg4TwQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
oRtzZL4VJ4iwysPsC8SXYCzXS8Fw2gtZTOskLcDV+1B9Nzn1zTyNtlo6lNICRmmK
ZRVu2BmCc2G+fmzynYlNTnSa7C0Cuel6FYpxCBlOuk3OF2tzAmLAuDyOH3Z1Yjzk
a0aHuoCdIRKv7BrZCdALt03JeUmXKPdOmIlkVGFl8yw=
`protect rights_digest_method = "sha256"
`protect end_toolblock="Jn9CQpRhJt4rnzZPRk+dOpzAubz7omckX1MrFd4p81o="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 9280 )
`protect data_block
gD6l00tciPUa6pDNTk/+t0OO0nC/UTtBwLB41d4inuAUA3i/ALrNyoJVcBnAmEQW
ptbcNp5fxEUJjnOxnedyZEuEBxWRieZFQnkRdF269oOY6ph5ZifxrqxScjDExJk/
QyC4366GIo3DwOFXNoiH0YU8bLHB30qn2vsrmnHvdnhVKuxTDXDAHoSYf+8QErf9
BnTao+9kqQbD0aVyPow6E4O48L7YgFhhqetd5FdBerlIjSyYQeL/HcmzvNGOGckB
5WWahEOFNymg+Pk73XDfzCSq4PERG0cTi6jTQZ55PkTljFtEGI9OZbXTMGgNKEGr
s6aX1McSx/ZI3G1MglwQmPjzUizo5Dp99bLzpqS2VfoCeumRuIRqjMWICZb8gt1G
OZrXdTvv6Frl76RwQtL9gEjJuXSd8YCYZp6CXHFSDdVLruaDgKWIDEInXqjlHnS2
9BWNnNk3g87061foz4Hhk35pk6LVGKxkWlaNPONGOF3hcUof2IuKw15zxfFUEjJo
tZpSrUTv3gYR4zOS6kuyuIlJYiRYu1mLfADNvfaonA7eAWk0AxtoS1eOBPoQPSY9
IZhFkRKx/b9ozQQZlvg1etDndrA/72Q6keYEVNgtc3bKQRM/rsLOKcgxB2RtfcrU
XEeG6YHXu8gCcvtJ8RyXqQ727zVklN2CjZt74j5PqBAihQWK+BdGHo+4r3JWJOXb
qgqlkrqfkS9uvQwVDuQVaqhxYY0FbPdZWzDZDpymmbSC7rCPrQPvJsXrSvXKamhT
MGYO6csHy8RYMv+B4M2OxtyWW6Y1JaR/tj270Ruxn3FZlCFGQIuVjD38njVFDCw2
ikk0UcjhUgn7iKdLVtcB5kGvqylzTg55B1tk4J/M89bUlWNqY1lEN6fEVq4IqSoO
bSBI12IVhrwei1fzxbBlBAkFlESVKtWbQItww8rE7RvNP92UktedfMKJzMCltO02
ER0aSi0/0GJj6MmV7BqE3HCgSja6lEH/NRJqm32IZi5vF3BQqzwWr3BJT1Atm8XE
2xZdMhfiSsmb+6ZJIo3Zdy3uQDwFdSVEaKLURmEZ66y1QVMAVyMH4EXLmYQOi6ZV
cPFNpqnCktvIX9CbRVUFdNnGXAC1hnZzyAvs/pdwoG1wMS4Hrtjy0k2Y9WGOAZOY
3xuo+s+pEaOHh1CMjxgtCIcJ4Udz34A5ybP4Fnqjjls5UlpB4RwKdGoGTR0Qt7Rk
Xrjh0qIl+EOVOxo5w9uriDgGBl67nGgrQ3cwBtRMh5Ri5Ih9tkzE9n+fbsaJuKsX
mOadOunuxwbmyC0nNkPjsPc+Kq5nAtESZuikiT/rCjNKib0aEiOX3caU0qmrnoGW
FyOGZTqg9lX9Lm0mx7b+E2FhzCq/KMOwCa4eg85copjz3cpbP5KhOtyJmYul67Dx
QxtjQWlPdECUclxH9gO9Hx06I/kaE1n89cgPrALD/olaBLN7ll+1zsdpO0FNJ+l5
+J4eRUWkk1QnQPoL+ntJPvg1s9q2czVXlJ1wkExxIbUvQMSvt6Q2W4RZluUYk41c
1mgESmloPGSKDtReES/j8Zl7N0G7PFvEhb2W7Kx8q/1lM/uRQYCiWeIHZ1HLrvN+
g9foCxAFGWo97wEqqGk9O7cdCvdI+wVjdP3GiLdMRYvGyNcPyizIsuLi5kusek90
2B5EGdSEtwS8TWDEX15P3EqleGv+SHphFp68wqXu3xaPe9rQqM5D/nog+LudxAni
rQY1TALu/p0TcpuTDvsp6AIJVnWyA9K8we/DMRIG5g0RK6cLKpfAFmD45tfdCDiT
INtURtKM4AEmZxeHo+fj4yMO8IJ72LV4tL8NsRhtcFxkbRIMigl9LelDSGt/fWD9
v0Yw/rTxWXoGeAWpEy3In9ndHksa4J1XgfAOeZNTrZGjbou7ZuPJDlc5nImViNHU
LKw8EWZWod1e0imtvhsVW/p3PjBZhVbQjYLb61Gyaa+x4JYvljO2g7Ipmr1qhsgO
TG8qa6rLRnDwMyFb5kCJqi3kXQVSyrmnrYlsBbIrxlfAnoQU8dSJ3urWnrMdffM9
00JZjXc8hG642tWO7Xu+mRI2UZxX8/YyAOGSLBQfBb1aHr7k66wRIuBk5XT1PBXI
udN+Oz5vS1TO+MxVuGbvnzc4kawneFpzRKMM4+geQnLbAxs9AqdwmOp7n2gsXUHK
CPP1i89NdwJ4ylQ9Qy8ElCQyPYs//vPuBV1eWOPKmdhqADErotxIq8CEaYBVsoPk
m/qTVp0Ai96yEgzTZjen2MoeLEIug1FkR6vmutu3Dx5DDU419L3TrFlNEtdlbSLp
J36oqTmOtFbnCJMi4rWSaWO+ZzR7yrPoHDIWzJ+p04DCENAl58u7OG4uq5UY2YaU
4Ar76UwG7qsnvp4hPDP+vt+QFUNIUUEh73nCVVdAY1DbKtHqDQADoFffavw9+V7Z
5ykJT1Vw55/zBeBwXaS8B9O0cDSKKJogxKwu5NiOUufw26jRjgB9/3vq2gYtfSKR
aosHuSgL9c1zWo/l1OhL1c/buIALzv4S6rG1O7wwsypQ3Ta7oty3bYsfeaFnbaTy
trj1aNazo8SmscUPdLFWA9eAcM27CsVKUAt/PpEOHRhMMJNNDbshEB5TEcl3I5HL
D2gn+KQ9n25r4lE24XTDKf9CjQPNBqo/PrKIz34I/h78ZBOoBi1rS6W9XbqyHc08
bqQoiFyZNC5CsSXAQ/PfIF7OzqIcylzdOXRBP6C5fYy2NR4JhznPEUVTPSwq4GPC
/ZzUYRxfXi7jGMEWRF7b8bYRC0A/CkAsPW/XyiQTcGOLMPplt5EUioUB6PdHDVym
9RgSjSDvDZPzlqhjzuweGg6lDkfOub1ctvOtFjTzc3zpzcP4M+CTdwpaDeNws3FV
yXJGJ1NPL8ylIznVv7U/lHZ8a6yu+7QG7rxTQv0M9y2+kEtOZcra14zG6Gcxgb6W
ru0KN2f4IvEGIZqZdCrEpaEfmI7h46Q90XRtW0Vjk8edvYcyLWJp3BP0sY2oLdly
pY4QjX1LX+mmZL+l10utAVp1LM/Rl6LeHUePe+0I6osKCSd+RUz5w8cKT6E8kjnP
IUO8emRLnNwTjaaI7SVPd5EAjQiHX1vfuNkUqzAgd3y+Mev10GDWYYC122mSw+5s
BD+vmZ954HLo5+gNssQe5lNgevmyGONrRNZxeoQs2yBYweuU3H5dkcIof3mLRiC5
enDjMn2A+oTU1WNMPoZ0p9flsBKpbX2qw30b4O9feJ26hJhldKUDDNa11wcpQgTZ
KGqblwKtxTWbd8VPuMhsHXlmXX4TSsSOiUr+rdaP62LxKewjgvCNDkKvLpEbgrju
b5vlQF6+WFYsoiMSbH0II+ahr3RvU762oR/3YNdGBrwkmmQfjMlKgJHmMGdCEryD
/30hwzEdmfTamFP4Mw2YU348K8Beg0ZrmNPc32bRH9gVgDkrse5J2NwxBAztTu49
/dDWTOBd8txm1ANdik6tqk17qbpqxYNJZ2TnjgCXWV8Op6uvUCsx8pHwxc/+E+0m
Olu48fEFvh+MTz5Zp/hJsDyJe4PrVmhdMhHY+PDtQk7zKIToDHcq4FNV1KnU6gXF
+QKs8OfSFPghphcaBMSW9pmvVoQDGqE8F6vuVzcdeKOHEVm2tJ56d8+vs22rgNbm
UyY26IjtcJJSpO+EuFznjHSbRRsl/71W+Jhs/NA9j5eUSN2E49Aq22OZbYxyhnL+
O8Z3sRf7OhsMpwbqgjg2et6WbRngh5lgoKKCdl3hrXrISZl/QQq979vi39wtaInr
N2exF4X72wfxsrEdFJQifyn6qf+CPMZRZj3td7gOxIkkX94/hkfvjJUH5awDxo6B
OJKrDzlx4JSyApFRi7jHqpWhCpKHH4ynBO4F9WG98eEE+8Y0PsW4KSZmniS2ZQLD
XHQhU5PUGPLjD3fJXAGxOt+2WcQAZObgWD+ubBahrPGMilNcqByX14drVToE5h1Z
Iy0t7tUSRzW5ZdeehP+vWPLIIKsum3T0+uCUUgL4TOBXhG3fd4U8q3sMrL7JaiXr
UBFdZ0d/fxSS2nvs9S5xvkp2llY+A+j0ry/IfuxyQGC49xQP7b6fkUaCPQsE+KAU
r6qYh/EaRUZaqopxsMTP26bGAjK2ZmJb9Izhs7GcNR+oFxHMHe/2y8kQbh/ia7gc
+1QEaA27J3KR+WGii6B5GuAE0gkOMkbib9+ETnXk57aFzYUaDIktBpEJXCn0FuqO
4H5gt5/y677LtgDudqliVadA3XABYPvHVhXuXjZU2F4vzkPEyQdgOsFZYVnRRkx8
BEF1pIHqu4EuzFSofG7n96mYt5FJh9wHnsgzcnu9ZC4L49JB0CVDl79FMEb9ZCxI
4HozXkQVzMi3Fh3LG9dOji6zZ4asU9KyfmTPUmZ9wzK+Y6WdlQQRcTe74/8IRGQu
h2B1JIJGTnJ93+QG2lYWu2sKh+mtosAcm+auHM9DuRt2mLgUAO9EUk0J8VW40GZq
4lXF0mWthFNRGQi0P0RE+Jqlyv/nvbQEFwdSYuwz9KsqiZzuxx4Zhb7sw1PoiD1U
7OX2bzTGGpNGFzLnTbKJ24KfncKaAR9Yn6/aHklMN6tfz0K0dzwbclIFqIkopPSN
RDlgwN+RtZS/tR+tDb26XRVpS929nglAbgmnWsnDb4fD8w2w6lEzmBdE7EBV8KPv
1a3jHxzPNKqr4nSUxrrQobVi2MLWc3PPJ6fHUTRdr9ZOLjVQyaq/7/53Ll0usU4s
/BIyUfk9aLFtB8EJguaa38mJqks2Fzqq1MlW8pFxEE0eXeS9EBpOtT1CYQzrJBhZ
No1YWeZCJbyRblpMRwVTY7Sx0P110bMljZOM7Wpm9mtLK6jH/VfK7wpVFjB6jKyE
ZgGvSyDHwvRPnvRiaO8XMnoZgIdx9nMQgHMMR3L2XTzJ0orPnAlgkvrnhwzqBs4i
Tws4bLjdtYz3TM2OmDYlks4fDbYjR7rCgWMRMl7ZkE2Tc+j+cS6KX1jPqHeknKt/
j4mINecPR155cjmI7Pzip2dBz8Z16kfL3DZ7fS6PY0YW7wweVzCFbxni7ODz5cEo
CdSHgSr694mPwbJf0jlYM3mqGOcqH2eTIbSiH1RQIi56v4tDG1BRZhFYq3PeQrMl
g7/Cs0ZitpnAObqdxqePg7CAJkCygobYbo5xccKDavJj0VrT1Y5bM1XVtuDmT7+B
B9kY0vn/c+J7L1DHuiyC6TEw4xsEcO8I1zLfCBkEVbRfdWa50yTgYN3Dg5vx6glX
by5kMpuZ961W4y/Nxf88rerhf5R/hwStJyqC43zZpo6xDwI0H6JQNqhaCOWD2uB9
s5hNkJtNX1Wlg0f5xqnP9AlG3KyiXguRCoAEnq4+dmssvq7hpp7QCWbGyB7g5YCw
5O7aoi0jYUbgXHZTNTGuBj0PbakGI+QHLMys9bf/9HeTq17qqBKJ+LYJ2/zqR/VK
rTbLi/7VJjObJGsVDrEFEgVU+01SP4MEFg1yRmS90IgTB7YqtWeIFhEajL+2aDHb
7VDdL0uIJVyxQ2yzwNfB4rotzovAOFHHBMkDJxNBXXaFDEzO8dh+0Gs/pIsaA4kj
zb64NkIbOtOZ/xuP/wshBSdb3W0+J6R48QpjSI8K/3o3iD1GQUqGV9GkOSAspRpV
wcw2xJhRFsS8y58mh09d6fURxE6HE/c8ZzyjXHIPNxTzksnGejcpr1ozV81ayKFe
sHYtlN44zyTwL8otggQ0XpfhO2ZX+gYiDDn41xEf8ygT2eyVFPtxwl+0UN2gjllU
VpJ7q2x0Xd1ZT6Cy11lsRv9g3XF+LKGjbjUoX//r6nMEO1chcadS2h1IVjhEsHqJ
6mjFpaKqtElDpBvM/PKSaGYHMn6VPFR6SRzwfHfuMTA0rwoXu2k/YirG/RJhS5r7
Udgu+CqjAPGmm8cQCfMnpNse9sYpAVYq7SeRMp1XmMZaxVeeHiCeFURLlFHOImMQ
A+i45gwIp653Lmh+w19Rr+R9lNA/wErbeFvk+D8BHr9P+OLUdKSnIVJ0ae4H+m1x
s5dJRwaWJFQXp8+KoYmbBsoLKXtS5he5/ufNjwUuNcZ6fwnqGgNYpyl+61KowNc0
42tqeGfQoKeU6WQmSRvJmAqavpnD1TJCH9jITP7w63phcttAA+80ID1TqNNTTq6g
mkRRxXIdZO59k1D0c+rXCg8TWwjEUSUzkpHEyUsZE0UZIlex+cOD5GenbFVn5q77
mRQtBjxbxsfXsig0y/Cg3VgB92tqNvxQ9MBVGi0tcO8sPGJfsKoMrEdoC/WzGgu0
5frdbV0xuZEGIvSDn4ol8xW/pNsSvOytQIWqpVkKB2xzXs8AE2pGBdbp2OzbMkY8
NlBin2SM5ciBJaJ4lIWl6mZWODuvjyzZJjUlQix1jPtMau7zPRNZ/Fxgkwv4roZ8
HuLxD0QducTjcrif7/zr9qFurdXoWP2YmBz6aYsIF/0FhA1rvH4QcNxrFeQ9nNrS
sZjHqq1mXkONhed2930sPc/F0/uVELNdIglXX9bETGu8C2DjFXpmqLXS37NUnOWF
rf4LzshJxS1pbSbJdnfYLAJYF8+Zg6qO5VNnF12aYptgJnSpYu0kuNgn8mGWjOgQ
FB+U8MhBZDR03Li+IGSKpc3GHA9NCc+8X9A/1Wfhai4nRrEdOWcJZr4bcjd95M+9
0lQ8/kvUut+GEf7R/svPVGtDS9rVWmdaTCxiy/01GaOUO3hSpB2FjSowUyg4UIkc
kEHV0YbabVArrwXkOS6ItipttBugr6AyXyClNe4e+kbzZmzXrNN1e/xi7InpIzRz
1Xo9aeNcWd0zy1MQ06sziSOqujhGzvzGC+NNZiTpKZOwgHiRJOEJdypPDNbCsCYi
Ujk+waDguIKAjSALY56J/wyfNdaUle5PnT9+WH6fMMA4n2gnMIsdTwb7mIvEuQpI
cNovueElXjsDHP2UsPutqsanVKJGMmu4/kWBfITvLJp/53t+NeRCtHFztPgCTTcT
+eg7D0yPNI5CV7crZSxWP8lQOoEP88mXNSVL4CwwCyE6yTonIdXlAlsY4BHZEq6h
srxMcd3x1XBQCuQXWuiDqUwEFjuGo9S1d8ekGqsKr/CXnuMf2qGatV8MyR+u0RaM
4xsTAiCGiHsiPreHD4HX8knn55NIzljPZzBqRv58eqyMFI5BL/tIPTqp2RR98LLQ
ZHbNunbeBG4gSKN9SnxIw6xHiMbwA/r8zEi6ADrBFJR54j/7ctfP4IHck3j3tE7E
oV3kYOBkUHTTMNgb+aI6JYJ75I6m5Ion0UaGhYeZnOyFnV90DWs6FzCvn6Y68KYA
Xg28cOGQjcVCVBYotr2BIe5lCmNUdMFaaxf4qB1L8iTVWOd3Hi9C6OVdq0QaDqzf
KW91DVR6ds6xhHNsLWVZxrH5Ki/89bOtE2QOSLnLRwxQPNBMeFbQVeILlfhsI2gl
9/9k/rzgfNaowo/pi+IFZ6ZgTdtCLIwMKHZ4jBOJpL+4XzkpjDv5VjUyL2iqkx47
AhCMRjXU4g48Tx2T/r5Z/c3k0HUCe1hGoJWS18uq9NAfDpIGuoBhFIm6w2hQbpZy
G4n86VfhtuMhlhpxz6CmJQETendq1WEwpllkXtdxcV8XD52hTvPK7AV+YX2ApOIr
2dH+dIAxL8a4R0tdvVkNZYxfQyusa4WSN3/dmENrGEqDQQIet8F4oQzV46Q32be4
psrkbBR29QZBhICIk4uGwZT/DwBHPvdmf+O2Pq/KXUICrgwOLuy4N+ypLh5huPdG
WlRyrOI72d9L0j7h0m0zJAVPAhbTtKdUmneFZyEw2gcUl5LTVkruH2doObxGCZFp
HW1c2QwRufBAyxUg6gLrY6MaChLAxhSHM4oql3IEf1n4lE41O2j75uXV0BtcROaK
cV2/zNcrDl3ulYYxHMIH5cx0OI8AM9NOhH2vNcfUJADN+ZXd/hRwMaGHvH0gIypw
YM3xuouEzqzmjKK04QUFOdXbvm0A3xP5AscVEYvn+IutKrS+E9gu4pkXmJAGH7QJ
hYXW9lBWcK934uaUZrxJsf5B4t4bwSEBSLklr8RYOGSssa6d+mlHUkjeyGfI5qnz
6dozAm+dqFaICt5Yas6ZTVtqvASt5N9sPAaShnI5u/Ak89mXVhM8pgozXjK0/cQH
bxi5vWKzctzohPSUcMT27jBp+FHkBapZrS1efgpMCx8pI9/7XJa/Vrow66WEMgB1
B3hXyLQqG0LnrYI2UGvmIcWjtX/s+6KmqisJtoB6L2lrcrjDxpZA5Nua8LREthuT
HyBBZbBHe0WFVzbll4whzVwYpQ15mI+g+pFpg4fDOUWZxtangSCeRYlSK2dBfhZc
UT5cujFhRPMVeJ5IvHhLMpm7ToSSajkrw3BjkqCzQ0lvKDc8Y9EaJlKYQxd8sD3a
oh3I+JAFToflw7h85mYo2j+1dwqsCYcTGSGn4fTOj4KqRdARmyFtqmM00Z4Jn1wQ
HMJxCyygwweJ3UjW0Ky3HJeOxiT8IdYs+uf+DlRITX8Q+MvDJR/JHrGgly64d0Z8
5dxVVW9uUKRLnzbMV36pronxzjD4trt9BvskMLsUshv1W9mI7LzmhKSccGugY5FK
ZmZf95zjTdVXhD0s3qXalEdWeXgyUIBI7EILHXe8CyYdtI0cCLQ1npwipR9mLul0
IR1J+fZ1Pdi73CA8RZVv/yNrDC/Wg9KdP+gFE+0f1C64+AjR9CmsoPcpLIq5r+36
PiF/KirtlrUwgIG27O0yPNUXCwSmjKM+YXG/r8ctnh0/SsvB+Fo4THXnVH0NAwU5
IQ+CQW6bOC7lttVEogM4NUj2bhtxc9fmwUsF+cQ+ZRcorsz4wJVEFXMWkwkNgsFn
IWO3IW3L/90x5AnQ3RPB5XOM8TpvIJLRntq1gFRpO6DV9p6ZKv0nD0g8HP5RpsZY
hLbGMUKubmVbb778uLhSZxaqIlmJOZVBAMeNzGFjwXgENISJwF8i39JkdKSI6q+x
cyJWWVL+iNJOYV+021K/hnSI4EMP+rzpPsHtrORWxqnffOFQVqTfFgy0UzD67Vl6
z+giQsnKfA5cmLeooubJ4vHe1y9m3A7E3hzGQ44sYvV3ZO54NDS3OSkSmk9iTGFp
ilPDhz0OG7UX/IXNsl86+RxktNGzCDF7jvk4AVfwtOhwYIB39Z/Zrm2jKq7N1dKD
cCG8dBq7iwVCMExEWBV77T0TMSHSl+7WBXohYKzpS6EXhIe/fg6Xhk7SLCx1dlUd
sQjdaaDfsqmxnqzLMciw2QSZfOn09DBsDDtT9jKs+mlb3uurBULeBv1G8TDhlnN5
iSxZc6hHTY5ajikxzdRv52fIyYTZ3txY4I6pLVoJu9tvFUNpD9JiTo5JRxWP6aVv
oJTHQcyl7HqqnlNQ70YtoH3Vyl2EDq1PupCsg/N15f+McUXWHVk8DIPdpRH+CZdw
pJzrGDlvOeAfD+5u85EsiTm5HEet+bY38Rl6MdpXw0II7l/YmdKdxg3Pc8R6gxrU
/lzgr3U/hpmlIqJpVPxho07nMr/xaaNTzBknaQe790zMp1Xq7Oai22PXqU3UBNDP
WiJ/bQV3XP5+raIPB7mlhafPPZ5x1ji2A8/k8jWKmqmXC4wcd7HEYIvF7DyAWTJB
nL9qIFVD9GCRnabxkZNu5K1MkQxpuNsIKeucJcz81nj5+AnIJGcpeGgzhCTmYcm5
/0ealWWyrpR1u8SHPuTgHLH/NnoHQhL4wa2dzADphBEgwgX6HWfcUWE2+waeqtPq
hKfhuzkoBCQqRFIEnSX+wixqMkUtGUNvj31e6gpxrPlxiCThL876mDk5D4ROZMeN
NKgp+r2iIOBL9y/7elaJs/n9VkIl+x435MsV+v2QI4oDQPfFi8yIB91ePo1tqih6
ugZk11s37inEGrN5N10ojjlp3VRTTpkHlUrsXs6JpVoJWl+Y5xfUNUSyYVvCr+gU
ZrRvPhJ2/l03y78bMxkVyKLUsvOHFjwSmF94F1t63Yzj4lVvNjWRdXSvD93E832d
Szsid0E+OvYL9DVVQqDilTpu9YB3jrDQcqT61293V32RTYlZCMYQnj+vfVqwGNdM
Q9ZSgnH+N7O+/ke+BYQKq431PFry/j/jC83M9uuW6rhM7r8S49lZGqRlLTXJKTuP
jLvAS8QhlguR0o88tt8hxFKytx15/aR4xLxMIyEZwBJUxJwn4NTkqgP4itiUUOhw
hsGeMnF5rYbOe9O3az7Rs8A0trH182Grynw4kzm5oesW8FcXXwGuigOqj1fJpjxv
Q+ZDOJloF4v2XPOkNmFB/pUwrgKyvrMfpu/v4HzDf6iBMAREs+HRXHscrbBaexyp
UoOViYhWk9I+Dk88bucTIM97ycQIvaAnhxUHS4URRdR5+a//W3eYWNqG+NrEIBQZ
ILUX2zfz7lqKNGZifqc06otTGzQLKj/4O6q9OeGYxugpo7OdRaDG49/ZtZf5r4r5
ZnrsWCyeqB9cmooitVYmTNYwPt7+fg5pppd1XkuBkmJZugSKOB4uzrKhbKREM2df
5eVPassFFwjry6lTyMk2nhw1eWBffI3e1dMJqPN/uxFwTs4L9qgyfjTM3n93H1fL
18GImaIC/9xZSQMppzb9H8JqUfKQBg1Mg/Y99jmSY17v4s6aSMfI9Jgwi0Ff8dSO
K1MT66vt0D9m0iemqQN7F8M1x21flNB5M7ig0+Cg/4MxRKFdCFdK4PyD8yF5Nglz
G64M4hLuCbBFTa6khqewWVE9M2HmbMZ1/Jg+0UOF3QLuo0sdy9HZEl9IUxe9qtqr
8hNNSG/VwpMhsdYuP0xiKzoGoDm8DRTk1N1n0dP1U60+zYc/vcso4VY5p5Au0jMg
t5nMKMfi6cgxMi++674pRO0kWBBqC5StdWp0HCzE1sZjAeolwONa+hYnzJ17cLO9
2JOjJHQrlLGo+iL0ZoFKSY7+M4HJn0vmQzrf6ywX/+ZRKNSfCh46iOrHETTqfAu4
TzmQQrF5wvKHk7apndcc+NQs47WUxWI913ISeFskYpeggENNalV5bB5OHORqzpWH
hKmlkgbwwl25OIFptGvRzCBeLdtsElIx7sRnLFpl1lqcPMEP5Lv356x5Zs8t9S6l
WfVoTbyfLTwWpjfyEufS0Rq/CpQd2yq3THAF9nX4uVn80XXvgACoscX7qWUKelM9
MElfcjc40eP9uL55/KwjgSNP7EfhYlj2sBZ7cEwsuRz3e/Ngu4XV0cyyn7RFRso4
51+8MLLXbPW4H3tZNZHl4rwMHWCwGR+MYPsFtEK3ccv7N7PANQ+dwPzhz80YXswm
ygQbKpuB/DCMhrWgbB4lkE15KzqxutTWVpIxbUzfx8tB5B0HZAsMGduHd29I9YJ+
IXVsvPHjXZ2Qi3QI+4199PnMLEkm6GeTKYAi9X0k0ZPlKqpZz2zIsoQHBm4N8z7B
HcATzVB96qkUuh/f9v2rRp1AuJvP21isKaZVQ7ezJKwRlQLPPRQGocpB0m8+jO2v
Cn+B5wMsQ4H0xISsbP5L++V4grzGY1aqYe2YgAZuZVezZsl6PyOTzIe8UBPeTMcM
+qeUrp7Su5uQLskl7nFAA99mh9s21Na+3AwH9Y0Q75qC5meJ7NhqxXtHP3ZHdWPj
EgoU+rjzV2ZSVhjDPeXiOkdkWCU+PIJpGOFYbDtT5XmxHWLprf59BE781q4HJU7u
j4ixF3CKNjWlbtDK4QHHt0rNg5o9QhoE7MrZKuAgbTpLZWxTWNmLNsF9EgVxD6Lc
NzTHMuvZRNJSVYDopNiQw52gHdXZB1nV19w0+ZxIRHyOECDYx2VWTWUjuSMVUw9a
JpS9IpYAmWvDmLJCxXbFRwLhEVxUM2xnfFUdhpUTRg3Jvv092EZIS9qPORHhHxbG
HDwFIwd3kKF4v3/U2u5x42PJ7Un6Kf7JWFaKB+ICejrjKIttU1YuNSiPms5ZSBW/
fEikU8DsW5XDP3VhWul/isnpJG03Ny8Ij7hKpxokFWqQbxiIUStSTUeR/ZtQQZFI
cgTQ7giQlPLUtgIQODmTuGY5WhWL6rRXHJuteKUeR7tpjL6VTDUj5vQQKCylp007
5rF2OG5mVDFmkNhMZ0GpAA6RJBZM2R+L/RjFGhTPZfC56PS2RXfFIzX9pfELjg/7
3JAF4xRWZQ7XckC5UD05Q9Dge4QDwliWGVrtUuXBblV2wbqI7AnPDKLuwqZhSORU
gDKNTqHaO+M31j58dxicbujyS+5EOzo+XKeQruxRnsJ3My71K9nsdyH3FttVacIL
t9z5szQsBt5+gQHXWnL5wDPXkXP0R5gzHDdni2ALs2kfnFsYF5QMfn9ZZe3LOjf+
phpz4JzdOVZKmEzMZj7+IM6rTsKQcx6ZN8A6j5LBMB5TZBbTeWDOJLoFw4mBchBs
bM6rd/PvbSgaG/x6Sfv2mw==
`protect end_protected