`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
ddtXksX2+yylW5zu6QL2Lhnb2d1sD00763mmSITNX595NcHTEkwn0zB1Dry37fOW
FufOhVzEJp80NC5qZ/+F0Vk7Ik02dIR0elf3clrjeJRK85K4e3Hoo4xn7YbFUIms
l/8VZSb14+JVGURjfswrIyCUotIzlzVYZ6gzoZwDXIi5gQIBf/gI+KxNXPaKV+PQ
Ufys/12rjO6aI/pPlqSm0hCvftmBcnezN2hk1UeXgOIuKZnogjOsf0iJVX2aOOWE
6pD/psybjbnsNB6kH5uFTA5frkzIzkzl5d9+YDm9OyC+k84E83I/7/j+rk4L2dah
QJOvksSIzN867/4Qt8qYTQ==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="MvBXkzurAa5VTw+1JJ70nePUfoQXBvZOku/SMmg4TwQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
oRtzZL4VJ4iwysPsC8SXYCzXS8Fw2gtZTOskLcDV+1B9Nzn1zTyNtlo6lNICRmmK
ZRVu2BmCc2G+fmzynYlNTnSa7C0Cuel6FYpxCBlOuk3OF2tzAmLAuDyOH3Z1Yjzk
a0aHuoCdIRKv7BrZCdALt03JeUmXKPdOmIlkVGFl8yw=
`protect rights_digest_method = "sha256"
`protect end_toolblock="Jn9CQpRhJt4rnzZPRk+dOpzAubz7omckX1MrFd4p81o="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 17408 )
`protect data_block
gD6l00tciPUa6pDNTk/+t0OO0nC/UTtBwLB41d4inuAUA3i/ALrNyoJVcBnAmEQW
ptbcNp5fxEUJjnOxnedyZEuEBxWRieZFQnkRdF269oMhoRlLmoHbyuUVhBmNMtd/
BaoestqHP7RYce9HODGkmeQWqja5zRv9TVt+9BWYIKeioGq+2p/HqhI6+GlZNz3H
50ZDYBmTWhcQ5U41V/uCjNzkxbmiR9WiDltKi64nQ83BjYRFKlSkQ9t+bgeGkWdw
ma4453gSH7xcb+dvF5cKvv154OY3taHnJVNeBVmmPX2/hZaIoxUbYO8/P8H8jfiE
EbatF+EJFyZ6DCjmDXNPCT9j3+9bAAYVtode/HjSt5pJ+gskxRe5aneO2yuNzCZF
F+Z7bWTEG9OBqlYxJzD6a73GwiU72xhORPjaJlTntJfakuHDVLF0bO8X48h0LonB
c/BW5pA7BNtNkIlQ/kqWcEow0bTB+Perdm9ChcZHEusrt9RgPk3FVbSHfHR3Rej/
mgxZ5nVAxKKry/SNlpTNqgHTK1CtFueP/dvxUHtX+frgra2uaKXhZZqbfIgELIQi
lc+mrmcCSN53mBtukvoVV2xN7BI2X9rK7RWH7war0hIhAtkxxEga6rKhHkr9Qbpz
VQH6itw8e2G77sYeFYxNbSbJ/j6ds/UKHKQBSGEl/LJsQDl63p8Pqglp3tVfZZ7M
Pw1K/Qe2iDr1SDgS7VFljEmaGfrUpLo/7uELY03fg9h4oSGrJCEQyvf5xkMaOn0Q
L/nRCQbVdut+qeH1iVAaIyEo44f2GXNh/0hwomlFdpZ+Xso8Pd2vw/tuGpwFwqGp
c08jOTszh06V8z1rdrJGBZMrKrqqALJNqCBF+D2cHKjM0DbCHoWFlz6HTRuEOVDS
go/T3Po/c1GGUrA9gnUIgpGz9LZOA0C+eSQaYJ95Wrj9FYEywx5Ch8M8MjamcWfI
q3QoYj93DV3y1EOXWDdpNYzgYUEFrtC8+rn1BDe84KjOqXvSHh5Wc/fbKUIV/olx
8NZR6Wlrcf0bgjAIwbARoslU9lijDCY9soTVeKOdrmx98urgQQa1tfW5/sGn5s4J
/YbymPPsS3ZbdHj8cAZ1Ya8GPyuYobolpLFhkJvoWte5TMLY1NGUHqvVZpoHbTDs
aUsXkZfzzhT8SKCCkhGmAmY+TGiHmmeaYVsEDVosSNJKhao2s7EARkVBdGd1x6Eg
Xl0R+mJuSue+la3i6HHF5SVA7l0V51DCY1SEmFj2+0wEPCRgdjxvjTzdyqpRDaYr
mEWAzXYQJHJEOusqz4zZTH6Cibr7ru19hfBqkDAM8N9vafrlk5VUid0Mt55Fhua8
rOvWwk0pebTPvxdImhse+pS1TvWsB2cSv1ETIzmaDN18vzcariVLJvovZ0hegxD1
enio/tOrzdh5klqXnUkiDftqEvf3S+xnlY63UUOMQINUO6Gz0J3GtQVKtJB9sbjZ
NsIsG9eQlUe2HEjs/TGyALgN5XBGqP+h0F9S9e00/2kBtmj+c+A5bp1EvebPMTUD
7M2j21evZne3vFsr0quBiAukJVlnIoxknl3v1AnL4iKdhPuyQAaISh4ivWr5H7wL
FIuBwYK/TkaB1WOULk4tf/UQuExytQA3Q9lTh3D+ZmIMl3f36ixCTw4/ZzgxST28
Bb9PGJM0PfdYNkNIs2Yu7I5DijX3+mBYxRg31CyjWldBlUgQnzdivWgX9f/m2TjD
W7MvnK72D+0pcRpe8M0XCmgHjoq3mkg85ymj3zNzggDfa81agNZraMIXVLeietw0
9tyHpLgsRIpmYO4xETip1W+v/+tJZtJH/Xm9exl78oiXCD1HWZU16X12g1UFfuN2
iOgKKxdajSnMUZlqSmPuHTdGqO8sRnzd8GhwHur3ZJ26umEEgiBOl9OUs0VjJfen
QvMDv31P/WTaa9EcXtqg5CXfx/K7ZxZy/YUDNjadC0oWj2PxTjE3kebSHTeDARF2
oqt8XnzMu/kSQvAFTUT30T+Jtur/1tO8IqZDqfHa+b/qP8sufeOVIlWPQpSJ8+0S
tNX7phUM8EPb1cSqOAL6/LHDcj0X50+ASvbjjQ8fKwaGiUMAk/MfyWtK/cO9lxlc
5TfOKtl6l1XSmbiH+YXHtQviBogsw76ZNvjq9wAAeEIyFpjvIn2s3FUP+8phYW5E
6I6XfK5QsDdFmb2VhMvj/F2JGmpa5sbiiJJf4npLbU3dExHuD56GmORW/RxUyhdq
S+4ZpjR1upEVLzB6ebTCVjmDSUsiQyCSktslAnpeo8CdIlUGG7f4m0nnA3GVy85v
N/FDf2uXkOc/4UouBpJ6JSRyMqrVPlMErPZ2KzW6C2FHS5KeJybJCr9xwf99xl2j
CHtbW8v/Eb6pHhdDgMd6R9l2fvmCRw28YfNYICXy/sHJ5FVqtHmJZSiHdZ90cBt0
tWQkZx8asl1OsLc+9SADMqtYrEKVHsUkNHpOsrGyJyvUZZGlBRJMQmGBOP7MFf1W
TXfXw+rIjkJnnOLnpo1CvZkiOF0QWkmJZELU/fjtqTJLl/u/n2swJOgzyO7mI8Zw
OCVfsM7yhp4Xhzk9yjDtHbUlOQniaI5SW05hdt5smPCT66Ois8DwYpOer9ud/UFS
wQ0J3o9VVeRtKr5YTnrtOxbGnbbFGDgZnsGwcZZ+r1Zkf6e34f1mWNKAeyur7F7b
HcqClRRPBT/uxJvkGJDO+2K/Ps165riZpDgK8IJGBQqwElXf2wxGXQ6VZmu62DQG
c1A2ZLKnVHO3ZPJv7cqrphP/mmMMsXbf3COcCJAeXHdwkEz3SozWDKaJk88Co/79
HUG4hIBq8foNW227CecTTngenFx+m6D751VpOhcZ6Ruk0zu0cbzN8tw9qMNMQql4
Mrnn5IJJHzGW5kstTEFGwzmKe7qneLn3YTK/PE6pq7ep0nTS8x5v4FlmfzanpFBd
dSayv2BGuo8Ts7ZnuAYjKtgfDs+KqEszUXtUYsIrLrtIcL88cefp06eBIXs1rYtS
Ruf711LgUGd6s0Qy7vM1fK2/1ZWr1P6aIdSVlvFAnkn6Cuu+WKf8WbcJ+ccZLagF
qe7rCx0Xo+Vrh6mb+O3disxeUVRLFP0w5ilMBs1bOoBLmQPfVSr8LL+bHCNefs0w
sRjuFHIf7jHxNw3i0BY9B69I6CiQY13xTuX7uJlIF0kPaTIhY3HIDszOxCA4Ea/W
Wfsj1m1sHEvI0chZ0LC93he3nZA1NdOipwdX3jA3QGpsrZqTG81jkZH3t8tkokF0
wgX0NxKwwNmy4reIRY3fj7YCxyhiDsysAQM/5BdLJhWhqv4Ok8qpWQTCthpE+Ko4
Xs6//Gey+KgXgZJBY4MmvHBT8xCVXz+unHHf0hC3eRfBSi//i6Rq3WDHRKsxjEBH
DSGdNMvNtxuzLPKhwBAXNKNi4cxgOB0ca6LM62Y96A+kTDhMcerJ7qAEOyUB+zeg
Z1598Ch8jwtkGYIAV/HNVgN+n1F/ETOblZMBHC9joOqCLegns0iNzPDHFqPoh0l5
ZtDEu7TYeTw6S9DA89LCgJT9hajgweYuLnF2mNVF00KqyY6z+uWY2o4e+2TCof7d
XtVMy+ZzpHiQIlKrhctfdQoXFjD/WtcuKGCp17WHHa8I960XHo3QCFnUtF3n/piG
FyuizMXEOCzKLYuEN4sulZnAa8Ld1CRu3mihI3wT9uQH74IHzfOMVXK2wtdAeIRQ
HR50DozGIAbfZxtFGUNBFBVtpK8q6P8UEzP142dwR7W6sPABacPwN9dfbyRXlAuN
UqzW5uclfIM0ra4kTimkLb/STIyIF0Nm39cvimLJzFqFPUoXn+XVcZQwP0b4dXXR
/9zalzu9GL9ediObvvqY+DYONJll3WnNvHhdmXfQiP3JmDEXEwlbWvU8MQM/AHuB
Ezb2DpLFHi00swHb00ced18ez1ISWqRXcJ0nGzM/yOys44N3T34NyoGRXNCiKvto
23EyHfv78vDUDOyU0wbG0n+Rt4dN+ICOgruHjISyqox6QzhYr6zETwMz8oqCkDn2
+N4N9e8C59xFReBuFb/q5HzIGVU433S1Mj0TOPEnjVMVFjocEHQaK4uqB1acEQJi
NUJQidTXjiSau2ImnkXXvvoud7hCAK0ME1e95A9Nczu9SLmEvccJ1xmiXIcMQuUZ
f9JEirg9NiA/DjaBoxoljT+mxS5XKKfqMG9rTFqxM5FF3Q0idyGzDoBVBiRdBqnF
ZqDPl1HOqkh+zY0tu3aSmgVQwlvheEELLZkZEE6wOsgj2DeG+aZgE8QYVdewD2Jr
JDIdxbTUE79A5jfCeSRM5sV473cmsqsvip0/Rw7fJEwRORsHcadZ1TbqfZUi8d06
/zAqZfitFaSGsNBm8Btqla1wDaAIeLOFlrs/GQV3IjRUQma8W7BNzej/ARG976oQ
AEc/Ye8XXDu/TK1gBBoPGQMtWyqLKd/09wynBfSTVUnsRh3YPn4wQoKUuRtuXqh/
aOcNi7jhz5xdiiApYOO5z8r88l1r2GyljxobPFTx4cLCRM849mFa305BQpQ5Mu3r
6coAMA2coZLEUUb75AqhSWJ593x1OfkGV8Lk2/y852CKC0ZFAC7Uw3uI6g3H8dZT
QFIc9cuAWfk0+Nz9OEuzKOBwtLNL7gscmY+vfpQPL2MO1B1NeFSPhHMxvWpNm/xI
WLYauD6zTIYZAXJbe70cBfkEp62z/fnoh4Z+W3QzRXdJ/n1JFT7Gz3OvYImhlnJt
yvHP/WqLFq84mCPgWoIF4wG6SISf63MOzxhGymhimwD7etlRp9q3sIZov8SEFNm8
ivTXIjLqvA4fxACvhz3s4+fRXf0l5veDU5MBLgAlLAMRW67mxaRrVIk7iY21RdgP
/K2yRRm4KUV49Zeo1FkkQsXzlGsqV+Rnvx+DZ3rniKJd/tL6q5vFb7mxDvpen2LC
uyu5yxCsbKwaT4ewONZcbVmdALodaXktE7TfNcWEmd/LhtXISGvJAc376aH5XKOq
KlGEffcCp6HjRb1fOe457ps3DSf/psgsoOYaZuoWwnzx7hkSmVv/aUN9Rxy5idBa
CG2P9/jabMDHmc+1iNdPIfWeXQXJe9lWjg0rj3u/EC1deBDGuF4Mk1fxHY6OE4hz
opAXj+4dNNO/sivDNn3ez3lztWut3VFYuGPaX9r3BcAcyMMPUdo+147esawMTeBg
FnMF82v02D/bS+KgKuBWQ89epvj8NQJWfiIVE2orpFvW/SGQ+cjp6z9uGH5AkGyl
3Rcawjoo+pCblOJYA2vw9jOPmNE2o+IaYuS7UR4q1ljGDdDQPGbpRUznPYuEfznx
fdDkuJ0DCObmuHoVn7zN06WvpRdw5MuDSII8hr33NmUfEEAQVE11f2TzwPJM8Zrn
erxff7IvWYPifnOsIyW3Pks2/aiSCHdg/kqlHq4b8HenYlDek/TrXwg91IXmyiBH
OJdR/LeDi1PvupgRKC2/VU35dCMVhSz3Wxs8RCuGUaSlBHRDL+Iti4stRpRgSKZm
SSauz3Rgb7PjE5OEvfzT9foFRlxrGJm/IRVMz1NDkAEpK1J4+23ipe+vktUtlV/B
KdXMghgVdIV3zQK912WyADURQekRxNVF/VaKc1knf7WklPLeGJRt7/JNCIU3px/y
6kYBgzVKP2VNQ7D+zTDUbor7mJx78P8aG4QLw88IjZBbcmG69rwgLx6L8JxDHUun
ZJIGx6AqnES09qewhEzQqMqwyzSl/MaSnCE/NZ/4n2kg0WwZCQOXH0XqXtZEMKFL
5j8hEHS4mWwMJmKXKej48gjCq8MuPIY1BStqr1/cSVcBrfcliVIPzm8pDTiprTlk
WMT/AUjTMFIWg5EcVcjGXij5Q1KyDo3BmX0av0arrdHFj0WYgacE8ehWWAvOGHFA
zqNrOTHbJ6dxBCmO4eWyLN+FYgcT7+MMKcoZEB2wRcLl01VWICp58Bgjh+jXq/G8
uqGy0pw6bYDBEjpNM58CO0l+QcPMwoxGo/EI/7pa/3t/QJDDaBtccYisjK+79J2a
CwYzbJM/r2PfbncycZ5InFFwIIw81BCVPVM9qpKOvNdEXN3YGLw5bGqlv8g0Ut0n
CIHb+hV9Ts9dHFhYtMYFXVuSGOaDodFQeDQ4zu64gpm5DkTMLqia5gufclc/qX/C
3VsJ87lt4C7bJTUMsmvsvRr68oAHeeuBLd/FF7kxlnPSxMf2SUENMcx2ctXZ/0P0
XJwc1NeFoWLyg3IhwgHsq98sA+R7YraFQlA/thpW44rtdPK52pROsl+4nFNHqDjx
4TJYSK7JH74ZUqrjze/JObrW4g8w8ZPimBMoGTqc33yGS4BwnUXjx4JYAgeFpes+
eTs1jv9yfzz6vcizb3C55SFkK1bzvx0wanSMMaBX1/YXYlzvTI76DmF6v4cXhLnG
Z+Sm7860uyHwLNYRNzP8+lC8XHiY4ME7zxg70T6rqv+8Q2gw+qhnCSFiGEwL1bLp
VI35mEM9Nfq9hnM7xz58D9Qq2VZCUv4NOXwnFQof0X1Bl/XRg4KNUo3UmzxZWVFf
s/JhKdfMHqoS5ok/n9QIyx4x1VST7dNOtpSlmafNm/yqu4P7szCnVLkRAnOQteN9
xt5qsytafqNnjgYbL9SPiTO/yHX8oBj4l4r5gyRsW5EtCXSqkpj6F1+/QhjYWliB
7EIr2rdGYqaTzzxrCBQMKA+WBJHUqp2qt+6aitYMML0ipuWgGmiKTUHbVu08RDPA
Oh9zb43JLQi1N7IlnalHOXS6iJucvzOSEcWLIXpaF19dCW+EBd4AOIsLWdjPDi8r
U0LFAlkisFKpT3otJh8duK4BoMst1XCKLG9Y9NrWkKEGYiWvSiXJY+wDmtMok5kB
dbNe5Drk4QhfPstGlTs9f5F8Hkp6CWFWvFYs3Xhuou4M0cBNjckZnrQus0kHIFMr
+KZB/6bPC+Ibt87AMLWpdI8pgoMIJgqZXnIXR0bpS8691XFJ9CUoUlBUlbGIObUc
qbZhL8DlyGhD2sKwv31GkVI+DmxJ6EgOGi471X+BXJtMrp16+cR5xJEtz5xwkl5m
J1td7MKULxYghcD4uZuA1j9ahdRtnKjdkOyCg6PwgTFjg1t+5eKbBFDu8ZhqBkaR
lQkjHteBkdtnDMHWun42V+mO/EyxMgzBbzfjg1KrFjGZI825isz61YzGZntzwZQB
zG1PAP+1uqfgDll2S7TXLhMMpU68HoWJiVuwWWZOYDmnbmeiGhAon3dc6eHkF/ul
xXzkR080abEkQ6YlAOhL9eQVEnk+rOKqU0kL16KJXSDAK3Lbnrvk/xV1nJz32cZw
EFMzeeSEpcYmEPk+A2ipZwf1UFe9sl215FmuU0IizBm70t4ipr14uKZJmYgIeOqx
vhLK2e2zclAVhqCAgVtZ8rdaSziEqyo5Gy7xSYrDCVvQOJPLbLE9X93Z2Fxo/pYV
tMc063/HFLz7wz2RcQQUYG9vBIC2xiNIYytO9ybThRtAys45BR7J7hek7MPPV98l
rgoPPSFcxnlM/kHJiNSHbXWS8dS6j5RMW6wduGl3YVkiXOJCKEmO+Lr9PiGk2bEI
G4hZkBvYtfROrcFUkPsE/6sB+3HsVdjLZmt7EZaBvD891SC9HSMZ3p2rTxBdS7WU
RiVu2T8Ixys98TNsWW3ccMZ6Yukw1c18+y4K5OKvjeyR15SuKCA3kh68n0kzfA0p
YBe5kBxU2XFW51wgjxcJYW1NWHGA0OWXtEB+xooobKGU+knbcphSwsT0xXZ+0NAN
KcXrPfl6ZYFBx7ybt9MrHG9mJ02/VSCb+vJUGWc7LFmTyUwpuMe/IWViYYCV+cgt
dnpSjxM/AdBfMuXPpd2tydtVW9K0HI1uV5Bm9msG/MCbx5yL0WHen3Tn3vO+s+fE
bX9EZtq4jfv5a9LlKkqn2W1nJoMpRMZTsFuBZWT9SlU/el5vQiaHdrFfZQ89UIEj
/o9EAPIzIvUQblRjMpdldxlKazFG6GiFGRReEYhJCy+0ogpEuaUAmdzA1cXNbkU9
CY3OiZwspVfVWFYJgdBLtydEbDOML+HDhiFUQsYa0jEpn0UPb1zyYaKZHIh17cAM
TV6kQs67ShLUtN1vtP6cbnyvo9h0isEG+Gq6Ueq+X4T/jYBDFxF+xHtaWzCX/x1+
Sj0RVgf3zdMPXzR4+Z/A5rgOUcqKnovuuHRoGoqhO8qXUvQcRE+e9hwbRzK9tIP6
PVPJQELnY0yZh1RobGZb1D14NPNcE44BBeDwAK6eWXwXrwfIhqPE5cDsgN5k+eoC
ZVgHont67e5NoYaV9fjgp1NNTCuhHo0ydYGAaerbu9RCgVOK+oULS+9Ch+rlPlBK
pHl2zpDRHkZMiQuJDn+tw0+35dCG0I/nFkqKYdOcjcfmBxYTCDxvdy3fvme+OW1V
l2FX3vV5cWTU8NR2h2T+0Q7CqAl4azeQoV1nE+xaPeGKx4fpQG/bcmJNmLY5qNvC
1PQWCG8yZGl2M1q9FnBRf9xQD2xlj5eWBz9swTMvPH9Jp+LGSlGxiQWCzF7p2H3W
KIyOv3hkTMYlCxyDBWnGyJNaetbtvIib6SXrFMSK5dyAGSTAuUl8f4vWBVM/V2uE
H6kWh7KK2aaMtCkIHE1djX583ddsaP5hMSL5mLX6uCTpXrySZgfJdlqx6NlpCNoM
bCzV3nnfxhiYSLmIq027Lfe3k9OZs9tWz7+CeCljw2sZ012+TrY1Hj3Sa00g3CvL
ZAiTm+zng/oQFdL128uZjoBQEif6XNVYlx64NZTGGlMLHv7402Ne3/aLapuW3C4F
OYOFuLtJt3YH0GW72vqhBFrlkI+KDwwh55xJeAfMWO8p6xhEzslfgVqFyKDDXU4P
xLj5XbYGHFDYDQ019bVrD9tvB0N4YCdif+3MBcmbLNb0ofEC7WoERwp5RxdnuwVa
dpGEGq8s/a/eebTcew/wToRWvNji/2hZY2fBIT1kTIY3SBbcGZFy0RSiIISYiV4U
Xytl5L3TNXSzBKGYjCLz6IW7HlTVqV9fc2VK4cnOm2/x8XjObAHehFBinOua85Ox
GYWjYgxqe6VFzP+pPqPQuKgrA2W/R2s8nYTdcRZE4cIuFKqH4ASY4HAU7dOECJ8/
GRY5V/IGELY926IcWLSmc3sf7eGTjKasNLxopDV5y+ESElb7gR8M0VnTHrf2HXkf
abCPuiS/QwvvKF8clxVRvIDvnJeOHiBuSILdh20W3lLoxK2rT/TsO+DV5RT/gvxU
Wqwn5BPK7THv7j0d4nZuzS74dNjjscZQ4GlHnwBHeQIiFjRcn70sf6mGS72JpJTq
+Tpi3vc8ib9xNBKpC6lL25nbvOdhuy5WqF8PFhnv0H6qPbXBbx7qYiwfgJVKQhlG
XhJZo1M8eZXceEodBYUWh0uIAhOMoVjxvcvnFmkOVohTeaItm8bx9lcA4xbrfUWM
yd2kNZKKpYgKYrkEnqahLpKVw6BnKj435IkcDevp4CFdnYZHIqUeRLov0zU1Xodq
U+JEeoffUNQKWnTL7E5oVhgxCvHSByeW5ZKOI+23+xDKCNBEmnFq1gSFHwE5+SHf
UfikVorJwOWvGjDuowYleLWsbKOhtUY5LpPwAjtmE/zZljynr8uEXUScHjLqTnxi
yxD32WlurtyA08xZYBGnXAcf7N029AlmwHqLeOUFxGF8OPipcHF7j35xFvMjN6DM
H59o+OzUU2HwN5QAja7iBTgMr8vaRBcNcuPu8vkDF7uwh3lUPte8Fe3Yi9e88eMP
Bc7lbjJwarEwNsIntb9TiDZVtjwGRwUYNCpjQifcRMDo1QOYW7BUiAlC0TO/Vn5Q
D/Ju3svFXYS9aA/uX7+dTvVz5JwHlTPqMwkU/JyRuclOOYNZlhFKJDCpe3iPB5/O
daisZhyERSpPWosnfgWu++pzspYjzkv95iAKlZdKLo81Xp17lxQ0kaB+KUqPnm3o
57N6QFYIqyWy29WkyBjXvbGKwdSvY7nZH/E2Pn5c9/nXo55Y49mYY0vsmobzt1SK
bTT9xOo4t0cYkCplzxL9kKPXjnzBO2C/ljvRwj4eEA+06s6KmPlUhB6JY/elJ6C6
Pa3GAyWK7yYfUGaR4CVoBOFiZrbkv5NAS5fvEdBcnr/U40TFrjNNNa7xXjD+jxVS
dinpa0OH8LyInRvOtIzrEj9daYzO//Il052+hQCbxyGRf9yMng3qOL6mfzf0YzG2
XobEqmTJ5tv71MvLzrAVb8mPuLPtTly9z/7RXvGdffEnTMcRDBmAr/kgdVCrWie2
zlceSTE39TdnkmqPUBG4h4L3HuvPewXWrLH7Olw0Jc1EbgzXqTn1zKY6dXJXul1w
TmHv33ohSv9if9hBvPuhvkGVHxP2/VI7H59QCMlJFOfGUYSA7WsK3yG9MQt/49Bf
R31yKKla1LVz79kMi92BOWRMR8B7F1ri7E3ZdACQTM6XwG7m5YpiitJIz/PL9Dkx
d+geFaCllQjxDtl5J05H6IZHc2+F5q02/4fUmjvIEikyLFDc5JCIsBVpqjupSz10
TCjcuIuY3g/5GyrPrck/1pOViKQeAjTHq9MAtgowuQxVhNWNvesdYIaIOpJUo3/C
F6p6JfaElGdsECae9fNDxcZyvXhXkg/umZm4KTNizDYDxny82V62IZ4WzqnTl6Ic
UwpVSzkPoEe7zMB6c9j6I3EQBmRKNv6yRla9O3HfQAqUv/HuT/ba9WvH0PwaijT7
kDo2ojRR1SKppusf1kBSVHJ2aNHSiAoYEz0qTGnDW+ZE3tg27ERz7rVZcOL8UPp8
5e+OAkO//nlzmUFpLRcWI3NIcc17YVMX/7UIAIp0BhvpWIQSAnkxmo5dIa9wfUBK
dfOwmq7eo5vME6slqLoygYF/uNwcwMgHSuN75JsPUhcHAkrxUUQdvTavrW8BbtEy
tqnd8rc27KuZfCZyeeVDZ4uK0yRpMVMDWe0/NF4UjQeNW8zVSLDooVhZGBzdmyqS
dZ7IMkWnrDs6jDgaJrVv/rXJqDnmpZ84pc+v3qWlJlsKRk4D4eOoSGqWXHPXF4ZV
/Ps4fmG20b2EH56zi8NK2ZejI348bIxSGhDPPlMDWVQkdxBdtzXTyXykn50on/p/
wZ39TEjGRlLCmYZdtcW5rh8+tep2tYDjMr5MM4gi6InnMp0wJguREoXYSj9iXlBM
2sqf0VCGyPUPEK3/aw0UiBHPKZAe7/t4i2jPUYb+1fkeN/SLUx9aSGdWiWoiUghb
oFjuPlGRBWLXn93sAp+ZyBUhm7qsvc6YdL9fAMISHVFi5v4zgX5OT3aGYf5SQfUO
z75i4oihn4UR8k8COkUhqj0bAW+kJ6sWLu+BzTu01ZxF6u/zyRiwq0LM8WjQ6vLx
f8YCQr9Vf5II7XVIcG7UkzMajvy44G2978ik2ORCmQmv6eJFwbXMhB6yeuy6XMKD
e0TetKiYKYmQR1qvICMuyxLtXYtm+51WvGKe8ppqsKRDvfbDHYxbVOs4F15zd21U
U0WarPQMw4IZDMvg6553PvMhr7P3wHtvZJ7nhae/Rk8f8tNqOLRlJnEx1v5Th7B3
CITzeNaFadRRg0zHn4xHVV5vqzzinub1kbQJvQ0q5v1RadmBsaSN6bT48GIT+CPV
poV1D+8gsPOBP99A8aOniwUTvQXInFE6MTVLjMnLmRjaZtibB2GAyzcIe3XB3jxx
2nfchpc3se82G6MqyNdhFruOp8ZUV0TxESdjIMNZrrc3EVK9ypcl70u34QTMvbLf
xQCRgodlZu2l4cGC6D7WAdnKk51UPGoJ1c2ytLAWVxJFqNSFirgPhjWz4a75ftvP
yHCMxr8tLoMRlcNlT7jg1TAGbFpkVDrPRP/ClI3OxlxGtj1lWcr8Hi7uLoIiiu8/
r85kwVJkRPK5KXYgZoPNNTCOU7ZH8TZ/vOENl+d86/62Wjogkj+RIC9AqnaWzpHn
fQKYvsMyJod2RfiTRAhW3txsRwF9mkGpTeSJT5uDi6Rc42Vkci/hkG4FsSevkQ/5
SjYParxvxs6jNwAEYviAC3wJdGadrrIa51Yu7kBV3m4Jy7TBmqHIVUUmO8tfCZD5
ZUKGJ7Z23547fR3sG65eGnC3K9peKTnTmwRvjoxAX4y5UO0ymRqwLz1d/tpkX+EC
2Xp3Nq4+2BXSJfWvgTXQZD6mqO/o+fpzFN98UAVb5oRppg9wfvWg+z+aH6TRFw50
OcCeUJOATnUr4/97nd9CWF/WbxvkSSik5DW589C39HPFoWs9VYyST8MVIqcLSfV+
BkMJRkfnr9UHR12COVLzIreVMRdoIiN30l7FoeZgfpiD51n2rBbk8p1AosLXbsPr
roZK6eVtfp4BM9nVnk1XQdEutIacy9DBrWzHYzfy68Nsq6ouyIjcPhIkWg53MkH0
ZYvOHd9sb2urwYZsQ1eoD1ghPn0UEAiKL6tBzWJj6zTiXSUAoUc0lcqUvufKZgM0
rqx7I7nuW9ZDSC2YVP2eitqg8hdgOlYlPQKAFEeElfS5CZwUp8NOEXHJaYoGOAsz
ZGBlxCbks7WFAKbYV5IQh2NuBZhJCK6gxiS2h5qCiP2QLORayA/9vMXidrW9ORN2
uW0ZXXHjbRQD/QyoHhuUW12r/iaaTXLg4rCmeAthOl+6dwOkAKF6JdZ/Fs/jNN6K
Aoaz445sBUd5393IoEeHCOHb8isBam6Tr8H6H7TNXSmh2NfBYSEM8YfEySjhmcq+
FRgj1hvV/xftnqjE1V818EjWde3xiVpf02PwM80VlQmtZduGjsbnk7uXEjLCdGA3
ZnVvwHivzIAS+gryNT6fH5bWQBga7FI4qrSQe5GDcbI2vybPYFcJZZaYBAujjUCh
oN5b8wEQe09M9S3pcB5dPHxFh7Y5nLrQlhWZ/aNV+hkk2UUtccdU7/ZQDDj+GQwA
j2xDxG3NQONCTFLSf1FSerI1YGHWPpfljaw78+/qcFz0fXgkzibqIGA+6nG4JNX7
n92/4mBaVA/Z1r/UfJ+znxm0HZC2LvTZsAwvmpN70Mvy49DM1ToiV4jvUuqWAc4r
C+K8MkdazfMfDl89RbQOO0c+hfAkvDFoqXqdK3u5TQnTPvQt2pkTZhPtmQzQjmRL
2OA3eyFEH2uc2aPB9Y5yYGe0Q0o8S4M+nMHqkkRQscxzoktR+DTNCwabXAEVDOGp
rEGCIApl6iz/tZoMXUGPWTKe6xfiaI5MKkclR3Sk+tTZvq2liikg0Ub4RDgMywvM
f22dZf4njom4Me0GFunJTTvKF+7nj+ItB9xRM5Gyi9/bSDt65oto0X7lAbiBORCG
cJK8Tk5E1VXyYniKBB1Y9C9F3K+XkCG467t/xmzFqQmlMSpXQvA0dyTvluvwbO/s
q9DRofXOo151v+RC9mvfcwOACtKmfMc4ejhLDtE9v2bvc1rrWrBm9nRSAi2pxFqj
cuCJCvbL2ka0EATZLvk98I4U0cFW/IRVpLfe/Viwy5aLZRdmX4NFVv4O4s4lAzbY
tIiQ+aBkcL9z/WA+CGId/vdQe9Cxa7J4K47ylaEEaOQR0nhcIeTXfOWh6qg2CPV0
fhJhb2U4leIydVfBbGvO57Zf5xhOqlcaxo8pBVSwaJBOkpYjGBe+AYKbSuskeXpn
TFzJpMTkfmgqoNk/AqpwCrxkHu0rZBQzEcpbcfCXMnpc4yJTjLK2HkVmINXIJ5/i
hLPQnjlMZHjjIduCbr0J75TZe7977WmZt9P/iVR3aii1njL7M0di3JXNy8EtIuPB
iMOrrJkHqmwdTV8auf3Doo+YPTt39mcJdXR1hGvTteeRm1QZrln6P8YC3CtUVCTF
omo24FWp4TvhrPHypyru+Oz64bvKqFjQ1nQqdfl3BxMP/iAttV6nrm1j/cDbCmvf
dHxqROPFQ1Bb3pBK8dydkH6V3wsjB4j3yq+O5GvMhhxCzQ8pPpCmOYvkcO+4msQv
bVTK9wLB2NvO6Pgf0nG+lQS8xLLiUcxVGiJcY9dBuvq9SM2seNWnfxpx5BGWyhMl
Ya/9wBlR4Ku9mInHJ5aprHDde5GU0JP/D8/gvYlfqUl0lZDJnMFGmPbTJObhWiVt
LyT8xPhKJvgz+Ngqd/PksVzC9d/v2DX8UOY0jUc0Cob4BX4AMTpRhNQ9UgX55dQI
j8CZAES4MoPdgo4GJLvqrSyuC7EwROPYa96WHapySCA7ptdTXkQIPbaKiio2CK3O
4oLC8VU8oEozplGS1h/IZCgTSoPh+jwCrsKIvMobGguOWDTQ6XhH2dRNq4KyYJgz
p2w4BPtAuJJEAGcSJXg/Y1FDvwdBuYhwq07RJv9XrG663TxqFiuKnytAWqQRedvU
zNMPD7b7xE3J4Vim0lcnq/GGuFNUBcVw2vj5/tgQx2BwvWu3aKkQqy9idqCO9o6y
FZafp8tcvn0Fi3a2Vo23pXzrqQPwHu1kN1qzLgkLPW52h45y7fjQgh3OYrKp2d1+
+JxYd8F+sB3hiRpRQC89js/ywwo3sENpwU4Qe2bYeQqhyfrPha1O8QecHC4KJdp3
l/OTrdQ7C+LM86TEGVQFv2lk0ka17UMK7vKP6/PBZ8yvejRFegzGQ+04/ixAQOHp
8c1nin4qB2qhOlz+w2V0vLnd+QugJ/4ocSQVPxi4TUNMdshVirk16cQhmU80JuIF
CCk/YFpSn5wT1cP62KDUqnqFW11K739O+/Rpu1dyM7x0OtFfewBUa588YjBjiyFq
DCWOtjUkL4jO5JQhOasHtiTPZfVibAiVsMOumMz/MkTIlRSIwlYOw+TA4dsabKXk
BahO4XpZOxb1Vdc9cNO/HMQVXFqvaJdcJaQlme4c3DhiE8FMjMOkVc8ckr8Mtj/U
Bmttohv0NPOBxTcHd0uzwLsARoiG+2UXpwzEh36mCb/+0BbXFIeSsrxNK0kQiKKi
5ZfI1q3WdsKk7XyOxDlRvjS4eEkuM81VglkbmV3riW3s7oT5koghHXI15atX0Sn3
MDQqGgRweKAKJNXbrU3KmZSRf4/PHhRDMYMiQao1iG0oi3WY+gECzJc2UmtJXBH1
OqsRCTAHm35Wm6xZKe3OjCQ7tavyQ3cI3W3lv8Klcgnl8xCSc53x59ctnQaK5Rsj
XIhyFVCtHYiiijRB9JNQDeJJpz+IaPYdVWxeLWHpC13jMnxX6HhszCNXFealtuLY
RrDxBhh/7AYY16qt8eLZd3c4boV55Ez0+JDRJvteqA0GtMtMsC1GbPEHAgqA1to4
ZVa/uvdZt7LST7gxFjvmEPj+dPX0YhNVCAhI37Fr3F0gNBtEdqU2amMjytBKS+rV
UEmX54pUXyWkDaOlSRtwnmQ3gU0s8TJ/JOrDPUiXGVaJz1zZIj6otKiKEabpiIRp
hJG/Osduo7Mj8WpykJBcoibPpIwW+OutWUJ07L3B3od47ncT/94gIFkfIfOweQ+L
3y4mkox7vyC7aYXG6acn5fbVoao3uoYNWm05HfVVFOrIpkE/AY4qYa7y/kXazKcv
x26Ja39UcTdGC9upJllaQ7O0di4D/OanqU9hLBSRNnhcz1TWj0lAXlkejBKOSDMz
R4M8CeovYK0dp0UrBczz1mny6DwfNftQsE3+13peHr7JqncCCmKb9cdQFXOic+a9
J3wFSnmGhz4e36+gvRUbx9csH0EKdigwXoVTfgG1uYxn0t38WcuNZjG09ez/mVcl
JlFbzBNZKC8jxVOCNp1auHSeDyYkx2Oz+w31Sd4QENeXIKuQuJfadsMFKRitTZqg
lJxtBnSK6zN5AHD9zyJgFOuGT/6IihQWcfAVphFWDtBKFQTciDfaW9E8ipN3fe0m
FvwrFQ3BzefYJuYgQC5U8CUg7INDg2ihjhN5D1wWkuQmke3K8f4XXoDWCO8G2rJl
D0ffchvkiYTgbvvu4vsiiJAeJXW+/Z9RceSWgQXGBd5XW3lcYNhBp5tw6+l6wvfS
zWRyvZ3Yyba2T0J1KDM4D9+Kdxob3RHpBaYzPWqnYASubF9iIXi01FZc0Q2FcPlb
qA3ggifP7f4zXGePZA71dD9blajDzKNe7qPIx7Wny+Tw2puXnS7MRukUj5SymJXc
1l+LYuOxHbsIoem4WxSX9WTS4qRyGHtLwrd12SpwzgHPwuTp6iRq/3WZs6eSkRgh
Zn1mQ91oWoCZFYiZcr9qvHXzkn/u9LdR+BR1FhC21JuLaK9ZI2YSskuxqTsj86CD
iEWhPYY+M78VnaFudlm9ba5MEjur8XMG6wuWeLiFzcxSAWxZr4ZllSkL+qr21NRn
CirRrYKggkCckzItwEWYkJULmdIUKnCaBhfeNikUYnWFuCo0lsRM8ZRaCczGBf+L
Cf/qkYaPH/RI2ujmjGv61nDXLeWVImgtlX7K/t9EbbgnKDyADg3TPRV4+RPFOcLh
knU6T/ThkuPzetQ+BHWOs9KTbKQSCeZkAAYupLab5BLUt1hFGK5IDB5gveE4Ze5J
+N7yObNiuwhRpenr2mtnkxqBJITAQlxTls1c3Hjp1tdk0YFaKhqPHjhMPsxWpWUD
w46gSDCtEh8zczBcQtoS0xymp4jFM+Jz9of161SwQvfzBGxgL7UZVpIIOS+H972t
C2QHXUZBJk5EdDWnZG/SklJ90hcmlTfWAIcy+2vpyLq+r+P5W4zxrj7edoC9CXs2
+trvqRjrYxLi8kpeNiL62aECxjKTAMNykAAvhjTYC7PC/04mP42kUBj7FtN3syyv
Wc1GGQfzI5qkH+rhDWbQEZgKdoGY8BZ+0QHwUckYJPiE+81Zl9KyzUk0a5IKNKrG
Dxu2Cwv+0aSok1XQUDdhEjzU1S1zUW/6reSttGj+rdq+jzsVGdI1dNXSF6+Poys5
0vRGVOWzULssFAB0s+b+pPCr2kSeozsgaNmxUtiSSd6kuOGqrDFLgJmwIddfOZAB
pDs01+9Xz3sonjB73YwSioBp/IIjKLpDF8ke7XLg5lHwzByxjWwBBriXD+5IoiV9
UwcgvsOeZ4u6uxbkawGiBZuKX9dL3mEA+RE96AyLi1+wD7idkXuJgnL3uTNs9wUY
5x4NwaVYYpoQr6n6F+DbzhNZbs96zDF6uKJ+gqyz5ocG8STML8D7mrZ80hN5XpVX
2mdnum1WPB8li6NudkHsYu8DGEo7hrJTzI/5VFTu343oswQaEpnXtt2ai9zSEXky
5OyP5erXUxVCPhZTF9VjFLdAV/kqk+7fcZEjPhDHSkG7hVuIpNdt3ninKxSpVg6q
UruldmmHxkoovMXpqDK+sibI2g6CkqPhhHLxlzRlOXYUf2r1DkgD2QHbdhDkU00F
BWk7M1Ea2t8yAVDq73aNSrlJCnmlpjGgi1JC1Q9xbZ3Ei4H4QkH7//rWIFn6QhY8
ZOyRhZENceMRCiycp4FAGaSmgW+Yx0QohdV2sZDzLHGZbQ1X85yXgIbb8IN0+S5+
KKrZRqI0lD/GYPX2/ZyzdTUUWGURRMhHHJ/AbY7wQqbAh0smi9/zm//wq2cJt68V
wUh6viYRgnodTmTnCTnO4i1stldQw0ao796zrA5EQy/sYiq4gZhYwR26ebzoni4v
g7wyhOKWMVQcrIfcxiIp1XPeBFElpku0nBh+Vd5GYDy92ogExvkQBVXOArc5YZA/
3Jh/6JsByrEOU7OaVqAJkDdtOk1CluGG0XPsU7WfXFGZ3gaYCUJH6XoacZltrfsH
fjnb/jm81WUTK7gupmoHfFvM8BtAbROFhHeR74+ZakpXTIf9irdR1HWJt2zpq9Jf
JR/KGEXUBN5HxbYbL8Qe+b7DbLRCxuCc52/MmVHPjjaoAZDGLY+cB631mnRbrx+j
ihggY9xNL1hmcqz2buttL4nlno5BF/T/JfPfkDaU4BzxLKCQ32beUWKyc27R3uvH
YDem9fTxpjk4Jz2K1tP2zxZGD1dim2c1gGO4s/c4h8zhmvsK/gZnGeV7bdHM2gAA
sJUTSzywdl6WT3qJ9WiVz+CzcWubd1KusMRgEOHtsB1fctuCyujcVSTAlf7xgXA8
ZdDQb1rs/2A0IHk1KaSAXrAUsBcGtnNcDyRUROMlczzuflxTZ1LwKUDg+Oa0PvgE
TL1N85LSC/2AjOKrY7Eiax5vtIIIzVMLvY4pEwvJpzxG29Op7Dxx3ItDpmoY41tP
ANQX8cVFcSWRjWNrFOPTZqK+IQBqd8TUk/omfgJsCsrm8QMvsZS4Pru1C0vS10dv
wttDNcQxy3lIK3DL2RWgjrYfjIVY1iXJvzSkoNpL6xjkXBMwkdF/EthrhxajwZKt
MtsnIHBN1pOVwVfUb/CzVLtq7qz5rRnyGem+lamwxcgDjRd2tyjZULvYMGusRJtV
PSkmHxyCt4eOWV+Z2FNx0Jq5Js/bEDipYx5KY3D/gpSjgLBnNeiw7YoBu0/teCon
xKepQjtDc+UEGP4Ihi20+CO8DU6g8XLE348Ub10Ibv62+2r4C6fJ+noeXfWwpVYD
/F8kXE5druHBIn0HFBUp8bIjV7FNZZJ32AMOtW3U3HwZdz3w41vrp6Vnhffl2ymY
ep58JjPnLhT5TeeJAVQIaDqutKFZTZibbXbYuXlIYOVrShEFfyyKzsWScANi9K/Y
9YQNt3QAdyavOJS0tgCX0isDxh+nGhyzeHb3EJM1QJ347+dzcdqe2QY6+XdbdbsK
jdfkd9TaCxNhHKOoKV7K3wJUc+wiRlLbiSoEEgxLEXuGhs1V4lXDi0o7ROvQOZ/k
plX/d2jl3VUQK17g1TsgqtTnD6wDt7+QjZc3xdRSVdDljOmW8agJy7jfmsG1hy97
WWwiNnkELdw2DfqtTDEbq0nnZXuayAgUE5RPUOBaY3XxHlb9FiqqIsD4sDNCdtyq
/ZXNyHoRqSdLA5Tt0dGz+siic7jhXTQxy43o0cyXngRQvkJXlZ/ox5/MEw6Zt/C5
St7kixXaz0JB+gKDyHXnNPC1RJ1JxWZFDs7I21Hv+D6J1bfSkPJoG/aGHMybBX9C
InDSYYcsUcGvGaQsVJmmNUTw1obQubbPk53Sgb3V4be7+BPQs3sFYyrDFP+B0LxF
TL3oWNhZIu376bdxVdF/C7s5QgABhfDSCIEKL4G/fyVM4Ru6LS0joNoiLW84s0O9
Sy/nbIX/Um6RuTLj03kLInflWIQ7mdAfyLGLTMmNER+p6uLqmjf29bnrVw8btCep
ioXdXYbPU70QxSPczm50Ve7/gtn6nOhDV0J6TDEv5aMoHDvOBmuQ+/r7jq0OJBjf
tHpJ8RyBaM7gDHsda+sZkAjjGFe6baa1K0rapTm8s4VKcgZ+4HYMM+L0hAyxixwr
hilRwgIWU3TcEj5E92juxTUoRHIJIoWMsAFeR5KuCeK6XAxFQ1Zck+d47E33/14V
2EcOQoLryyuguiaZfuBtW3dU+nm43iIvtaR6sBFfWf5Hx32vEISnEmOHECcHwm0C
HYu++6/jNIR1VuIv+fcyJyMQzWaq+qaMwqXJdCknMoTUppPGmg8NRVVJ0jv+YBFs
hjHyEHh03odgaT8Gi0OPOMIBfK7X+r7AdcdbOFfa2yled6AbMjMVHX18BAznY/xv
9Vr+QiYtTeFkmRGTaVXDT2xx9kifnpbIaacz/2oT+scE2lQx00ZVlHNygCZW4JKL
1me5PCm6HqzeHQ3LIsoFpqWRr3kqh4t/TVWOW1EEeVUeDu4KqRLRdyrog9FFRhiJ
9sYgzHsH4p9RNbkGR42yDM0o5u2mIP+cWqEKUDNQ1Ns8nNgxOUMliWLegmV2umKU
+pfB0glWpbdQL1A4QU8rTjT9FohCp1ecF3oEp2pBQCse7QVQeAMHS6t3HtTVUhD1
a6Pd0FsT71ciMRwJf+YHLpHvLAGljfpfOWURukJLdAc9P8I7PWg9RDy6c2DME/7B
T/9uO/Sf5qF7zxq24H/S/ppumG5MqICf8381UGWx9vWEUsU5qvXlQ1wUsx3GEyfa
hhYJWV85KT8bB9v+aeuD2nCEDt6+NblZSjw0QSwxXZXMTAMr6Bp1AF8DORzWChd0
J9MAH147FJKeHGA98/9VCHBpYWOcM7mCuGqxG+TIZ3xCEa48rz6mfJ1JbbWFgpLc
iG/vif/6iZyOZUZPQ8MjcGAGa5mkSDUsT5ybG537k0cRlAIiESj9+PbRvda5U29o
VGYOT5jexsQN8Id9gGVcujrFvaR80fsGm/v9CFmAdlA3kJP000bNKUtHxAFUkQcs
WryijkaKtFRLM6sh+NkXXNRn+AXnoOetqgMlCgKebx9DCINjYYnjyG48qUwxWHEq
hwSZ2aixTFQCKu6QWDQTX3BEcn38ih04sBaOgq8inVWTzDrvoboHqIEQleu0/7WN
Gg9cVTJvU6i/VR4/UGvBPMHgVJzvVUI3WHNnHBI/MW4RlSFUz1EBQQ2btT2uOqpz
IJLn4i71uJSmgLfu8vvuf8djnwHOsTR79QKgL+dxg1/NWEv1KkZc9C9F7EAK5JLQ
9dSlCHi+6eV+4R22moP/Iley9s5VFuRr0pXQoROB1imqrzvqpRTXWykcGcpPSyN1
9DA4/JusCGEqOMBEUnE+/4bV47fhkab6rasQea7d1jGN6FSQXRWDg56tcf7BwaY3
p24Uxe/EFGomh0SjGQHjim1I0SEejoWCDO7aqQUFqSF+1wBR7cw3ish4IUT4bmv6
4UCe5Ec5F1OSc/YAF5xeZSJO668TZv2JHI1oSXGFlAeZcAZiD19sarYXS7xmK8e4
p8ld8GZwhhGNuj5AXm80b2JUodMopf3weAgjXY0JrOebB/VvtgbIGCFRc+fJsnuH
ub9QX2quwtalyLSxRPUt5Q6kVb+M1Hxo5quie6UwKUT00wzfj4V0GcAOIwqXgpGA
YWZLvCcKHSzYfUsSSIYTYQeObcTMaCtlW5VWz5pPTAp2XMmzRlzuIkYpQfEfi8+1
yNE6ASdTKmuX2ESCtogP9Z61KbHx6nkq6cD76jbcHXxBB1zH0RcnWnieGfG8Y430
0i0UWeg55b+8eSkJwUsZf+8rFrxWoIkFin94lkOXjZxutCZziYzClqpfmDw4fmwb
cydCOzJ3z7RBO1LVD+dWIQ7IiCkCwNFPbMq7Y08ZXmvwVL4cVMmp25WVBwzCvG73
tGlUinGP11d46CXRcwKur73DF4HdtynVr+c+pOx4dJbHL6t2OED90ehQcBlWV0RK
mUvUJ5PeFiby448gO8kBkgvINqv8Ipeq2t2+z7wHNX1QkijnY+l5iz8GTAoAWS7I
mh7tFM1tN/M9QG8gQ9yGzMzoAmZGfmv8JTgZMv08OjMEsfo2dqlwU3g1SHUA2Ik8
2cCJBcagERo5sfSo+iGoQNGGdG42v0YRVLTMx0uCbnyWPAR+HU34RgDxF/uqq8aG
4hAIVcz8HPOfp969FE1asGYeRQivywsv09s+xiY7WDV7V05hE0Mj3rzO3b5O9Di8
LWn67KA5oVk96ctSa1qVgNtSNFFUI+1PQsnHGZMaAoRkVFnidmMzqZyGbyulO6/o
3nafgWQHQAxmLXOAx7wKPuTGo3KtwNusI0LJEL+i2DERYvrcChOPy4UlC49u00DP
9Nus63G7/g95WWTy8nOw/ZO76warg4TNuRMAGBcnjy4zy7q0ScyuxhahWgv1DNEZ
XGhwwZtt835vFV4DWxx3B+ZPmxsrB0igIw7/iSdoasUF78RQCfDazDLePSDfKA86
eHYiThbjBeVmxH5em3pD9Crt1ALnyb5/lluTF0Y8ZTdNkfd8NZ3PHjp002g500Qe
k2Dk0H0gHiX3inD/9Fhj4SgnbOGjl0isITmjqNxBveBwpamBJcVL4XzfJCy4yRos
Y/VKz1+uT+2huP6xnKi47u0Zd34hgXr8G9fj2R9lVcFtLKtU9oBfRluMNYpXsjrS
m1ENYgHQilrBzcS/8i52kx18yh/PNVfnwwsD8IT10tdYBDhHG7OUInzbP6bMaJiw
VO/Y8yYWg7FD8xCu5xC0eBk53+AjFrkEo7djxeoN+wbkBbxUOm4A42jK/IOASOka
jQC5Vk5K8orCgab8M0jU9PEQQ75UsTQcX1BlRpuP9zSNB3yg+ZfPY3VrF2IMI6B7
xk9D//qhiZNQFc71cH+2joT2ke3uwDmRNcdfQJbrWhszmn1mmMf330t5XFVSiCV1
xI7MQ7TIKlFbNKu67gO72gdUsjZ5C8U7Okwg7+HRKGhU3p9UAPDtio3GQIsIZi2v
hU1q1S9Ff1BVqh0Rnmp1QUzkR9x/N88AFNJwhwPA+GuTsr5ng3dgJ9HnBRLBLAUI
2v5FdHujedfQdEPVZKg3Wv1TvO9lm0O3KnPcLltmnuEuJqyvZUPa3U3csYMmHMnB
iZ4mgQ/Slu2e20v92bbzGhhoIFJf9YzEbog6Drs6/B3fHULfU2SLdEpxYz++G1Bu
NlbLlIHUkjyddH1CnPGX2UcaWgDjU0pg1WcvEmbQEXFsENPcBEXQNHBCd66FMbg5
VmyoltkXeHdQa0TxSAOymxCHgFxGcebNJe1RKiYJwk/fxicg8yxj14s274DFB+Op
VfRIuPlyNwPSLtfFCcHQWMwR2jGR5oKXyAUqrnbhCATaApRTc7Tl+nU7BM//Hbez
XsAjJlZxnzKFgXeaSWmzzZf2Cv0dRXIiuzOJwxJTIEGH7tcVwo7eMNwwaEI1Kp00
HD9POEDSs/0WWHkLPxkfz5nDWdWohB+Z1MO3T1XIKFAU2XvvwZ3WGke5kFjBzLO4
JA2OonBfWYT7mGvBX8fcYaIgQb+5wUxB3WxgwWe6/Acr2iV9lAIYlOXMJcpfVDg7
pGaWAIXUM117vvt1rNZlIowJ376oIK3Dd9kR0TSRJbF7PpKYsJC666qybzovgOBm
DFxURvMaHCbLBYImbPyfvPLzHHCba5q5f06F8dx5SC86RUE3k/Sc8rBM4lMPPD5K
UvX9wzk3Xamg3YQxWIXO39DHd9tffOPA9pkSBUHq131oSQKmiU+0eLMbMZPJUZL1
wkXLmS8b6huenMHiftlc0+CF0U7qQXhJo+HW/zbUmRHrSSpxU+AQOiLDjpXOCOkH
qd1N9riPnQ5Vm3hIhqzKIZYtwUfYZCCYmhOmKo/eZ7kflONvFTbKTx7UAp1lv6VO
m4MliZ0Yk4J+m2r0jlim6EhDlQ2c6xM1t3aGWfvNItI35+GJv2n0G4r4EPNzOsmR
MKWX1Y5psJVTWTkzJl3tGsA36GrZ+I1Qdnykx9h4I7fWOe4YB4zmy4cw9WISO0M1
PnGydO5EvfnqeMG69uUcZJn+Qa41Jo06s0SLln/4Vy8G1Z0Luc77UB9spQrF0qar
sSnr4l+JAv+Vr6c1Z3808iJmST5piS5o2ySglFfDIrM=
`protect end_protected