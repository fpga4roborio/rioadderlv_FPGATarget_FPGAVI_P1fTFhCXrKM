`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
ddtXksX2+yylW5zu6QL2Lhnb2d1sD00763mmSITNX595NcHTEkwn0zB1Dry37fOW
FufOhVzEJp80NC5qZ/+F0Vk7Ik02dIR0elf3clrjeJRK85K4e3Hoo4xn7YbFUIms
l/8VZSb14+JVGURjfswrIyCUotIzlzVYZ6gzoZwDXIi5gQIBf/gI+KxNXPaKV+PQ
Ufys/12rjO6aI/pPlqSm0hCvftmBcnezN2hk1UeXgOIuKZnogjOsf0iJVX2aOOWE
6pD/psybjbnsNB6kH5uFTA5frkzIzkzl5d9+YDm9OyC+k84E83I/7/j+rk4L2dah
QJOvksSIzN867/4Qt8qYTQ==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="MvBXkzurAa5VTw+1JJ70nePUfoQXBvZOku/SMmg4TwQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
oRtzZL4VJ4iwysPsC8SXYCzXS8Fw2gtZTOskLcDV+1B9Nzn1zTyNtlo6lNICRmmK
ZRVu2BmCc2G+fmzynYlNTnSa7C0Cuel6FYpxCBlOuk3OF2tzAmLAuDyOH3Z1Yjzk
a0aHuoCdIRKv7BrZCdALt03JeUmXKPdOmIlkVGFl8yw=
`protect rights_digest_method = "sha256"
`protect end_toolblock="Jn9CQpRhJt4rnzZPRk+dOpzAubz7omckX1MrFd4p81o="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 7648 )
`protect data_block
gD6l00tciPUa6pDNTk/+t0OO0nC/UTtBwLB41d4inuAUA3i/ALrNyoJVcBnAmEQW
ptbcNp5fxEUJjnOxnedyZEuEBxWRieZFQnkRdF269oOplPWLYVmDrUt4WuVBjZ0w
hiBt+zFf5yOp+dJyWIu6FwOaLUS3W2UbRzblXl3dsRRjzwWtKmmC6uRwRT+d67tl
fgrdZu5Ux557BU1F1E43ZtdJx+9P2sz27EWuFr8dHgGVIyCfyGn939SWYjoKEHkZ
qPnJdjl0IM6lfk0KhnkoLmi+ngZqAOjt3V0PunBE/Ci4d4uuNYCPLMNwXzYpE4ot
MrSJXpSjQ7zmSVVz7PvLot5KH3lc1muaEMZm4iCTIKEDdGkGt0DVdFxJw+wBdTc7
8BgSg6agdLyEtrkonJUBpPAVPOUANRArqVLNna278LiEy8ucecO4H6xJD2Lzbdb7
wFNQ93HfmCTQqsHwNQm9eKJajQmgQy8Ptmdr2hwNCH0URb/4RFmACNl8JrMRlakL
VgTKgLscuriBV++0GLlUP+qrJkobTW12NDo6oBJR1EpD+ql/X2VlNDBaYNmJJoOV
3jZJ/vq1Q5Qi/C/fbWKH+rdQi3+yce8hMxdMbA8sjQ/lXtLO0I2abE3toHa/pbJX
B2dSmJCcL1KeddMKCXc1t5NCvwSwHhTknuAwVxK1glGszmX+RQ1Tb6ypkZkerG3b
IDSejnQDVKKP6t+z9Xvfd72SnVyUXW6w+CbHM2sNyZTP2s/pGHrnlZdPrpjTBZwJ
MRZLhEsjdVTTb3wKlXWXQrByPwn2SxuNeZwbzQ7gc7oR3ONalQ6a16R8pWUxrn9P
8p+mcj7FlJNyYBgU9ei6uN39tjFV+TxmLpQVdJjlTb0dQRQur2AGQ/EimNBLnKSo
U5y6/FcFCFRpMTcLtyN5Them3UcVuE0Yj3GUAoLe/Ixto05MuxSkXend+bjGWEQ7
t+vIutbJX2OaZH4BMi4s3znWnY+Q5FduSEaME/KCdqtBMx8eKyKY39tw4ZZcxZGs
PKIwS3mYIGy7QpC3uIMm1IcgGT9nhJWJSyhiMHoik8/Umk2e64xRo7BXhj8P76ZA
6W0/p6jJKp0S2HYi7JL05PbTet2zZBVfsOomomvELVqnkmr/aefYfRyM35e2v/Ve
NcoC2w0toTq4Jh1w+pWgYtWefs0sMmOrZHzOaUp7VPavNsFnJNNwW8+SCphTcY7A
S77nwsHzomnTy67eZbX+8Q+9PKtsUl1pwFeDdEQ+3GvZgDXumXU7aesLqH8JTveM
PDsfiUyVHc7vGpPV8l1PukGhRQQE9EiPdP9EStZ1u1VBXKMxZjUkyGY2EQto46mm
mecreouSE3FLmoa2rQsxRpPBB1jYEXqvC+jJZiev3NmETvT9/hpH132RPWIarxU5
NX8uOkajwZY1easumAbfNbNLTHVE96x8qRI4OE0TdHD073Dh5Zn+qRoY+CJbzSY8
gib7Wb8KhmRIKdkucYvuB75qrZgfTImpO6rE1jbpbSfvgWGT74Ye1ayAObRpJJxK
6rkpoi3TTjqRaWZpAwcc2vOV1GOGcP6sjgHxohIXPTrVI8prVS+o1ccQP9J8qq55
zNB4FWfQv26z0RW+GP64u/d8BwjFmmblS86dgOHvXS3MrCe5/4mws0IlFWYLf7uE
qRksAikdmW+YR3U5+h0C15eXxK//5uwHruvGcWcRHfEIPTFFf2/nYh3WCP6RQKjW
Qj/Ba6KQ1f8meQHvdd0ZeQTEUMnp6zPUiYEsuwBxYkLO9MDQ9PTTO0zF8oMRbYLP
7a8SYl1NFLpjogC51YWxIkCXERVymH3WsZZgvWVh3SdVmuiJmVxMjuMiUTh/AOqe
6A5udd79IsBe24W64JhFaIKdjaMxFqFNd/SMkjgXiFl3+uw5RpXMCuNBmwC4jdJO
Ee0ZpbuuuUYYqdRl4DP4hZBD5isi8JgZtinmAqEPkQ87+o4+We2JOwsO+UJJzV9V
fGd5Rtx0W8bn3BSBC3rl2czsJIxAQQy+xUAvuLtqaopbqf9Cer1uWEpl1F/Ld+5O
x9Nl1mPmh0ItAadQakaTEYsPwT9MCC6Sj+4RCCs3gndz2bP1LLQzK4G6fdmw95s/
jI/x96vGpdUcP11wHDVpANWGi+M8xR/YeUZgj0YE57apQH+Uir439ZZX2RUDnJ0A
a9jXkosQYYHdlrlAk3vzuPsloFPSJRufdF13ySbSn5Wjra1y4CgAfgqE7fc+ewl3
FG/fB16QGsf5tLHODPlk8oiXRSNIyfj0VF0LSVUXyjV4qcRf6g4nUPoJ8Wwj7KZr
LVL4wryZuOEaiouRY2TbkDhsIUi+kGnUbpWd+BcFnuIMA9lRqwzrJ1RWUSirhDkj
qvKhQqOC8TcxuhNP1nyXS57KwJ8sqPlk2DLWPZelD1wOBhmdHODYOVa9X7d1qx60
JwkwrKrmqp+ugOVox1NVu+cnXgr+9i0FmSffE7nbPJah6p5Uql6ZSKDmGCoJpaKk
dLH7th9RcN/p3e5UFvRgFZxJwMwpTIZCuneMsWKPPZ7tScGX3dl6M2Jx0umcFPEy
FPPHPr/SC0UkYuQOJqwfkwA5Vj0HdDciHfInWn40z8CniqfwgDu79hzh0HzKtP8H
UVAtGhRDI/ePoit5PH9kL6v0fqaU4xW2p1yOgSW3IV2dSA2ZqBvzTVE0kBKHorci
XguMEkdgJg6JFbXRFnMwnqA5sIojQMhJa1f7X+zQn9gLuQXiiRTJjOgzFa6jdlis
fuolLUbrxKQgC6bbavdbPyUlCLe5GF5aazStvvqpcilxbWZJXXoucCmVecWMfLJC
mVgepppDscCvlCh0ofmcHa3ifjD6YePlwDQAqgUCi6HKsaLuvqNgIui4GBb328FE
dqQ5KbH1IwmDIdCCkELgEktGo19abUI1Wl2SGqxpsS6qQk4USqngrJlRxHVRjWTU
NHYGG36qPv8UmQmtxONMqOJZpUy44H+SzFI6qTgE0bSBTA9sFHj1SXXY99EMhRCV
Op5Blw72kWyK465bSb944LvWZz458gs1QRp0ncyhfninhU3EBN/iMKA42G735P49
KgpZs+8O5cMsISLw/u4oL+cJi6AjyrI00KKbtID8VQWjNnFmdZ4YrCTwB2+tNGmF
hjzVafq6Hm7BuDzZj9AyBivxJ3Zdm0ia9guRHpq/r1uZOEVO1BNmR5mn6stIrNEL
M46GhqrhpUo0fmBK53srHy3AF9AYyGRmiSiwDY+ZnCFh8MCAdxF6BljyufFfB22p
7e30E7ilFDrJPgtdXyiH1rUE5SWgl0sqckxApDyOVMuf93c1dIdCu2lJaXvZzFIY
SrWem4V5gAkdT+SxmDriOFP2bUEuv/q9Se+/Z4AQELXWiUU1hPeEnHJkzG5ISRE9
m/icIu4SQ1A92DOC0wtAxTcZIBPVonPUquLGO5es82nvjI5FMnJ1Fz9dFIkhUlL1
LrTVOMAMOjmSCwkmgTuOCpMY1zfflIPH4k4NHBS0jemkEMKHZ9wz4D39my/Ryb61
wlMFiQvc602ugeu3pFvSFPCUEfUSKbQBZ611IQNSW3hx07Rs6gu8u/ZCD8A6rPm6
tJLKlJQGYl/oEz0g2188Hpa7b1AUFWNMzwwbMtoe4DY2+x/v3ZK/8i16iE0E8rs8
8QwP3Wy1wpIiUZUNoxm0b5Czx0NXEDQ0mYU7+0GOQLLCXjuy8S3EQmsMghbTOETP
FcIn7sGKsbLTFkDYDIgiAV9xe0ufBeVChIm1e7i7qLfWfFfym2eNeuoaplUOHWKC
Rhu8wgqOoXyTbmtmEJow1P2HEbf5w7TSWaCx11hn95QG4BmLbzIOmIOSKQ/zd65F
eXkLepft0xAZlEJyd9YWJCayaRHuaNYjoA9Hz6dwim6TXOlWh+5D72q+6kboszqK
GaT+uSqtS/3S7d8IJBDbQKXDMAPg7AVZ/gC6gTdc8EZ98xakvwY5wYy4bjEascaH
y0qLn8gKgLv4zh/ykwhWNBpE5BG+W34nDgbU0EoX2mcrWAo1+MetAlympNU1hY8x
T+7J7jYdKIp8QThWBaPBz4IbWgz3GErLVDcUXASG8hOAkf0mUtq1ibE6+ZaxklMY
Lu3XfGL9DppYPVJ5WqtYca+p1mpI7Negmj0+k7mQATrIWzGG4YvBx0Jow9Xx81zA
3aHo6p7TjRsIzQEkIf4EhCbla6RE4NVGNq2IO5IeCECKcbeDXwHCF3lQsiNHdC8x
XmqbYzgloQROtMG6DWFMBM86xbtV5CC9BG7Ao/VRL0K0EKt/VgKQelAhPN7JpWv8
92yuiRLuC5kj8694xYSARWTYzRooENOHBZy2qjmvHDMTPfbt23ej5Un82+Zp6Vcg
FGGgfJF6PrMDF1Qb8C+1xNQpl6MqECeLEyhNNiXlsakWwNx0aTmcvHL1uyU4o9fM
Bvs1znC59q9Ql/aGPSAYHnCVFdy7ZHDFRHhHJuwVN7YFhOAvB65YhBd1kmH4b5PK
ZrtfmtNz4T4kX0LJOnj3T/YXo14+KoX3ZX1gh0YR0Zby8vn6motvzUD7RoK1qpat
EfG4SltI2YJb0c4UXsU4ZXV7hbs2kko+7Lf1+gQ1LScLphHmZxFiDBz4gwPdLQDq
zuS5tDEChnCkknW/Ghj91TR6gfbh7GL4dOZwBCdmJ8MKhIGjs1aqucdl7ncl8Hco
lrq8GcKTiN5R+oer+bhk/jj3HLAfL8m4cvRs/Y47WlK404T956fI9l0/f6K7t/Jd
/4fc2nrdyk5+tKkWu74hX+YqZKg/gzBWwixQAFRdr43+EmO//cC/yt/AcWIPVSjh
tjFuI8nTl/7J6pOZewWhnzR7/R2XpHeYPPaApRIWNvLEGM4JK4nnOHZo5k4JxeM6
0GKZAmH88dV83GzVMVyX5pbQPuDMEW7w8STC08jaMidshIoIgxe/e5xCnVAx1Y2v
VlpOtgjiwcBuSgUSpF5u+gHjzPXK6aKUTMvhgRJUbTue2by6dRoVQLynhYkweQCL
f/TamER/tbUAXFhl7zzzak3VzQVAc7IuOHfsTFWjf7DU2Sa4E9xZtukSkiZPdv1l
eP9cJG7Kl3rBGorsb5SArFmTO+UxDRRcf2waFmo77TQe4CQ/VsQeDDmo/QZ6q5AQ
Q4QJpRtQPBiGB6zvG8pKziMYA7Ax0YEBMNl58gEqB56PTDHujWSOYm8FFdqha020
/xfjDoc1bSF1l+S5DkmRMorXtjcYYM9Zy/uhcFe71K8CHP/Rv8JzJjhLCYmwL0IY
tERkZHVErn3XHVLLZ2nuw3GQyPF5ZC0/IQ4Oe43DDKqH6iJWvA+PaJl/03wt4C4m
CxeFCiMigGwTVWMh+iRM7GA9Vp355Qn+lGK/PRtUJD5sOMyGgdwhwy8U6sQhbnBg
h3uv4Zo+7lsijkmnvpmF15WfBe3E2KJITzx+0vNRYlXkP9a4C3lunF3BCNc/4bBm
vtsdvZLXwDPrPVHSxET4XHTWsv5IaDLyOzMu+KJB3eZZKGx46EEHwzJTP3M3BacM
7zARaKYolW46QkvhRDNT/UBWwWEPfiDmEA3VowgoEVS/q3jHj0LOLcUKpWu+8BZw
4BDIwolw9bdJuB4IIZCbhDriJgvbk75MacOSSRfEgP3fSVlNN1RGItUejSUxwLHV
bb6QOgL7xMgIz7Io+GqhjmQ5X+X6ZOW3uDpdmps+sRvbk3rsGtSLl28BTVzJnO87
LsKvxvrSV1wjvjg4hQAPpXdHbJe+wBTL2MOfhjrVmRjugDrMXNn1cgiUlG3+bugp
cP8HbXFFE9qPlVnDYCpFnC03dLoUF9aJkoBhgoR7o92Fi0PeZ3yWELmoDbzw9lZE
2Gh2OQVCrhl1b+AJL1pXKhqEyh8H0PM1HWJmJxPXMQf7pNjHl+JZMB0pBndk4MVN
0JQ8aFqZ8/z4ahumzhCbogbHJLt+rQYpgI2Pyf+LJ3WR6gE+D1Bh+FHM2Pz7fhKi
k1vF8mgXTLDPNlgG7liWtwtI2lflLHhf0wkfbQzUI/7pQYKokt2eiWj9sS/6nJFk
VC2fWEvcmsy2OPcND5HLuTre0MMuhVRYfU3oZYSHqXzX5/le23J9wn5/qYBswAlh
uSrkuYV20xJi7m5M3x7O/Yd6TrK7FhNK7bzCdZ5MG0SlL/LVLtpwA1CCfBV0gfbU
5orYiFmkm5Iql+Id0lcbt2TjKblH2lnL6Rh0FQpLpxlg0GT+YuW9iaEij2b4HfO7
vzd4YAqtZ5IocI3ZEIliE3ehBtimLaluR5+yI41+9C10FzmtZQsXInB4EpAsTtZ7
xPPUR8nujE6Dp25knVS8SbywcFcswQHmQ+frKdMtUkr6T2vpSEmhON3+9q4PmX5U
lMGg1yiikxRFodxlmzRWm5H8T/QnHDNUh4wqAE66CWbJTBaa1MVm7M0kR1B9AG+E
9ZE3D8XXo8jswePswVbAW+AkW2GHVgH0NO4BJ2pUg1f4TPRVYQ17BiufP2PrHE0v
Yz4mOb5KDlj/PCYkZ4vlkdFbD9u1nOm8tQDIjJJbMzmNpnbCExpIGkGp1jpW3Wii
7SV6Wq45FXHzD5lUzDh5wO57QzwivvXMgrPqJIOV0kHaLrXmSuM5wkXQMDVfhDVf
CvNe3BECywO5d+90CX3qXly2RKFyUZQfa+qoqhvtQ/1UhJchWE2y9BL0nr0/zZnB
h8I3MZE5XXvsYiWAUlVsSs9T/5Mq835xXC6CEGEAxeAIH55KZ1pm9LEpi8X+eRRY
N+wXnSytleu8iLztydbijam/zawJT3mLSfBAqeK7dO+q34fX5QTPJ01BE6rPPkDg
4dUNh3RXMR4mhSIhKibEzg9naHIUqJI+GGdvMLNP22vB2bENTeqeTlsfLE8EReck
P4bq2hn5D3fEwyah8kNQpr5J/pWxIm1gkf1Lpze6KEZiWHQazFo1XXqBwI//XAWf
bUEee0jsIenMm1rZStBOlFX8Wv22uVYXH2nKh1gDPt6e5kckgfAqOXghEUtKt/Cr
U8ZFlFW5UNMHu05DYqBufqkjGiU/9ZpVIRQOIhJsv+L46HErvzbIY7tpDLsvqUbh
6kJC3oaFeBANCkgsSsbU48Vvqh1vSAv7oJ3YpZDwd8SpjUOYVR/nxR7+o2T1jLxk
nwjgy4D8RjxWwtWnLjKWIrKmr5WdNz3o3T0MOdgE+L0e4wSBHhibW0YDslB0rLOa
m1+18xFeSgkYaz5Eo6c2ENwpe6fl7m9QzktBMQkNY7CRpATdGGMLpD7ENRlpY77k
/7R2e3GHeZhWZOQSDAR/qz2qE8lN8DhdUGplHm/S1ckBy1OHRcQDg0wP5j80W1pH
qlgxC1LYNCrAAhaOfJG0BvEcPqCm/+mcL70Y1DqRuIlxqfSAW8hrZ/i5jvhY5oy0
Hghs15rIq8o1ZZp6GKxPcxQN7x2vra8Yk8aZXZl3pkwnv6WHocBF/ULWK7mVqVnm
G805UD29iw5WKwu0H2/q+DQ/bftTCXRHco5IkHI8m1/Bd6rbXznXmrOrdMp4Fh4S
EJ1e33A63Z2kWMu7YJxgHhCkzeZxiVTXXnFIPhFnWNMNMDeNzST8AJJtou2UIfcE
fTXoC0z9bG/Zcja/PIWh5T2BY1TZBbJDtGYgb00YSwXBRHR7rBmWVuHPdgVcA3w5
Rh41l8ir6Cc7QAYRv+NcT/RJssoJYFbctd1Tj9t3ML0bXUKj75D/Zpv3JJ2eCuI5
k7u/sjt9ro5aPefzMwS+TbQR1LMAJ6q3xFzCZCOpWsvumK9/FPKhH5vTiWwm80MQ
0DxG3ztMLlR06YVDQNV4YnMiMOnOOtvTaSCGc+214rL7aJ4j5UM9mMznzWin8Ndf
wyLKHhuIjxGljckfLOiJcMH8MfrTY4MtSxhU24P5b8+/GSK8rPNYXBqMvezPoHGp
haefAnCX0d9QC42KPX260FQ/ZoYejRN840qhjpp+CnCov6WZ5tKZXsgJjVt1MzuB
MPwzOz2w++dwacm6kKa1pSKWemC20gYHvGWVZ2BJRVnBlc3KIOde92T76E2WnQuS
gx5jTL7cicR8IDVzW3TUtlEdnqzlGpCdivm9VSLoQ5IhGSU7+nraijEO9E/Xtr6Q
038Hwr6ERcq2Wi9SgWXdVbWKbEvh8xTjc4ZKB+qkwdvZ6mmJrj14cqRCHuFiMhN9
XZi+migRZSfcJsdCi4FRZkNy1U4zlen62K3V9uP1Tl2nRL/QzpFmK0dNEKIlxEth
uajvFDsY5hqaFX7RYJT5XDz0OXdVGtOTMfkO/TxH+eGTD2N2Y1JHRO6S0N+bvAE7
1VfOn+D67usG6uuP3u3YONAC23F2IMthVPewy6Bipsqn6ohXDDGdoZ5CxUuhsWOk
p011tfajFYrZ3L03fh08Fu935/nuI8Gqc78ewfdiroKfMYwrSU9TvkAsChiACmsX
ldRApqfwzxO1KvqvBkYPrsi1q6E8aQU8eyXJAVCKiHuNHgd2g5Y/JXPWAxeqtIq6
VGTF3u7aDiErsNrxbCLc2I8T3yQOR/bqAN5XiQnkQFtqNN0CdPDBGZwYCP2o584h
4/lXe1Wx4IzemdKzxYjvP17hN3EfidFYG4mrnbPw4G38o49hqGspCsTtGib92I+j
OzL2LCpzJYfe5SJAnewdwU4/vSeuc2tpBwTPQGPz8aSPG3fXNBaT0lXSFixvdxX6
MA0QC2aRLEsE2iWb+2PKiRMSdwiaCnfM7a27E7Hlrlfg8SprEh5ZQlPI+6BZuYgj
tF5X2Y2ktQgI6i3ddY96eZDkzck6VDdASL2SyWTKiwriyUFwvCsJERaXjk+yMjOT
2D8YkP+dibzsk2WRFmjuAAHvQodCXlQKW3zOTvErsEfgL4ELx4czuVXlqZtxgglC
NHgZW0bH0Pa/IsqbPKxw6sPpbMl3QHSPvWIreQJKBKjcLw3NUWrKyvXWGUiEmPdp
zGrzNqDvkqUO5hetLg0mAF3cieb5Qn23k7Qc0ZGbEk1O9gnox0pNCUhzqMquB99X
2aG+Ou9MmdmX7skPl4HBeil/gnM1ydPchZRxd4UNi+ikrZQGNlHWrEn5oFK/54ga
TCwpN7pmB0MNAI0aIusgzoZod6ndh8AHBKICDKu5tvy+OSUn/VgoDFK0mcghSjIP
JF+nN2yX/g+eEOo62+A9xX7KDJtLO9KNf3URL2Gz+m38MqitccJfhZSaS7+rAhei
hS8Q2cOiOhFN0bJjnsZ6xJJswtCLqgFVpvvsAoRYMtq9p6IP8+g1AeVIm0BBsk+L
4C394+/vBxx1BW49MrapQw4sUwSJpFqSTBg1G1r9VUgwf+zRPm62lmpZxqtPADrq
jstGLnCd7Ktms6lUqJEQFiW1+PZEyFTLOVK5OCMdU57MVxfwaobfmyhLxfuWAE+K
4UfwnAmKBue1WQUpqxIq2PD4dLGjrqbwR4IdSZz7SzYUIdbA7FcP7R1eILYd+7qY
vsRaMl9c3fuBd1FrmdsEBvqoU0PYWP1uF4t6IDFBniLAEJiR7nbCoy4Ddfb+YnKm
QNWvFVr0ORplOQSeCJn2E7eZoe8CmoCSMBuvRpTOKgXjL7mgo45LGetSekfoGb9H
jp+XY9iXsM7jKeU7ABjQuyM6fCkppp3AnLEQ1VUKBedwGNyGkljpkjRMlr1XV1n8
GwGQLcLGTNmSWDpr9oQfgTVLbO8jxBwdiFIgtyiBmSrzUevzcls0VLcFpvvs4/RP
h8dAS+XMi1PPXILru4JEIsDcbkS9kwPHtViyT3H7kFR5a+IWDcnyI/pYuh1Lajru
we1ASfW4zn5FA4yXmjj+NlzY9/6HYIEr2WcjoP2jNKqX76c3Z1inecKb84T6EkvR
iur4dYv4uEJSBEzbmFmx0Y54cUJYHWrPOCD2sIY8etRrue8xiauObcPaVFkNBoUj
asQ7gdayWW8YCfATa+W2ORDWDyIe9OnZKhBJgVZUQQSsPmhid+Ln+moDykaIi812
OLa5g+0lmG5GAzge7e34IeZ0VoKlYcnJX/2lnhYsZMmq3ncaz2JytRVIm2XWI51E
WdCnL3F0RfKWT+TWEXqEZj9V5OvPIj3HhuNcqDvJ62GHybaiVLOkQexsCtp45Oqp
eVik08uZIs9R3OL5XemDXwLp/L96hfAUUW1apeJrGR5BTOgoQqb/6XQHdo/2X+HD
E3lSP5FDE5JwBdbTDRzFKZMOyndwEGE0dxJTI+eDhNr4jM4Op/Je8IxDtRjzVHi1
fzEwaFsRMY7IXz/vaVs0rA==
`protect end_protected