`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
ddtXksX2+yylW5zu6QL2Lhnb2d1sD00763mmSITNX595NcHTEkwn0zB1Dry37fOW
FufOhVzEJp80NC5qZ/+F0Vk7Ik02dIR0elf3clrjeJRK85K4e3Hoo4xn7YbFUIms
l/8VZSb14+JVGURjfswrIyCUotIzlzVYZ6gzoZwDXIi5gQIBf/gI+KxNXPaKV+PQ
Ufys/12rjO6aI/pPlqSm0hCvftmBcnezN2hk1UeXgOIuKZnogjOsf0iJVX2aOOWE
6pD/psybjbnsNB6kH5uFTA5frkzIzkzl5d9+YDm9OyC+k84E83I/7/j+rk4L2dah
QJOvksSIzN867/4Qt8qYTQ==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="MvBXkzurAa5VTw+1JJ70nePUfoQXBvZOku/SMmg4TwQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
oRtzZL4VJ4iwysPsC8SXYCzXS8Fw2gtZTOskLcDV+1B9Nzn1zTyNtlo6lNICRmmK
ZRVu2BmCc2G+fmzynYlNTnSa7C0Cuel6FYpxCBlOuk3OF2tzAmLAuDyOH3Z1Yjzk
a0aHuoCdIRKv7BrZCdALt03JeUmXKPdOmIlkVGFl8yw=
`protect rights_digest_method = "sha256"
`protect end_toolblock="Jn9CQpRhJt4rnzZPRk+dOpzAubz7omckX1MrFd4p81o="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 31776 )
`protect data_block
gD6l00tciPUa6pDNTk/+t0OO0nC/UTtBwLB41d4inuAUA3i/ALrNyoJVcBnAmEQW
ptbcNp5fxEUJjnOxnedyZEuEBxWRieZFQnkRdF269oMzOOiYTKBE/TxysmcEF8lX
6cRFCJrnjgkJxIpHLdg4S8bkA9UQkTqYChmK4NVAhcrMlX34wOub7HlgAmbKEWzn
4ScFF85quglcIHqvIV7epYgr9oCrw5J/dlNq1m+IFJBgDChTtxDVAr3puddGb9zk
w6i3Wc4tkbrY8XWf3vx8v6KWwPHa1Sjv5gpp9QHURRASPdhCBD83veMgDs1Gzw5r
1yXC24nkJ3PMo26mu7YZyMtQeXDoGw7awZCcKHFKHW6XoQbS2yDYrcQp72lwb8xj
EyUWZgjD0uOk0Sogow/UwNa9qAPj5tZpjdMQlawEa0nz0WZqtv67mqfjBoXcRBT0
V5QrbufG0t4XMjyvcDOTKvkdSRmeeioQpxq6xZrrCJSjMCPlVRkcCnhadnkdN5i1
JQ+kAlYZrIEF1fL7OvWBqS5qpg4drEgCKFUU37ZNI+cqKtE8Fh4HT+Q6gvWVjEKY
2MXJfboAtnvEq192UAxy4u8lvRxjIJsxiujb8OGquuAhcrSNaZet8DjnkAjXuYM9
eshPzt6oZITAh7RWVoCQgiNo9tM+w0ukfjcCpA2TkmnsBcYqL/zyZhUFGvs4B/84
7dYOt5R5m9fDO2GKNB0LCICnvw76t1Xu7SxchIqIump6DZpqkgxzh3KkxuznZpvg
K3RggtCKf1tFZ9kkMm8TvpYjJr1vzEkFUc/OhIcLie87NPmnX8T+szJXPWgIzKa8
BX4LMiKhSUee6NkVoIaORlMBDDdCLIffI9F5nTO7bm68ecjGSyRmBaQQWQljnl+G
twd4HXHrsH3SkdT/6tbvs5SKDr+wT6QaOdaig4AeG15//5bSNU6d0D6KHqRdZJm1
T2u4RXV1+/cfdWc7eA/d2ZCoBHQHR/poRt8Dj+Ky0LJF1FUPVbSyZny8UpTqjsnJ
2S1HF7giLC8QY2zy10J1nZ5XTjrAvYpsBBUGokbbg+52toOKtVEGc135suCFv4IS
ndRtKAfmDrwWep1bVwZ7TaHQIy6Kc3O4q6NA2tFNedyh569gzIjSxajTGjyuUFTS
k2pb/autS4bAz9p/5MPSh6KwV+w6sSnXV0Wfy5oPLWENsU+O0avVy/cXABDbvwgK
x4n72uYDsvoWpDLXndEVDI/ZmDOsQ3xkZwvFQ1XV+njnkDi85UNwvWXsVt2PiIIt
Fuk3wFlhL3ZWX7iY+W8+bpDqEx9ij1VIj6Y6IOnCC+XUszW1j8Kh7n2t0O+eWKMO
dZgHKZDwsWJCZ/V1hT47Nzu3nj5nI3LfE3RTMVsU2OXJVhxJyl7UWetF631nYBNJ
K/Z+iXAhY/tDLVZjDgLiDIYHMawzlbf1o5GEukYMr+C9zwBW9FN0ZgftMUYfDwRM
DzhEo4K/Jpph4NBtGiH+/eKhuHd36ZQBiO//UBAdj0Iikq+zz7kfruErZJUcG+TD
vvAl5oDl/VUKnLhCItItPKQ8mWKpCmHG6eOYWsWwE/XTPDbvZBL+9lNa5D8JwKPx
5rWJixLRRDkCr1WiXeLMzRtNbWClivRVBnOf5aFB7Cpemo2T/MAw6yFunohH53Qx
ntbdFzWMKcorSNefo4m17jv+t4plapomhM7/+HQ/Fl3XCroYuCU+6W/gFLV4wnF/
en+ziR0Je6vsZFdoZcMFjJzduPm6Pshvkp7Nuv3/EcAgF/BEOTb2n9DVFVGgs1MK
pPm/vg94HQx05PHLMyHWjJ6+wab6dMa9L1bOoDPdWE4a63S/+CK0J+mht9kuYkSU
djmdB663OS/9jykzT8OiyjbUB152g1XNrDQChjGjAJgxoP+X8WFT71h4OgIkZpKA
SwmSOIkmkuaLg8xKSs6h/+PQFXB44y27t99gtg75d/nL31adgut5g6UK3PJogjjf
3xLJHchZYzpVnky4cqoKAFixLzmEQ8nSAMFK/NYSuBgNZBoJS4Ttx/39X5MSFGjT
8N66Bfj8O581XS1WI/tLd1l/Muzuxz4ZXZcPXxtLA+4IdD8bfyEVmiiVNKkdeHA1
XnaOvaPOzl7JrIG4+50pT6tNRlsq0kg1j7jVm2+IIMb7A1roMQOs7hPeitecJZ1G
GvG2gIPOxtHpVlmTnZqYRd2CS8CgYYDGtxtfBICdOO2uoQriAfjG6sAmPmogvRCR
kjxTx9yObVgCMM63rF9HbKZY4zHWMs61NorAKljgMKkr0hWSl60JqqnbhkOf9koB
ku16se8EFRZfOtNh6yMe+HsgyTbzo5vTf4N7tz0SDr7EViq0+VajganIbK2sjVhM
3ZxYFfzsp2LHNYZvH+y61eA9OFdl8Hg5vWiftOXgkTFoOhlEz+bgw0PfGlp2j6gQ
sjTikY8oGCJnTMm82xFCU6RyOgPAdISLifCH3xO6plq71CnvUWmwseTCudrfkzc3
5ZeILM14gaU8wiDVzNmsXsiuEAiac2uEYLGz3mdUbRzw6/ywmPo21u/q7T19ykJL
DFvD6vUF/95yZTQ6sOVWvULD0QiUaMU0bDoO1alIrrw96WUH/skb59Y4A/W5N3+/
X7FYEew7FllelKwkieMTy85dI76P40VaJgAw56Ek0ViSqfMCenkXRSq4M1RCd//r
xIp9QyPFp1d3T61VqTHcXnTTlO4fxYl5aJygyQ9egrmkKUsiaTzL5wh+E+2N+yl2
e+Mb6SjEvBXkHG/pWz4LjjKCzMHOrHQrMuUb+fL3pxL4e+PsR0n7rIGyuLTcMjoV
H5DXm7hMOyRekfdEdo3/QG4oE8FzeapF9R+EByn3bywMKuvmDsZmwFOuodNyzP0c
yEf8C8agmU5PJAhxNaB+Dpx++iCxIafby9ljFRC2tsXCLZmmZo0JmCKNcgyBJTgv
d3wlOHgjoKGlVBSVSkMSthurKzP6BqTY+MM3xknQEFZrKQvcsatM+tm4t2kplFPu
4c2faylhzJuVTrVxhjBH0/xujiWKtdxXz7thiJ3ORbyyg+ySeqngyqJsZNaJ1aGD
EfGuBJvHfsMdlVucyMAYxuGpgeRdmVi05EX8bqmH3k2lHksFd0OHHE3jqDEgmCb7
HttpFEzmZ67M/4IQXxbitfUxgFn9y/W6cKX4lhnHZLOOPFzzSBTgtmyiFlNGxcUA
xdiAhIXa8w99bu4EqmQ7HAGhKzJmosILKPCeBwfhDnMCIMpxLeVKLoq+1ajfhGUN
yqARUngq69UW+710jAUzS/v0k6QqTHfcbFq3AIwLWd4PIzMYVkIZUxfZ5wC/ZAGF
Vfy/YFjcPRBOlEPWV9bzG6KfC8tCq9SDDZMhC/GNAuJniwPs0xM7lLsWbcm95BG+
LIxaUk6Sz+GNK82Xs/EGzlcDvF7QAdSZUfjR31wg8fgjppYjhIgXo0J7IZiDLq/0
3J+loTNRNOh8W6ksUisrGq2CT585I+yU1iAte28BqjbryBfDKOzBTQPfC0V6YQQ8
WzKii0Je4U6nLt11P+CLMzLdWlkbmu8gK5vNNe9otnQPz4Jl2xhBPiv6Qc9eX4as
xEXVIeNwJnARQwX5L0+CgzaQTBYh9vEvTbuJL3BH/JggDJ3OMDKZ/e/02hhPFqeU
cte6FztZ1QMWZuq0gPgOnBCqQCehuQLyEyMPJv8uhnWsklJ77dutrjsVIjbyaKzl
H78cAAMrRZcgDKvZtdGCcSWHd63uNc3V9khtakOPrHAqcrakQZ8/GJ4x9RprJXzr
kuRaBOslLOz4mMWA+CPpCZ2OWF1YpXXu/Ylfr2X+z1q0Eq+EATS4B+Ih2jm5MX+s
W312XNE0e/D+DE169a4DF5DblhtbZDl1I2XaNu9MkVGjmtfQHIszZwi5Lr6N+S+p
iDRivQbpnV8ipkve1xASwUEJcNLwcORq6iF1AuD/z1bGa4KHs98fEeLBSMpO1+xP
ahpXhpujj8Ddt8uIpcyudKrbknGDE3IrT9WnczyT4sGGJEb8BgRmyi+d+MqA5bn1
bsEvKfmMggehkraap5UR6IKmQBdDXybuwp/zGHL3ynuxLheUhxN35CgA5rglK/JE
cft/9nn6YZgFmQ/eyI5YFvZeWO4ouxOk0VOIz0B2y7UNBb7hOFjF7g3gE/dgUeHh
rF5A6dkIsLK02SP99bybLlypqEMmYCHvyyNN2CBLu7Ryer0Ee9/Ss0Yj0LC2MwKE
YhTU7ZuHixSySCZFovORpUYhrjgxM/KXRujnRZR9ix2+eK8IUrAI9X/4Bf9ee0Ff
s2hs9Hn/ArGsp45h4edJoY3pQUwOyObfEWDKcUVCO/SzJbi9hK0ycG6GZHDradhT
Iq1ZLQNGpMJDh1R4dgSgTct2ObgT0/mayvDetSbUT4g/C/n+DYrG6YrVTCM/DvSq
cpBh5Gg4MmZ2vr0HeORxEZHfkbTok32MD2Hl3lQnsF732bAMCNfJGFd2NA/1Ffka
fP64PY5bWcWDtmbH0ehlVJ6dIJNKDlPMoyvubajN8OnyrQOkNvUMGOVgZemliyhN
o3eNmxM/gUwlW4eRVIBSMsU4NmMlp4flqjeljEQpJKUVjkjKVe68SaWqy4fLCKLq
e4Zw2hzCykvudtXk9317ENLP8rnNwowJbl9sqGWzy6hAxBPEJAlYwTttZsFbbtcn
rzk9c3okf1bnRBBEpTfNTf9eN9T2/RcMY7tszahCTfpyqVv2H0UXvmihruWH3CBX
CS6/r7nJYadDM7BPHUCFVw4T0Lvu217Md5sJSoHEKdah2zrPqnOd99XznWVkM1YP
QaWIsttMO56Br3GgB7wAYcWZBmWUzlR4tm+2NKhtQ7vr+++BemOsxvqQ9/TpuUe/
9AG2kpZrg/hBn72fAmdfftg15h595jXCifhajLzENRkrzZhWpV0zcNtqXP57K8cJ
zgVrh638Lznz11wLVxvU5IRJZ+IkEF3vsmrmW6SpO9ldFAUYb24OW4KtWjuzjAHy
SrCphAfBDlnHVdJZ+9jwvTnQDcpCkbhW8RVnwiSTMDCea5ZX+NqdLT6e21a88Nx8
MmBbHZa6KtfxM2WDMYPvB5kgcSbs62zxZZ252NjP08PBCwmwJxUzHIm/EaYDVIaq
A1QCQRlNmlztGf2joHHIn8eSYPXz4aYs474bVEG3p8M7t5zl7cCJ+Xrb7ry/WeDO
LZgmhgJQS+L4L+9YKG0h3p6fNjxyTBVGxWDnp7qefGP27tW40fAA/CqI/yd3zM8D
n4y5IXSXBcY/OHmNn85+d71pTXlv5HiHL6nUhUaiAhEtN/43lvAJWjXuq12xEmhE
+5BHM2WnGE19uh0VceuSnMckOpIPYiXB8lio+8xT4YHpMMop6oIiE+OKebQy1qJ7
bO/0F7n0wlS7Yq5oHTTFknpia1ZQg9CZ4nW+iU7MhHVFfEndIHMp2WMoun49epax
pBhBzSR7KraGnAgGdRB73JVvMLYJZuIPJK9H3E7c+PT/NobQBQDWQ/he4dKQh7OP
be1+lYOfunf5k9Cp83WJxqBjkK+xzv5usKfZBG58/Zgjbu75D+MugphrxxjrZwm5
wmte9oiuWuJC54mNjbItF4Rr07wwQEZJyvSoI5/N+HbwI71wl9fmY3/nlWeRkwJ8
lWKZP9wMXuUxOz8r9B7P2ucxusICrIPFEORh0pMabO6EXLPXI9jkthEmjQ1yvcj2
k2ziUDAaFTykITyiCWogxNmoeYOq8ijspQRlAs0sbNuuobe8JvdZolOlVvdVh77D
YFYqkGS7KNHHbOiGXunKeFU78NXKe+cm2kClUVx/cGV8asJbMDcB9HJ0CoM0nKv5
aB57z98HEYfi34tSwzaJbCV21QV9czj6K6m5qtf7qNKp02rt5hJcc/f0s6SvYn4c
mK8WQCLvUrxhldog3nL2j7vQ10i8PecyBIIWp12cOuw0zVsqhOQxn4f6aTM5HrrN
QvjFgwPmWdfpPT6tFXI2aXyGgUqvZSIjDgiVN3gdOLcqjLOswjv9EtHOyQEBLZ9a
TFVjIrkuNJxDvQ6zJzHoHCrxHRAzYIRBd+gGAZonBYNokecF9xyhAQku/GRNBZiT
JjQIPIKnO5Lxq/A+gsvzdAM4GbhVjLzBEdaZLSkiyj34hxg0rH0tkpcBeUZLCmpA
ggYv0H9L2tsxYyXPDJbVcRn9HKZOiUurSEqMQ0ErSq3YoYtfbaPQe1QXDA7ba/K5
yHRv50U0CLh/untgHWYlCXKjTbHpWVXNKpCDVytW5JAH/SoBMKmzF3deF0fqOaSA
BA/2gl74jxV4sUIGu1HlngN7FKUHyavIKgv30E9GAO9KMbM12NQCeIu4EcH5i+Y1
y5lyKPBscI5qkmQ2k87pgFzfKLtcMhzJnHV61+FXMj1cCo3WCt2avisW0dQUEV9k
R/QrFJWQtK5r/xjoVY+ekq9AvE1sKkKsGZLqGwDOcBb9Mt1eFem8Zl0xsLQgwdZZ
r4qOVDLNT91b3h5gMUkgldE12ajpnu4v99QVInXio7h8eENzWR1Id1+0OCBEdXYH
VOFDGItcCS05x38urVu1mLGwUs3Inh0kMc17BZJ5359EPKMcMkc0QsCcMJLNaSKk
IRNWzuXhxj2VZpCZzBNlDEvo0hbP+qpWr1/79NdfaI5I+HAIdrI03em22U6ERj8b
VyuW64Ewx6JtrwSlycCx+hwuZnizgGQJK6BvSjVzgu0pO0diTpuUYhsK1YR0dkf7
iKc+fHp/i/BxD+fgZOcC2+u3WeFk8eY2nQVYvA018t+YTcZyovQAg7bya5kBFQ/C
O5M79YUyRrZig/P4fEy9peT8aoL4ZYVXWm212kcO7ArOeiRtmoIHRIMFFr3IHkZd
Gg/B9AuVb3YEKctEVC8KT2o0CdMvujh+iiS4aZ5rXacMoK/b8ZThMOC1/bn5v+ga
qJzmrNMapf1GKKPLTuqquV2E3Qyffr64kShZTtExEL9IM7MPpCR6NgKGHwTUoyDI
ze8ke3kx64v6SAWdcNoUNRaQOiF/jEFCJkVCaxv6HFYvRqoA1lT4/NcJ2vauaCl1
1YgeJpPyIt5kjUQmgHRshq/iKhZFckBsMlaRK5MJrGTREQCSxMhknVaBZJj5pyRy
yScRBKhHxTwD61S6JAVCfezTBrwU8LQgS99yopiBNL7k6Y4mCEIMg8Uv+UAzNQgd
3ZL13VDbBpnCX52UntnFFY5C9lOMUVukW5nezG7f1YJEWW2Qt1pf0NoKMJDZDJMr
VXdi96aZq40B4AUeG9pf+8ySuMh5GnVe8Sby2lirq8WiohIOmfqdQ5miezwgiSun
BaQJ6+jeFbIlx4DtFbH6zWlBEAajikMAkPUOHozUCeeklCX18Q8yIeeyM+AKRtu+
MpBJsHtn8gjNJUyCTLlfzA04WOii2XFb0svFyRbGppt1u09dUC7oa2qk18iLM3qW
6QSZK/2bC4KbmP9fqhInnm47P2I18j4wX15qjRraxHg3y45pixlwS+wflFdl8Z1I
o53GG+VJVK4/spm0JBwWmtD8uiSaN2XrU0KQYz/6qdo/k/B+CCZzgJI5psL549af
Ooit7vU5oKQ7UJ9xr7+eQid3/NucAUlXYL8nIrPdNSsSGT0BgGAP6sT32gYJaS/3
tCFjFY08ZncsjPIvyAIXVxf7TAKabtqcphu7ZlhZZ3iySoPiZqkaIsLpLu4Uugu3
uWDXm9L6/hocQ7o0EWuvG3yIxrQN5B2+LQDDCPkf/4NARgM7esJsyXuMm/Fl7L26
70Ioh8/6Os9ISvHyOwvayrqo8dvMr1Jt0JvYbZpNdN264CBH/FCvK/WbySSImGIZ
GNg6Dyq9B+M40V4MaOPlo79lDfHAjx0UJilUbEkSqiVJu7Ca1nZhy4X5ZGq9BcZs
i2RkiSL8WpNzG9/vBsINpRXpKAoighquhJhv75PqHBz81y/QN75yYcyZD010PRfE
KDaycovLs/QOw8M+eMX4j1/PL0YEeAS4SePfgeymjHr1DW3t9c9Wt7F+odhVo7HW
YzXJ5OYbqxSfANrt07MUaiJv3VXYw9LxqDwlY/gIFC5YExzCABrJR/n6Sjmn1Gz/
SZ4CwISaYOHM14iHv2QefnJBc0H1eeOpRYTe/Lo9+4UsCjwuojaDR/Ku3pebiBEK
He3YtTO0MXLjGp3AQ8TUefrzx3/aWwym4Cwj3FYIvVKpNSx49vO9vs+Xf5B3QSqX
obl5tD5Si9p2yneMHleYYwTnyBIXheNWQOUJpjnjNvLNyedEHm6TMhkI3c7rEvfl
6WerNtW49tKtQqlL6m7PMWgiGohdpv9Z6w9OPP/lPyG3pP7ZK1SQ2IhGkRt+2Fug
myA9u/T9w6Ro8ebFfJWAJEQZANxvwDRmcky74ggpQN7BpGf//P3qND+QuQiNtZbd
f8Uu240sFvCIed1zyAyClgGWzbQseL17zwEz/Lwb5XFn2hwN+zjmbQe65xkadm7X
TobR/mLQjd0KoALr50AVmIFTeqNSpcCooG2+eH+r4GM30YWKeAThxVkwlhP4eEEp
3UZlDcgf5zdzuPLjGFXoB+1KKdiBjMccU3cLo1ODwTAwwfw6f8Yudtl2FF06TybG
SOvQGzlrGh1x4qJz2k3IH5aO4hXCc6HlGxMBzQQuS1Q2LinF5HVy8HxAqMUJNGoD
rQ6JZxPE1A3PCczILiBdiQan4mGT1KHSDQ302vLk8Rsjoix1wG0nWvDTmVIM9opE
3MFhwbnB5IDVBve0nKeH2W/F9lC2fA5bVeeceTmEUu/xhVnElvDbiZgdfJbh1Pyh
GPVDgMuV/KbMqxBObiKPeGA5Fg+EekaKH9j6WY2Xl2vyyPwYdTZiJ9ph6OZtsy0C
tD1VJJ7xNXzY0VGnvWvETu20Rpkl9w7UDF2FQ8emACCM/KCEFAVfCAfJy/e95hPq
rE3/YEkJO8YVSBEbQiYbNOzjaaVpzgXnFzi7LatKuie7fFCJtmbUoZ/nan737VSF
6LSOGUTPb5ofd1tpPQUxYyyPfpZHN1zvRCZ8VJkvSG5/IF75Cvhpsx/hOX282Fh5
n1rxpVwHdL+PakKx4+AMPA3Jozt2pTvS5ocGN6CwYr+68zhHf5BdntE1/5+yyMJN
s8cPiemAZwciEJzgj37urenxseqS32H39dByis4sVdE/keUQgxWih7ruk8op97Ct
5jRUhH+tIRybAJ1CmfPplwweoo02tM3zl/dpxVq/hdjfiGGrhD8r9GkGQSiBmilr
untkVivixx6HBCpULrVyn4VGWa5DcF8tKa3hkgyHswdeUuuwq7XomBFoXklTewp/
XpiHqfgLr1K5321aG7w1l4GjJPJzbZ1g4UCqyJJuZKJFv7o2i0CwMVGbxdETkUma
1qR6C+6REEg0FywGhda5wx840g6wUCGhj6jnBEKTPC189YGUHtgTrnGWP1Ed9tDc
eLgnBtLthZwVSg/Q0HF9TsrXKEBE7lia2O7EFywRoZVlA0uYKDu401Th5hRehaB3
1AG/wLkxmWwyziKZKr+M8i6NK0q5ISEnZgleaVxofHv8FiqAB9r1qa0qxhrGLyDq
lLsqOkeXPkAebJhhJnuRC5q95dNkrdIylbHVxvQlNxlXFTGXIIxgnMlbNJfHteMF
ozDd/LLDGDkvSEyGH9RiwZJjDN9vnkn+dYsygrhyYpoyTQ30yvfAnm0Q4YBKWHJ8
ig/q9G5bzdhLxNuCimgfzkXPNivsYP8cyhod5MCg87VNvqnIkpTug8RWb9F+g9fK
4tpty9ZV6H74BZjZJmqsZAO8reUVSJenaZUwJaVLBt1ygU2glcHPtl724RWFN1cP
KG63T6ZBYXHrlqh0OaJ2hJ3g42Fh268Kg1VYGvkUOPoJ7Csi7cNUFxs+86eQI2UT
ZWbBi2bm9WEQeMIXfb/HIaGRpRJmZKb93LtOb40yF+V+rClSS9hWFTEdH+McT/6P
5i2uGvlHgY/Hzs5hFlWTCCPTYRrBA3jEjin+R83CheIojjliTkJdoLc/+2ZMQGJB
8JzQettGmqpYXtgsqj4zEqriN2PrJjbMgMGme12Gzx4MomBkMv3u9Nl7eqcTUKWg
+h4DmASIbdfnoYFayDYr4A9INfPgkz6I9vHhuZKmhTbrMGmvCY+pGE0IpGDMC1bR
RWmezPP6XbBY2RUGTZG3FhbDXsvTKJO/d9XBtj/Zx2xiRTCJWsgCoMh0/RLHojR9
QMPq+pPpxf3F/6HTSykdacYiWWbS1M2R2rku50BvtoM1lWCWeJkpnUAHo95gL9S9
AGdLm4C0g2yFgyacWqBCXmez0hLs2BQkOoFvTKIMr4An0tNt5dnJ8bRc7TRA2+K/
y8zJmgSS6Ed8mw4kOegojItKEL7IzONARK1EYWGyKsZsX7/79VgdEGN1qt0vulgI
p/7evcAdvrqeMCZWyZiUe12hvb0lhZGwpwqA3m5R8UhCdXbxKn6ZAJ+ZenIu2qbl
43jpoAp/n5pJNf7MjqywWnToOWHlnZdqJcLUGVR9bmXqQakeXFSAyLKxhEbdVIcg
k4CKenRw1jltAs2CZSX8/YYH2R8rdFhDxTEkEStPksgG0P+fBNXbvikRAveq8soQ
IUQdZ4W+UQfHNrNu6yT1AZmkOFoKJY7sE12UpArf4HWmJPnleAY0PPypewLbTU9n
tqSLXxc29Qx0wX0Qjvf0xyVZDQc5HFhEm27yfZvt4pxpeLns4ll7ud+BMEfuBpUD
wfQly1svnZLSWj37wEks845Y3GgJnCy3xXTEluM87Db5PdyyzedZj5lFJL8IvDw4
nOgwCEjqzlHReXzSL8vhZ2cbVDEcXGaTXrM/gv9kL9V2hKaBisaO+FXultmrp+GU
Me+cZh46NZmR1GJgBaFFTkfR3EJCr8Dqx/YKp1sd9BPI1rMJ+lMVIq7l4GSFz8sb
DT6ucSfg3wb5XnDGdBDb7eNG5CQro13Oag6LIA8TJGDadg0xyKX6FYsvudCIqN9H
K04KL38+0edjvBxmRu3r5c6WeayZFM4jviU6Tfy/u7PXY4JMwetq8d/GRJEUvq2J
Jm7oqQGoRAxbjjAoA0tIh9gZVQxfj9Wa/ADiXrzrSscLawGvEPPUYweTmjUdRZLM
e++xP3DyY2yMMug7EqkR71JzCtVfopgA4qWwOqIMVlMIKUAY87nMl1ObwjguY7eb
meX3yrBUETvIQaib8nOmCRSGRefX37XBMPTH2yZFTg9L4yrWaxwi2yV0HXm8cls8
59/UxWhBsFDwhvqgqGBlc2qxMvbeXsH/ProbdwP+tFlJkw+blVgkjMBdVTaMLUJb
lb80ACq1uDqKblCMSouGKgFTE6jXjRjSaCspvYZVojPWc4bTdFQ5MqJ/yIdWRtQZ
oNJtKquCqpo4MHOx2uSF9WPhfB552M+aLFcuCAe8VDmoqECeNdJ13mqwhKKxKb+c
Sy2YQ61CeGvRfG0Mkije+g2g3HMl8s/uElF2jX4Z5YO2yDW1Ia+o4j4dPE+J1FZY
TwN2lm9wZupXAYLWcYDNT8mCz5682kdcw1PnGO0QhF1tXUmwgcAz5ilvL97NIawt
CPB+gir85xfXffZrBpbKgN9qQIMTKdhfnNuvhSu28vvZem6EUFmblRxck9eyYGWs
zsdocOXPJuPyLOcbTLIRMhztG74c0reOF2K0N3uc2BBmOibQD1KQE2uWE5cVeQE+
SXqORysH1i4lpABsmWcQuBtEKvUaMxLnjFq2o3FDu3VdavmKKi3lbtKjxulJOGCU
v812Dz1WIz2YclBHfrNfN29sfj5soRVNzMjQ1Mvh2wfZMx8UjNrARqgHhdylKnHl
+5/vz8n6p+N1nAZ3pWvT0TkqLZXBUfgGs6+mgkRfnPwnmtCnnFr5mYu8tJg28DTJ
q4Eoe4mrLFAlOa2ry+EJcirIrie/Qmi8nnURzor+YNnO/n14EJPWNcUcJ7W47aqJ
ajOnz6Jt6LYdg7NP+X8xeBU8d1YvIKyvsdVAxOw/Y6t9cM+hW4wI/F3S8qnfDITi
l21Zo2D9ruaG3RLiHpPyuS39huB84xg9gNEm/BYfNwBPJWkjqCabNmpdpJ2TTas2
j1Kq6L9RA4Rc7R8hQBjN3Z7SA7pKWjyfrP1Okf+WyOVMEg67rO6f4ZGn9lbfy6JX
FpC4793Awgyx3thl5CrEC+qJLAEa0CZmkPWndeJABl2rfBly4pe7/DOjT8MugIVC
5T4Huv7gMzlGJH5tOYp+VlYwZ5r9AVz23CGAWvZySwhK0qy5Brn22o8TjGFBjdMA
HRARA16yn5g2VujRmqdnaMe94z+tifUAJLGMXkrEncTG2oyOXnsEAFreNmuOtFTn
mNW9/jokVDsxE1WLWg8OObEv2ou7Mfto8xBIuOOioFngtNz3oCqCcLPRdYb/SD/c
CV6fFMQHVIBJeua6QJr05v5e/nLsVXQ0GNQ76vuiK4fTwSEMvisi2v/Ih53fu0JA
xgHFHOj2rdVWZtBdua6/1qx6ByZOoiLSE5sRyFjt+tBVDt4XHbER8Jjdv3nG5auW
snulEHPy5S9+Pytr/RU4kPlCzh8wp+doNvhRSPXiGOyrx4koHEreGkt3+L80ye1R
5ERGWcbAUi80Hqtb0j1QiJ+Yv7L918mqa4Xt2dRS0L6i65PG4CEXt+j4gKDG2de3
JOwQVA/eK0qN1wd6qta6ufPymOIEsYSahUxcaExE6nDZx3dpkfFEHTuWyS14qAEG
Lorq3DtxonpxJfimV7jeJm/YvA+ozF61ZnO0PDzXISK4UZSjZwcvw3lOBqxoaf9k
X0WXl8s14pmmMSXP1CnwyAmRp1Da4rB+hMdJ5v2coaOBjx2MyXyaRLl47WyYdPXV
0bV9zqAFCATnQwxCV+HYsndNXgHY4aMPUtMc9I38mIEtNOC52AhErkZX6PNshyHV
WzOMln7w/TWSd+YPub+4J51eZXO86ifrljzlTjMQialG/810fKsAEOCkzu1cu65R
oj9HUpN3Zfqd4gHT+q4/Smq+mHoj71lfdyQxOMaL0N13r8P7KXV63oTxfxH1ASMa
Gw7LFhEeisYmqdxcYpP6lr0UT39A6nPIvpcco4sgN8DLGtnf/AZ1sgAbp8v5hRtO
Qw6W+wM7aywkvwWCISzFK8m5Mg8WsqLMH1Om3wOAeioeCVTpCptyNVzpnnjU4RDE
VneZtDS9YeNbMlUUqZ3V/HNGORnfsHVfxFMOo7jMyYPyCYwSEUTiF9XpUh6QEBqX
vu3k6SHQE3GDtp0ol1wk/4G+paS0Mwfk9t7SbxXSN36qxfvZKfqbnjA7jZIz2tjC
zS2sjnc5tm352kuP0O0lfP8mLjUuIfxI2lU7LI+4QvotTvpUOyAs6LbFceiAZpKn
rlDYPM2mFH9HW75MFbQPEANNdaS24Hv/5JGFU+JjNlt3JmLVHHsTl0FugNmiheAy
vCazeEcjDi2hZvanhsJtOV+NLrzma6Lhhb7ZWkGE3caXg+a0qK7CiCQ4FIxGuA6S
TzHsT1byhaCy61l8ksRsqITGQlVljBTVCIL0gUuppX8p3ad4GKv3k9BsJ+9NjApW
YP97OsTcks/8gYXvEMe2GD+yjWkB4GUWFGtDM6ExfYbgb2Me/3/eput4XxqFUyRo
B1/jAdXMCbNfPR+HyEaei2SzdOtW6cJqgod7TV4QJXiVI1qSEbvqzO82b0/VsGgA
x5J2b/1dOHIZNvgUe9kHNRvnUYBM/DbRK8vXSNtbLqya+eC9ODk4uFXIaBPjoyrn
RWmYYgYR/Hr92pvs7+F5b8W29EvA3Q2H9eb08eBOEDobnlFnnkZ3vd4LaJFn5dyq
4DM9XxQtRAGl5jJNjVraucYHRxQNUZ2QUr6ulMBKhGj9+9BofXOj9IWAuUgt+uSI
5OwikzzDOJ9Q/cR7Lf7eRdqLJ2k/nieV990ejcCkZgrJfYBIXhEVQqYYzfn6OONc
qkWqvRnqqILPC0B+2YNvdAs8FAoaZYnMp2Gqo+EVSAOc80x00LGChSNrISnmi9Bk
Hehp/eetkrUQBEtSSe6fPQUR/91Xgf1lSxI97HqGxIneU6xEAcOOYA3lTtzbKvGf
VK39yeqXPuM8SIYyKzc1sGUi8FdxxJtcauuUAGlwiwq8dIg4tmgJpx/7la3dxGBY
CnbIHwwnwr+Zryxc6NfOGULTnzQEEKqeIgfrp6l54UljA/a9ekyedtLYlU6V2sFt
Figqq5d5q7b+yWnUX+r91b6vKjVWjxK8es+L4kLPnvDoFEeLK+A5LKhKRg/TrYPE
4/Kz+5BZiM0rguJEc/Nrtu2jaFEQSEouVrwzz+kAb79Vj3vU/lB0wSI55SknbNGQ
7DETaIywPrzwWNW8n7yVn+F/IrvZQwhVNLS6TZcHDM9l2BPV0szpRAWQemd1QeWD
Dd7eknjRniHbTXEiU33vRNerPIhLXsUtMSeX78LVYHW0ypj9ug6owhDaCZJvNyQX
24IrwSXIL3oslvhUwyjHCb69OJoFf15MZWA04R5Zh65XsuGN7B5QspZ0jfdvxuX8
o1TLnC7RzySd+mluxSh4acDLF9kR6qnfeYT+oXM15dIrU9LpikmBpc7y93Zn/r3z
5R9hQQ/GUXl5SsU4DA4LrlQ3lF0hrtEfzEOD+tyobM407VbLg7Q3kur1Joqyv6G5
g1h3NRGK8/f0KQgG3/CrZYBkPgccF/yO5JVyMuuBKmtF+ASfq1Lp+eipTQ9ihINe
GlAa5GHuyVFWh8gLq/NgUA2nF435v6Hwmqfa+3p3HokbQrkbCihSGdmEE/Gn59CL
l+20SNOvetVLh/CtmxdubSxj5ZGnvKuUUKRCteD1FNyuiYjVtIaRubi+mybKMFTN
05WluCjmCGgRPzml5znZRLqex9uRFq5mKdu5A4YDEC5XByoLK18U5fQAwtZaiL/P
ZvbX6oO4O3Ya3/32S4UZfuz3p9QVhc6N7YhWvyuPppjc5nWGUt81zfO15Mw0AssP
IkKeqkjnLhPkcavLixhv0KCVzzKJG8AWVU5wkcGJb1c4bAlMs3P9pWloUuxLfKdt
765zaVoQZAq5WckRtGyXd27kNFzdX3txe52uVPjKbxWf75rwiCAi4F/bWmYfbcby
uBJEcu5NdmsD4KR2gFkjWWY2uSLdlsdtFXPsJY+0jRV9jx2aKQc6EO9p3YPvFoEc
OK/eIQjGyWhR4VIVyjGLO1fzEJvrUUPMYhr/0L+wM3qvdiDD9HX+lDhfc9vRxZrJ
4IGbSGT+cfz9p82nYA/OUjPLeiXNT6fdkvSiMPczaPBZJh3/nFPQudYwA72ypPEm
a+qlFhvLuvYGPrC7YR9rhxQMyukBDzbBoWTwHYGM21bpHqIvE5t28NdAe3o+n2a6
fmohybSGQQ6FwaxrMZTK/saZ1wwfYhcttbFflYL8mmNzWi8xSVoNgqdX/2B73tpM
nb0Gidg3eM+T0Kh1J/YmjPYX7PBHu9RK/GyTminBsJlU9vrbhShqEllPbHvqTqlE
8Os1z1UEc+rCOKEAhY7ora6QVyVsRRZg8OsWzYDUIasjj7Kd5uzGd8j0C6LQRX9v
SXup2IIVyPiMiMXgwKA5Kx7k7jXglulCGIA21XYdu2fwKw0c81ynG7xgrXaf3Lfi
T6AoVeQdmJsYEEMt9ifkmqBpgmOTLDDoYvEXe7ZGCfkIYsIsrCos3z2JGKSCsN9D
Kgouj4XFcJzundMZ18j0KpC4tU4f8aY60mlF9r4hpHRomF5CTLumHENMc6VTLMYl
LBpZrS9P1bNRnN4HRhIjau/10/GumQ88XCpSevZlY4LpNNDfiuQVtWQ29MfQiqW6
+7M/Xi3FYIoGUTYVYnMMZA+1lSIgvn4MkzARO+ruZekoXqt6o/ihVxh/HrmrXqjS
aaf2LQfL5U1lLmyDkmQVOj1ahcBqBYiDbVxecr86vLg9A5bwCF5m6pbgomXuEkIQ
Ag149xHvcGLxMqJwnQcfPoIzn/5u3MrQZLxIh5yhneGSH3pIa+ERrok9y2oqTYOY
l4MJV2mfLOrga19XE0kmIFQ2lj74IQmufS+ZmgRljsImO4gKXyzOSMyaVmt6Ac+G
0d//bgcYH/vWsYp9puzBirAij027clslA6G5G3eux4P9rSDJLufmUjiFEGvmsGXf
guUPSZQ6tTtutdMA2Mr07med3Sk53RdmMVNIMvlOOEWXONXk3LJys5HxvrSRq5qM
8QW3270nN0xxjmdue1BlTq+oK4mRQ1GSCbzQT/jdP+OpKEDtIw8M6fsTwQ8O8+gu
5TVTDNQXTvtfymV0CxsZQySX9deQSyhnUccjwpaYp++m6D5mZFfqzTjIwRs9Nq/H
8MkWl5q2/GC1kC/1B7cGDusqAf9G4oOLP47Hu4Kwqmycr/nsemvsEByrqptBjZ3z
Pld24F2NoMpTEsKYwELPlyjoIi10hAo3XIC1G/wqYT8IMp2WJ99pReoXmJo0e0sI
nBswcDsBybBKxPuhc6GsWEVU4xiLW+Es28U4vXj4T70NejbOrU2LXQhewH+Fiey6
P1+I3bXnji9tocVuwliY+cXclMtLkVd1JX2vwTxk8C8YycQy3aIjxVDMIvRDjqem
aUSSou9bE072tRXkTknC1YkkQJAqmGksdO7sr9tDCYzCtOS0ZPWtOvHWoxNRsOxQ
hSOTooHNqq8l8wLDkGNq1aielAIBZKQSwl/C/jJWC0oCSI/5+InHQ3chf4x5quGp
7Zv2jX8PLUTP2/wZrFe2UFuKsE16EPE+7t3+Harj1D76v9Vua5rygOm+rQeW7QTr
TEl9r6vwoXo/RCoZgyEKPhWYDSVMlr44ecWSRUerYlbyTAJZM5lnIstIH/WWiWlY
cM4tsaRyWIrlJFuaSstvSxbN8jxXrUQ+I7lXWpyPh295P8tbdRzXGRnL2fMkXtXx
1lodR9F+zmhXx6viCFVvH0MiyV5ajEoKkuY8ezXSQL8Q+yb/C3bTwH8d8hU08IF7
u6+LlLcaxg+VQxRdrDB7d9SJq/RHhAwk99z1FQ+5Xvfo0m+riRHNPaOZhUOlekOl
ZUREbhKFpf2po4yeelh+1FiwVRXZVbBpc+22QnghUwstNirMCTiBGEPcwdGgjhW3
dFnu9fBY+k/3ppvAAqPb4i4TvnbsfCikv8Rd2U+JMCRpDuXKAnLPsaqhcRhqSMot
eHEI1MQoNbYisQ4oK+OwM/R6cn0dF+IBlAn06qHMXO63avVFrrAtcN4OHn+OhQlG
CFedkkjZxGYJ/iXO8ZqhFFDbMAjJe/hqVsHPyXZSpoGTM208aU4GhWE0CQMJxsIm
iCz8lffJh8wEcpuZ7/pnCnH6Bm16fI8xsLqerC6D7qkME13gx0qFYdgDh/hGBGR3
H4iUckOIfslK8rj5mq3dRtvyfdJmswzlqA4OjUPhzgr9ZfUOWiwQQsqyVkK8N63P
FTN7BhEpmBZPLvqtHwRWO8lnr5+108ziACVHrWngLpJnxTCR3AJ00I6TcJ5LwMfB
KIHr/Lk/s0IaEsxbA+QjJqx3xQv4FtgeeH3axB03tNeRs7v3IXTeCPY4D/HjugJx
oHpfmsDjCnuwy0LbOKLTX5Y5/RNTrsgAIOw4a8FMh0UmvIvPaMU9u296BdbBEN29
uFHGG7z7tKpVBSZefqRSk/GqohJYuSm0yGLki1nw3dIhBkKH3CD+CF5Mh9+9rU1l
fUdDcLYpbUs2QtevensDIxwycVC/1f/F0odDr13FKgVOsYIACKDl6HJgTCEvwvKU
5+YQFE0TgattU1JpYpRLTrYkwZcUFMaFC7PO5Jqh5AO1WEfcJjY1XrOrdPjIwm9V
3FRCMU3JXVVRcSS3oh7DRkpuQLeAwZ5qxDpWmujU/aTUtRt/DyOsIIltUxYq1y7O
z98wcyYaE0h/TfguIFz2mQqjwLVbIGvaktrKxpM4t4sodjtOc//lAMyz4X5dhbVl
canXd3PMvNYN0QYADnfrOYmp7aixXXZu3LwPK0G/cCHduwDSVeTk3Hv9rlqQDUNa
ROl+6MZlM+btzCkBummRg1x/QNRRzdil3anp4Tcy+L8JQhtnXcP+dru2RK+b2hR6
XjIzzSxp2w1zih2KQ+sOg9WdXuQcWeXAgIED0MI5AqoSCeH+BUKIph68tm0MbmyD
vWvCdrnc1zazhWgP/SMvZ/2psO2TRTS/40Lu5WQojo4LgVP0qhANMXG+pSndYJ09
bW35OGH1KpfWdO84Ssw/hLeRhZZR2MUlp1elMpufFnBCBL4G6I8WNukVEZ2eqzT2
6dbU/LqfKJ4Wri8BmgpmDvBo3CgnyFQkVYQhGDnVE6ugW0TuWA9/PWQwg/Jwnr2L
hBkDUlifNFzTuphu5po+irM0Fb3Y/JN1P5E+t71Lxu3EFajG6SPAieZXfGHg3h9h
PRE1UVeshWWTqxe/nygX1qyTil0SE6hB/z5D9OC/uOJJwvHly1DbqMS+jD7giODW
MNUr6f6e2n5f3ADsfPNrHHZNMBGiD3uoBkQVjWJBGYQmztFeOCxQemK5b1Ot5lbC
GaCcRAnRzi2SL7cZT94xWEz+qNh8KwObrcCHdv5aGfkPc6uhO6XbsHzRmPaaBvZJ
T4ksqUmKJpIsE6PZ0s6Eti+jCbZ5R7MMqqBiQah590vEW+PmRHArbAbZmOv0Iiuf
Y7ztHE4id9g1KShgwpTQBCW5B86Zs2CzL3QCJfZa8NsYC6VKu3ifFZ4IEYbN/hq7
D+5VLfeqOuSvH8XsqDnKavQjcsg20m2eUqK6dajPpFWc7TUXb8NPbfJxPRToJkPl
koCbB5IWDWBPo1F2ZV0XAF4wI+wLhGT8RwqceTpCc+yYLFzSRi0C9jfHu37zDV33
nT4iQTucR155s/YDdZGSnuZzZLKknqhZXtwifIAlAfQaHJ8Ayso4UTlaULX6Gmws
NibF8V4sgAvtcLVvIuUHU+yfwEleOWhQv72miAlgePjgaL8vCzDdpoJ7DlxvcxIg
QHDgHYYHvORemaLIwHFKGUW4000p16PP0XH84FZj0mEUGVWbbTkMrOC0wq0UvU0d
9YFuSb8feRH/fEnFwqwoRLuXGJQ0gf5NvTf6O83y9qEE35r/SvVYFVaWi8ZtUrwj
TrleEOy7b1z8475KcQg4K9XtJ4iwPPUviXPBPNoQxzoONocCIbim21pCOhmujvJ5
DQSiTqyGuAmC5HHMhDVxrN3eeGMqXPlsckZsPtdTg8guSdA2OZEsrzdF91bD4Lv2
LSVIUkvG0XsD5so/+zliTlMb/gvVKwizV36JICU61F/7F47BTdoUqtuqkIGj1tB0
MSENFpcg7dLtA2hYQflvqL4+cekc8rO5SZBjWb1Dw1cb6OnRJhtQ4t2IpGRaNemD
niePpfnC6/TDcI5awYlzUeh3VMiP1hyoexNI7eHQamRPqZtTOEHTzbuztLzSzY0A
Edd1/5ByMT7zEtgmitdS5wXGJlXQrlB4qssgjBHZVRgttsQIpmd0xGtu7AfBzkpI
Xs+cBAhF//c+Tfc7wN56qe6pmTYPX28IK2T8KwCyyi9pBhHfQHYcTOR64ATSY1Th
yTHXd7VQE9U7d6qjjlOfhXD0YHkuTm7tShYKUiUPZXgMzRpcpgn5f8Rl0CYsr+aM
huc49rcsN0cMZkxV5hBlFIBR47ts060QSV/A90znJbZr5jBG4Ov9fnuUpH1vjjkQ
kYthCNBwQ+e5d5K3Y4FlC6jofnTvjqVvfuVKicaQbqeVum7+/CZOOecrfPHQUgSU
gxWflWiLpw4Io8ykn/gf+PQkGJMJKkbKnx+9dVV6UKSSB/cwc1REAcb/1hIuGHSG
hqiiVgcoGrvzYy1qvvhKHGNNuiFWASTr0uQc/okZrFu+ei1bKBiXrhHFLz7yWJNF
SKV08PMqzW7ZYjU9ONeofNv2fsDQONaJpG6pJsVthkuCmV9XBkjJDHUDjeVefzEz
tjoPj6h462JcDiH4+cYKufsXz622u+4gpTRULFMERU1iehQvNGBhKrXHv6wKULSs
GYjhXlSUcsp27SUYyp/xLY1+ZYjIRF7NAjDLOvgkmJ3pNgS7WNCCT3Mi9QdKrgN5
lzmDyzRaYHOVisi8EtcGu3QeFCSpUwYt8crQ1coUZyG4rPs1mv5Z/kpcVje6wWBh
VKIfndsYwVBXlRVM5w5hgEEd/JgflubC3K9BBKqWS4VBLkN0FWZnKW8uhEkJzV+Z
RSPRHA5i4v/vp3V07z9hTQUpUur56ogsb62yUzKBAjr5//n+Zbm5RcOrfcMvIMKp
D45nVb+bFpYw9FxF9PnqDJtnB8KhAgLczKcc8bLaR26hqlrSR3H8D/FYWqx00CEo
BmVpIfekl6hdwFqskL/5svG+Il7QspyIDj4/2A0ax9hmItv+Yvyik1ihxMCbo50L
VBaose3kjsKEHI2/aqfp9HFVWBn16m6RuLmErq9KWSTH20egWgoZeDCUnq88EF/t
t1IK0mYAu+bR+k1pN7bbfEkX0+yak3aM1JWMMdbVrRUxcX3eOrNdtsFtMyAYxhaY
dmyBBAi+xN0BPpOTFeNHeeiQDpDhFnI4hi3Dm+e6OzzHA4PAaeh1DkHj1sqAxfrt
N8SEbp8xIkZzP7+iRD5p+vRLphqyzuIuzLsG1FzK+Lua3RtGj2LGccHWypjEG8YD
0CI6tY5G78tENz/3XqsQK6gQ3ka9lykzqcYjZ2/YhMFxmufBsgnjnDPVbDUgjfnJ
ql8/BTh98E931GY7vekOrrhXkRWwEi+SZi9HOWhSkm77C8pQDA+gGTE648z+bU94
J74gkcPlUT6GQjsHmbIy0r+GmLJ8O4EeXmPkDGsG4SoPO7+1fvYs47MW5IbEZOwC
AggO7hNiXxNXdeVNt9UO8nRn3uqgv0pEKGoQhq4L+axrQQ41R2UxROjrA5Sxgrlq
Xo5yujd3O7p/PiQOjCceD75F81gohfH+SjAipDSGk90BUMcvSwxcnXnCZk9RqMvJ
TRLiM/yg3QZSQEAd1PMd/3oqeTUBixacrteOJ1a4Ynp0ad8jB1RxTEI8aPZ6G+tP
L8d2y+N2eSviuV4a1ejrLB9NVN6CF8XAxQ835VOVL6XKFvdIclWiZ5PKm8CKmqxz
6LTLThBWn2eHESqdkbeod+apPCXUY5z4j96Rfv3vTipQZ6qE502Id2VSuwlmSYjg
wiNeaBjmIWLWclSIUl581sY6gIwckI3TWLbOiOMRSWNaDXKL1xFGlwLaXUybbWY8
TXGRb0K07D83yO/qNuunqMoN7YEIEbAzjsUg+KJxi2ueRO8c5n+kNtFViqmYjZUy
Sapq6uAzCEQ293/PcI8tHT6FqjBftzrn//XJ3IW+4xlhvozqvOhjJJialvMwev0U
EKogC1AzLOSx+Z9zssBQcJ4Nze6ISU3Z3r9iLNaWU+q0/rNJx+JZnZdHFN5vYZKy
JUErkf8u1ZVHVsUCNEQRnprudTeVwasOjb9HDxc64ASW3aDfHZkdQrsT66xaa1oy
8edf0BDFlik72vx7tWJMv8p78igqPxSYycP4Z6Xf2F2L1g0a6urczGsS6tRAAxwp
aP/pCi/wjWYk/DluWC6PmkpqLnu3JZruHyPOTYJx7fAaOviyaYSXw0+rmJM3CuAF
X7+TZ5YK36p0GKf1U5J6YA9CwsslnYfgrfRzBsMa4kzNveyd8zJgi7nsSIT7ZKGB
+HkRNV0IVNRaWBjFio8RE/kVSxGvoJIFGFvmRkl7jR0riplXm3nGBIE9R8FisWKN
E6BajUgPyRQ2Lehv2GWkJ7GlFkXS3Clo9FyZoOAfEXQxG48KEc315Bc8bqYoXfEW
2W1BK49AGq+9ML8dhctfYC06T5PkXtWc/Ai4CqEW0ORIkbh16H2UPL+Tv0LXQvWB
vKYEiAnnJlv+NM1f/VoKbHvrdbKDrAfTpmYnWovZOVt+LW1useDljrkVYlOwwQdw
RtDGRnx8SfJaQFfGDXRdqjNhY5BTSRXNQGA4wFc4szTMnbN+Tws2Z7cZ/017/Gda
/ogjWdsAr1OfP2/t/UZ9ovMeHPgJYAVByTKhxr3jr8iGeHrDgJNarKUelc22BNOI
hecwpKnz2/wE/n/TNIFaTyIzY0+87YriZ2VK5gjmERx2HZ+A/qcMVQAZJ0gSBBMQ
9C4Rbryv3Lu0SWA6GMuJapH3ocAY1cRrccVLcWjqsMqsvoVGiyQqWrxmk09SWr9m
f1iaDKd4fE0EMep4G7XWHTwwyU3PxSFrh57CW0kKxmvPC89y4IM7/FsiFRjYfMBf
udMWWc5vp6e6Ps//fTnt3rHw1R1akD2+ht3BpOhBUqOdiQVMFOPIGHZ8UbNSix/f
4V/jCmn4b2ixxALdoTwPYn5uz/VVxwiyaexDLqQLCezLqjdhoEX1CufS50BVGKN0
h2jKWR29JUzMlSOisvAW0xQSeQMoIsZU02vF3sPDnaTxsjwzBfvgwFF+6KXbUjJv
pW3M9WgHWW0nQDP4rjeFJaRwNV3z/eGtl5YBxN/bRQYUg+hPvlfJKlTGxxvIBQu5
mbgmFzsmojRPLdk3X+6B6E4WLNqM8SYvaiOd2+mvU71GJOhNQnPRxt1AlWaWyQfY
lWQWXPRQ3hfTA8dtyWz+b3hziWiZBK2G2dSsuJIzG+eYdrJdZgcqN8THGAyfShTV
F+grk5OxOzg2IR4al4UpeLdHgOHD0Q8E87mgcWCaoVzt9diho74rTHFlSjJpc5wp
beLSTHbwKpj95Szjfcv9D2T4HwZVhjMIrNp7WMhVgKQcqr6lGgHMQGaKdpreNY+Q
iBFwUNbgvkCcTvMZVTkJXUKztdNA0FRf7d2MmXc3fwvjEVNoe9YKt0Q0sdKmoSeq
dR61B6YB6FwmKG8VgtnPnyJ1d1zwyaaruSSAXGw7WfsrpZZEq8B3QW1oEQMeYpNW
11AMKAwqfUigh6KUr+ag9lYp3F205x0Lzz1AUx1DS95pYqmc2JhzuP8LGI0X859b
YO0G9SATMfb/pS/FT4CPn5fQslBosFUqJkZ9I7Zvdbi8qvf+IcX1Ah9u1Q47h3W9
N0ZQ81CeA4qRUorEMX5iQ/Hh2xoC315AgxT7NAmMiZDj1AvUw32iTvRchuK3Db4+
GBpzojSye4dG0gDUMHPNph0NMnY8t1NHxTQZ/RF2C6Fd7maIZg2RW3dtmprxF95p
EKVYEneYlCzFBLzXT4hEyzV1sESA0z3VJmJu6Zm4US5p879jjHTJbPO79gF2YT3w
66upge9MYz2y1kgGb1P7RcMLgyfyj1bsO8ZZ5T6UzUBhYbyVJdKUH9wXIWtjSUe1
XXEBnnWE5Ww/PcxqLDYmTf2SXCexDVPjIJmO1oXUA+IFSyeF1fynBH3hGek60R/U
w6IyXPH2oG5L4VHJvvatrGonlsyN84mfOCOi4qjkpV4Jo5uyazoI4sZiPBrb2cWW
5JrqvIc9RVOg5cKAcFpkIpiNEQh4PJw9leX4R0sTAAFgUg9xEU8ZUe3Ro9pyWa6U
cqFAR8yTcVW24oj7nnEvXz8zYHly9+gT4tzN5cREpj04pOhkFqMbAGXhrCEvuXND
HiDBEU7TqYRp++nhJGkGH3mIAQiEIdil2kv2HTIWl6fs9bvSsc4pIXHFef0c+txI
L6EyrQSd/kC4qXM5hQ6PnaaGbuAWcOu4o3HFE/VmWGjD4L5qROH487lqYMX66Z2n
rronvCof6tqk94067uOUc/TT00UYkcnw5Tm7h1lkCOe4phW0JAnFSo+25UVU4G5j
+Nu5MPftZDJ6lWD+RMvktpWRvNt7cMhdtTmBxeBu0/5i1usHPS7nTXjTAdB0SUxN
PeJ0VeSPOS+jTOXl81u5Fa9iwYzgW6kfkOAAF771GwwpNevGMV99c3PPfwV2K/rU
51PCM7PK6s4w+TB69wBS3s/YbxfUmK+3tylphLUPpWftxWQRCQILpk2Ehit6iJ/R
5efH8ucNpX8F16ggJgmho9GSKOzDl5hQH8MThpy9d8I9qTCPFGQUvHxYPFkLDqFI
VhNWkFHIuty0PMSzqGj3ZoHQXTwf37oZX1C7SPy/f8oaRd5hXfOcMgQ1XWJt56vP
uotacpwwqJ0JMc9lBG79Dx+UWr7umPFVM18Dz3uuBRkB0HSeRle5K5dlF0XzRmrh
e0oMhdecNuJTc+8+r43n/wX/SU/F5tSfacrZrmCgbOf6yQESlhVasYk5AelYtsDV
DJOQdrM9FE6pZwQQHHCUfSNL15hsxB2NqTSxte6HaZEdDkSYu5b6zib1uf+GRZff
QtmJZCB8kAN7iksuK08cFfuX7IhMWgJ22gX1tyBP2bJVNNqi0iUJRFSul1Xoxw56
HizcJbtr3CdO94Z45/Zr071/L/RPRh1KxKHrX3uKWxvuOIfot/nhpeOpN0Yyc8t9
WtrR7oJjGWvwEVDx1TSPgiPrcEd3Kyk9hRR2ofhis5mh6Juo6VgirXyVCcSxEah4
TLTny2/OXjKKw26wwjxkId6HUn98IdpNTem873a8R+OEJjy6c9VlgXIb2yBdB4Ol
khd4egqkAms4gbAtcjZQ+iZvjgPGLAwwQxAqKwMYLqdZmHy7t0D6oZqkX9Ao4E2V
wbCzD0V7V0XP911Vrs0cYrKx18eboxZQdTAmpQju/1TJ3oEU2Kanon585sAORaF0
8W07vrsC4hHblHbXXUj9DRPe9RLD9qOqbe/+lF0stYO66GOLG9vE2hF1KKgZ7B4A
ZWJVkmSgYr5wCffkWKSXo98JGhMk1FjLUZphXIZYTrnkPY5ymmLt1IeYRVDVcHu0
TSfnljiRlQ5+omys1LClXCoknAT0nqDw03yTkmqxvCc9sdJeQGSmqmD7cJlHa7Nu
LIN2DcYhW6MDrHTBdanEfM+wqGhNIxOo9Yrr+nj5oB7aJHnfdrmIOSTAjljyP8fR
aPWdms1+ySMw8ESbAV241g6Fqb+n+wm82qD/NO7UXTSNuMs4XhUsp3zU3dGyEslf
NlVHh/B2MtkqOduC459eN9YQ5nMXdlV7rmofmyOruJ5v/wqNNUplsRL+/ho3A1VV
gtFTw6l6/SGDmvcl51G1RLlLvOKtjrNfCAYD76Em+3wERTUHxQdr5xUueCwexdW7
PUDF069kAoFAO/WkC/kfqCa3Qa91fepcmvx2R9ytMkvNBJ4+52eQYwyydBhpUo78
9ZmB0kjg/rCER6m4fZhX5z3atO59CpmD0ZhXHEdHek7w3m4klTgFFjx5CE5O2Wtr
S8Lw8PVN3iCqH7FAyGyxs50q2hdcG8i9v80HBDaFmaCgOSR6vPYeZViWL2TCZSad
VQb3/kjeRZh15sxf1R8AiLmsfQKlGQ/qCz84K8YO85tRYGjMkJy2gtv5umpXqvv+
7I9xwOWZiQjfbPxhsfRTuVp4VYg5tVY2/iuiSTiowtnNv810YPmgINHfrZ9YtbUV
eJhj6lOXX0XyNOQkza/hNiDWeC75Uiw21UqyKmLu4sK1WTym6dewpwc7oIyeJR4e
flK1ojr0Y5ZkAk6XdFO36fdI0dgI+Ry/R/4SesVMSCBUEFTl+zHLCdsv8L78Xxc3
rocLIR716QU1fbwcK/NCPx6aPN1uS7uXV7MlTQI1H/SIqtZtujyzTfrvY5lSKCiD
hLDlpckn4JqilNPqyOPzeSslwgPrxjgxswNSxiC8gGFp4Vf831u6sEl/ko5WXrt8
9N6pqkzl4MuyB7I4wkdl1xD8IpzOyDK3HeWLiVofwVdEEkz0glO40jQeC++KQBOA
111J/A8SgRKRg5jBwRanTuKjCdjv6VlN1u+oi2a83kfOFNOlJSS4Vlx234Jrndzg
JeN0qTIcMjJ9jkXdIAemaDustwIiYtWFvJMEbsPb29aWUqdD+Zf+mSD3+HvfScz9
yTeZOhWzQw7Rh6Df+oCVYZAMwEuEJWtbecy/msXhh52tV4HT+XC3D8kJBijjyVen
lEFUuV3PzKEejKU58cDSnOZuLFh+/4CU+uBe6p1A4Jfo35i+XUhpnAhud3OFF7/d
vtSm9q6q3ojFVfFz+njJzRgq4VhwDPBhdcRlFfo+mP/U/Fo9GgfIszXIGwhdR+Pc
EBFG+LqgluyMaxdxUmzwrV0+7XAqqo9q6kCEe2hawNBK8XZLo7a0ROjM5UX68+fg
3VckMepCsDCVyDytSRztv/3hHAuu1eBhFJvkNOpjOzVvACauv4kdASLUBjmE+cIL
s5JcqqhVXiNRAOrc8NqD9NPCPBGfoDq5teURJUPKSJdwO4VD/nAqiuMoLTtZF790
iIvMmLur01IPxb1cVAgA6zCCY7wCLeS3XOIESNLExy3n7GQPkb2EFkVMB35ePFZp
M01nj+YKIhSMcCMU+UTCD2/6WVCyC9ArkEbhee/diXeGNyVDOveyinMt4HMVcn8n
f2gf1peUEPsZuZKYSfgCvJmOvJDmLwgtyD0cD1iwyQBqRHUgyt7xF1uUVFiTEbNG
75S3JaWU85kRgONzPBt/9//jChx+7P2FEGQeIuG0TRG1vRVWtwFXSZNwD9E+J6js
6rJWXO7SL+P1bLipK9mijnaTMR3cK6ibCHCjVeONVIQkN3i38R3Rmz6Ot9FIsmEC
4B3w7mwP76VBb21ySwRNIwlR6A+rRqwDjrtAsbh4CXvp9LFzTBbYwbs7jLnFqNhF
6A54SI6e93k4NJTCvIHRxfENHCl0U+r6uxSGHo2xuu4t/SFenXqkbuEJi019Ql5n
rjiBbP4ftC9yvOUNH7MAH50pIEQ7N92z54QqglJiBkvG9lZ1lD155YZVidRo0dT1
rEvZRYCfMHgsBJ37q4dH+0ct0H0beHViUcuJBAP5M0rOI17IjVbDCTeNaY9H1uNQ
0sxm7R5pkrS/qaqoalclc7+mWWDs+5BBEIWOO3KDclIM8Rwt2x9SDJzxdeUrQopj
HOevboj/fgaHORRpx0ZJvEPb51fZKw+EhOqcgqDLVisZ4yB26XYJA1wpFapDt0q5
JJW5agWPIU47gV+81LbK3eiMZQHgsb5Wwug9n4O1RZyYvFuS63UDYuyZpuzwIHch
iK6PYRhKo2GSgeLiJUSeSyZCjozc0L5RYckKVTOtW1sfG+mnoSHGohMCzxDfH0yM
2s1HuwFmhsJt4qNkq+B+CZB5XxwtxEkWjQOso/cMXZc4yE4/RbuM7PQpng9So6nQ
dgPrAZRcNEwe1q9odKLiGYjfwQw7PnXItGVmE9ir1GDbPEYiiGG8hkTQH0ypkAKP
rXoHHiHqAWY8zI4c3nQ+6cjapln8ijwuZRoH4xAD3q+9J9ylcDjRb5l5gsoIfnwT
DenGA3AlPyX0fNk5S+tLAiH3EnF49oRTs+M4XGwVko/doXKINz5UQ08YxUp2wKft
ATdueSZmP6HWDFPo8E+sj0jQ1QPIYXMuLwHMUeLYIAxMZPWAAHtu+9K/cGzhxXKD
WnV1WEUg4zeXvFlm7BKr455n48uqOlG1rV1K3/0kYrEwPABfFcPx0Pt8bLBAkh3R
nb3yRCfl+aWhKZGYFJAuZANvc1dSTMCif8DgeIRSysaB4yiuCm7nDuM3lddazthI
/wxx2fGXMEvsLo2dOirWosxU0b3NbIaYS6A5MKP1M9b/Q0PgXFGK34JPv+vzszn8
z+2zksJ2qCJYHhCR8BRGcu0OWoPnUHA+kxlw3BwXm64Qx3mtrBj4y8kqj3qPZI0H
CbGzcVkfGuJ9n8701BtPe0WKrUC6UjjRyPP2fxeuub41rITbx4CD9AJdFXnrQMo2
cX4ATExMDzkzDgrm5W8jVO63s2MgWR/mlsB8ZWWn8NydFQhDZ3vsHKWxmFE1u61t
buTSW6cKfkgEdvLtfHFONSLvbUbJxa0q+g/RhH8KGgw0fpFzk3LuNU+4xBsjEUDX
Q2saE4jQPDRiExFQkZnQEbaCRD1va094FPeUs6ouuT5AiEhNCmL8NU0xkEf7qsGk
22QcsaUb8MfahWtPZ+wTjtCYVO28Gr4Tx/vdQgLdEO6gRZOVm2Fn64oNESwR/hm7
WuyN7RluwghPXZ8o144gMKZOjgIWoQOMfMJ04TuThlGsHh/pQRTQ4zv+7kl/YNsk
tJ/9+TFyQKNOrGexTGZRt/9D48IvE05bJkLIMVRQhZlXugjBNojqKAlphd+y/rBS
pTjFlHc65KxIDmzVnEag21y1Q4shRAzGQB64ZhxyFjLX+2dM6x5E/+a0EstxFQgs
zfD59tnWiey99I4qASk/uhkaNpxqVZeigRrrpUBveiuBcAatTs2ysqCrPRPL7gZD
JEULQw0PVDyeyNKO+zmMq3FJIGyp/UqwBKTtF2wuZCxq+db5SaZlgW8Qdn59jqN8
Fu9ltSVYWMMKka1lrSdGS3fjh11k/KoXDfQ0A7cBqv4UWptgB/LUFudbgT1LXr7u
hj9pOAlB9apJbQpMigCajBRnYlvgPrU42HVpw7q/jU6zI90HH/I1acnXGuPUQrAs
oJGjTFcehSUZuTAgniRkzEYiMrWEtOiwBHAAYOdSap11M4HvsNPCYIfv4qA8nZBg
glZoaPgqCxYYI37lSljX8nuktl09PPGPlalGIufsvSpjiXUpbvCUnq6iOCusEHrT
aHe2iQQXSbefJwegPwgSZ0125aESSeEUMhfSXy4QpzevYMioUVD+sDDLsvilqmYJ
qpumYG9iiwLEfiD2m2eBvEH+bnyDnPUjOxbGQSvVKm+Bc6TDLYP99dnYzLqc74Oj
lsVOzENl2ILrDS9gM4r6E5F3PYtMxfpNFUGXsa0N9AJxN4ecSuV7+MibFO7cYpL7
we4oPwzRWehNrUc6c3o5GoaN+WwCTPETjGat/d38xK/1+Oyzu1/D2Wo7xDxmFA1N
EOT8u52Xi3Rrhd9Z26x8a562ziMuFJIPGJppy9dJgSCAWUiDDkYceqnNiShHWiSq
K31sxs1tSJkixVh2XYlVfOoMjEwgVs6qmAATtNnrZKUIz3PDlqQhNnls2f37Rz4l
kXE7pY+TQFoNfdKLXVdv+lMvl5k0xJqsaYqFoRU0QfvNumojGrdL5f/d69j9j0z5
WnyFDejVZPpDXUFfdhpQ4aPerueL6S0jTcJe40aJxUPZQJIdW8zZuHtJG87CU0FE
WA6pjO9+2dgSJmvkjhAHn60pNMqW3iMCpS6wt21yB3vowsW1bITNW375VN8uqVR7
m8vepB7WtPKez5Vklzu9KWHlNaTseyMtMVs1iK3DSiXgMoTHJ7YMeZs/JNc63C5x
zVD7E+x7c2dLVy2OrDOmMkpR3g9JzhIHgxmgDoi7/2pHdUeT3LaF7mtRJFTsq5jc
0aoen8d1gZkc/jXbITCwA0lhVIVkZsymzW6+G2092MaTun51saFYk+98taugwrT0
UEQXuDHKwD6atXojBvPRI1rOpd9ek96bUu4EzuHER0I+uytuhGKi1hNbtKpQG1Zz
TJ/Owzm4sj3wqbaq9eHJKEmxHCH6zn221PK8xmfrrw5dBvwqKeWsdHLVt9+jKBZN
fmKtQge+LsnC1KPbSxIeZjzHnp5fke+O5gmnIVhuPvlgLL+Q9EgmoO4unUL/nnP/
fiJsNjGWTy7BnV0jVOzZI7hT45ohWQwHqhJkv4QEVrunI/LUKw1hfbCE2RcD9sEP
p5tAFRh3jEBUHgrcJnDCMIp5f9ksx0Zz/dRiMB/evqeP22nSerpE7c0zXSOgyDas
6J0KX/9gmPg7pKEeGkZ6x+7h4+O/za5u+u5WZgCQhl81bbxbjNXGSSWmlvEJj6rA
gmFfH4HqZ5eWpzlD80wPjUSJGoJWdeF00xKFs2EMxCEuYcKZzjKPFFuMJtmEJaeD
4sm7FYv4WjF6BMw+Xdw/2MULH6oqD7/e3WrqADWejW+EBwmCj+0i5uHa4rsqeqQu
02xUgU2uMwIHaW4qPV3YYPc+g/DpPE5GD/NWspiuXWuWa8bhm3Tydm9zvnyYPnDp
dm7orB0KV259qUIQBjp5F+5MpVesEJLja9XoFlhsNlUIe5TaS50IJ/7gWfj+xZaT
ehquvvEBQsyAqRVqPDNjFyhexaEVsavHaoLkOvDmSjcv+0DTcojj4DKTqmVJ7VbV
yPHNmnneNloH7ZdRZf06I2qIF8GiU1VmYCRt6xVY2bHHzMSoq15Y9NLUb6xY6SBH
x/5OBAIQqNkrLAoXFV5PTix/Z01A4+3VNdeTHZQ8gd051qpEuKnuLE5X2sURn8zt
73hH5slqwrO/olsXmyAZu1vwZlQDDcEuCT086dfoitT8OGFz/ANasOn7SetGpbj3
PKptjXm6mwkw5bVQWWi19IWnoUoyyMLFc8DrrHZ3F2qtT2V+6c2wzDxk7YhSa473
f2z48BdsvTtb+evypstKXwHG0o+PabfSf221V/r/5nvbNr0dYE/rsmSUuVGj7ArM
IXwTyYZsliHBHmRIw/jFrYlvOPSvwqS037NFKD/fLZQTwcH5iXjOKxVhIvBK9XU6
mu6GncQ/DVu3zxmN0hxutf1kpCK5EumcO6G5cc/xHRu7aQKg+KN6FgMjIvq3sa99
A4JZ3Aj8g70617O9J8cbBnLBk48QTniyVi9eTZ16JBdvPXuKjloOlk8grJnMajeR
zmfTHb3NMrGxsRudJmLWm6Mq+vknL+BIprL0l9rO9cYOTYQ90FCBWN62PJJmQijX
oZtGEdoMhZkKkwna+IXaUa2iznqdEECrw0z57h5gV4wFnSP3TStIwGWK14F9IK8w
ioZPMGrVJQsm1SDQ2werPE6BZjI7P00p6jIxxSqEjTnZ9GXTMalH9V4LPAuaHQhv
9gjMRSiByQKOG3yK2j4K23mQ/5Lhj0lZxfplPac43OUvvPzxhwygVnkBjnpeXzVL
lOx7tq/ACCsS8OtM16rn7veL2w4yF/IiTUlNz9OJW3IYU/Ow2c/H3+Vs6c+F3oN2
0Fnqf856LMN6eIALkg+MRZnSegcXTsxHsdKjKTrDjrFqLxjyibW+dI5FnTuStB4t
9Gknk6TfPpQYazGKLg/3/JGIoj0GA8J2T7G8EGbm+ZArgvGpLHkiN+lAm5rEAjEP
MoFbiWN1pz9YaRycltIXKlclTTzfCmO+dqe35NLHLFcyBo8lJfI14jfR2MVbobEg
a88iIFikbRskFYkcL7gsoGa5b0uex0R6Jvaw/YkYbkv4mpspYdtiWrKQ+ARXmLxx
Wr0W3V2QUFFDeYoD9lxHPtOYmN4Y4jJTEcERf3lXdHMKKh79SG1q3tgMSdUM260n
S8oN1U24beXmLzZMUTUkcDMcQIlK8lMtwe00nRPxT4T2RbbKLcfJ9ieXsFV7OTn3
NpLWA7bRSzy8NewvLPcAs3rirehE87RGVAxQHtICv9W4OZLTXDK5zPtxzypNeDi2
j5bwcb9nYyGx/cXaJD9uHgpj85mmwbSaqKiKC8niE+AX/rF2pMGk7mtac6pcgJKS
F3f2IUgoPihwD+U3+l8g4jNZ6apVsb0DWH1zWhqpW4JgoMYYnMCqwlto8B5udf5a
AovEsDlUG88gKPcddCkYqInckAaH62pbHNgZD+CugnNm7HPqmsAcCB74dB4SArvs
H1+lxIDUY+m7tK9GJuhrLawozaUTrpAGPdQAMS0LgIxjNGE8sW/xOr2zum74cS+B
9Uvyg1H5E3lo4w7u9Xpa7joDV7mtr64zZPg6Zc5sQz0Dew9zIpL3cKeBRPSuOG+i
Jwienc7z3IBTfGvkS6NqRSJuG80WERcxhF0d9Fs3HL7Vdsd1fyyj3DWTME+MVwDu
iL2VeEYlqWnohb1B6y0rWZM0Mb3/SkUq75d0bT5RB++03I7x7+KxCSemaOLM5KCG
ZMT/nXBLiojcB+iZjSeOzwgaD1kHKc0VdHRzeDnDWKUWHrzMAR8qnUT0KxNzd0ho
groJI0Oo342od7Xl53mDNJ9y7dm5doJvzFNGPM8Dvp7jI4NDCzkpsXK2xbGW3+zV
VentX9djs1Go3WJOWmDb5DvJ7dV4/UedmhvQ1plfeDvSUlaoaWtkT469+oRj8i5a
n5F2F3xFLBV1k1YOCyQmNmY9eAi+VGRZQfNfwkJJMB0vjxdS13vuIRwy3zVMrXbS
N+R8ALWr2ihWAj+7Wbi8TMDuOJJNDUXSaEpcat1ANei1s1rT8SltE1LBNikBvj+C
8NCesY9QlhcFB+U8NzZa4TNqmgiNsSBvl1/AhFO/fzbAO2ACm4hSzlsHA3ZW3REu
As1pP0ZTOSQLVE/JGdIUqbron06EOGy/j2LIEpNVtyqFYdN82zezxF0qQI08NWLb
tvuXlhy9JHYOVVHVLewTgxcZ1YvEqMivS6fJQQeEEHbE39K3dSg316nseYaVUWWF
hzocNV+fSZE0gLMxD7Nj+WMGIKrkGVTNL67Novft2+I1rVRhvQpJCuNf1sZSDP4r
nSj2l/kkPcVatYqNrEJv5UqPgqDF8okjZ8ASBnY6SWiZ3fTjQrg52cHgVGaWAQYE
6c+oVJ1drRPqmeCX62Erdqnbx/IC0vrz+bWH8JQCdUG/CxymhYZejjT5V0w3AvZP
eu0+hy/uH1nCH5V9cYM7s04swRJJr1QHzcHqGkalgA1KVditnpORjaskf2dhjmvB
bK3lVkr+U3P56wuo/d7dSnTM3B5siIp8j6tJmhuqNASpIr5LlTwwkd4E32cr8hon
mV1Entw1MlTsnF7FbHnjDsIaN/M9HS4HfTF7Gcx7vjrQHhh0Ot0VzXC9gb2S/OkC
ObC+GRW3YgXfOZTq65yfMVOU5H3K+NtNg/jBhJ4emo6F0FocwiFZH2AjDyklF5Yo
HMD/dxRPOSSporfZMZ4fxRrM7ZBxJHL/WgSzQBN/MmCHMFozCaguRiNa+ISoepSy
0bWTyBP/OfRly90Qcfsj8sUMtLKwWoLigg8aXZq+euCBNQhcNUg7NlOL/nLi43Xg
aTJx+N+EPYM75o/IKI9rN59Hl1VwIG9kqmM2Wc6VlcT0zaR7Y9HS28ELyTxetoLo
fSk/ukbCC68yQzoNxXNJJu4tbY+Fpl3MqoJgz77JkMSpKtnjqZIYzsdNfYn3H3kz
vqGmWcgjeiYSRr2SKrjNb9VkIcq3epA19VJ1JDeDxbyFLRu98DonemFe6Wq1Ybhw
OJ+fQNp1bF2zGKWyB1zUK4QBusxGbuysBpcm2mrBvEZgqCDnSXxbO+wBMsPpiTpd
tCR5nrWC5N2yARmZgO9sMOfc8EiNMCx4+9tDWDODUT4D/+XzabGC9zQuhcr+qfpX
QMKpDJe3zFcFpiYJMMsQL63Ji9BBMafqYrCVHmuXz0xzaTiMWVCT/Q8i4+8rIyu1
wxTvaUJo/He/el2xlvd11aKTJVa9ONvEo1z+4fgqhDQdQ0SXdX7m67ftdsCVk71J
O4kST+UU9B7V0Kw5X8RGFrL2Ol0EOIG/JnBlvlcrJhi3dHHytOrrlnojTlq3KpR8
QsioISwQP3RfoWhXX40dxDOEKDlBh9c6XAnlSYW8/IMZfP07cIAwhdJcW7EJMY9G
5dwwjTztHD4wNEQ2gf/19O33JoJuXXtK7yDhnbLAfPHEb8FWRmxo3VtdC60wzJlf
z3/4smHRYvruOSTN3dq4InFlmJ1ZasGtYUjqjTROUF82KQTYMahpy3evZmOakdtP
fM4wH27bNJD0VxjZ0L7WDnwyvFslKbxNq8+YNKGq4h+jXi3azOj5easU8odQ3lOQ
YEVWt2YdjuaJEAYnqgxxfrdfCOftWAMKHp+jDWP6OC9GNFkxGoyupbU+dtmJOC2+
z9ciZce1fmji5ktXNOBMR7PdcBdN0VEvHVcrPld13CiKec+t4PKzIsfoqskhMVmb
mbeiyLppWjrgB0KiYHZUzxUsbbexw5YB/lz7CXisjXC5Jl80vIFmd2UscZm59kgH
6UCygh2oap3gqQFWZlnh66aBgBV8PK0i57k1guNknEYkMBnk18JIy4veYCHmHHXm
JgbKxyULfCuTr+76HGcdUxyJHp/0I0RhVrgI4JolSAhw3lxMMybEvHYXOFJDQGMd
OQc8P/FlpieU1hszsRhaK4T4CYiaRazXRlmELhnJrhE7zVaJ+P+KGYNhPgnOtKqA
sZw4T3bCVaNzMJz6MfqzXo3S7WgeWoLUHGcZVrJJmRfEVQBTNW7OaSvrL7MoUBrE
INYowKhIzKm9K5hfQoVL7Leu5Z4GokZR7mY+OzaDGCF+VsrtvYs5HOiIR6ge5Hxa
w01J58G5uo8P2xRLRNnANQx97CH8I4yKeABwZAdgSXXpGrCcgRV5Xe77Rgk8vwkv
RHDt6M4TjT0mMJWjp1umoJQ0SY2cWirjPQfvcPLvnV0/HtWFL76dPhtgAzO1HjtL
KS7tRju6T/RrHuqT/IbVhB7/UaGI6ugtWU7frdK/4spVZwvVjl9ILDfGe9CbXon4
xQfJEQZgV4uFRDoW/kSYt78lT9I1vm01vbrER8CbHn/DOr/Q/X/BAIyOESJNIwsO
pNvOgBQVlGmfkmh2C8Xu2VLY5IKc9EDO/udSYBkx63slOGMGS8+aWcByAjtpIgCz
uIzZVsMCvZwwrIbZI4wgYy6uf7xWx1WoNQlpUVFjdUuSFml67QxAvUz5YXAAROCQ
RGYgM1uACQXXJ0I49Nan+EYcOifc7gNWfKPqgmf3Jg7FfdwFIVN+nudbttZhxSo8
TApEkeoAhyfuUvDOP2AhQfhJ5A9Jg2Y6UGjDqAlPFBtv8DbBt4ZLZevqjbib5axu
+Ul8hRm5MYBD+Oswl8zDMyeLqSSIdAvbifU35IeLgK/RWiZO+fZ5SKXMFl0o+jnJ
zcQFzh55NxBLE+fgnkIW6Hy6EGfl8Inb6ayJ1mEjyzT1EGNoETNOc/7xVtox5bqP
fQNtvkpiQwnTiqSjd1q2nJWGJKutHqIxd4opMNnN5Nvr/LEvI/uvD7E/9UkYDHjk
T3IAzEk3ZabQTyZaKc+8JCRpWgxkQhik51OlhMGKlQGvhRMKiocNPEBqh8t1vwko
wGSQNnAqbCYySsfyS/FCbjnyrCRr/BCmiBpx4XBCpshg56oAkw2CDlPHj9d/ZiIe
LAMRm0uW4GfJnjAZwAluGbTSFVIoUs+NVn4ko1NFEN9n9qhn5eUFfgLg8Ychg+kF
yfhYiDoEzyuBVMjiYlGYe9nz4bewr+E0pJnTH2B3ZH5EyzzhHu0lOIkIbaYWRjPY
FKMKeQ7bAigy663gU95XIOI/+vzaBsNropz2eeGk/A/3snH7fb8OEgFPVwluQtAt
g4h/IC2Rduqksi1iS3UmSupA8Oj2ZUDGN17iVJDjaklon9EBtzdSEArNAsu+FcF+
dzLUSkG8hggANpq6tQU4h8HxJPxJ6BtdXcQz85JCYP8sxyfC9vj1cjIqE9gRuFz9
b9ZzCah8pgyqzmO9RVndO0Bhmf6o0tF+bF6ASSfc2CfjW9GXblDWr/z3IcgxxNYP
VL73/I6y2kHEXQ68AyBXep5bcWCR/QY3ikqsxsf8ZzvQJPMD7pXMK0GCjbRiwP8M
vLRcAWD22bW5fhBIVezLVgy9nQk8Zut+p/XaTzfE1aEU/WFgFvI4LBG1VDO+l1hM
IR88ZQEsnRpBLd4ltgldfppIQwDZ59xkXaplIyKrsB/q0Ij7PqC4HEFMQQ0IZdFb
DWjPI9HMPph+j8v2DRIENiYE9sJzjbbJloFxDTWzTigm+v8+/Rz3ZbP0pq/yvATE
Ai7z/0RI0Eede+H49jhUu+tQrDpP/uuj8bUFa7fCNFSWeCWGfbmYgbw0hQpuKBiH
kzu8Lux7doLKElaIberkdrtgkvNYflT/we3xO+sBpVqJfjrtr8mZYjYjM2CwjJ3J
kq5ZRD67kgCybuvXm8yXzK+2fprL3705Y2mqW1mGm3oRLa0qt1jOKxlKvA0tkM4K
1bR0YOapes6Q8V/CDX7bWgYqb3fXu43TpBYlTcvFpVp49YN5nUeHHbyXOaj4Fiz7
5vO8F4dIw1zs5CDQ/xHVM5GTLo1JFHDLD40fnjiRcIGHEZqi0W+xJItTalA+dzjN
/g4qUjRN2xxL/tblVbfkvmLx3yTtBpoxETksZ6kXvHNYCwDc6aQS8vS8MgFVAa7l
c7UZ5mPLUt01bx75jasZtZAuiON54hY4+U+mE3mxQeJsmSDa3vhU0jRqOPIxfIoc
ntlj0NO3XkufYI9yBOJPlrIHxyuounCNJ5VJXyBKC8G4PdbhhwktUM5icXMFRrhe
Mae5NWTh1gzqg4Pdze3PIcyHML69btyKYmsWIJj1+EcPctE9eiq7hNvkk3yqpc3H
qaLjcO7QbGOmBi76F+4Y9Y7Lx/u+C8FMY9RdN8a1DnZZVIdoyXwAp58ERJzIfqG9
IqMQFn9RyPSbByXpkrjsgZvCsKZXt0FVL6l9sat7o8+PtqRp5yupOxTKTVDudWdw
LlC8R3fWsINyUUDHif13g89QRDwx+O2DJENM0ALWrogLJpq7iHv3zEZy0oZdXKde
UDIpF84DYBbMoIejqQNWIe4/ruPIHMkifLDyoAa9RbrbRJMOmj/1HlMQ5sjz9ITS
siA1hnjgtpShsw2h88NcN3awUSaxEdP3Pj8+w3mpsZjRelK1+EfV9rqv9p5TWDrL
s5aPrW5cjGd//MZgjsu6FB3TA4CQb3sZ+3vvW75SzYDCACPrma+ACICDBFtjz6WH
PUp/ndSGlsd5GiJvcbGpHVzQyJhv0IyYHThtbA8f84EVOYVi0NaYtvsD9LnRDlNn
M2pTOf99aWkLRzwcC4nV9oo1CMrW07BnYEa01wx4YQhJkNK4Q7ukiSoDHgwd6g5R
yLKXzik747coIp2pVRGdK5tdjAvhS90Rx8opnziQS+BvpSQTcfhzkE1nylHJHEuu
zxkSHlTVao7zrnukVboqJ9qWTzEdMwYnJr+7wJjnrNc/pxoWmf+mR2nlhAnebMEA
/2di/aIaLxImJwnOAPwfGKWOl+lEymyI7iM9QUr3uXm8F7CJA9pfaGFZZXF8FF2O
p0Ljdmn3dxT2ZEXKY5o60gfZMt95vKZPQ3F6qrmYeV9DDugS+KEAZs3hkzfdcQxr
8IjQXkhwTNP6Bh4je6d76AfZncaxUCOpu02wxi1q63+IML5fKbt6O+GHu3ThLcrh
ndDHGom2MNVOoE+8MmdTpMee1CbWk4EpQzzSubWTHN8CJXfkE5v9SXhKgfoeLBoH
93cqpAKWLzwd5FpNmAHS8lG0MPzE6afD1T5VxURHn0wCz/KMJIqTlbQao7DEBalR
BYpd1BWli+v/wXVoc2MpSzw62rsLGOJheQoiw+H2ChxDnPg4xngZaDvfWLu7SXEE
3FOmXoIeyP+9cdx+IyX4aK1L6MEfT7V1YequnrhM7VMHh1HyWm3QRnBCcbUG2Z78
6ALtxTSMW1sdBwaZbCxiLYX+KYD6rBGku4Uz8zrxiblmnmRe2oFMaIK9+8Isossx
pXF2adDpH/u1QYrqgxlO2nBB0mlDkvzAic+ttpWIga/TcnXiDnM27Bx05Kr7FCpe
Q8dEfF9nAAW+XF4jwxo0/6KRjRVTnLqDJZlf71f3X2XwbnzhozX9jrYbaMUsmFa/
THgkTBVjjZQud0H/R4nq9Coz/uH0ilqXU11TGMbRXK2foxqTz52+/bdTzA0i5zxM
8h2DXL4uoBJb8TKdBzEWbOe7PRulctrvRxGCs9rOR5wBHAbvIYDV4YGcojOsMDIi
K2vWAAeU3hfk5QKzEmdG6gNc6ra4stNLxsUEeF4TwAMIrnb6tn/A3EPhwexIAi1D
gHlLYs8gGUTvYaVYf5nTGzJfuckOppnRur+9+PqIYN/E5cC+rJ7d6zn+cc5aY9EW
XFaqnuv50EPASSm0i2mQzp2QuZUwj8vChJBgJQ/XM7lxssSgRXboeUQPcFbOOKhX
ueq1ftrBygouSJi0gSvwVaQgS/UzFRkPxtx6o2q1GPU4y4b/ZC+iVDgoxBl/Q643
ju/2xR8WNMPAOwcG1XAsznyEJ0ekITO5wbJLw1jHwt6nSR+yATgfaWzwcnXgycW6
C6esHiOCanDfH0UlPhU3N2yIjkNhThrA3cZlC/Q+6i0BxSn/jPbktKUH/ficj2SK
0yEoXm/qGCGJFK5YPTOvhOLSlLx2WGe5LyMGGYWLaNoAu93CHMivKdqc3kdWr/xl
G7y+NwjAmHDgPQcHKErEzCVFrA5vCQCuh6PWjOzn0bznyLMPNf2yMdREp5Ikxe+4
aYu6tYFExnrd5wO7AIE+FDbJ6AyFzVXQpTGwBFNkDHlcV2mSGRLaHp5qbxk8KDJJ
/UU3w5OSHDZEclj4mtsqX6QN8G83g69ip01LiKkCxtWwG6s9IUm+il9LJM3czU2q
rKxLtxIZg1CNHEsToK7ORmTZ0ldaj7b81nH+jShKhWeEPS6q/MVCaF6hdGwiDmMc
jyEVAWBUb/uZHl+uC/FsNY2ap8W+96gRRbqoR6Nm25mHUdd/iDyK28iImWsyyjdA
79LkpcueaA2HgQvPhGPbml5RVChNkk0zVCLgw+acSo7cc88t7PdBswoL7WLXifHX
6Ux5tbZ5jfuP7nzY08yzmaZx+7OQG8TcyPR41UUYPBZ3JJzGEgCo+j4BtAnVxBfQ
MuMtFZAKsrIYebRGxnN0dOUICICKeV52QkO5bEha8JzJwz6EWugATGCH6v1HGcAH
2/nBkA+dQJHryajLX/MgWvZLzbguEbU8VDy5lCVKoj+8j+Uw3p/5NspjWBKfBjb7
jpbeVLi87iidXg4YkUdvs5IWzFudAnqjmUQcayb1z8c3W9QsJ2tntoFPT91nMZMp
vzxR3e3Lu4hiwrRAYfo0OYTXm7+T/1UYg3GXdJ/tYsg0YyBwdUvXmtSGVeH+C8/A
5RM43eULQ3IN9+0iaNLvh15j34pvDdWSGZqoBd391r215RZn1S5CExTRuPONHF1f
i2ZyApfwHHcKrYk5Sga4PU2YNgKTsS3j5tga1JjcxUuwc4+XI0DBcFnPv4etNGON
EeSRIGsqmPppp2+eWRJLQIK1T0mrCwdtCWb+DVh5a7RzoD0inRhH5wNkMVNLwI/i
9I77p75tJht6JoGbxFOBB9f2l2U8KKYkfWMYT2r+CaNjMCaMflbjF6n47zpuFIjt
U0iQmZMTSoPrInbFrZ0YGg8pzbci/ZcbVPdvLW8lM99QuUUjkHE0gn6MbkJABCtQ
iLrAkIur79URNdaPMLuHRvqjjezp2Sy1SmoYwlmtAHHdx73AUemi91wgmZbrIDSH
IVpEMcTwy+VUpFuzAD4qUWB+ResEWty/BcQVgpKqs7mwrulY2RXe3XGLeI6yEVuH
rjfyH1BJ3OuIDdE5Q9aZe41jgPtQyUAKBO/EAHwVi93yLVD70KMlX2SWLdL7LDlG
sLapUP6BvDTtkkrwT9j8vMq/ILMvBmdnaYgW4GeNlIHvEmW/zy+0A7tOdOfRZyli
3DolOWNpDl/tyvbIvyD9hiyVDd1HCv4OSIJa4i3IwemF8fIxKdCWk/Rv6Q0Cdfwy
M1DR3azGjke8qT8lVglsNVjsMBo/f7qkxOd4BIWaQorKtEYGYj70cWkBVg+Bnakg
uRsCLhfBiyagGUky5eu2b0vJi0Z4185w3v51c+NRC+BF16a530PBRxO1Znoen3rL
/KGB9I0VENlpa0FUeEqS08kFIF4Q/mOEkxrj3Ia0pn0hBpmrRBqyS5gjtYi8u7SH
ijAofqldBtfQ7SdSSRMTkHmkdAF0fIG4vuRh/CX5yDwPIH7yyrkQ9+3G3RKOhGHY
Nr0eOuiQCwMPvkLRTpBuVhg15aZRDULmLXgbd5jf5MnXNVu61/5+2wdbaxV/IJda
zrBdzb0nKXJEkr4fSNFjmD49u5AFOG5Rd5QUVE4oSNkjkmil0fv9zg+roFzLSf7w
9aHwSU+j4Cc+Qgko6KOFxvzA6OaV0j1fVQeEnsxpA/S5r1NROPJe6zDGL6IqmCu5
zsauutC1nUTJuVKTqrZ2T6d5oK5kZrsts6imbbaeymEBoFZZyfUQonuXgYccycYC
62oiY3It0U20nnwMcEBwRoE3EbG3+sFEK8bDVqDREUg3GfScOWgX5cmhmGMDPpS+
q2n++mRqwJz+kS9N1oO2iAsMWEzTAMvvlnsD8hVLipL0ihlH5LYawADfdHQovQGm
S/7RpS6pdJuiS8qJC6v3zA6Xjsp5W0Iq4mzdTWsS5UeUlrAdFjGg1dvS+hYOFoOw
vRGKXj6REXFleMD+HbYOdsn7/rizca8dDNTskbdl97UTVNm1a0E7OIMzGN3cCKu1
4fvGB74AA/ydsBgxO6zjTBaxzMn37WcYTORdQ9SlipVykv8wSG+EG5lgYTqP0nzI
5SSS+d5VtTz4/gjRU7z0A7g5Osg5y26gs3sixNR2DMv0Aa+9G2eK8yIrDXCgQxS9
oRUNJxRv1Hi5IvA2YzyD0zrcRPdXPKvVK6mK3tuR4rIYAVvKxTO6WnqfGXu7UZPb
Tz10OHlB82F/o4xCNWL1v66yvC3Y/BW2sMMa0w3Es+uuZR0Woq/WAkw5/yBQBXys
r3/CSo7vOdW4XVRW0Y2tOMrCM8Skpdrkgmv4IbH9pil6t8NEmWZvKKQKlB+PsyQF
SywHQDM0D3bEcQikDO/UxglIfh0lLmHHEkxbbV2KgHdgit/3JvzMeZ7/3074wBXe
7AjtxKAJsCqZxU0HpoKZbPXc1tJ4J5LQ891tRS9oku2bRx+hMZDhm9JJZZzQaD++
hfJywIQIXo+N/LJU2WFt/T80u7dPuSbKV0Yr/dOQEh3VhK/HfwEm7heXcgNMXd3a
4AjKPR4YSMFaMyFuuI7j2f4JRq5xxvWzYK03Tv6CXPG/5Qjb6i30vPAtjS9lrEfo
cIkSwN1HrVRUcvkpG/xpVa7y2JqCA52YqjcPiyLOhZne7AyF3akjneJR+JmsQBnv
x6ds7DVIhv6uTSntZIj87V8OlRyQWgGfYxGwc3lnWyw8CNIu5rGwUBzKOUl9dd3z
aUeHU6IrdXD0UxbXJyBWGqEXAOtr6tbKazxVPhGhxkjqwuM2aETUfra1ufSkU/Zl
UDHT3HlukBoEutMF/OlyFt8d848WuhoEnw5SNWdznUIUgAdnyfWvTCmxbzkipLL7
AlCT/PkcN+3UGo3RAxk87C0/r0T07J9I7Int3/gO6E0ahU9v27lNs61aEXhV2vwI
LiqZr/55InDAbVWwKFA2xwhp1I4J3FmIcjAoCjh/y4MpOYMgVzavoJ5S7WJvKJy3
rlt/Jv8KCIBY+JjbnV3zGQ5USB/e1Hrq4UJJ1hLCMCqrBUVNiti4CtLs1Dzjt7Xo
DRLfNeF6PQTiXdrp/0w602IYinOQa8McbvKFhtRk69Xl1KseJKpGo99LA6UKHGZA
F99UMvBkxYQiURN0dAHSREeWp8fhPhnYJsVYFrKcqkd6MB+/PgT3eE/CCZ0vXhDH
e7eQyG6q74fCRcxUNNjHKeghcujBZeMsZOP1rwHXExenF+OXkoL9Jk/ZjBiQnj+c
L2E2oRRqHabEVcmYgX+dKHvIE+Vr+alZRsfRa/2wCxycPu4r0fhVx1kaPEu3Duij
vWZv+mGN90owNeQF7XWJmgZY4Cy80mLFqGB/BAmruL4dmA4/qGd5dnFx9rvmUTkO
8PaECEph8D1HHFWRs9tis0CwTy7ob0PJ4gy6IKNTL/emx+fUQTScF2UJhkAlU9Sb
p5Z6QR+bljN19TJpUBPX8ip2GZ1IY+PABYivivgmjj4ya7CAU1QMKYDNhwL81V/l
0S66ewLwZbdtFbhiMDL54h5WHBGnoLgZNLZl5H7+euYzcAGI4JtDpXwzZ3JWZ+N2
RnW55bhMpmuG3ogp1X3Ww9rpp6aBkXt+twdWWyZInYoiL/F5I6RgaOyuPLAtBAch
MSFYpFbfow663++hVJLDgDosetwV1KLD6R+HVzhOAbvO2d46AW7QDnbz29Q38ZC2
wwS7QSY9/YVPCZFFKZvEaCmRNeF1Cl9Z7eBEyoCczNFJqzL7fJNBrP4iBzcOXBTn
GlVtSI04bPYJi7Iqqbo79vgEQWLiH//7lQkhxOTm72s2NZUTV0n3XCnN0Fg1jyL8
qy0ZeBzi1QNeYYF8U7x+YeaYV+RQb7ZJmBJfUz0lujJzMRIhIXuVxbhBks+0XQsA
7cVhtzYYpu2e8dwa5o5lq2XN44Ci/mTDb9ofpHin19QaBaAouWNI9d77wMgxDy8N
IqzjThkLo9KM6mDphkQjpfAa7NxMoXG6dzMdnvQCENQJEcitREOr7JZqxqeZwpFd
hFsDqR5UazuIqiuESnSZPRYgF49mVMrK9TihYYpnybwmiH0QDU/Mi20TzS2rpNeq
KiV1lY61Aqyuc7hDJiLvM3bO8xvRxUzqqeH2PRpfqsxTrpJyb1lkdi4tkFhAwbSZ
vveSyqTmH3fhez7rrtCxkwBx7rLXxmFMSoxpgxnwHB+uOcubfoPJJzL82qDiiH5V
mwuM7Hcu1kS59cNetAlYuIP/ZZ88TbY/NgGqMt4DVQESq8uatBFu2MlEv4MQOYsx
QXhAMjFTaHyTxxhoiaXoS416aN+gJIhM+MTbxJQTw4qddyDznaQRhFeL5pryABIH
xeZDfknfM9TNvUcxF7eeTgp/S9wmOqHfz7tJW/aamwph+gWwSpSEY10lwUG+LOS8
`protect end_protected