`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
ddtXksX2+yylW5zu6QL2Lhnb2d1sD00763mmSITNX595NcHTEkwn0zB1Dry37fOW
FufOhVzEJp80NC5qZ/+F0Vk7Ik02dIR0elf3clrjeJRK85K4e3Hoo4xn7YbFUIms
l/8VZSb14+JVGURjfswrIyCUotIzlzVYZ6gzoZwDXIi5gQIBf/gI+KxNXPaKV+PQ
Ufys/12rjO6aI/pPlqSm0hCvftmBcnezN2hk1UeXgOIuKZnogjOsf0iJVX2aOOWE
6pD/psybjbnsNB6kH5uFTA5frkzIzkzl5d9+YDm9OyC+k84E83I/7/j+rk4L2dah
QJOvksSIzN867/4Qt8qYTQ==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="MvBXkzurAa5VTw+1JJ70nePUfoQXBvZOku/SMmg4TwQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
oRtzZL4VJ4iwysPsC8SXYCzXS8Fw2gtZTOskLcDV+1B9Nzn1zTyNtlo6lNICRmmK
ZRVu2BmCc2G+fmzynYlNTnSa7C0Cuel6FYpxCBlOuk3OF2tzAmLAuDyOH3Z1Yjzk
a0aHuoCdIRKv7BrZCdALt03JeUmXKPdOmIlkVGFl8yw=
`protect rights_digest_method = "sha256"
`protect end_toolblock="Jn9CQpRhJt4rnzZPRk+dOpzAubz7omckX1MrFd4p81o="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 6752 )
`protect data_block
gD6l00tciPUa6pDNTk/+t0OO0nC/UTtBwLB41d4inuAUA3i/ALrNyoJVcBnAmEQW
ptbcNp5fxEUJjnOxnedyZEuEBxWRieZFQnkRdF269oNSMJ2WerVRnVinFdk7F/0i
sZeYdbp1g28gFbrcD1oXRQFCW3g37XY/4i7Z0JxmElVRtQJhWjOrSjbT1jStl91h
tEBwwTZBGy1ZDgx82/raanJCTjNcxodJwlctDIAZ1Hh1+jgsbR2MTr4I5UYoVY0f
hQHaXaJBDIRIY+y82gGSUyGA/m0aMzCb19B9AJ62l3VqolEwBALqg1kJJXEzAve9
a/GeBmVlWENyscnz+BF9BODsXwiOVHgyTww7hyTjrhSY3C5gUEAk+z/iflHIbj7I
o063KaEYgZKJLVpD1S9itbhUArfLrvi/5lWoTi9d04YA39oaHCfa9xErt0J0ytDH
h29zwvpGDReZpal1Wxe2raNZR3xqClWTyh0yt8erGpEYMfgZRhlGM/awc9PmnahI
kgTnQU8wAQoxWlAbb+RPR//fxfT6FNs7bO1y1KAaMHfwK6lYQOIOOW/K9XRYVZIf
L9FrhVefdlhCGa/T25sbj5wJs7PkwhuVeLouM564wCK4BSPo+RwTDjoIiL8MR4bq
g6y+p+24PItp9jrmoFgr7EywO5u1TSKao1LDyw0wzevDIrniissSTz2FuZqBeNR/
XCleRUajwNk7731uhoER0xpmI6iaR3BfZtKKe4Yx3ZVICutewQ5DFOpBz+zNTsyO
l8jnXO37mMD7bCrUNlclqi6bqGZO9wALeMuoWURaTXt8jnr0BZEUKxEWFIbvTFI2
YtF12RRNugJfV7drGxnOkFyo3E3eNJDGI9z+MlBDj79h3XB/K585ZxICFl/+2TCS
EEloJr64MIkAW2mppMjgVnVNxrh7Q8vcaUsoY3vsyhX43cMuxRD7+4X293B/KSHu
Lh48oW+QouoquOk4lBnpwtNj/F2k1i8ng2MASYC6Suxx0/BsKBPAStJ9vjLlCCfR
bL9Zep80idD6HXYckIHyLy335oe1aCDxvolDIovpBR/TdLOh9nd/kenGm9MRL7bS
NqDkWC4fjrgIB50JLnx0jDi5Fh350w8z125FJ4Rc+UjJdGtxxbSF+wi8DQJiHxJ6
EtcksAFO+IfO+J/Ef6vbvJHWfVPZDki5gUlhZHYbhCSrvCjC69QWb53CyCGytZqV
4oXFfRqxwEEldwNNGcvJBqSBn9UZ7rVJfHsFad+slcch9ivVp+8WdIxSZv+iBD16
vDtzQNPXKxUXe8sjonrWLEVTXE3nWuRlCo4QSSv/fWKXK/MDzIkBQo7ZSfyQSzuU
OVvJG8nt99NZt1hCkAd/Dmo0QqVvnTvnwtTexrbgPjxpPXO1r3TO2jl89kg2m9YZ
yj/VhtyuwzKfowZa+60JdF3+4VVDzdO/g09T8B4thCjAxjCmNePjWM87WYKSL1Hu
DXPuMJboyhYN1sya5tOE9bWLOyPnELx7xzRXBGUlQ0a0K57lipEgc2aPEMgqk5ZR
1S/OvjlYGHkG42NJ+cI/BtW+WFoOG+EinBkGDcit9IHSIG+88k5/+U2YNKUbWeoW
Kwjwu+iaYoYIsol1V02vkZMoUbims8fmxN0VtN4Mx6NZK4v2KRsgom1D6lZdp6he
dvbsSeEgUMiD4GjaYd8+e/6OKbdijVYbDwfkf/1CdoDBNmWnftur7S70j2Y4Zo56
/u0R2l+Vj7OPeYWZ1xSknNFkzwTjjk6y2RG0NO5T/dyQlHbQ3cHMSN3QMgiQdT8Q
7Ungs34gjyrWfQ1Zddnrk3WaOXZIwnclM1/ybdmV7LxvfjE0K3dOFrSKEg2styxc
wmiYeyC23NOURRCc2mfDQ+onO7g9yE636QwML4b4IdxoDk4mTUIuocJWno7vjLaJ
IhX00gIavOJcOlWhJAWrcrf7unY5nO//wnaXhZewmBsaLNe/a5x0Ks+a551KJVka
1hYUt44SzxpSzvwr57E8irWWbiZk4cin91Uh/Wjo+3tk7iLx0QxN3QvQdhT0jkbn
+FrWIo0Tfj+XzFI2GHYsUymdMO7vLVFJwxP3PJ3nMwVJQvyYLj//4tSDmr8nroQI
nXZ4eF7L440G073rzumWFhj9LGqDTuq9aGfhhW9EwM+PzZPFn+Xu3zsyZ/4LoE/h
fRmzEd9MbBnmGiTU+vpBlxxT7XuYLIJK5c4h2SguGpd5VM1L/PCHycmsOkVeu5LS
nRbprrsOKyuoFBqafnRO8tITCIcT+Gr+bw22hGcPW3yCa2Sg78qTVrRqavufIFrL
3A7zyJYfB0Qe2RVjTah7qcT4onw8HdlAYIZpVMtCCnf9etbkJQFuW5PkHrlONPg4
uhE+jfQq/vBTapPTAD++t0oizVWJlh6JcS6ukPmvftWdjtIssuN6d/uTAEOlzZzC
L5gY8MZVbpPNk8HQ6jt0Y4N6lr69qDJUqC21kCRe3Sw4dcIjWvwqytB0Jx6zK/J2
Y4Qvl7pSocU669gk4ft7cPrBSapPGKXVkV+ZTPWTjy6QXlTLKbjOgd99LOYnZBnV
QbLylJHJlC4LSU5es2C9bjXL1a2sHtLuy7KYvf0o7FSvLcvL8TK1hSAcDuFWIXRh
6979kKisrfRCokFBnew52qq0VGWGoo7iuAUzOr42Q75HraroBbiVewfC49kOUtLX
WQlhIMvG+LVanQTY8geinCcl06RceFohQLtmpI4ppkHeVqhaszitrE1DIHyP52is
+oBf79GlZV894vfwy5k83YhnT34+b5ZTQGtTjwBFeGUajNT2FSZ7+bzorJi7m9Qi
vX9TwTZIRbc9zQ+N42Yhs5r81xrBsmwZMn5F7tz9SCs4tbPkJ9M8JpUq/e7nQbu1
ufpyfWzSQT+vpUUOSJoGAYOjUdBwNA4xv7ZEvANeK3imYlp0SDlnyeFmyciI0bis
JF9toaLsTRFc6BJ60uDtO8oXfHTd0Ap5YvsmhqjugJm84zv9ubhkNde3ZqfdINrs
rOGYsHjnL6ZmmjPfO2ktitwZkYnOcwT5liqLOc7ESSSlT2qQkB7lGV0AGnIXPTtE
uuNaveL2+s8mXj6kjSIPs4g8POAqgfQIwdIwqAnORvvKl7+8R5+7pxCGMa4jbC2a
z87kXxfHtvLR8B6t+mJQ5iB3LZ/oEGZpO8/12/U5CbNSVSIhQPB8DcapMbxNgaFp
Qrr7Gr7FoYJlGa77DbWnPvA0natcdNkTLeTOzNh6P8aPYRQTnVVmLe+6yZh9Rda0
5eo5jwwxl0TxX5jy9y8N65rCuyPJ6vviQlOeUOx0vY2LTnXTj1KWNCP6pKKuwZBw
23bOCjnh0Hg0Cp+6fsNH+8xbOTLDGU5nICENe0kaVWrGE4qAMhprG61Y8oz+Vb1n
4vcncNr5b05QNPIPtNm3W2diZ9Bw/gbpGe95afvjmhShVifGmboHpkSCLVHNO0w/
ibqJl4cuNFvlO1u7Cv9TtxCGNCz9vzVBoB8f3aOc5gGxYrW5Q6bbfN/OCBGvuxJ2
6/q1QdqfS20x/xi+psl0i+TGxLaw7kSf2HWPsf1Qxgr50CzwGurtpXO22MH8w7rN
ZKH6GKsINLb5z4d8Dqp+L3Yd4graS2FpID5X1jgsGqROe4JzGTRrgp5Mm3W5nPzn
lOretaTCgZZbYUR6MvrhejPaFskazOYR67pLBsVL7REPAV0pS4VukN7WWaFHBNZ9
/ouLLJDRsWH0jTqOevXqLEVQbcqkZUOFG2FEC+WBMef4xjK4F9W4NEYeeCBFLgK3
cDUlYidrOGr60ZByA/jzBAGipZA9sn9JbOKyHLaMxeX1k94JJfpelzeDrP+UfRLO
1wKUhrmrmcaH5DohXuEBZj9Cz3Qmu6vgd0QuJnqVluxyMdFKr/BeR6GvtkMFcziF
awpWCky5hqb4h5NwA1fDqnC8z6QnJIZELIc/CcJqjWvsaA/Cl7Hwvi2CdZIF1HCk
j3M46yVUUbodOHgdgO9HjzrKMiQEyQpxJyyhuY1oXDsnjsza97KejqJoigm0ssEw
y1S414V+pj9W9Wew7pQnHzz0uuh4a03GjEFKz3sGQUaIU8OWHyClpaVXsJcC/2Ph
5+akuLYa9dn6iqP21XLWY4HzsLsFkwsLEjtpEQUqbrR3++Qr8TJd27SpEz77UJQu
kAcd+758FXe39uahxhZhbT6THQujqEjD7RcbW2nc4FIXX0rWiQEQtbYW6OXIUFW2
WFqCPQxwfabw2ZZ44xRTzZUYx8mYxBw3KeldkyGhxg+1S13bvDbwUDLLdre7WAi+
oXvKXduOk9PjZ1cxWAEDikjV4jf0QQJrCpp32wgJgvL5u66q+K26jU3n1t6Si/Qv
OIcqmuUZZP66cCycVPmB7PhCDWJxwA+FUCwYIqS2mi/y/L0GQ5VTe9RL2uH7VJnO
oZfFKF/+MWbbu4NG1SpchrZtIHTBHhJhRoxQ0ZZtPf72tOA94ZLjZ/XXiP2cA6QA
lsLYlit86QgEAgJfsAPjF7AfowCpAsmXp14CUyhXY2kMZnigZ4H2a7aYIIQUy9S1
rZ9Z+gX1m5wbLI0/ewf1YXsANQSVGUuFwUemU8RV4ziSUktZrImfaMWwMEBSIY1M
ksHWo7/efOKN3adIvEBJ7QpbMLP+IEoRLqFDJT5iY7AX9DnKqDs7ojYZ7rgzMNVf
eWsdT3OaDtUcYTPodsgMktOTsWEg4WCURQrCGjhh/6cPHrtumRwYbW0S8Pc+VdaN
/azGp4t8A6ZA6c6OykRs9Sk/Ne379Gs0exHb0GSvfwBDlkVxiFg1nDhNbbu5W+TU
wN8/yYYzLCUIIMgV858jWLM5Bx1AioGsZIll4sYAHDwyCAjGglz2yHbQ1JL7I6DH
aDLTF4DL/iEJ6lkLem4Cjx5Wkl9bbfNiSzMGwgRlB5Xc7NLwQJg0plGBOgOPSO7/
cepepqlu9teNuBIG0TtK5t302uazGbsJ4y8VHkW59nYoM21xQMQZg2GG0b0oaKWA
s84Ta2YFo/hZErAo3pu+g9LnQti9OJnOvfP3JrL7mESRX1HpT/W2zdZfvtTrkstY
M7NG73n3/WFPITYoOQshUFVXB43iZwaoj97p1EfkfyP9hoIZLz/Cb4xtwiQiMfe0
vbyeT1J5b4qiV88xyR14od39T8MxsaviiW1hPbrQIu8AD9toUJccZTbaxsGd2byC
7UOWVM+U6EnOjiRQfTaXf6avfVLEJivmi/zwPERWWRVHDYfbSj7pd6qKnUPpfA2P
En7THAcpJRfclUHAZPcLBoCgABgiq8/EkzHsO262NLA3OVAAVEtU4GMvTLDS733A
tLq04ZFqKhR3kWSqbnI6fnhvtYD0RWAlhV7Mdg2anvXo2aUB8XoT6S4/0/E7fa44
GP+oeGjdKUCSqIc8Wy2AmpZDBMFUaANgT/t+2gjHuJWeDu5ApuNm1hZKFDhn4QFY
lX1spO+/OvqSELpDR2/bkxVhfUka+gO2WoDrTbkFhbixAvP79n3vysFk5HZyKsF2
xL8/tJ00XjBF6UdhHvEVXE2fZjR12SoSHCaW7ddK4saZhWSJgYirzRr7GYj/pIu8
4ORhiyGPm43Jv9iboA8ld9dJGa5dr4diTUJsh9KioSIK/oAMvKvrLyWZMN+hSUGu
pD3fO6SrE0Kq4/FuPOGA8yL5FjsRa/ENmp766WbLm/Vo7rezFPUre2/7KxnLuUHf
HXAMasMkklL5BlAhF1Iv04O6hUB77x4WFtdjbzpRTb9+hnpIWMOVajf0tgRmmcMX
jF5PHged2H0m2lK/FAzAuUEDCQIJrUmmjWeI9g+oqL/+UAm9QeAxw7r89sQqgCIW
p/AOZyicEkSwGyMgJqmTvDqoeyjLbIkyThsZaIIzQNMinMX70Do4gcKoeY//kvq9
aDWMEhOoAuo09OahvY6TIEJfocvOHs4FPKNg7riFG8DMVb9jqiwGb0TUcNC6AYdP
zdPahrPSy/78Y4CvD0PSomZOd/50lpjGpIl/oMmhOKbKblbFozXvrUce0oDIfX/k
hx07JxBy8Tb+Wh85GKn1lBq6a1eJqN+ZoodGjsYf4LHuB3GcNoOWeTtfPQdqI6Bt
LvJOf8a2jznTAUEaQzLoqGLpEFOr3jjRxjQ+hyRqMfNgtws7MB2keJKiIkOxB5k1
6//qco4BDdLYnpKj5IumKZ52pFH66NrxR8ybO9Qv1aJQAXaV9ckTSlvZLbHisBnc
N5lUOs5M11sZTqy2PhA8S5y0arVqgOkRfDkBM9Vt8M0m3of6ThU5j7IdhKNWvA9y
FTUPLo7S1y1Bb52bXHYwv3aLOV90z8wZ4kAPRL/wSF+mRRC9lJ1/ktBkszzVHHcA
VRAFeQd6ZlJDJOHc9OeF2OTNwsi6VEuvR5zg34f4pNVqPtg5zUS44YITEhOhmVVE
eEYuV43/LQOreDn/VieWVqRBrDAD3XWj126xvyoFzat+AX39nOQzYjRlsnhKXbI3
ExLoiwuOhiTvgnjleVUGtwUM6cPDsvWNZamQg5O5shGIsPbD2ddPsqpZ7TtuXuQT
fnsM1zwDao8r2PLabnWNShjGQSXt/9c2GtVwUOyoWliwQ8iglcgoFyGRkJULq2GK
q5dFHeXcpz6AQKELUnIbNkgyNmtpQTslFX+LkwDtm26Qo5XaWbmKYh1me6YqzcQX
BdnrdfuPiqZL+wNrYp2Ji0NmJyLqs9wyv5cY9EZxbm5gdPm9mq8AQKIgRIou1kwe
1PG94QvpCY2nNTi2KB9k8kL57huC3CP5YQ1hs+m7z/qDhtsXpSXI6722WGV6IYEP
fZlsSKMDGeytw/t7kXHC0cuNtW4Xew5gtKtifR5ppoecyTznPlbKLj+XkpeRAt+6
HNFBlVTJiZomoE/816ptWVh1v+94crYxd+dzyHSdkBv+nQ5HG/zhzMwM/nZ3tF0B
dV8amVvVIt6CkfgsdEbQ2LJ1GEdAPSrl+kYE0twICXmv60XA1XFJVC3SidCtwfMb
JiQMPCgApQjpKqB9WZwc+0ZVlFlszml4QzygZeLfStRzpRAMDZKPpO3NAq9tAuAD
gied3qMkq0QAsmeY+mhBZCaalnHdpwWqwNyZE10vNlkR/J7m6m69bTcMgtsqFxUO
GQMFkcJlkHIafqajTavFG8idq4dTZTSqYjdoachwr80s5qSeWIDCi+Q9TuIcB0x/
GxaiitWlrXPgjYFWQGqMbDnnbqzVBbSK/sPj7g6qdj3zKi2H0DBhiYY9YTvZaSM7
E8v4FLRYME+kE59acjdkLtg525LGkhC+/uui7GurpKWapIorHTNMzVFxHsalnKD1
xcmE0Ow5Wig8FN22O1aTB7Tlv4lS3/8x/SAittYy0sIAXBNCWBQE6KR9Lyt4Dn/F
LK5dThelfEDWc4+Cas3A3ARO2q+TsTeW9BSixmsFwOtkc7k6y7qrbqZ3xtozescf
nzFedBLxS88N23MdwIIJkpW4B+IGD1+o7/5I5kDAaT8l+znsNNYhs4/6vOZRU0o7
l9p3nVkN5ECdsscQjabXRVDVHks85n/MdlyZ6nQPzBJFpimJEmSJUzKSx9J0Gyfi
mjMm0g00cGgG6Awi2VN8CpbaXbsES3Fe/ifdvexxT0fhjDgjlZEZgIG5d3I7HySn
SytYLjKqAs9hkPS8fIeRjS1dQ7G5GSfBimOPdlNVx2ouV07xdx6RQz28HtwPIB9y
wiMOpSq4ELCt25NpIjzNGOqbpaGJ9KMeHdpgBotEXY3+3LApclZxf85+ndazV+3z
o3ZJ0qow/icUQumdSUv4tlRT7rn647v3SeNWVvM/byDwtLL9ZIsZ2F+NIhynJgpI
G1WkhvmVUehr4BzD3zRfP26HCsN9wpFNVD7Iedwp++LmhmxcdG5c0/F4zf5F8bmA
64bT8X1QcLzFdihLhvRfMwdQB5CDMDTjLpyCNWzfxpL28OMKOQ8II+hDt7z+6xlB
prJ8SYiKgOgWnBIIhqshjrX5p/AAxEjAfXeSjm6dqBFBemhka9f+z7V4KZGVdN1W
Lons3+u35cGXdrygQNj2U0//fD9Ho7yx7xtwOv8NNbJD5kKy3bKKokrqjQg6Zu3+
ZZ5Sv7z/NBjI3EBrfuYoTLv9XKImNQAO3r3ydw03x/UlMYF/tFtNHpHiVOnXLdCK
kIXlHWvp4jgXCaGgONmNzqOPTXm/hPGJK9tOZL8vLVMt6cALxHlq6fckmTd05B4E
cZoZUCQ82rfWAC4tx3ygzEi1hiceea7D6k/SoLY/00rIwLbUsVFEdxcFYT/gFHwQ
1V9zVhZ5OsQ3mwtcvJxGQ94D8GKU5fGcpxtYNViot9rS+yBqQ9iyHZu3ORkEn+9F
BMS4pMZ4IZagVfz1ZG6n112VdAH8q6RCOPb9eS8SqGGOhZeE286LZsSfldwvdp/g
0lspWh7v0ru9XlfvOfTSbZTcKD5aAjeGc+Z9Ee9atZRJFJVowr94kEiEPtLQMvtc
N9pMwzyBvyQOtRSmhAetcFsRCbQ7EFjlQCcTbvjGBUDEcrItRjbbMpgXU+Fi51N+
7ZxDtUR32vpcngbqvrW5nGuNUKoG75OB/kZr8qJv3kGuU2e/LuzlcvpncZ3l3BOo
G2CfPzxMlnhBB3inWFQ0sxUyst5fTv3G/uCnumWi16hi/wFEIkDCsu2OOd5fJBat
ZlXbJHGiHklFk1wOPVx5PCjVZ9SMxGCq34XgO4oHLUlaWX7SKDQ0wW9VhA9FLhg+
kSBsMKNcbReJRxMF8XIkJUOT4pgrz6GH0B/bHzY97zEapOj5jQYaZftMCwYkSkQj
ITe6M2LfUhg1sjXtiZVrRnNp7G/ERJfjV2RpK2QEiPQwUnZrIFJSlw8ZcmqwDXJ9
PM5RtRKQi1WebWtYQzYfUK0k93LypFwad18ADoBHDjPha5/i9cV1CKP/LUAaHbZ+
xnpzVgUQfaxr6ODN/REL7hoAXW8y8KPyMDaxx16QwgN6uoGjDqR8h7Vyrs1nkAoP
lyRslDaFJAjmWeRXHZrgtEleq4Fbp/Wg+NftPXCRwDs=
`protect end_protected