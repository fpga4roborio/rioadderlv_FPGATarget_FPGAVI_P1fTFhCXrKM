`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
ddtXksX2+yylW5zu6QL2Lhnb2d1sD00763mmSITNX595NcHTEkwn0zB1Dry37fOW
FufOhVzEJp80NC5qZ/+F0Vk7Ik02dIR0elf3clrjeJRK85K4e3Hoo4xn7YbFUIms
l/8VZSb14+JVGURjfswrIyCUotIzlzVYZ6gzoZwDXIi5gQIBf/gI+KxNXPaKV+PQ
Ufys/12rjO6aI/pPlqSm0hCvftmBcnezN2hk1UeXgOIuKZnogjOsf0iJVX2aOOWE
6pD/psybjbnsNB6kH5uFTA5frkzIzkzl5d9+YDm9OyC+k84E83I/7/j+rk4L2dah
QJOvksSIzN867/4Qt8qYTQ==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="MvBXkzurAa5VTw+1JJ70nePUfoQXBvZOku/SMmg4TwQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
oRtzZL4VJ4iwysPsC8SXYCzXS8Fw2gtZTOskLcDV+1B9Nzn1zTyNtlo6lNICRmmK
ZRVu2BmCc2G+fmzynYlNTnSa7C0Cuel6FYpxCBlOuk3OF2tzAmLAuDyOH3Z1Yjzk
a0aHuoCdIRKv7BrZCdALt03JeUmXKPdOmIlkVGFl8yw=
`protect rights_digest_method = "sha256"
`protect end_toolblock="Jn9CQpRhJt4rnzZPRk+dOpzAubz7omckX1MrFd4p81o="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 47856 )
`protect data_block
gD6l00tciPUa6pDNTk/+t0OO0nC/UTtBwLB41d4inuAUA3i/ALrNyoJVcBnAmEQW
ptbcNp5fxEUJjnOxnedyZEuEBxWRieZFQnkRdF269oOtsEi6w9V0QqevHye9BASm
04Tp/mmkRsUwGEQX4sso0Q0a5Fzs2/zSs5WiSmbIApSVN5YRKFSSlERoK9gfh2HE
1IyUH1NX+BuyzFbA4CzrF2LDhbelYoAoHZWJYTvEweWurdb0V16hRVz9Bb0bU62e
N8TiAoOJ7sZYPo4iVBr8tGl8PlGnFgpSR5YC9FUjqCSOS3QE+qop233d1H6zDuj3
8fn7l9S2ETp0iEvkGDQnhVxUdm1+4qwYwaR0kbM194Xu4X9dS32vuGx9C9C9veI8
LBt2p8GGP06lfMotjAxjYQeGViNKQG13GwYRKqXruGUAngab+ZiSqwIkRMw19dfu
f4/r18UEmq6ux6U9TcjE6vGawQhq22qSK14XXlZafHQs4Tc4md2rxOWly1QjpDGk
xKcOMIsMpzP2VsQs3B2z55iVZebXp9Qv8TS5m+fAULsGD7Yf9azvWbqCj9/yO3sj
F3Xn0kem08FFFLqPBVILaZCUcS9bjCPnqi1MAueknCFJjg6yORcBPM2LbUt27wT+
p/vQFOaFkZ+ybpmgql/YB4tz0iQOWp2hWPUw7gYuqxEMVLEh503W7OG9+SNJbf4s
kKX2rdRf4s/LfoEo6QepLJtNJQMunsC6MUGKDg2c+aRdCl537yB+i+ZrGkdYSGaA
BDhJTWknHWao0XGdpbFqZ0DA/VeVBTNzat4PYNegxnabXzPg/maQj7HdNG52qA2V
L0UR2yYoLpTEFcoNenFVPAsB+NWcZjoUqRiYHmLTZ1RfyETXZMbcSs8dJ7aSdSsL
HriBh+EuCbwQt5acA8VV8lO9yhzji5Pcobv5lDGVg2XhTEG+ZoE52bj7LknM7xsj
8ajb570bgU8NrfX1g5eGm4cBByFkoqAEX4LP5arUuiTHYKDrkrF6SZmjtmWeajpL
NOgfSNFb8VrXwRbUyogVObZqCDbfG7bK9T0egYl0iAsL8j3UG60xQ8eI3nd7GUzV
twbWPF8In6XCb/0w+gqQ3neWv+IHDUOLGjgYL+OXPbXS9RxaVawz2dx4lNZ0/q4Y
sXW7XGIvLeNkoOM2uX8w7vDqLo47LPNmjDaaLk2N4ke/gCsAC0Oh1dsm9bofnwic
LfEr/PGqj9HO9vsIPLUZRti+bFHSswH43bQ94vE8UQVMUo+GJ7WVO9nGEOASdv1L
w+k/df/nT5PV0p8igCKk+Vgg6DxPI/k0Q98gKZrtGoCJa31cruEITkVWhKMzGoO4
wm5Q+e3PfUPXuXj4JnZryN1U72exhlWTS3qNFaiCEUpOgpFN2IKh8PkuFNb5xrpV
mVLbVBitPdwRHA+3WTpk0MI0yXA5FUWkRMZcL0+UWmphpZjMkzdtYSNiP6MOx4BQ
X8idSNmTMW+7D3J/2gLDCYcjN3dWsgIHDNXQgwsjY0AQ/X8quSQKNUSYPYry1RdC
BCkNXRZIiB3vdLWXx7gCbEYcT73JtGmlj4NhcP540/kbEwDUNk8NBh36A0SZLROt
eg7PxYRrumtkWjSUtrMBeISQcUZxjRLANk6OG0Cb7BoADUelkvniHO0DYHDJeR/F
zw7uC/qxt4UuDNPAGni4EYb7/VbtSVzxPF+++MANe/zQxib0+7/1w58jF0+87fYv
SI5s3+acJbVDQPmzI376G4JbY7OuQQ71TU8JnRloyks4mhmJlylU83y4rtsO/3kM
kOZ26HndZhqeFGQsRvEmENn8bYZcw2qz6p1a693WheIgxmP0LZ3J2O4U0oNZzfLq
B4/Dfo5XLC5TPEsGo43wnOc9+8QHtNPwUzVDFzQWtoDUK9BfwRCdAPT4dZrhCu4M
zmn78ApniaXXaFH2hXJT0RuikJ9uvAbSf9NPQV3eRRFtTZ7uEz1HaFg7iAFOpVNR
CFkwsS7S3wbuj585ROVGjmnyug9dXKTLtognSWNdvYlW5uPJ7bjkjlfl/EGbc5hs
QfBN/GeZgpK0biqn7Ru9xOMZHm1id7PnI8Hmin/Nny6tErGa3/ebGku6ge4hp+HP
UTAEOpNHhkN8c9z+fdeHhM57MzCoHNZb2ajT7pz9DJPfTtBJAtMDWpf2r2L0YDXp
GETH5VlmVqZystrV+EuGqcVSROMjrz+dno2eAsi9iXm/mlXENyZiNXIFd3tkWSKD
JKylvPFjlLbf4uCq97R/zsgBB1brHstyBSwaXW5qO8F8WzOIRBS/3nJo9uFxvCIF
Tl1g66L0JyfYWPfly22KmAPFSc9di31/4b4dIzDdMAkn6vj+s+pcEJvXzcWYQk6V
miGBZAHmqk3JCZAObRph5rsTaI/8xztnwwrbsxFh2LmzL9DKPUf8zC9/buKs6P79
scWcwCO8El0Fy1x6IIWD0m8hhNJAamyXJIsSpola0FbJIN0bkOV6DudTaJp5WKwL
X4clvoq6gI/5wgVUnIupiqb2xkR77fzNWRSyU1vOh5cBr4ClP87CBeLK4VxT6Klt
l92NvshpyD/VPK3HNqcb1SHvHS6l+snoEYlOzmp0A59f4kpQVVcTaG1bD9eU8cbK
TzCAsbQPbx7nTu3JonN4PyPGx20/JiMhVCGUVGQfUQrvl+kEHiBeZjF0B8nQMjyK
gygDSfrNm1UkCD1bOtWKhn0M+uGYEYnhPPGgnE5VTqvQUKuE2TL5DfmdT3UE/9hX
N4pgGv201b7ylhD69DKdIfoqlrb60OQ/vrLvOMqBZYA1RPCF81Z061B5RZs3WbAQ
I12l7I1sI7xv6+rcmwId1f8RwynoLuQAiTjMsR8ACdbzUvq6Hf9Pn+OX6kHFenc9
R/ze0iXZFHkKoky+9tfo61YNxw4fPn6DIObbg4UcSKtrWXgBZbf+u9j+dTxOFOuM
vR7ox342n3FBn0PZvtaUsQ+tlPY9T2DzArGZxlc/jNj9Vv2WbEJYxREvlUHLirxC
IlhHRFSx/+XHGz+Y/pwrNvpZpvxXXqjEjxoWRDo1tKavOxqLNjzjwQPNqbjYfrFG
PTzRiJ6wRJtTtUZnr0DvFtW12DCIq8LEdKwuem9wx8mDg78dQa4WvB95RHArHAeO
NpDggErTwLJqNnATbAigjUUcPirbear4B05CZPMYsEIGoDOPTLEuJwY1mTMpaAqH
UD833hz0AJNw+MXrpbjgAjDhKMGf8nEyKMkRGL1RP3B1DWykQ0jGCgqGWD65idom
iHqU7vJqP9CKarL9cHC1OQZxFbRTcH3TPa5Q4VXxixt0PIlzS8ObPFiN9u2JOhkl
8nxUrxjQgBnwx1LSnjPlP7BYLUcWUjYJrLuGrFwlBUsF18qaiSD4vJWJVfZZbLLN
ZAShUt+F1LaRpszSHMQIrvs0O8dME2wlhw3fgO2wofKv5QUD0Un/PU0Je4gy3D1K
qAL938aUn/XjamTwyzcntN331RE0680vzKkvjLgEhChFt21OJZgKBXXVUnvgPRkf
70ubGDC6fdskeCSpPw2Fc9VLFjIY2RX2isA3XKaK2Zc1QQQCQopv3STBdsoQUlDH
wFyUpZyMdCtLx2yLO2RpsVRenjX5HERf5+9p/QFtInjuVuZ7QnRQd0IXULdQ8mzZ
10RnYtMABVdV8batKPbrQgWmJqkYv2F2E44r9tsyY1x2EKut6q4aNE3sWDYh9rB+
+0U4YjGPwyJBMqkOVdJvJVyg/uUXKPVI9xbEYCtr84IwDCqVTOaWT2DhUtFioWvT
UeuuLZNy1Fr4/2qHVhqkGy7Us+Tng6nYd2z819j7/4goOZxfkHhYjwWonLOjLjUD
76IRHq6TmWqZhxc65o0CL0ZeMY28Uyzg9KcqfYQIZteElk0BCcVw4d8AjSh5+ANq
PZimPVugJ/YeFbN02UpPNzIwev4yWuSKg6x8qSr/0HDKPu+QtED9X8Mae/VFd+ua
l7gsr6DX8jaqPaVUr0xtKPTiR/oTT+9Q6YuOJVuM97XECgjgOsUHIfZfBeXFKmO9
sLnUf7eiYhG2ARxkn5PwxNNt8s6oNpVca8+k4iiEnZzVwVZ2TBl8/49PT+PpWH9A
TDMZ2pek7jPmoHcHUN3dd7tkZPl4s5Www/KLzcGqbWm5a5eXqApNNBo2luWh709j
xSc+lc5ta3z/zNaTS7AJBKdah8zVkyA29J3wGcD1Q12FpNgweL61TGUMihiyaJLG
iJvZbsz2aL/SXKTO36fRvISel+OIlgkceo992RqbMFc5IVbklAmZXJaoeWF8Gm01
YRADCa8JyH2nLDxv5nG9fHeOIwxrTiAlt6KFPu50bgQymoYu9/X+kW7xuGvIt3WA
noR2pO7UfqxFA1+VkSgKDlQTW4pr8iqH2kpIXK8XfGNfkDNNssOWV6ZzG/7gF/hD
QQ3hGSAwouxZf9EBiaUgynUyNKgIvjLynAVgasbta7rMA+nEE0bFpbvg4IbrbN2V
+EiNTnrhLq0qp97JaLHIXtut84v/XgF56jICfawJ7M29OwcV8GjIFhFAODBCGWjT
AR4XbR5w+vRd1ULIjDWkQU3KGpC8204Z6NI/Bs8cmDgPS8248vT53Z4GKKWy9iL7
uCSSduKhvFBvvM7Iy/Zv5DCWs4zT5ZoJ7CzHYe6exvHy2gm1IwAqfGfRUT1IfOgc
H7TH9eJ37T2FC8mjJ8qqc820K3bj5fq+0yDX/NFDQxTqcyzN+vUwBN/GmfIAxT5U
Ab2HHnBiu8kac24pWibhinrLlFkd5Ug23A8XfK4WYc52I8UYSanf+wINNrMoZqaQ
UCl6g6CFJlwkZq0IfVD0KXZjMlWel6W2MfIbowD8eLqO9b3fRHd6eccjDBtmoXp4
eOHW/SBq3wESTcY7MdcQIXo2QiPAEBOuNaBIZGVczB7WHwhDEq8kgd0eGPRe4EWa
2E9LOpv12SyEqqfousJOIgWRMgeVZCrbOUtsp7d4pylkGrlXsT5DG1LwXncfdRlB
4macgfeZVgO0jgwyQgKcdTCVmLHyg7ia6VgLuqrlfGTYhHyP90aAHXVzrLFlJnD9
lULgTaN/cYg8QIGLIPEx615htOKsytByEDrbmnno3nrJHHoCxYIM6keuirkEIPMD
7rskmJQsWjVtgmOdWTtPVQCyKObMX5JSs7k8mZOhWTcc1zwCJrmHzEb5udPAezut
BThrAN3mL4t6TP31/X9CmOGBT+wkmT2TYYjHUHMorXIrpamHJzpEl0RYUN1e2X1K
PwHdHjMaoDGltVyDa//9gWegHd5TmW1oEUXjR/r7L1tXhfVQdHP6jnjYmGQo3x64
06OIbjt4TIbQzAtTrpe+s75LqZDw/+TsQcoUOWaWZUwuMpReW24BACKig2jV21FR
KO3Q1tKcEPnIglyu2xO7lEAPQWBm45bUzbR3SQ5EjyyCAJ1MLaKAOdkDF60dYyOE
QoyQw5Uv2cY3kHbPmxSwzjDHh/V9/mj1ASavAk4vk+aUhtI+zlV+fPuqZ+14vT1z
uLW55Hp0tLYmO4P/8w/Ct2xCqfeIQypG8325CVsNOW5cwcTVC5OOgQRHAY77wlWD
sEAZWpYnGPav3v3i/gtaXpWTcfl729VpVT7GbBxjWxVUxG2Nc31mK35xiTqvj+li
UNWYBr2xfVt3u47LI2GLbqLF3u3FsvaiG4yHcIUKh1e62kj6VERWpdRRsP0udibW
ZiY2p5hEeRikEl1EnqknPQzWI+ytuExdWtSY6weL574damiTz8fNbW0mistw0Dej
5DYbod5YW424a1qMtIAlIC5agyYCwVqQjDYwzeUdsB/hzc/wkvWNykF+VfB/OSBD
kxlqHY8o/bEfC7jWvnFavkabFkna1uK4AEA7wokQ6iGS0XYnFDO4z65NRGgQNg3s
IN7HkyTqZ/9kMLT1ythUUOoVPCoZkOMEHB2lamE0b2lNdMP9clkVJVhj8ocLKb4s
hw5XGamHD0gyKPpnEn9ODy3MivF9bZEslzMRXFLVXOmvq099PfFa9qBd9wndhhiS
4xm3ZBJRbVTLsUs+bTejnsTafH/Vgc3yfEl5NnKDFSSlUuW02HSYdDIiedGvWDPc
Wkt2NXTZUQDJWUcMdCuIjqzgo0DuDVQEocthtJORaQJKGJjpzWWPCV7GHuXdeAc7
kJNUQIE42Jr7OvKSd+plsuvLjO4XaDYkj40Hy3l0j+o/W8Q1Ys6QN3dcagr4piAv
dqotpo4yHUx5gzkMf9I2zzAWWrFmlg4cvuIzXoB5VVN3xbT7Mddj3D2i+wxZyYJo
Yp11/R0EYBOVXB7a2D2W6BGZu5z5K3jJ69qkvFeTsMM+5wONJtUQHj3rBj0jQ2mP
hPIsswVb977KqhfnQgwO6vVYF20xOV5YzuPjWJLETeURuyDiy1b6DhD8Iwnp2cFz
r2ZY0oTfF/8Jn1aMBR2HJs8w/6lZo15OmVMBaZeHYmpucme3WZFsqsnpuASRuZ3U
SwqSl9LsWxiTD8EQHjrjcr4BOIsoaOoSQSDuGHlZCHLZMzzLHq+27G3UtmUR+nAh
lH661+cLa1vgqsi42oe+gpljxiY7rWgLzNNUum6Dl2TlBR7mVjBmhtL9Ce9dm9tR
7tb2IKDodjhKWQNRIIeWt5OoD26w1KUAng/imnE7JOPtiwUDUXPdW+oxWz9iaNVR
HmVfFHrb4f51Pn/hRyV2jCVbJ4UVwDyH0gqJUhM+ryv1S6OEtdLyvaZSp6HJQ7aU
KsLAmPtr/kOmhLAX6d/QdRm0GmmpEgZKAYvFhi5zWzMuq4i1G//ALcpOxonzJqYU
ORxkmD7FXfhOVDV4WrEmMFXiZ612g8/EDXcqBT/Jwl65Ajyp8JFdQ8Iy2rmCUTA8
L1R3b184AM3rBrTMTpTVTjNAP3a0kDXBaqy8ezee5G48pC57SIP3WDk2I+RM7tIT
qtvgvOvJ32RnDdHpCSu20GLrSkvgVzYaKRCk1zb1fOwTOpQoy/CLR/RAD4Ygzaz+
YAPHZHbTtWSXA7Yzb5i0dnPOV2AR6t2MqnUV1+SeLhBjK0WFWHlpha8KXF5Fh+B2
/j+ok78yUzWf3EJymlYmPYnyLAEZb7ODslMfIhV1mIhmVwYRNccRjjUiF9PajOfP
2B5QsvhVR/NtYGdYL3wEdH8kr93CszWk6OU7r2dyG4gN8yr+i38Bz2K7KIq6KfJM
sy3+g2ly6Ye/h2suVqFDI8GKh1B1Ol89oJAnL/6g5dKDYa9DVTCCAL1P8hgXTbP4
2a81SXgaH6XxcyoIurEKcr3aDyLirVZnyfnHBMbNpXdANJFIU+17CgkmvIh2p6OU
ZxZwyRME2SbdBPDx6FxwVb4qLXz4uCToYlEs8WYdzd9sbOjd5gmzeKd7uHMdXD3A
qqye39UfmbQV4dr6emeUoDewwa7lJM8tEOwWs6zKbH21AUIuZJXtaa9/RrLGRugh
jSbpSujK7VFdvRXZqKLNkZ8Fbz0Jj0oMqODNIAmm2zt+tzFaFRp8Ti8nAmKP/gWq
D16WPQwtWbEgiG977Ul3DArAC70TZdwjGLKXd/p+KIVxBmWVYUO7CCaotQ6fQs06
3D+ZccRnLJSjOzokmXvPzX1vUY44l8k8iqBMnRbOHEry8jp8qetWCfeKAOtJicki
3OB8NfludCG6f4yUGQ2P5RrzRpd5gkeg+H6Dpqasc2II1oEASJjEaV7NN7AIwGHO
uQgsmF8VkVnnNyXZqmV+cHV5aCll3rbS4I3LW5MwA9RU6NSb/IcNR6IIGcT52oni
4HpRMsxP5xDn7ZxOMyZYRsm+nhVrmBTEueLGO2mKxyckgK1GwPdmPDtoTHVFjbMX
6ye89kXVbMxeWkZKVFaDNM2qLMQTn27XjgRRhZgJ9Cu6h+srtz/m0LoetQcwhYET
OiVrOh1X/DzhUfbq2SGTg8aDfpM+IJ3t3GcVB9dgeApCdQusMgFB4urv36ndRh62
uqbciFYmn9lfblqpINR4kwrwW5w8sn15WAgU7hYn/PH3F15q2kJ/2lucsN1EzQPD
iSf9RSO6QteVRl50Ic/dFe4G0GLjCAKHk1h1GYgtzyNuVQNh+srFRh2aONIv8HKJ
OxTP3QnJXlrX/AEqq4WQbue8+aN18oVo1vpSpveBD48sVyxa4ENr4gCUKNXDZ3OZ
jyskMEzyAc4XUnxaLokhrVWxyhIUj4FWAFVQyTSZ1huh9jcbN7nIjGS3iK4fFIDT
sPjaAW8PZYCA+Qjzcbo/Ftx2mRj2CTCroonVpxRw17kkjXw0J/3SYtrS3P/4hRsr
UeWqr8CEYRQZFeoIYDQeMv45cagW7ZlvwPlIado3d+r4foS3P7odNFtHz+wuIf2L
yhhwxsN8E0xdCmBKH/4dzvCBEAquFcf/8OPCRpanjfoN714u6LLXsUAN9JdQcomL
htw/Uaxu6F3HCVEuoqcPfD6HyhurAupbWd/Puu5eBWrTW/AZP0Uf6gMsBNQVN/wn
ndmC82mzbV/8vTJXX1PkO8Aumg0zuVczIcO150fQu6lullLt4SsunIi09AvjZ1+z
3J7MlvVdKjMzAns6KG4cVkRwaMElY8JdDNqv33bvMOlrfbAHxpcK2aWsE8iYArI2
tgm3mFePvXJrLENibs1D3HTWvhhChbiXTysXRyO8OAq+0CdmJ2kFaz3+a044nQZM
S5z2NlRmw/sGVLnpjZD0/1usioRAXNoOQlhYLDS/NQPoEM5zmF+ryNKGLMzgU0T1
qeWvzm2Jp95NzkyeO2W/0URolYM/IIrG38LOzqxqgFzKl89rO32MKc9X5Cnxhn7z
yMthJX0rQG/qdDwjqhR247cdsS80FgQy2J58CAms9my/lKhLq4SKZUv08VN1Rl2p
wwi40MT2Egg5FIvCuVeOD6UR7m2ttDU8kyjNH8FoUtuUPe+z+RT6bQzmLqFdptop
2lvtNDLrmqbEGBnJD07+lHPLMbcKDL0B6sq3d9Y/V0Wr4O3xfWIQ9NCIs+w8D0qp
l+w4u1OXY4++gT+JkR+e0Y+H/mVvpufOv6bANEWAp4L47MW4qHFO1PZcmMawbdKq
qOmZR2gzpzW9z/AKMYGP15UeXuBPA9eWGQlY1ZhLiHzdBTOpbeWx8sEUfLvurP4X
y806zpcnUXri2PONEscW4saX2yMQkVvBbb1luG1xtGCJj5jvcQteY8hFSDr+qvme
2fewun6F2ui7DOjTQWtCQ/99gFYWg+ehjERkzmuMwtg2Y+u7pgdl8wOIMazD0YBQ
Axcmv14KWD5hzo4LEkHs5prWiOzECD9kJp/H93DqBlc7bNx5THIfWItfNFxo2kYg
M0J9q2Cp4bxngOsfdYVZ4NMNZql4U/Zrsx+Ad0NQ+Uo+9BZqxDau1suNtvyzVOaP
wcMtn0vvxZbu9QO67qSzECYxeqd3ulP6heJjRoeWob6Bb1Du6ENTD1Nufsq3MxSs
g4R/Q759Jr0W9dGKVxuy2GkCoutwBog3U4PC72MJkoAOOmIy1dvjaD4ySpg+iYYi
6vvNyvW1I5kLlig+x/z/ky+9sSuOmAonEPFXWAnxFp/UQq5ljdU7WAW4Qs9WQM23
et7MXd7POtND6LGsUh35s7o66yLzBI8zsdKYG8BauLh83sfY8voJ7ijmbilBHYch
3JToVhJhbl5XHJRT6T4oizBQK9H5QGqTCzgnEjNj9MWzoS3Oz/J4Xd+sFMNI1XDk
dqOg6pmH2NxPP20LdpPqJqrfH3HVOK8Mg2Gz8WOktUmX4TYu33wfNIogEco7ZXta
P7jppN/B46ImEYUxxk8HDcNjVsnu99f9kXQFk1UamIiALo/MCBhMjR5Hbt2e3YBO
hzeQPaN2epayndJpMV6fOSu5v5AzZXOZwUONCJj2X//QxPBzoYuPTb7+IxRUfqs2
Bv205fe5ZMApJlRB9cxUWmXWF9miMNAfM1B+JbifmcPc4Ffnk8ivAfNdyOAHNUqh
3MvLaFvDuatzK5qFicSuhpK97kTCZp3n05Z3d3mxTZUKXUu5v4YotqJRg22mydkB
I0TWCb5SfKb4dLIZZD1O64WUvfHvxRyTYfpvsjnET/P1PtyOwO0sI/o8THyWZ4BS
5eAXYBQmDQto+8u6BKlgibyfStclTUxniqTsGzzS0iLpUFTmebvefaNgXg2kjBJZ
VTYWwxIHX47S6SbQ0oL/7iyIbIUrIdZlWZmBEXDikU3avAncfQTPMx7sScEe2196
8ZvInH8a2IYuq5irAaVysQqUIyUEEx3zq6kCkefMPbFFeVRPntw8XNUbcERnOOM9
XIDqtgMfHnXlxO9pNMFzhHJeDUxULqhvOnLw3OQR75kOX16e4mPyxIqWGBSPWqLK
lfDm2rqc5ZlOzLzcJTNkpRiLFEBouwnwOiisOBmigM33DiM5oL5XNDQK+W6mxU+9
/YYBPJqG1wEgX13GqF22mJwxQ6k/6qYGb9EvvuhiMDhGr3rvotzd7wP+BLc+sxo/
NF8S1MLsbEPlZlUWNACByBiOaxKCWh7/279TeL88bgSiJ8WKxC8PO90Dqm9e2fr6
VwzcIFCYkqFY2v9Lk8AR3vVzOE5j11PVpK4CUYNhJZc+gkb9eH3E0mWjoXlwzCJC
2L9HSJk2l2dNIi4E0DzjEVrlsLEZd8uj4WACWMp9FXMXrXgmRLbB6jrZAKrZIq3d
ydEWu5/4+SzAtB/QgiA4Na69NzHEOFNSLDgWi5YQBy/77k/YCyUpHrwAlqCYv32/
VLGG03MTTKdBrEjqknnZrANj4kRqteJwhbX7xlaFIVp6ReEJ/OCvxbAvm6FrAJmG
sbaengiJXyK1aR0CHdtk8qmKv5GKz0mTEKqFkPi/vXq8Blx/OrXwP5CQBdq/zF5T
gBqFlzUGcisbAKuq/D+9OiVZUWkD8qlaUIJjeVu4tc2YFg252PLTpnS692bgUfSE
F4S12Gh84QT34A7WjjOKB0LwaiwEJDYx+4Dvg+6VuEeRzmJ4ZO7KdvF9f/GlUBaz
HICOeqM3jo7fG4fjAJHnxUpJIxA0wri9x5jnAa+/vUtSrOa84PS+LSSOlESzZhBy
1muPXORAnA4kFUJo6v4sCEpooKA7rh1OnE2EGyKTVg1qhCtus95Cnyn27fb/maR1
Ch/hIT77GhSjmBd3//miPurzXbssr11fXB6cRBxAHJGjNhp1RPXRhlnY2GVihw92
0Jla5MPazNdRsDrapvyMhjZInIcfa6IsNRM3we7J10LNhZxC9C9lhg7XgySQoZZn
ZsXFW+XVHIyPH3LOBgnqgi0pXcFiCNw87UABmJcCbEGZS4S2PT4YCAx3iwtgk5Ch
CCskWrq4FR7Ep7J61X+ARjLqVueOXbHc6DyeopDUjxPY3wa1TI5O0bn0SLnqHPqm
xP1jrA8wpp816g69sxq73h7mViE2iqBtcxWAFztBrfRuA40G6C3ki/swyv/tTWg5
WyrJVm5djYKN+nWLT4taRTo7QNRs4aL+fZCB+y2ZI8FQQMRX86JcjaQOa1Myzq5h
TtP1gUV4F4hIGShu+UGtYqEEP/MJhai3wMDFDZTJ3t7xd7u/n8XJcHL0QCJzmIWU
9iqoZsRUyCrUfC5ox0hJOn3sCBTuDYlbdFg+PTsUV0BmIeD7OpJFqBYFuDapvQe5
df26LSTK3/EjbrQuR2i6AGa7pfpzsumWQSlIIn1zWSmMnRm6qS1At1BA7riRbM7f
ms3NjM8Cu+ahQRC+NE0DUqEQ90t/uBCF7EB5dzJU/nWtbf/36SOJXVWvlLkp29Fe
32yEj58fREiMWedb0XxNmT0ErFfzS473tBohEA6LiTH20lI4Z0yxvFM6Uh4LxRmL
z5r2mabKo2cpkhIC+dGT6SDe9yCU0gJfmjbvECW8nifi8s7ckJk2WsTdDY/xdkPa
0+OtqHwbeZflpngty4amXA6B28HuqEvZ6+1FDdz0AgIrc92t3o1l9j6XR7p76gYn
TgOnpGxydbD4WD7dBiR9ar+qg4hk4ROrXl3IduI9BRNHduhf0BD/USynycP3LWUf
ttHUskxqh8yFLzmcTkLqy0Vvu8w6R8NyPZ7k807EduYgRtqQDnzysy5KyhPSI05m
znxLBr7XyqWYa1As2TvTYDQCqlLnMJlIEI0XCdQ6o3qc+1nyG0aWPfYPDGu6sVV3
V4RA/IdY9qDQtcZFJeaHoDUjzJZFJf+sm/rHgb0k0U6M3+4QLajAhqMJtN7nw10K
Cj8P8L3pfs7/BptFbewKdPkNiXkBQknHVsbONB85qJmPAeFAVqBdfrL9J4bDf01v
ipFnWzjOdPBSpy2kVwyE7ebZuwxCl2JwivKElamcNGcqrKJQBjfWgRwpZxgVUxXB
VlNCAJZKKS+/yCT+enwmmpykQaZV4SM14TNyuU/vHJbKF5NA/iuZ4GXaW6Bp9y9X
+1Ggqibj9Ngeph8D8j+Lq0DleOHywLHAWjVdlrywH9OeWJpcF+9jM5wSZ7RWZT0C
u3b5SA1iXym7ygYhicoQgbmiFBIasvAdtcP0IKF8m++u+tzuZMl5fRBX4GlmL8Bc
hyA5Ne2KkLG6Zf+hTd9wOE2waD/JyfHKJAg82X+2KYE9cJrpZkvaJvIDgOSl0FeK
zsshduSS1FQUW2YqA3zChJgMJEmLSCDSpnv/egnkxa6S7qT8DJppiUOfCOsQ8EOO
OAMpKmylFAFgTawhWXgmLiUHuc9RYfnIrR8KpKcmfO6thUivMWKMIa5TEWyMwYu8
gHSAB1F+KUoJ7iKg3Uc7RvAOsJYb49IGEXK7SmCsWWe9Yu62lDm4QUIBxLlw2cL3
OxciYIpQQDzmk4qKGtdbyr9b3YemNp+Cc/mG1m+kAZxeVIeN8TR+Mk3OKWsxlxPr
u6U0GsWTJv4RHbcTUplb7saTSvm8A6z7gptIzTb5YyYFEm0o9IT7iEHAulPwXFjC
5qgitIVMWQWlVJW0j1kmEe4ZzLvMCYK8dVaQXCgv8+0FnaSrogAi8CFZOBsP8/Lk
j0hwS38nZiBRcNPJY6W4MBANywRsIVwumyDxmeVZ9WtDqqNFPOcSSbloQcYs3ykc
z9Z9LwdlhywRniLLqDI8WGwPNHYK9RhSpfXWVDYtZu6Gs2RwvZNzgRlHnDANEXD6
NhUzvAlfuOfCAl/jrATg6ZI0wUuIpyjKn/6j2ljrZMEryzvDiWE5GgBL0RM0W4EE
OA42dGsc64W94A/7aCzElkeoyoUI4GXDy2Ol430uBl440VgLl5gg8zdf6X3qnFqT
BjlqY63dkuf5Cktq3WtKYz5XD3JfzaiNn6cu0tLqwG2imMu/fLHlxJBajP48tj1U
wINx1caIxTj+Yu8YoqYt7JxnD0xNt9UfCTQHagvJ9Nsun2xyt3WCY1jkfP+1Cw1H
pUMj7q2G8Y34RFRCDJ5aPV5P3Pc7+QCnIGrSwhr06AicUSzfESBbDWoOcTMOm32d
1dNeZ/hBhPDW4W3zYeBpYvEsA2tgBDX0DUpPxVFM1ODfXnllVHobvU/oA20Ph9Q2
ks7PaYpB5zJ7+sPjF1BoHquCcZw+zMjGFYODzXt5dfcKDtJA2gNAHzxknOc+VDKh
8egFW+AXJSksN+khnwW3SS4Y6nQXmwn13vKK5g3lmcbOnxYgGrSOAyk2Ns5sJ26O
xg6sARXhwHOQrySr549d3yBxAnV0yjHD0aDEAnpGtlsgehVYQpY0BUC/d/Jk6mbP
4YSXbN5XTU6rq9q4lc/X7F3DJrxSmcgDQQoMZB9IJWGNe+Kxvn2lJr86bJzMCGT6
V1FPrhcxPcIp7ohik6HwG8FPernGGp8BjJ71W4eFzxWy/SpT+NcE+pxPCVcsBeS3
HKWh4GnZmIU7+OPEqaCuosHKYpO5R/qQYnFRUJoteI0N3vv9kmlbmUvgNT32xhAM
MYQsZfiVTserqnkYRfDJvZVrXJC/LQlY5IiuT9tCiMnwOnX0prV5nwi1Hhb40p6q
m7q3ZCtxFd+rCcyFb8+Ynls2F7azSz7IYvE+CSuAOj1k6OGAovHtLOn6L/V/XiZH
un+o88kvhq/ufJVuH78GMFp+AK/hQgOLL9yKBUGwx9oOaQcJfuTdhAnyDZbElPFV
La+Cb5FvKSigoKkpYP4P/861NKWuCyAAiATFphVKOGzfmcp/KSzQYn7URyQVUfqj
euwV2wHBvCHqSL002iX9IJp3Gk1lXJnLP1rIqvfuKa9Th7uie0H2b/fpGRXDZ/+P
s0SiheYT3WH8C4S/Ln/ov0cWALHAO8E3+f8+mUcMg3Wy3/Fq1inXF6Kxtwr2mOp9
QfJFlp/ARbwL0zol7XSVZNJ4KqHFf4ZkFjxruazJuYzLeL2RCITjkqUtOl5XHvJ0
YllCx+bJXhcA9R6fU+NgteslFT+XGJ102Pzn8Q/3n0pmNdENSK+gltQAK9LXbi4y
I8YbP4Ce0Ahty5iP1IaVoCvjHKdtDe4mCyjg3/apJeTc09JjtTSof1vEASaUNGRZ
vMcXaDS5Y7u1e+MbYKNyjLDjms3HSRLubCRENeqpLc6lGDi1DoycCA6Lr0KDNLE5
5R4MxZ6i88P8c8vxDxZmFRlR5b6oHLlRVK40MizRYo4tIdEM3BPLvQgd49THmlas
yXFfz05kDl7TFsZuPrEcnGanSMtWoUeZD2gKdVYlTQH1tjaNoD4fTCmViemwDOPd
tf6U6omRnvVpAdgE+cEqnmvs9CzFz/uw/GRK5Kx4L3YuRdpSnCF6WKMRJgccJozQ
IaAjTJ0PTbEh7NXTEyk5P2rIGQkmq7wSRLhE1ZwbP88wOANYYqztVpjczCySGlS/
frQICvYiOCnspTPnCgSoxxGO8Qg29ECZGVTb+EB4RoFRTcTkBBv1ddK9ICbdiW69
c2uTRNP7fR6Id6BEE152XDRrymQw6P/tHL+zRoqqUgGzej+aBth6/UEaYNvEHPcV
IIwCVX3sP1NXPggbmKVBeg5cc2kWyQoq99m6zkmCQP5XLIn1iBB3FWZ/ZNK2T1Wz
H0iSqq5spwP4UgKzQb69Ppr34LcshuAmLON49kSZNM2qiWny5+a3vutvwzFap/ND
9CwDQADYa0jMQtuNEmLOL7sJUW5mBbsK6FsZZHM33UI3g/q1K7kGBxtbhGUqoFGc
DHO6QMl5vNjKC59eT4GK0IiHAhnbkBkhPTThXT5fKYUb813FcWWvGqrpbS+e8avY
ejojAncEaMhFtgsf0vS5F7pSLHG45VXGHuJLBG85rxxEcFiAbW/fIIY1HpJlX75+
MSkVeC/tURr6eBgzAQ2zVzVPiTA0yVYeOcWb6uGfjKSOqjE/nPpFiBR7td15lcL2
Q07nZ00W0K/1QAVxfrlab/J1mi1HTw84CkYR04i2fpMf6kef+CCGF4SwBN3kDI+H
HkUj0oxDNIwwfFlHmr4YLEvf70SMv+s0ApV+se0yjtcJa1kwrJcQWv8joXf1JOfb
2pnYHBLfd471vtYEL1n00iBURyf6fMr9/PNDVrMC/Zmsk2mwhHRjvM/mHhDf77Ik
nbynbF/ggNuZMCpU2L+WCRAccnOqruc5cEetdz01V87u7prxHyKS6GwJswCSE0Ir
g5scwanS/YcS+WFPQXGt64s9q+QnVvG8Y/vSkx8/QsBFuRNSnPYM0NCBE1Luyg7N
qlSNOdtG61JzlseMS4V9vsPnp6fINMffCEhlp7bU7K1ZLJ53w3Lg7yviTQn1rksw
gHIq1MG0RRt2UzBr7E96t9TsI6Dh6HpZO7LNpjIAuolr7GMTawhf4zco860alXlY
sgBGeDBW+2DjKcFoBGKRSBOGkyIwhk5tFxSeMxCTWdSzAZVVRkScdGMIH2R/8Y7e
iRhwfDkRInKvXz9mqDlBg1QSeDTxvnXgo0VYNOWY3sRrVEBow1U3Ra8eYinL1ky4
okdaIRj2cVjBcgPgSfa1HLzIa5fzJRaq4v1lifs0Y8Vwof2ycKR0EMYS8oZqc7rV
NJUDRdBUiRmYgGDRR8nrS0/ESUXlPQ/TyjHT0n0WoEG/BcryZl2DB58RT2Vc3FRr
n5vZtVudDQDV8DIepUkSrsZHKDGHqLcSlWd9YL7/CaKeL8lyxWJSFkeAVTdhbjGw
gjYZstBUZ+0IUOa+xJoblCTlv4uqqJkF9B9MxWYK7BwklG9P+JurVGu2y2CyobkL
Ejfp+6akWm49ymv2O1Wq8H2FOVbsaqKBoFh4ATiGFNZEtHOz+qGzbT2E/I0k/glT
dtprgSkWrftaFLW2anRhNRc/Szz/3PbCF2SpcVYA6bJp3JCUOd1bUFy7xoEdFxyx
aG5dBihNOzouNMHn7HG7UTfQI2mcB8FbYJ8JX0Jr70hGqPj6c9D5gHzBzbJo5fuy
iH6wc4gKeCsEx27LSmAXSdBuBVGXNPSDD/4GV++b9n1YY3R8V2phlR8dvNrWiUC2
edE0AWn2TBO0Se+Fcs8Te5iwprsFb6DtkOGY88M6ecNM3fldVfVtVdv54j5KnK2I
WiqEGeUb4rLtiI1H6v90mfbqbbegxXNmymcKOp9YyjmQUGvvRB9FxshJDgb1ceK3
sFuVgzage9dHQRR9/y4VpZZ+dCEkJINgFV6TPNS1tqhkK2drY4TFYa1pF1tOtDJF
BMVqP+mBb60LkY8hGoFvWpMaonOAsGNYc1/xmV2YsWUJgNQfx6L02Q1wnEFsi82T
lc40v3TsGXf4Vc7W697RrNkwqtfWJBbB+Fh/8qgl1yWtcpnt11wcA+URfBsWfG/5
mAuq6YbQl9HMJfgAf0zhsSjzTY0OgsZ8rVeecspHLbMYgaigIRJZ2uRaNNNQQNs1
d/5KFmvMTbMhqmRp2uCR+qUDDpkik1KS2bLg4BVIQtQWizJ98asbKGxulOWc/4ZQ
+G0JjfBzZuBdZyeK4mDNbvypV5LdBT+pX3Q98Bk6mlXlL2BFjO2onh6ve4p8rMPv
wNxLEo+tVoCJbM7Bm0vrksFHCo7rGnZcxOVDDqe+0QBdeG6AYZjdyIASQjaTkf/G
PdU7r7DdZ1QYYAi5Wi8nPgFn0aIno2hIZWJo1mzSYtLShXeX+JwsDiRjt5DDtpkm
kzMe13nAOcYixfLCy24dpmJyP9XdQkf0BjW0W5wG9CEA/kcIbEfOxUDht7bMnJEU
cpIL94jYVzcHW0ybjkEwWSkCRbi8k+613x8hn0rgydEVLPtGzbdjOEyI9djxuK1G
LtChr1DoxwZ1rHWaJG4s0cVLXO2pV5h7AuFzd+2qd6kqprIxUc412VrIfrDmtB9s
NWDihxlfAkaG2kSdsiuvW9ZlHCytnQNDS3e1qBRP0Hd7hC6nRrv1ethtIelWAzYe
OInwwblw/GYBkLqjqDMWHWl5hM5H7Jrlyh6n0RWLTPJMi07DpIVJc7kfyoDqjYXj
ibWII+ldjbaDZtR6z67oSq1vW9jsF+yAqWp6hHrlF5eqsfCinJ8RqHkY2VpgG4jC
0azJ7id9/8HEi4wpacVAiVISKEm1HhMfzx6XWeP6/151FbrUqvazqe+m6ksNiPra
znzrOavFG+beYQm+Ne3E1z1iZGuZfCxgYhB+fEEiOBIHjHpxs478/blzQA3coXA4
tOL45KLui565uogzP5zJf/OfG+xtBki+gL7iUrnYYLDe2i5V306eYOSq8ZRs26tN
pKnV1gpG02G/sUPeVcwjl+zidhzMz5VJ2hdoQ8Norze3s0S1MdyYAIyeKXWYr0RD
vDh0MvqG7Mpu+EMfEsEn1Ur3KKlnF1vWKo4rBd0d8fJTx3XqxrYQNBY47TD4YAhb
SheAi9xDfsLScXf4KPAuzAEeU+XA4lZ6w6dzXD4M+F8HFTuZo2Dw96snYok1k+w1
i5SGsO1g5rIdn/nSLjKtOX7qsbZI8DavcJ0OnawCSXKR4yhiWfGiLyx6Orkd/LGX
AZ/hhlKIe2mRafR7sqJj/uEINjlr1Mjrf6AjW8NIWUtTBxxqzRJOzqZ7N0+EKw6v
pvXs6jTrMPYIvZmxXjjakvMFERxcMTfs6DMQpWy3Dbc40iwIKueIJEXzEGn8wFFh
oNhP4MQeatl2lOufjKijaAb8R6Cr2VDNZJmG4N1koPX373NVxw5qQuKVRMHJxNzg
eHsWlKxfoh69S1Pdv4DdH3l80f+h/tkN5Yhf1fyK7T+PKvFLlNaBFgQrhnLsR24M
ZAGGvcAW93WwJM24iueBD2VOBgzVfp+m6hb7b7CQ+SmQfJCDMcFHHHA2xFW47SmB
jsZcsUg1j9W710OY80GrdPgqrfnRE8rQkr7c5FI7+6Q/22mEF+5VZC02cKFaB1ev
lW7ghx3DYSXRevOFK+L9FeavH+k/BHnJY1GDXgSLg68rFOnrhWDAOXYG/PsxvpjM
uocAwQ+WeyE/H5FK98Z6EJwvhFjUaNy3yKTOxwH1tydWIlZDT/ucc8iRfafdgHZ5
l929cK6T5BcACI77xAn76jBSQoVeQeYGT6SXSSFI2Y6kS7KA9AN60gTYR1yJfaST
tE0ZlbVzXDLESE33xxZZjR/b1JwppPty3sYqZqGRRlxUJmswaf842Vb1ab2Cl4/f
4f2lMGHNjgqIN7VyG2J9Mz3PbAQ9Z3LiPzVwLu0LIbkzEaq5lxOY/HrtGr+HzziG
oSmI13XuE9JG335w2vuGr6TGFflV7uz/BbePvFCclvT9apVB6QpecHGEbhZqIXgR
TrkzeAsSYWzrgqXWf764oMnMr2gNuUc02pOZsiU+7LaXFfCgvej8bXPXrtCzao/K
RaKTzQeB3is+QV8xuzgo55kRLStIiBoSQGbqiglRYaTxmB6nJOPuVwR2RXyRIf1X
qnrlg4IeHvOaunBHppjKSuqgnJveAQnuBkxWwG8sBNZVOe/vuuw8SybnF2BijD3E
dufsQacZzsES2YWn7AGCfHyQKOnyCe+GFTAd8AmZf3B8v2hfrPB+cH8R6VWRv5TQ
9e5Hd6i0AnRb+L6W9foUNCnfwAGSOSgGhdf+aUvm6H+On07puAl3aG8q87rP2TXO
Ei/asEWybIb/9f76GEauXsrE8xYBfEjzHExmeXqttSDSIlXjpXVNpppuios3fJnB
YAmgOr0ROmZa/aAnRrzmSi7e2FXViZ+BaG9V1DWNOuRwVDMgY/L7BIiIOp3m3kGm
CUSS14RzDtyADFne084S0cN6gl2hOfdzixi4S3lO0/1HBKkcV+DNd24dvHgoCir5
Dy0j8sWPotB8baA3YVvQZ3kh0iUnya5+FvXSt5DifSf1f/NwG0pAjc7jNlOLw+wL
+y8pFgqJx9HfrgeKXCnclZ9lEbOzmpo7NyREDngWlzdLnfwVqBiKa4c/vcJq2zLy
XWQiuZu9w9XQ4mZH9eAov0wF2jnZg27sMdv6hKmqiAkvffIZtytYbjO45zwJKpth
5oXDsyliI5OvicrP7xQUPpJ8T0W9ddy5yFoA4wwPHJs67zDohYQKL/Yy9y9+Pyxy
9R5apguTHI3J0AIcspTubTEZ4kfRUGfMx7iHBQZWcQLATMJeEEAqIA8tvzEdUf8M
GnySjfcBsXpsqYU7JF20OGb+uA2uy/zcNMZ0O/ndIHorK1qQrWFqkSoFOlJ//LkI
zbNv74i9/JKhsr/SoAwyCo/2/XEU+zH87cXXyvimXt8IEnIEIoU4DM/d4Y02SKXh
kHdy3g58TxaqqIpJmdIUn2dazMy9t30of/bK2VNxkEqXT3k76wa9xtvsAYmEJ9L9
xanYPWRlGTcr8pwuRFjwr0ViUCf1LNHpWrVGyOEE1T5ToeCbXgB69WXRV66BrVHK
OHUgEsItf/UqBDn2ilOar9Dv6Fe4uDB4rZ91trwKqEjl6bcIVzD8zqWT8kuF1Tze
7ekQCSfJ05N4juL0tKrfY1D7jLmU4xMgPVnn0gb/9NmArbyX0Wg569Bmm0hqgyuH
uR7O4oPXJQye0Yx1cQEHLTZsacorB9YtfWl7brfunJAylW3MpFI4Q7Dq3PYLv84C
zDWEjVS67BWqqE4CixI4sfgMvQNdYTuB2nnrhb/hLNMVevFjXmUwW7vqKaZqUYYe
PWb58XfkiptlGD9XAEHR2KIDWHGUyrEiJvudFRDN36/BeO2OQd6PgLGu4Hti1LBH
BGQMfFRIaMmnWUXsdIyjGO7L/y6gX/nK/uzy/KGw15MB51ESC5Fjt3JejOq7dnJu
PSMDxFeNsP4OTDeEc+s8gZA05pYtXAlRF0v+VR9ud+QD7KfaNHKSRsyn2U/VVeDi
wNcipWCufpLYCyZPvHMX6l9zX4pqjIG9Z0+WBW7xRDKfHGEvB6KiooxO9kIXzbzq
/c6oiooWT2AmG0ahyMzKrn2U2JFpTfRPHy+yJK9GxUm3zpIF2haavUM2d4CAG0o9
y8WEmDh/0vFdxHP1wriXa+hXmOMKXhyI7ytKlHclgGuz2U4VAW0mQZVYUwDm6ISc
M2BLIOq3i62V7AxvHez/cAV1Ff5JyaMR/goSq/V88tCtyOTzSxM3RM1laNOB4uah
p9Iop++gJtK7zVZhnKo6VPy9weZ9IYaBLB66V/xAVru1PD//egSpAaT56lLZO+ez
YsuuroNAh9K5z52cIOwW+KcOJtqfz/g9LKKXFM24EMlX35ZuVZpCUxpbXWm+zUA4
F2OLBnB9DuaV+hY+Orf/OkQW+RIbnLal4sg6BeNloSjsM+Mh8eVYoqYbjhGK0Fzv
h81g53Pjo0FfDvWKPt4uGJZlLBfi9/aYG6AVuCH65ylmtMnrfw8gGJ96zoBu3rjX
pI9XytRkRhAxescmUodEVgcYjp9HiXTglIubXZRZYLV/J0ZpWoFzD1QLIRyt8DuF
LegIVRoG5ThPR9SJYiGkYdPVb6zOlZE8kwd72ec5utGQSkf27cTBDfTy/Iiwq7Ns
dPwTiqyK309WiIL3euLB6NUUe61VQ+eNxn1hxFP3QwxIYopqvSo2nliGCxvbVFyX
1sGowd3AJz+2g6qNIGKKWbsYtBOVH6enrvlM2kSHwKijCFbL0VJncih0gnGkWnGU
8CQuWb1kW1nPiXB1dST11sTk/N6OLmtTTldr112j7P8S86BIk/lXcaIiNkyfzuDG
VR0/dfnVIybQwJdaqcCRxny/c0jsdH5pHKTEhz09wNqzSj3r9ytyCttsXrQEQNJi
5aA15FFrW3S1Ph5iBcK0QGbS4Leo2aVHMDMdhRAJXAncQvdF37KJNzd3caGfOpo+
zdmU3d4eBYEjJhSmnwjdPcIzlHZZxj0eWBpcjEWHhugtuOpf54KpBxxk+0eByoWq
jCvO3JxxTW15p8FjUcrofek6SPoUVOINyEKFnGXPQlcItVmwnyn+avh5/5ooWqNE
ppXlaluf2Im3s6oy2fp0y1BCpWfZzjeE3OgS4fPqRvwQHp0vnTfUdUkog8HoI7h7
VyfflcwInNjMnqhPJA4e1tm9wWaKYvnK3occerN8lv4qBwJNLMhX8pGrxQ3D5dsc
TyS8E7x04lgayriiXCs5Hv7AIFrBG1KtLi0wyvt2R1Of77OeDxRI8qGLaE546aWZ
xjxN4pv3MwptpxkNfv3M/7zMBx0gevYwRD/Ry777T+U6+oiDs9Q+xQG/19gKkUV2
Z4lnILHHXwUlj8xGzenNy6Rq+mFGZfuvuKIlfBW045JG3HEQ0TKBgbHeCXB7rrsB
rDVwKrY6XAjBZ6eyYqfIvmupBllD61tiiks7f7XYguFR/nNh2nSj+RNd0F9tJ/W0
/DJZ6N0tajTDYynfDnVQ7dj7RMuE053rLAgQ/CtmUg4TnW2P8cLKPo5kIqActZ1B
EknHVMK7T4ZMnwPb2jDGFHn1evKAC7otpAqv4Ntqa2jW2Bm6TlIbxY1A7wTjgPkl
REqMWajproeoQv/XRaJde1KyZDOhDH0T9pNxQeTvxBCh5fLCa+cXgYegpx0TAuPN
wCMZw3ceyQ4ScTAfpGmxP99ghCq4hzP3NMFfHN5p2sMXM+6W+x6l1S0y4SUtjofg
12JqESiVXwTiHH56uOu6uaz7IWwHorvfujceaTGzsZpFJSgVJ/FSsqRakBuKNSOr
+f5aOY33PoLDw+1HsZXKUE0TCrOZfZodu20gy9O+Cf+m+X2uOWRj6dViP8GneOfs
aUt92botJNEMABjYTz/X2g+0mLcJapYHgG4kNixSpqHh1SCv0Pl1/+hVo+VxnYhk
zYpoPkqn2gt0t22Q8+g7JY1lonFdGy7BKaf5KIpG2zpg2TGGTXO/yqi48LCpKmEb
p8NuPXKExdccIhH6J/G8RW87vOQ8GrwiYvkohjqB8h3Bm+jnNAF7dbxLdgpQOYht
GugghxBl6jGAoksTtnEjgx+WddB5NImHHCCGzB4icTD0fZONhcKQbWzL5PlT3p2/
IivVpDKYY/ifceberWwASi/tFOhTK+lAM6M43rx/doiycmyyx6Qy6z6SDvhJPx8e
wuHYb9MqJ+QaDuCLwtPQm1Wz+ypa4VsdUguZMYiacQr6aXtY8EzKPsIn+ZrTd139
3JFtwSdHQAwDm5Mvj05rqm4wpVkVuzlGUp1kTxddDNxiC2zu9obysrI2thX4DvVk
jGRJWffY8mDal0COiJ+iiNzcexNASNbrv4Z8uCYDEA1l5OHzIAdICi8e+QOjDMc1
obAvwfSTklodexzEI3LeFzRtUR/ruhJt+gFxmqyZPJCR7/5aTZV0UIB+5nWgeFlk
CWZfZwiN2cu1DVafBB0ioa3WxkXIb2S7Q+lBvuvhoLkxUKmowsQybB0kUqN+D8YN
Hkqbq6o6pixDlXNibVDEGNfTi4tp03S9cgJeY76KUzhZiRVAxeMclhH+7aIXykUE
YC6UuXclbu6kUplbVo0l8WcqJgNKSZ5JN3Z9FOt3TybHqai5F75njPHx4VMNBt5b
c7eGRBWmneJNyJ4bJw1XLCXa8nhNubaZSqaSSE/tiVS/+JA5V5DXsxPJu1ZvcUTR
Rgab2EGqafkFy0QthE/zkIlij1iwoPcrFuHryeeiVH9Z3SecbsPuKPF0aT5DWl9h
gkyZX3g0Ehuqrs5bL0+wvEYhwwPiARdapOLYaXcWRC22NmO3J6/OvTk1JgPJ4CnP
kFizCyPG16q+g0bz7V/aO6wVeY/5Nhc6WkCrF5pkb0oDEXrhI4J8ya/NOCtLX86A
KH+Xbi7Xm5w9vQKt2xpFi34KfrpFHrS8pD/dYstWD/MVFeeWVoGMGuJtiMn4S/tZ
7QgADMJuMFXlWCJgnV1HWjUlM57jlozpUa4Ess7IPhkaQwOoTcMVOwZvXhslQJmK
8yXqRiUEPSbfz9Ns8zhLOWQFJwBLxKT92cO+VWSIUI3rcuaOU53YHo6r5c5vQhjP
7dzBXZNKXkBNxKw3LswdW2cFZ+9K2+J36fnLf7vYeTZnQpo9yCwUHUUUlRk8WFA5
A+ER/kDREBZggm7ALB3P1+kuzuKHQ+RuG0o4W009uSMpY9AUMJT084a/eJdhP6m6
zgwJJcJdfj9goMRjckDI1Shr/0oNQ0EuZtzudVz9GUXbi5LV27FbaMLV+/Jbgy88
wEaV3hVkQquk1F5ZiIU8uuw8+ShZ6R6Mw6ecRARdLOKe4TcvAOalKeAuVJCqwC+9
KZ44rPq/52EgHHBh4G77ZoLCrPmqm4EE4EmaftyWf6kuNhJAzI1o1XSkm7SxrMSM
nnyzIpozOoD/5pob/0w53GFvAhOIGuyLf4ObGardQ0w+8p0Y2jRdkxkjjVa+58dJ
x3sF1tUsly5cZo3IuVEGD1F4ZlqMbNBWKeMExWdgco+hEiFnZCilpCXJmsu4qWNt
scoAitSa6GRVHVJnsjaJjkC111YUjVO2Wfh0dEtlaDwDiMVSgVapIPMb47S01ITm
4OQ/4+mTkfXuKF3JzXfBH0zD2xJgd+Uh2DO+3MCYrZASP/sYljJNtB5twegdSFqz
AdfxnByu74rL/BcHWJpZyynTGIKhLBkcGGKPuABcsoZF7Ps2HayIhtQRTDMAm1pc
Wq1t10XFvJz4+e6XI0zA6bmMY4JWPJkD81rr5aCh0Ifl0aZUry0vr7MMLvoMXR4l
6l3aB2Tix4Ukp5OTf5iCug+hf0o1d9z+YIhKl4rufvRCYw4DRP9FMA4LeaKTI86H
kn3/BD+QLIYUl84z0kGv4OZp55TP/vj6G44kpsodqf3WhqE+l0+kUFS8TrmmZkTt
wAQDhC3Y6V9wPILluXHJBLrr/IgVmkOgueRq71GkV9mndaAsnFg5EDA5WlYguZTx
LlLPKPpPq5HjYkp2QNWHtn3+KTJyv2ZkTy6cLqCm5n38NSls2xjEFEv7vAOqiVUg
NqzYA+PX2keQ0HWChuxTy4rnpyITsQPYv5wDNk4sGeRK4DLeMfHC5O9nzJTxxs2q
G2jET+ahIEjT1tA957LM9vUfGNacERbj1KVZrm+9S9PHvef4IyzrvjMonqfzQwru
UiL0C03jycZIeyTEmDMC8FdiUTgck4ty1l2WKlsVSDTaq6nj5FqS+lFbJRSmYWJJ
6/CRDHfkbMrCSk3VBkKcwDJZEA4YwacI+8NRL6xAVkRLUUa75ERvOLjV6Q9aVfhl
mqWDXpKRcn91UmeWRyTAi96NNiIfJyM2c+5FnIkjexIOtmjFPHdOyVUBz5pJjcMa
Tj71D/hTV2ScNpzBqhDAWNe4jcc5NGlLFyIa/qPi52bDviZC2/27GQ21OxSaJLYO
Q6NNjspywpzCEsrH+IFuKjt6YpvWfk61wrYwp1KdyFvoGvOJpiw6Mg3oA7whS1Ee
uV09sFslFVvIINpbaeU39AnWq4uKhGfiqW+54fk5q0hrtolXGeD8ZiaiWgGCTx9U
NcLZMRK3xR0WXmNtg2UHQgh3ieZZblVRsGpFa1BT7dXfslm+o4VCdQmAEegRL+aP
89rtO4FW2+b+x4SDqKbT/dwCHqeudyuNe4iCT8ay3aRSVPUc1FYFk3c1ubJKSMWp
WcGD90iiC1jBdN/rvlZ8ZmhDJKL3v8+yOPSCYOE02Sf9SyHaxCG4Cyj3TKDegwLC
QB7vXhEUT6wWiYDw0sgfmhC3YhRkDINpvR7gpCvBLkcgS3ooftF3P1nZNYLkLcbv
r6pX6ZIjFWwM2y/jZX2Y5lUUL018vh07rsKr0n56JXclcBAk6d+8nBHIvNYI2nXK
raxCd4VLSrUv3WitRj+jWziwPnMwnLyGpyr/DsIl+LGRJrFYX8Ne4BBHCu2fKfTr
2p8lVcSfG07brs4tghv8i+YJyi5ZpZzVAogLMGzCj+PODeNejWJKYR8plRsbZAa8
3uxGtVcEtg338iFncuyiaINiFkz/GDwZRwiYTAFl2s7Ag6RKFRr1ETGfo9yMXica
zMA++zZgKLxrY9lzXhDw8ysVTPBdOzgR3rsYvAqjuzWirbapVATxmFEle2zaWiY7
QEspe5LYmVTYpV+GtXDIhp+6XAtQv649aReVRRmPi1O0161y6I+MZaWFNz1/LWkt
nKw4vw9983EiZ/n7uBW077T9Ot6/RY+dwVJo/k7t79Ha2LhekPJQhZU6+SaVb3RU
W70rRB6wEFY2bCK/dY379XTyN4yRNe2MME3kiOSYlsOCn8PF9+AbH3o/6BD+mgK6
OnHDlURBeDXhXgjNETAhwRO13ZHTk3sJZybKahuEY/+uCL2FWq8VNGr1C6cxETR4
H/F/5ZSYuRNUJmNLaoX0y/3k5A6NVGunRahuVZpLLq9lr3gzBadSFIE1DeMFo6NX
5C5oJtt7kdexgyvV7etBp2J7pwvYnPERxM/nCEzAz5WmJvNC1zUeb01Jh5y7GJDv
CoLoS5SqFxJB/XBOB/GFQvZ86U5+l3qApqOtKMAGw+MmHJ1Gx/XFo9X2z+lC0TvN
MQArXno4I0PwDTqvOWUecq4FOCkDBLai66x15yNKp0jk2goVYDG1sqcCREz7bm1C
dD5mh6l82fnkHcTC3ygYJAdsxvGXSp1VbUDrD8RSxGUjT7K5dbxwDyUnzHuxyZxO
PMo9c0dM9S0HhBgGE8UJAUqJUJguT1Gup1j/YV7wKxjgOlYDb0IO5klFIghVtWHM
/ZvqiqBmWRFzkOyrQ0ICHEuZ3eBKTQYyflQb7ydp2kvLwbl6QNTdReKo/ThQwybV
K6dQbUwv8AsT7fgGXvP2Y/0sXrIVsThFZ1j7JgqSzpmaMQ31ZkzMlfvfNmLeEYwq
aX2Nhxd0Nyst/+OS1I5yMTDk3f8zwB00eQSkqPOlPy4WehChudjQKnrp0VxvNE64
Bgv9n2xk+dQ8sV70ALrBn7WSwXA/ReDm4q7abio150MJJs+rehyyB+kigYvPp3lg
vWEFo4e4LVmlELo7DkAB98MyIl3y2K22190P/f6/pR7C0OYrmULUZ3amex46Lr6j
tSVKxz9Ln9tgy5car4Ed9rIN+gvfCYIF9XYHxIsc/71CKCY0CetVi+3fId6uux2Q
wtc1/YOw+HVrzB956ox8baHf0sJCk+bUPLxkzVbJfcObELDct5qLcMFhX+7geFo2
ug1MyjXJpgVWwOYb4Qkay7UeV3Xr8fsRjiiCocoWloZoJiTgViDKHNdEReLTPtoC
nQamD+QuPHTkOf08GP8JcLeIVP1Ao8f0Mv2UanutfLu6+drGTwfxMiNcoZ1yvn8m
jkUmb0xGDzEItnULVuTEypHxWEFaQnUOXO7/I7kuPczC5I+fkcUnqX/GF6ghkeNZ
bh048oIzx6XzTpzJ0c6AbeTaJy+SiS+DyzUJfwxgWfYGy/G797LwIk4BlsZ1dO1y
vtSjIWFGODyWSuf9KxccpfYAR70hxzqaOdMgpiokS1VFBgSkS2U/Z8tiitkLiFZn
YBVnO7mWf+0hLTLt5TJubIxCJQfH13ilXlSaeDO/HIBkIUvR445mw3a9E57PxyXN
5hT5Gfe56OV3mCwVy3aDQ6GTTMkSgnWfzK1d8geD0uiSTHV5oOEUhqCpJwlH8Q04
x/A4UPuLhdZttv+M7P7h6NNQv25BFblkOFxozmLu903lBeUNSOmgXrzkSUF6peak
TT5LNBOmwPzgZAbWhNwqJPCIxryX2g2BHSIurdmoXteO1sggNCs851gl7+T8qfz+
iOWHv4bNjNmy+TNyllHAFgpf3apBX/xp9Z/3JIDx6BVlHf/EEqBKTsfykoz9h65a
z5/kQ6HZ20M22+tCyTwKjxzEWeq6CgATsdz/DOFrXtJ6yOWTbAGYMKayxYhtXeMr
XwvrpZX3Py/2DnH+vxbBLhMp7NN7lkJvyzvOvt2NeIAKGUrIJdQRQmUCekzi62N2
02Y0qYPd71b8YFzhozMmIEk+fLGXcEw+El60p3O0wYSycqxcptgfk0yTmVBmuvrN
Mxcc4/jNgsvWmhL4slS63idydDgBAIXpsSyM2qjCvD2bkjx5jwFRVSA0vMAhkWD/
oD4+d+4WMdjqwqjaZdUHo/N5hq0W1vGnkbikBcyYfwzJIh/wpccIlgbNm/9g0sRn
Sc3fWecSaZuDaCasKH0V48FCsGthIG+fcDEvuMQdyTaX1h5GRUnb1Gr8iNzigNzD
VscTc9F4y1QfCnyJxH7Fsjzt56kjMAqtqG+Kk4pMbVQHd5bmMQomNI0Lc/Y06vYA
cnB7eB8W6DBNxu30NMz3r5TNf3V4KThPoyUWELNnbQJlfx/GMhMidDLWs53LX5Mw
BJODm4tguSHSQyF5OyacJNEY2TI06XQ4D5MnvHEhfuiXna9YUs61efuYiQHx0mmJ
mpgS+wY1F4DE7xun1Pv4O9sYVPWj8+cvfBFuIUe1YjV5vUdi7XeTd/BLjUtY3Yb9
WQ2PXy0bLBYXQKm/4Xu1Fo0EguOJQ19SzImXmWVtxEa5ZDjNyIC1iH5DWwldP4VF
fR2qHxfraxcHpuNK3g+JWRyBRrSZvbLC6aEengbaiiZhTUW1sYyXJfRvDt8sv0Hl
MbRlSJHxSpQxmVhxFmSkyi0vaAT5imirvqsa6UG5r3TC7J5xzsVQzVZloGUh5cNb
tGk4MzU9YReTwUGZvSc/kAU/48Dwn9V8x8W8JJUnZUIMNwvUO+AuzL9uv6nLShy9
wcNraqB+TptSkJKhIUIH8I9/pv5//DbQRH55lWsFoj1p5WffsaRwfw4e3p+czdET
ealUUnJIjA9IN/A0kLcsRwe0CTQyi6vMhqpeVmO17LjukvvoBSW5u247D4DLaWtH
3XCdHBfnUih2XVrqNqwvph/IPF+9ahmewwSthcCKPnBmfLNsVfsYPi20KAnlMPVR
FUuyHm5IBTCTtVxR2kNmROqwGHnybHmrqTcu/DTnKVPIFBsRJBZY4SOWa5dAtaPq
28caItLNE2eeQdpc3ohMe8CT8u5qGgvtAWQwwH29BJAlR6NX6qRs/YXagvBA6QRi
+oRfBR12vsESJ5vsyCXJMARsZeFplHeSh2tSU0GIPtgAg/XRxpWwirLjdO4fkPNw
K/qumjBbJAxXiZykuPO4dFZhBI6CRYMzi56cds8UjR5bru+OqUo4ehiiep5EV7tk
RP7Ex8iA4GdEjVSRkdryggGmbE9FBdZ7JIPJXqMYv5xnM8UVjleU5PziQ5icMUtL
W+C0l9/ZXMGlVR809aF0FlgtMLWd1gxIaseyU6TqiUhd+p3tm9envrB9O/4aUjkv
EsXBbRYkcrAREJ3YKR7B29y2oVnKVgYzJpiHI69+1qNJt+TXV0cDVHqtyji8XpFZ
YxM+PJzIHaGw7qqHRU2bVkpRVBw8GnHcZpx4SzqmDpYxHB70gL1UDNmyQ2NGB9d1
WDFTLwcQXQYHi4f2A7qfbOJAPWgFHeVclO+0+hK5LcfNhuqxzOlKlChJVsO6PzID
l2VNf2L9JNszi8lPxCKCbyD3JhFtsa5G56Xww6yULL1ggDCqXginMGwlKvw87MVR
4/cZOTvba5a9EobvtiA3QwpPUK9ujT8uPgkYPpsCHUzB3D1yVSdmfqfucKXeoIEx
8LRvJUIX8QiDqHApZOHyKVcVO67swDBaXm/iwhplbfAhnjgZE7/+eONGo4/hiQkZ
1QDA2M1+MzrglblmbvkvvfcIBRFlrEReNs/2d8xKMEUhewKNutWEru5c0O3GR06w
cg7TlCgTGprpE9jRFRn2TRf0bZ5vZdHrTlwvgwa3b9VHDTePmC57Y+8LRDIh5v1u
jnwH4fXasIJydScccgGPLHDfFxV3NT4GYcSrbdj25z9qKHjxyqkK/Br5UflRAgy7
MnEYFD+AprVy2tSxs92EKPlC2KRbtyy8jY0Yt1yXHCqhO8GjUSu5mWtJEJ1r8bSh
7dwv/nZHWExgSaWz50pKPnDQnFxVzMWgb3tWmoRJAYZYO+CuhqBvG3ttz0mtdJ4l
IM4F/2W25zoh1N8O8OzQTxWnljpXYYAYRlHoJJMKuAIu0nGHKtrKvD1vIe+WBGA0
9jBrVjU5cE2W8Uikqt3uL/NfXJ7RACWjy37TayMJRf+qywWp/MOWHkqicpG7LjiB
muVEOdJY4hAoXxfLkckGU++myAlRHkcGdpPL9ZF7/nqGI20DfekmyjcOvqQVc9Ai
vaghGXqBjnYZxBsESTr4Us8r6XPWKshfe5TSBC2cEHE3dSb781EK2MmLuZfA2QqG
Pl8jzHkN7WxjvmZtQpkSibBXQLET3p0Or2mnOOmiRzy+QB5+1/7wuI53Il6kPkvj
X84FkID/6MekGZ9Bbep7jG5D0R0m/CK+9v+Q0thLniE/7nkYowDP5xbz4HHZwWCn
2FrwOezWnNHy5At/iZIRo0M5PIIz7FjFGvUaics0lX3UC8xzAi7y9b0Vt8440bdJ
JJzRymX1Uxd3rxMdexUZ7VfwQyvRFpdGe2j0Q2FMF4BnKpv8x9myDRSh/3qCo+1l
hn8WhR8cO+UD0pRuOFgPrzDpTI0jndGLog7KC2d/EaikuHUGqnNpOsRIUfrvR/h8
VXIEqFqb6D6o/NlL1yPRikQwTHFRQdBvjqIb2DUyGBQVIQ6kIrTk3i5MFwjXmUta
6MhIeJ+ifWSlkqQkWhK5htU6mjXeBeApMe7IHYITm16v2xLmor+UwpspSeiMRLz/
h81xeR++u2MWkCnKhIqnf1GJo1h+grmUK5/LwpqI2m1OPlxnpyrY12VnQcO1Z5hk
sBSVKby6UiPZiTpr24K1x5xcEyiDchCr+fyUblzVoVNtxADtiJxRvVz/Fam0AinH
TkB7IpCYv5tMAcXbNfS9dTvNZ1t/5bZXnmpt3/ZRecyPFDvS0jH3dAhFy/eXy0Xh
kWucgiESCvTVO1Bgw4Iz5LHEhBwO6H51WrTYhG1McYqh2P/WeofJHxjx5LK/nhCP
+8VvMoJC8d3bdJWVOSbienuFcJgtrT5KQETOrQd2KLKB+grvnRQe0SXpGDR5XncR
mEBvxwr+r1Cy+iRsDMs8VSSVyZQbRTyGTKpzmVc91wTi8Kh548OLxRzHSHu8AUhv
lvAIgcpDDqFcsaZxPoSIi3oakmT6NTBAa2LjXq969sukJANUmtjUlHz5aN64B2Ww
PvdMnHNV/R/uY+P3CZcHqv6N8fhzIV/R/OGkchyLvzNEC67rg6qpG8TTMaO+X+MX
oT3/0prGAwoXnpCRsIjvD+TBW5Vzw2TtiHYV+ZMNkcCl5fzDtj6cb321E3cHdez/
IK2nw4TEz6sXSU7Dd5jGssWUpLjwlZRc27ZUrAYefw2xVtKEgaemwNt8L0kFQdEo
NwZ9JWVTK9t9ws9O2n+SM2UjfbA7eRCH4AF5BbkByec9avxI0jG8n4CnqpLYeR1d
yetwt66OcMQ4wM2rU61xN3738IsubESCAztRbyMiUOEi7r6Jn6PoFSN/TrrUPvRN
2Iiq/3BHXV0/BZ1/pnB+CXZlvBgYjwFLPNmXstVxLP1tA6LbQHqTH++m5/N0PQc3
txuELx6u4mruqEVGQDpeqIjDvXgRD+X1RJtRk3flHeP5Rt3Jrou6iThWSfMzvFfH
8sOJwHiSrs01jNXJLG9GlYegjjJRhXbCFsWtKOgDYTS2fvHWata6V5ghsrQOP93A
KuXrUZiu2Tq85lGkETADMvwwz/J94Kvysy71H2ZaAyXexijQ+tjT5sVLpi3NN/c+
vtZvf/y/6roasl//ndSHyouo1WifoKxatc9YSztaEXxPIWbyE4BB71z2AsSgf6oH
2SJnahqo4OaSRPZRmV/jcZCDvTifvCNzXYMNVGtzdk/0GPFMXgqcjf9KSlDZt6nV
7K9s6+GhrZpiZkTpluDwQvViZKT2Z0PcMANfALTw8kD32VNkKLs7HtL3I5B+fKIX
V1vOQ2Gu0TwYND0LRdpnNtjOjAsscbWAhjtdbyUPmghMpkspTuUZgrbPyn0anT+z
NGAu5gPDRs3BBbP2mGRsvFmfs7EnEginCni/RWECukv3kO9g8HnUMM41WVVfzzlb
pxl56XmXes2DgtScj55ziMO9DEOBIFo8RAA/06yFAFqYZHS+dClX21J8DpXlcoAk
hDOCUlNaIg4Z1csl31RmtfhcDgMAhmEgZUOvUIpV+/pUc3d8J6H4Mm3VD24+rVCw
g/7hZpatK9UEvQ/CYmlGLcG4F/FJI5AyAqXcJMtexTjOKinDLriqHPDs3B7ViAdq
FY37qRslFoE+IoI8S/f3UPyDjsA+ANezWHpge2Pm+eIfExDW1ZXj0gprtXmu4/ev
GzzAqJIUVD6gbPYu1TmNQVmMn9qltMXR5HbqBIkrP/x1PBC8qsry4HA6ji5KDGTc
BTpegZdHhhzZUmEQbFSdE7M4wOjVqzJaCqsJoXSwjBV6zF8rcgZjQ6xNgIMF0XSY
wW4veCTPOPMzWyog44wLWbocO+P9LK9Iw0N73GiZ5papSWflGNKtr9dYBOLHHu4y
0Gwhz7/td/EZ4UBe2KMuojTQe4CyYk3TWQbaP2yOjH+1cEqWbeNSc4geKj07FmNW
CmPbFCH7uZkUHIrMstFMZg/PZ++34RGw5qqmS6U8uj7NGqRpeynBcHa/OfAZQqWw
lSJrH/BhLQg3W/qK34z0K2+V2XOq8gqLH1bucRVI0SpeUlEJ2p6tCYcqVjNTtPJT
jNeaDYXyTsJMznusXC55u48NXeuLkH6mIWbwyZMHVY4nsPP1OnFnsaM0NtPH7hQm
ZhvtTdsMqXodIIGAPVNmCVccMkX1E/csCwyYfj1GTDiOvK7CezUEGQhWhr5oL/b7
xZu+omaI9qTOwQNV/Pr0tx5LZ2+ffX//e/OM810xc3nHr+W3iIxzyUmLvVbAmpwC
gH5mkoMsX6iau73kQvl0xxHbOqCyKsnllTXPOVkz8ivCAvbMqJeMjRzrj3OhlrWS
DMI33ZuLWN+HXt4aqdN62z041EO6us5toWWsyDIrQh5YuMmlWXnXmK1zcJHaQvIQ
qgGblRAZa3kc8krOivjdsmxD+6FTCtEjCX9GklLgk4cdZu02FeuAdZDTqSRv+6HZ
XXiqNbK4mAv4to902+QE0NDPQ8olFMVAA/e1qf8x3wfP5Ulz/LuMsZol+beiuM1k
KE6cjN0Ps3269XzswciCi7pwA2JdChORUb7Y06sgbSXc/2kP/SDi5+E7kBzRvMob
CSeFRVn7e+5oLKa+Y2BibB+w4/clSr/P6aBZ+QKt4g4LrRb5HJSiMaTOvnBFnzjt
9iAtGr9lq4t/SCmY4EP9Gbl7EJQZmCnbFt+Tamd0s0SoVmi7+JfvdzenBlABC3tz
1BdLxpQbnx5uBTktukjifB9Dlpobk0kf8JbUZs+2gJY+Qq2hj7KRpUatat4+Fx00
SvdUcikeG+THje9s8xzDxI4ijC0qsWtRJq0UHgQT/6J4YYwKPNcse4KqeuA0gzBp
hySYMyHV3VmzI0sPNjbkeonUrd+qMZ7CBMgdMWmM/SKtmC8WjGa8NN5Firk22SVT
WAFrHg1nk0XqoZKwsro+TLeqD4sIwqGkoWeH5KCIvWOujfdJ4I6KafgQFCFqGaYd
jOFNcNiOp02sxSvDK8MAN68searJItByi7oZ7pvfKGc+TARLy9eaTyjU7Bky5g5G
1Nxz8B3HwMUQXtmiwYYAY7P3Y7xjwoJslFaTJGvjQW5qNyrVWiTHOfIsx4DoAMC9
+1NCnlJ6XrtXmc8cocjgzeBhkAv8kfoga+2IDKqM9xRkEV+gId+/Rjh7chqHNbaN
blTrfnsAg6yEcdqoDIhTLepjcPl8i0TIHthVOpEpH1eFiApVmGOzRu4zDlLaX00I
WCXa839S4xP2jlYgiMfGWCw+On3sEcTuTxFHHY8xTLO3BlpaYKiiOyB7RFzoA854
qVFkloDvjGgHWNmKBVJW+r3TPvSdQp+jAJ8gIqcvkOP79S6U5J5cpzQfq5FVQENo
YctEuvHPpRpSCkmBju/OosaG7NQzaK9c/WDneihDfnV/kKnvyQE7yNIXnz7qQPvi
O71B5j5xmpIFJtrDZZeP+I5lUbepxDZ6+VWcDxsQebj9AR8ASYjutngZmBtN/ma1
cLGj+8jmM7MH0COUECsmfzyTwK1ckAmSS0SC9u9K2sX+4JmePT+evGLzhO93xDHd
i8jIld4fiXT2Hlh27mCNviuTtJtF7WhD9H/vzqAV81FRVJCZURrL65IgBD8dFzk6
kJWdeMFUXKDCnzVFuhxhx8IuR2tFuqyjNBNZXXYU/AA9YqvGZtSBS/fthFnB7i3A
ZXWIL34d2My7fzByIqeJS1WjHBhhhoj7BXmJp8vGje1hc7/2Zoj8CS8Vnl4rRu9c
XlL31O/QKAE1ByJuyjYbAO90luC1GCtdwNhfz5FL1AtATMJMOwK/aUhhaamE960H
ku5Wb8vpC4ufYeUJGkF9U0d1NLPuKHDKmGvRP4Tlv5y9uwPNDSrQcs4hso3jesRX
rCco/EvMVdDRXkit63r6LoaNiIJdH6MZZDVwaSI9cQildFq21K9V1nVWbSpys2DL
xugoiEqlk3FEocMA43GR+O4ARN//dV/n2Fzzrp8PQUut9oQRk19DRqUPlHBSm6ZW
hBL972Y91Bs8vv2D+fbz68QFTyGj6t2uukGf8nPzTYSb8ByFtY8qHGurGkQxxtJK
KEmTj96OJcwRSh8llKYHvjueKAPBU48SOC5TlZ/xZfj2kkdyJja0Ff5SvN5X6CJS
YUVLldNd/Bh+yDCdXPdiOpi9b3FnuMSMO47hytNfNr4r5pJjPS1034AqoTLTFNby
G23M5R1PzMCR6W8tWZtAQPF3g7elTTQJCZQUmFN2swFdQwmtpq1kNbg+sAw6SUB6
rvciGXgxafepIN6arndyxI7zc9n6AtZzwZRDmiNgvUV2TDplPrmOGpdKyIqF+OB2
lan6JAtSx2qFdLlY/OpJAjDIM2lC2KPdNCNV2ByVbwXnT9Fkkm+jhNgZaUa4PKCg
sVx2W+fHMGNy01itBq9H4xCCl7WYf7mBbP+iorEvcS6hwFRP1DCCF5xQgVAlQq/X
aCWPfZsj4ysVtQzVS+klO9an9gvXT2j5VmZuYUxpGhM7krDdn04h06W3RNZRdNkq
pMmvXit4YGW5MdAdnZtTSeUcnaYI/eJzG+JmJu4+lYQ8ErhLhY30adLpzEu7A5bh
vA+1qRwjlVxytZThTG7BtbKH1IKNK8g3Z+rc+Kah246dSoU/x/mrjmi2ovuFK7hG
e55FKfa6cvnRI+58Pl/A9wkp9hmY8vOhj0WyixcugBvmKn/172EP672nejnp4yJu
loMKl4lM5gqY4cPpt7sKiGdTZApCuxtceMQZTngJONr+l5N2mQqaX7rZRGzhvVAi
d6LB896qAD+s04bdPSN1D/Jr1ePR3SuN7Tv22FPO9fwDvQ/TokZuj10XMXT70rqT
i0+9izdirUN3OBdjdNetd9acaS3saJGPmOiBbeYt63mw+xK3vyW01HjjbSB0Xcs+
l4+x/ined+dWGRJtgQaQqYOcaf8C92rdACJ1lwcLd/3/cvY3yj0xs2rZeUG/ajga
6h7UyE5QskPH+jc2gyxHjagViLBrAeVAS7TEwG7E94zOw7hvGiTSk9Oc5YgrPgfV
FU4MCIARUEwTVUGfa6m6isiUYBtnvk5tT6o6shy89OXGz0//r2Cs2m66QDbR5IL6
+iFfAbUrER+F6b2W1o+jL7j2fh+9dnJZ2zq0bio9d07Jb/BXrVSBWDKbYsugJmxG
D5k5jZFRVIGZJzmPCc56ZJ/esjLF1ff8/W4O4Los3ZTOgyfFHdOz3w3U775gm3S4
xZIaymwzaiobBPSmtjpi1TQGlJzyIGdoL1+8OGyWBOauJy6nMA0vgMfcqyDF0Vrv
YeN1rhA59wr/owr3BWzbi6bdZGHr/MPvLC81eZiI2f6y/+nc8oH+tXrwvvwsnKNo
h8w8JiVgOaLC3oCoKJ1OD9KpEBhx8pqRdmvaMf+m3P5CDmDZvoqIYrhxlsc6NSAb
AKJ/RVHLgQMp/PqXviZ5qmaiV4CuZ5J5qWzEFO2g7lMq6uBf4I8N+W/z4zc9m5I7
5bJ3fVBTrTLpPwYw70jG9xkjfZH3ZkunIwGWaxnSzVsUjr4icEGWYwaV4y13352X
OdCvpevxKVRF9QdZH6D2u0TmPEurt582SF5PlJq1d15Mt1fgljZnf2l7d0BdLFLY
iTWZd5r7gNEAWevU9mFynbnfmxY3LJOss2og73kAnsJiHOHrADtQHNvUwe6VdLeK
gxWAkoM3NlO6g2pHv2xObtlxNyDu2GAZF2h8tGpU7q/imhkhmHGZOh6Sp1LdleOX
sRG+m9qq24ff4cebQd6OJaTbAK5csWIuLDdCsecbcZOSQSoD6BH1DHKsINh1S6/Z
CDeF9fzyYPaakCgPREZFso+mu8UOjJkOXNP/kIABWFamTyoWVO3WOf4MrtkTY/mt
vEliIOa+dTjr2A0Sfe4RAlf3dnaXW1aq1Wm3dvvWCqmAngfRx7PR3kHRM2wVS5f1
HBwhEmqse4rPzRZqAv4Gcgduuk3+fk3DEVGGViro5MeDQUHKqnrhlToxZjiBlZ/I
oLKgh8BgmnSXSaodCIXEd1bY5dsjixwb5qd0q9i1W3vxqHzk5Axk+ayY8fwMXIBA
thLzL6f2e4G/xtHgTB+N4N7m6/D8mkHPm5p+aYBKKFBx0NxyOfdzX3GdGORVEjvK
F0a0LmsfqKNjHUvI1BuOjywGxcdnhaXFVXXl6JWTZnM7216UUwh5egnAP8qZiQC6
xNnrfev+EJWuWpj2522YkCcbg+u5BChNS2bcCy+1fRaf4ib3ZNds8Y767OPNrtPZ
g+S7+Pbs2KwoaiuBfvcJyg3GLd+L1nTPocS3Cld4F+AY7OfYuoKE4C+KaKrsbFG4
ZRNb2oinnIQgeZiIqqX/Inyj6Wb7bOYOmiHMCkbsy87/wwniwX5izgKbOr/r09z2
uxVzZgiMrr5+mnlf5TKx/vjRnF3K2eA4O4zQLAmeg7xZ6phTWzc3jVZaYr432aU9
zjPGWY+yZkSCp0+elpavw+ZNtUNGAUUnd7MILxribE0Si9bO9Oljwv1Ax2Vrn+8K
XtDJwDW1lW2htBREqd7CJEVo2ZfHX7EyQkNCq+A6G/tI5bb9fjs5FuhxbU5qJkiK
37H4mPgU3hP2Z3fWWuLNJjIpFKvOwveZ9OaeoRa2+Rf7iNLrliBMAntxyHp2j1q0
f8DHbHVh4sFzilX7TxJfYlQ5ZhgUvm7Rnye+14WZwUKaOQMChR9Un3e6fwLm01xH
ODZ3MQ96zNm2jmIJ7Bei0EKLkjpuneVJRVfyoJ696zUpIwSov8TtedARYE/4aLNJ
GpMJCy+val5x8WZ6LkB4QpBbQHicxpzWReFEs9xEgdTxfdA1J/k56VcTRsdmwLsk
a202dCEhH3NGVqt6ZqlvJIMx6gEjT0McMj8ikuziHcknGtVdUUyKyn84h2xYRkP3
Xpdg4c237dyOmbSb1ut53DqUZZzThFA5xbykVRCSWQ5sg03hlfNZsfRFfxjfMBma
NsXsAAwPQoPIWMiqicDLl+4+fwx1v7qQ4k/7BLOTF3G6radskWcVcEcOZJh1PQMW
5uSuvEcw5xueCAhvJKglF86HAKjWprnnTGs9RG+wjrwD1DaQhajxK0psTCoAigNl
s1wWl2Arh4R1XBfmdsMcxWPHToXz9QIXMBvff6mrpv+ZOaI5B0O6/98cpjyK6PgF
YiK2VQH7VVMM83MdzqPzMHyNOgjYsspOOzSGmI/zTclvukFKKYJr6yLQqcaCJYVa
SR4/y8q7IZ8iC55vn0lbeo+d6BpzJoHs7ImfkHPGXgABQ0b3V43kui53EajbnkYf
TPyhJ3r8UFFqRbFb7j6jo3s46UpWK3L5/v/bWedU/ysRIdPSC6HtlGyL2s2BKeem
9Xc236RGyZoNhhJ6xsovoKpKAwY+5wdvp7iSuqC3KAP7m17B/FSGifIZkBUqDkko
ZvG8i7x/mB4QYp+i7bkRpHuRtHXfi7cas0mrd71NCBnsTYDkhQ9c9Xpuc3BOwtuJ
ld3nZZFQTI391y+8e1gN7gXoSJ8IXzJfKpsUxBi1kcc5M38/lDxWCYMZt0ZKHfPV
FxNx/IYQDaZ81CJ8c9fPIwicdKDEXsjNYixWZPKRVWZ7dTIhWPWNyLyit4+ps1Xk
dxwOTwFlOj3ebfSH1P4UutgiXNIkNXha5nrey9HOT4dnWLSIyzttqWKzuOmvKSlf
NZRzf5b6iAVFHltk4jv4YhLtbMgMzqzsYGldXte5M5Kqjv5ZuxTcCwZZ0/4Jztyj
xjFg4uEbSEx1dXyFY6sYBvGz1yrk47cgNdXW/FtoHp7ibBfpi3qHWgWROakEE+Ty
llxTvllVC4gUMpw/WRrQQpt1fdvKLpXD0/k/2rdaHQpSP9EZ7dTsn7603rqcyV0M
dhbtNl0N5ZVSv8svjsg9Qy80oDY+iuxPCLCg49T6e9DaFyTlZrfEgLAN7C8P4u5v
OaNDdfnlyHyfNpCwz/+wy+YcdoH6rWYeg/qo6NYbKe9hXAKNqNYgxasjQINNUPcY
XZDKBnpzsowNxZXp5ol2FsOknGb4noL/ETCWjSauSln5aov9jMX9McsbMC+YTJXA
jtFEgPL3x50ekohle9CVr+i9UrXGEod+FUfHi4RyEf38KKPiiUW6iYVJ/grfXcbP
9mciHt53mEkHFPDhr1uetNlpO8i75CwJH/jzGd4tc27md1uLEEqcKxVgWMT2RJ7r
3z26Utub2HS6ixM5t8P4Ykdt0be9kaqPzINeMC48BSRgClDGhf03LlkuKXHHRWtG
s3puwV7RLg73+cvNKD61vYiVi85tVpNymqY4u1Lugt7jzpWmgwKTTz3uodSrrw29
iYeb5fFDcEuXEUuQvANtIjabEAhOSWWqJAa676ttAGqsnfrnymogQghF1JYevZZt
oor06iKpqi6WkPlnVHYlfdP/8vIp5ZTFTqstBkxcw1kjhnMxh5PuDsmOF/0631FQ
iwHp0qVskAtuTvTjge2AEMtgU7aI/Q/fKWjUQNpJilZ3paJpGRNAJkcNt4mqLbe+
dy/LuWW56R8j09vaoNgtaQWOAIDWW4iuwgFweeY4lC8OOCdlCwhCJ+peZCZ5BDDX
WD1V+J0IM6H+FaWXyLbrNCGwR297YSxGjC8yqp3TnZa7oxQfqRqyxmb55jw2XCAz
jKnM6drAFhO69Vh99s1IVafA7fg6z4RQqzWYYsRauG9ekqevRxIzkTuHxMW3edaM
u6qDCoSOuXqTYI21/r/tmVntyZ0oDrCFcjotOpueWCRyQ1OiuqWZ6VoQ9p+YGRLH
BK0bzBCiUjXuvXXr3C97Ouy0KNwJNAzeS+uMYarkgacvz6EPYITHy8ynxgXbTGS2
FyYpG5jLuWUdNINUMffH6ZazVIefYeJcqGVxPC4WAsWjxLJqgE7s7tFQ0xLGmCzQ
nB9EA0Y5a0VFcHNIZ6JsjHw7lBjrF/PurX59kjf9TXhyWHTnB3xF41rxWu5p3v9J
2JCXDaXa+pYcCaFr0pSIdIsy2hWwZ8UhWJy56GSLQwDo5wfRk4t++dGFa/qY3AYO
yXem5q6lJn5exqr0OVUFC+VU26OamhKPjqnzi5wQJjFzuUsaV5e10X+Wll2AuJzq
IGJDpMWBkV03vmPdIsBnXBbKNLwSGzYuW3xR0adXb+xgYp/8DRfyks3tVp2cIWVo
zChm+YUwfD0eZALMG06BCo+tFx57jCAdTD5rfc78JvY+aNLEBnlDR15C+ZhsidQF
00zCZ/VPZIDa5XY3h5yfoAqvYHMp+vRaxEIsyewzTNJPrzPhuWvCUtsY5oY6e7cC
iteQeR6gfsuP3lXjHSiBRLVsi3nR7Z5K+cz+jcF42vOqAknCzP9+7lc0DlqJYrAa
3/s/kzFnQRQSjvk3Yvu8pKiK6Z4jD2X+b2JpWkL3EcJmIxuzJ33aN3QvofrMfMcB
dp8qbWoRy3hvZuQ902wCw8aSLQkWLFqSPcJTGGnRPuqjuVwPr+v23UNrY/0IVRfp
Qs4RMx/9yGI6hFMEiyfaESJPC2JC4DPtfI1pV4yqb7qd9MHTpch198Qj2XX0+siD
ydT9snHTRAZrA+mr8nu+E2WQyhoomN1mGJqbUMREufop5pCeEtOxm9xST705Ia2w
jJOv2gus9qryGkznvKsxuHYmObjngEyI3MMRPqIohmuvrSg9PyvDtrDUIQG2ZK8g
EzpnLiszOgZlKiP9oLRhD7mLVig1zPsfZiC8BsWUdNF0DsqypCTjZxpgYOcokBu0
kz9aj4RD+DYZVbU95J7V8Qdb6UyueI4Xo9WuMvj+X4RfanyVjwbxYn2ovNJqnDJy
RNQ7kEC5Eno7qn+2Ez0wo0zYjAcxiMBSYQAsKi6MDaPA9zEYQtPo25QGadG/ChTI
OHKCKZ+zHPwc9t8Spdb+6UyvOY3rGAPUoPaS4bmLGwOHjtbPJuYRfIzmc6d96ND+
u+MM+xL2tIRmllxdx4Lw445KVkjXk42GYv/CKFCUntMZ5LcwogZlCGeSj7/HrcPA
adiUKuspOnfzeTguxzbfZi53hDYftsvnW6p7wauYW7reAJdJRVYtmAS6qRo3+H8B
ZjzKfNc3KslHBk97Byge4C3Uz+e5Owb/lQPfWHHf4sNL/u6waIlXp00qKnkzWFum
jPIob1SlFcMteYhLB6bLme+4GR4I3pc+HJSnn/mZji6afSZx3/I5i42YpWPcGyOT
lxxx2nHqz5avBtKEEqimpJMXPlSJ9mq9QE3PBgcDc08v2MXUVIigFVcar1t5UK3z
sZ6NsDERFlwqjw8YIJ10Jdnah/4pzV835d1usE+Pib6JoFiFls5AWasBySaiTeS4
gscFKGYJFvSoc95hjKNdghSJTw6qfnFCtSAMt8iFcSEueiKg1LCFE/jVdSS2ICOF
fg45/rUToJYAOWw9Wwvice7kCs58MY4Xy2Uymu/sSG//Y8sOZHfut5M5z6N51ySa
cewYBeBy7LiBoJWtZ7djPMCWpnMVc+mFi/krioCxkXoyCxR4KcxO9lnbX6DLkxXu
a4cYWxHKv9K9HVq2E/BfK+Qx5eN4nD1UIKDPRFOSTGkyd7PA2bbXMv/qrGHqRrgy
L3vM5Lw9JGQEV2IqmfWBR91nM5PN+YrAQLobg57ve5JDpAA65Qa47je48oVFsJKd
CGkv7mJD588IRnJX7PUMhx6xc1zY2aYeiNdRIOZ9X+nkw0zhjRk3nYJuY9Y8QWOx
CCjwP/P2kMrUiDncf5RKB0Uf+WkkE04qDKmWgEwMiahxcvbCtq1AvebBVne2Wj+U
xvu+ZRHQmJfLGjDvU0ErdXwV2HovDnnUHOznrygdq4IBfvpmq18i/3cBh6lIEuGb
apeSwcCecROW+6FNqos6zCednJs4AkR6Z8i4xrBRhfFcPBvdEsrSfFku3/ANWWy+
cBvGTJvKhpCY9ckfIRwvsPI7UvFV1G0ua10n0nR+SPGjOLBQ8huve3QmJExKRdDX
bOdPupuB0lc4jpTZccwYcnA2xcMub+rfnMnsNntxsY/RqKS1osIFfh4xk2QjX4DB
h2XrM0ypIbAwaCKfLI2T9w33oZo+15DK1vLiLBcTNO80tp2keajoXechrSJuo+gM
XYTYFvtkzsvyf9K6OUWPyb6Dvwdo1sforSroL0uM2CzoTPHaFkt23WfUh9d+hbvG
7JduTNmcn2YaKekRT0NvrJ2rMHAF9pgYDo7ZsPsFa2D/tThVN2aapRTCTRAWKVYM
MfbYvfRtzluDEgHi9BSWZ9lLQVsZrCLfTZNg3wtusmT2RwgW5y8bzfwEsE9+xnbM
FkOxrZv+U8DajatBQYrQ+x8Ael8YVBTugCMh0YlsjiJFrUvwx8J3TdIk7gcsYQo1
/b12wBRXnZ7dkCmC4LYz+kIA3+iWcSl/2h9wIFM1IhYtEzZa5BMNF7Se1fM+5SBf
kadk9JQNZO5XR04z289zONXjlWPpqALApr3TrB6U8eCtUMYeO9V0vFRKjN6caVi+
m1P+CT1EFy/DU1z210FN6amO58H3dCTeRV5hB/OgysJZpjB8doj2RXuNrDjNkaA1
gRS3ywvhru1RYXuMlVrp8lEXVlCe4P9SmIqwTfdzNCq/sZcqWvKZVKcWqTL8rrWY
3YwdrkOKDT9nIClM968AZJSMbI/iHyIi+ZC4wUlQe4XlA6CVA5a3ZdV/Y9NNbYd1
pUHTo/4C1YHWRlzRnTS5UmieqfGfr4RyK6Bb/1FJOtYH4G2Obr+H146qSndmSctl
WJ2PdFkj9PDuqTGfXUCILSN7y++tKG4BmViH6+9V0xP+E4FNeZVX8/f5mtxCJ0wb
YvjAklRIfwFdOgQr/HxKE+Te76iOwxcXUQR3qRZ0TnJrgKW71yCBneh7TTwTpuo2
U3OnqEP7iWbycIbAR3uOxXqNOCHGVY/eWXUsRzEyGpS/BuskQDA/ptG+YDFruxtX
c5bhAdokP6TlQz/N4dofvWtvEhWescQFUejxx0/ouC2LMGhga2EiCfQFGTb3IGZH
IOL/yk6M0jpEHKADlcvpNJIkdNmVDhTXSB4jUMLm1xey6rFLeMmAt/sMBzxcMfBw
+X03Hx85WNzmOaoT+1ySzR3zCtNLWC1vdfHM0fPyXLPkOXjCiLUhH2qIM6grX4Ua
ffbxgDb4E1wSV23PZ0T6k05DtZF5Ixz4wmTlGLMcsi+PxpE8MzBb6I64fNSaTA1I
9jLbhDnjxRTUbm+tIZ+u7gmL+Nh3SL0cBTbfFnaWYs0tc2JJHrvkip57Zu9BR0eW
hHGigpRtE1np9Dcw+HEiLt+HlCLnevjmDCUjwSrrQzGJKQzrYxjKKGP2QHbKtMS/
lpcnWoebfzRgTQSc1whyoTHPYVVGouudPlMkOd5qL9kyLhesSgs580jeT7j0Amou
jYK+vM1adq+JsbZ1d2mfDo3iugPkhmeZat9/wONEUhJS8+PFNOVEGkMOiq+/GIcR
0E0sPTQEY5LNXh3CGSQp8ktrj/fI3JRHIP3vHgUZFR96Xg4Nk/pImSZdJGVvlvh/
E6+F99Jzcq90uYnViSdYSakKOsOGNqTojC9XfsUfPRrIbF1F7VGEVAZpEdPni0ID
CE02HzkwUogVRBM/Om8zbmHv805KOQJBYaF6NCH5iU/mns8Km8HDFmx7TwKT2JvN
HK4UC8DP8VZ2Ygk3PJvyWX3L2hEEvln8vH5JjjqLb+XD9uYyKQNjEuQ/EGIThGuN
gpggLcuzksAOHku7kkllPPmCq4aGrZpslbLzqCGHgzMVD6TmBL/wj6rKk49TXJsx
lFOpiywipXaQ3fkbh0F9UBYqwx3ar73GwPqqepuLdasnWQnh14Hgf8OeYOQ85tV+
EqET3kc+nusm87Qj08yVQdTLElPU2qB9ksarg2Qn7xwZc+Ne87A2zH/91zq4EbY+
uiigGnTkyydqMNSQI+YaTHw+bdJMBTnrFbN0qaIhl8SBUb2E4Gzw+Ka8ItFqsLgB
6xdzho2KTmCp0ZVoEiMg0KTmmXpuel84b2u9dp5Uidm8lSjck+KdLLA5MOqSGTrk
PyESkJqPccXugVERYY7N4N5NgIi2bLfGkvpuTEjT3tWAhJm72y8EayIj2GccmJYm
WpvA6K24q7U8gkcNMRurSMcpjFuZGb3FTha8p/IleMZzyvNLidOBqwSCYqDpgndz
oHKvB3/AAey1USTWLcTw6CO1NTe48EdX+qDDwx6iWM8Gc1BhEcsexv6pYcR4tVa1
kyu63c0RzosJtlOTqft2B7z6m/5Xz8eYYSIK83DUaoD2WWBW/0s98ksShVWvHlZt
oa8NXDdnlTSV+wicXyackUf3RCb8hDOl2Q5u7iqRu3zM9a3OdP3Evt7nzH5ywoIT
k01OpZViBNKnaWuJsmQZ/FVoacjoFjrH0TC8M5AEq31PxTRFmSE02LQQMljABuye
GWQdpqRHhW55HsgvVFf3S9x/gEw9QNWSyE8vWe11aZBQEHCmk7s8F4n4R5PH6OSN
19/GWarb0q5hRjkAGqBb1sLc+SPvDLlwlkdOWKlQiD7pUEQEgI6Ih+FZ4U4NJo8u
5z9La4K0HEVWh37RznIXwXydUm/UtsWK1nDokLV/chFkub0AXJptM4WFVex5KSl3
cRNVhmgb/8BBSC38gibjw9iJsx9oj9Tt9uk/Chd8mTnD9aMPNDkfcrkD3C+T7pm6
K2qkBpLwLCQtYB0KaDcYQpDhiVA4uFXv+9qWTLmom0E9LXRKiouwl3rzf764fM+c
2tHipYWGyAYDq5yyBJh/myZ+RxI0ZojUxe8VD7hSGjGlTOE7Cfp5yfE6dqGU/+g4
2EKMICSNfUblvXxKnrC3Jo8jgv2jMaBEw7wLkPsYMBVn9VzWtUa5lJ/nAwphPG18
Rwid5mDOaMbgWgZ0pEEGMrQfiAKgo32KT6iqJxGsjHmeOuQVjr1hmSr/IjiuFNpo
ZNO4SgxYKWxyhnzIKFLX0Ghtjk9O+QW0ooDpjfc9mZfZjMEmZS5KViKSkGFTGsPI
IzwpFIE2N4+UorDq4XGAufMzMd1e4V3MWYIHnv2BDLpKF5KfpTQPAEC9SN1oHKuW
uFdxoKHwqENldDXEFudb6LsoGNaTKQGG3P75TGo7R3/hoGFIhKR1+pWl2bMzUiif
WFAUP5b2KT4LCJd1PsyA8Sii5t2zFVbZpMux6Ng9VZV/1TCN+3EGC1AdEpNi/JNr
6uDgvb6osCkVOmA2EzKkVkw23TvLIkclBfdFjMkjXacQE/4p1yjFhsbT5bhb8tZ/
yuH0vGdzjyXtGUcATKWDS9JFvh3iL3BGaR/qTWg7M9/U9Xzsq3unYazrNi+lZ9+D
mu8Oa/BbqS9K8A78Vej+WinDtKQdw44gKoGgk/buPGsBDPPs3MYfrcBqCyf8ijsm
o16PIGizn30TweoLpE0ci1hP8/NMXv57CBL3EjSFcBvWdWGrPqiOAHcG823fEGIf
FYdLudEnqPDGH5pdYqMwW05fhBJvCje4rT4P8mV8ibQ8qYtSSjQni4o/1Or95LvP
P9xn4traev1Oq6ML+q5gspGnidsJO4WLLtJI/c5gDLe7pc6ouSBkDWpKMNXce5yu
88SCgly32H8HMWO5HJOp+qRDcYAxQsFAi+ldbzgTumwg+/HynJICqSOL0/BM0Iz8
bn2rLNsniOwaeNYlZvyWfw3tD+CwhrfVhk0olgP6SOipjH4sc2qGc1NMAbbuDRtf
bV5aM8/EX0lbpJO/BbJBM7hYTc8t446nGwodGy8qYoCADhwiFR7SgkvOowCWeyHI
F08HKdDfWZ+Miv+UEtNGsJEDRh1JkSurSeiubukIvaZBrooQ04gpY76CTG/u4wsv
18Cmnmq96O/BlTyldaPjxwQmloPLegAYzQ0++WLOTbclaSThnPNb2g84RUZuUZY2
bmehSn5An80g5ZMVTkCzZHR5Hs33FlqFHxud9e3/uQkuixegfpybx/KxoiW7u9KX
D/nX0CneMPyUaxRIncWI0sU7S3EaIX9PlGtfRcJ/aWYRmtOb+lXDSHD283C0Iixg
rOWOvWmUY+Do5LxQ30BeJSNcQM5GS/pfriyz0v3Dpo4GwydZRymW4dAcSlbje62o
375WLZu9JJ4JeyeM3Hdem1d0AcrfYjVEqz4bLF4BvuMdDgB4IGoUPWLwdmnFkrcx
0AdEeJTR0jrphscNd7sWu1zDErmT1EivnZKsvHN2YliAWPH/GS0Hb1leZlHizMhG
Fy8Yi6cWUyFFnFFMnUORp6Y0BWnIGtZLUO8PPdLkOBJ3HzviKciuLi+YtemQpnG1
Sjte/3vA+//r4kBhHaMI2ttn+KqBb7DEwaJStv9WOnCLEC3so8samZGUSgqieF5c
v57qtAv1IGEfUhjX1bLFPOTVRPS5uiWFmLaXHEFy93uM4qx6TtHRIf0JCyOqDubH
+gv5z1/ukg/HX5/jD+0nmyp2lIYXHDWetcEviikS7k56hc0b/AwRtKWFOEWUU/9a
6nDjXmREEbSYC+xDToVDwLFY5z8TrXYa95PTwHmMEPlJLYt29VNJUVymlsdtUikQ
jod7RZQRDkk0r5GqQDZzgsnL7Hyzs2imK2oe83Qoch023OUIZLbj0457ytO1mbAN
1EuzDn3uUHNziTz7ilVZjLUVz92SMfJ/CRgY6jjS0fFVfuzy1pj4/526nDbGJwoA
ScObGGinZBejnNQzdKi57WFo2vKxE1opYdz1rJ+pq0ewrSW4gWVhq7kbnke16Tya
2oHeS867XfHyU/V6UadAODnsSq2693xmjXoqHlBzEiKZnGEv6Wzl9OeF0i3pLu6X
4X1oNh05gcM8fXF8xNlQwXGjEobtqnybTGB31Jb7Q79mN1q1vP3OoxQcUEwkEFsx
QXSfRNC1jZKImKSEkC+BmFccteLCSQ7CK8QnS/MKaIlN8UrGgLUZZb5J2Y1b2eyF
agyvtRF34XoC4qpAhmXfJ2V5W4vegTmHDZcEnCxTGLOM7+mfjc4Q2HPwVizr4fpv
MNut+C73yZlo6R/segna4zt3sEBhJIgsYvoHPxQFjF527vgI9zl+R/+VeILdnEMn
yiKV0H60DaEeHjigb8SXShKCuqifFpIcq8ft6oAfAxdRFQzpREbgtxWLy5yb/Zci
qr/AlpR3Tx5YPiEgKc/mtIqZdkfgvQFx65kuZD0VV8ejwb40o4tzAwEN7vrGqgDx
ZNvpFPn4dk98MIdmhwPz/kvNmy3tb+QFqLgSRQAOX0VLXIOfPOYQo3I2PCeAf5ST
4OwMVDDF9kXoMaJVcwjMYP3O+8q0SlZxOnWiF6zYfSQPqSCS7TnHq/TsdNOZJ7JL
iqwKMBRw3aWp7kApD0dJ44t54wTaYPKuElfDBmJEcGaN70uc9kccWe9cNhIvCDIE
lFR+wyBtgkmgN8hzYjPAUUki0ve/zfmz8a39o1Z4UM9lO/CtKqS+8MnH0j2KL+l6
/Rz+7txiEQHl6Aqjsm/vWgZw8b60rC3vf89L497yJtLiDvK2CeAY3FSCkoNptLsz
NlWuWMEvoXko7RjWnhMPxeatXJAEJ5ODVcqobditphH5fe3SQJtoiQfHvE/4O74c
yp3JiVAVQAziCjn3fyZMPwvwqkrr72gJXzg9rZr+UYmhW9uA/JLx2MTGFrt/QQw5
ldsHmPITpsL47fGpJELUCvnW5p2ctoUdooIVJpyCdv2AjCGB53RbSVkNVRd1ckjq
nOTYhQIpfzGi8vMdlAKaIKl2duqKcVT9Ue9pDVK3c4Mt0F8c0M6EH69iHruSXPbp
4h9aZMx3xtPc45MV+f+oFoYovxvnmvztjdwhDt5vtucznnN7A/goxN2ipOZqRyWf
qhkiyQRKykGXLv5donFHvobJy38i0B71geRkgPEqOZHJsdECCvWKoK74JkodZ4eH
fE3dn8YzAv5El+t+7HdpuPEBrdUbIPfQjD2irQ0JB+pnC0zKv8qKzEbIdQUIss1n
AtNZefOph/n1v4LoyYlvq098nxNjNC+B5mYLhoYW5IRrZSSAds4MVuzy+FJNE3+F
PTuAzXMJcEOh6xqZlM6UQmTKLVgYd8yVFZmQSxKCIWruYOoLYvi8qFR9U/0Cq91/
aeQg+ltL0CiURUJjuxmae6b2V6lEkavbq9pd/J8wGASfBZ6G9BEnYtAqTNxOIBKz
iU8Iu4TnrrDURl1LMwGwVU/yihrkYrEVHc7kuddidjY9ANzzg3E8oYWmDMfA2Jni
WhABOUsbYevSuPXUpN6+ODzI9NxulAxybmqG2dVhkj49/lGwVAc+TOHYt5MC9lA8
6h1ID/TgU/slfijmsuWPSOiDoluPz4Qh9AwDgTgtt82Sph9WV5mBlfmXhfDJH3se
QctvFlkC7nY1hISKNdHqBdyLTfY6pX30Nl1m9V/bC5Dgu4+uN34XyxKMkgw6PERi
S04lM+P6A/n0HQsMVStSnVJnvbYhgOtzKOMXhWZ6FEkkymrxJ5+X+YGPzYtfLbsO
27UFV8uUaqTKfUQ7rd7wl+kyqV6Ox30tGJOaCC33DwbRT1tcKyKXJcsypb2cFkDw
acDOmI6Gmj7G0qh1KKP297Y/9kxFc3CG59UUFk2+rNbPup0mGrp3sM6ujJQRgT8h
fElXdM5lv1Z6ASnjg0wL070C3l+72HY8JWEcK9P6d3+/SPdpEd5Cz4xtG+9pHA/F
RXXsPBIelkcrSuosLo4ALOckZPAe7/Iv7DWjLt2SvavSgnjUP923q/UPJJFjxt7P
svNDRFOk1SB6mADS8mpACzbSvfd7r3r9l8mmgs+e5IvWyKxTmXNss7giXqzyRHYk
1FuBkKO7SszfZ3J5Z7KUf8OJ+jIBMULtHtBNgBXmfGiBGCjnlla6hqn/Qqig4uwR
ZG3fOQYfjtyokn1htY3Ju9J/+qZ+cpBMeqFycVtyKpZlIcCSKBYA5Vd+BUi6FQvI
HEbFV5QrHCJfPPwm92bOsoW9uW/odjWnL2ASf4dCthRyeB2wxhA4r6txfayqFiA1
j4jisph5gWWZm4ay0cEvWVyOFvCHUw4wSJ7unofRNL2+g/YwORSZYDnrtZtAfcLq
vJ9ixKjNIZx5aKoYEj1E07wyR9Z53B5OEpooFohDbskn1uSxND9DANxGr09ttqwU
PnxvUExsqA7DZkUoN6a/YfB+6W8NjNVItI1+AhYPXIjuzm6btcXNepK3dun+uaQz
p38aIzHI4kwZYZIlu/0Ie+qNbLHQYfE5uz7o0IsMltOP73SKAJRu/t5Yq7FiE7BB
l1EqDjRG3T5A/pn9fB0ACLZd9X8beKKnsKVBtoGHMx0BpcIBKSNLb7l3nPSHZnLc
Lvwt9AFlbWpOeCi4N6oYYCWyc+MZ/PtNJ1QXEbn4Ss/XCOoOPtHVFg9LPcr5sYtZ
lr9eCr3Di5nQvI0YkWFwWt7ClMSmgYz8arjKHVivY46MUVE6A6mctD67rR+v14cx
WTcWb20ix9mwn8hHfRpBE4WaVkddlJ5nOmGaAr/Up8obUAboUtW2AtGP6WC9CKz5
XCMsP6+i9up0+wH/+i1rmblvMPgqdWUbdwAEaLIwFH6X9KKirFZcPv9EPG6a+HMO
SFbp9Jr2spwSoZNsTbONZW8jK8bsYSPo6cihP7WeSmb/ncOmXiBgL+WR/kcQ6cBr
Lt2oCBGGbH7psNO2Uu6nsMDpiTR5k1WJTu83y/0nDJYtbHUgI5S43OndbQIZBy9I
/ibcAEYJ1keL8TZDqOFDGML76GlgKOnNj+ySmg77loDPFHxjm9XmLm2jowYjrqpi
eO1AXxr9xm3fTSPg81FE2X7lQNPLjga88bVB5wo36WcAGL+3SX4eeVWx3i88n0RQ
fpUTEXoBe+RoZ+04KcJpXmpTg2MJwMdHF4fwDXqAE1768xAFn+KTB46Z3iUcX6Km
wz4AnRIbVB8IwbAvS6GXCwGdhCxkzCXAf4HTMfJuBJ0/LIQXiLHUHkgj+YWfMW71
g7APsjkb6EQq2NHqVro2+FUxKd0PaFN6p2e6Xqui/Cm2gXQJcm/yHU7vP1xwqo6i
K/vVlqXxtFUXhx3DINTXVMp+0QLLUSCd2wKhv3UvEqDN2qQx6Fml8MInmZErARnm
CVB1aIOmyPexdu86a8FoMtvS50XjT0bYj9OGAbba0547n8qq1lNb7fdFvfGS0nWe
M2MWE7Yw22k/9IJE+TM1S0XxZUN5a4MwMsKwgitDH5lxjYVwuktkuGLLf3wryM3j
dzCMlp9IcEJlOUZ7m2PtlBMTguklJbKXHD3dWuc/XrW8KMCAz/CrtrrwQNklC7qq
tgfu5CzLAi/2dPfBuMNBmYtvpsQ5cJfsvlFqauxoqVEZscqkhOALc7RCiFhnrgJB
yNwEqsCb07oFlzYc3gipJEXUE7Sf3jReQNhOUqvhi3jcz4nQx76UZyzKvgJoVpBy
CHbPdsXyWNNpr/jnpuaByTIf5YLxCSqaL4BpwxCFWxcGwntlF3LsWk6lr86dZp3o
Fs3h96fA9+CrGR0n0Xo5Yy8U8B5QgAbXviBKKPROdgSyFZvOFXLxbEeZTfunEYnN
WNrNXavC03Z8aOfuPp7a/dpyvUUkQCxdKVyKy36962jq8HqjQBu9YLObgOCWMjdx
5BKiO8FC9DSc9O0rbajLxGfahnWvfGM0aPbXSgX1xob3soPUyp3CUhMc0mVaejJW
Dr3DaNX2YwKn/vs+JulginTnRi26s0xV89OCotMsUIIddFVyiAh9bG8ayEwAQr3q
dQpkWVpR8R84yvy94RwweqZsy3C3qIz+2ogoHN1c+RbRMuZD96WG8N9ZjQM6qUuJ
VIdJOSDUObh5r22o62dBu9/Hqtlkh5wv2/senZrgI4XV61QEUMOKm7NuRZiJEmxI
XInAeiMpoL/Oy+524hwlrbdqzoVW2wJiTWRj+H0C4QJn7Fmd7oobXOq+66AbM/Ff
bhCH29wx4LihC+DsxugwAhr21ftwON/IP7+6PFGqxODKhkDzaKkLz/5tJ7ju8m/W
b6bqnTQm829AAoszm00c2Fh5ZuSd+wsGX+POnG/UIdYno/bdXe1SzWCnhgFdLIi7
IppDiOsdaHfnWz4pGSAyqUgbNpoizsbfYWbN9KDJHMvAxvACMZifhI9dIiDDC4Jq
QdbExDSQ6jZKuZ9BW8LADETFOiY3vy1aZh+TgElLfLH2ehcxUsGvcIsgTd94I7Vv
JkTjehxeGzkUnlE9pnntR+30yql4AOBXcuC6Y0nd3HqKF7l3iBWSH9uQd4Y9Ku3S
pM21Af8HhOb3c2QI/uQ/UOsdpmTM4EFEXe5POW9TnYTwuRhGcSw8F8q7i6bu4IRy
gN5mRw7MQdBVjgDmOfmTd0xYITehzl+zN+8sv9fBaTuUF6CotUniCIKeJNt8c2Xm
HAt8pc5WP8m+fQ3cCO65D2RRrJRxJ/aznvO2d/jPK1XL0XA4UMwmFtPzq+IqNyOM
nZr0MI+L47DG6vnQBpqy1Fcrz6dHvpExXSRye71Sansb4oxiLyhxkoxIIX1YWxLt
OBVFy9gbeV2LsdEoL/N9RmO9nyndSlC5D0BzvzovAZpEyp915A33tHzi20Pw+QUt
Ij/Tx6uYIUfCQ3AXl+z6DXG4VR/KxO8n6YDodMcSVZiaIBQogPqMC4Y/rVO+Td4I
8Av6aM4G4l3NpUCA/LKXWCxgQi/5p9CTm50tkyocNZLPaRpOBYSgebYK0tzbk7eX
eJkuPmzuj9GsADeAOHfhb978BCX6ya2Yjsw3clvGVgKwrZhrET3b+wfsCzYArImJ
+kF9d7qDXPGd7gauhPEEKfncxUO6YkiSYDYlLa+LRy6h4ERH2HgIlOjy59GK574N
/Usu8BeN7CUK2lo/bDt3YQYTJHkfZ4i6f3t+t5AXmMiRXcobxnRaYJ4+UjhLmPCH
3cbCaaQu2a5nx94hvENBgGK7+w5n39FWOpXAhWQKgmwlkyQrof3Q3pvWWGlnBy9J
A/PehtbpF3vZ9f/pTQdBjofxSqlryqxNAPxk+Oaag3Gjh6JjVKil8QYMYmP9BxVp
y51RvMxPp49Ep8zd4OxGJ6ZjGGUWjjx4wBPK61u6CiaMeh9v7dROdcjCL08sIgjz
VMuTUO60d3ezjGKP5YP7DnS3OnRWeGLAw8zTQiyVMo8e9fkX87OtKUVfIcGwg0zM
d3FbeMwt+vEUwBre5CVzihzgeOiDLEMF1vui1svpxAR1Xvb+N0WHgcYRwIAIrdUU
KMZmaeai86YfP9YQMd8Bbo3MLIgvgXz1FaBdbw+OVXLFiAOi1ahI858qABQeCGwD
l2g1YQqVTHHfY/N4HhbdxxSEx+QBx8fnQqm5GN8iL/f4uJ2NFuFN8k8I+Kj8W4Mp
hzYtcuL5agZzJjKDJeGHMVNORs5Tou+8BTjaqpf2ztrOOAlBDQqRq2YLpxOdpExB
Fp39yadwuEv7iQnYYSeOF3TDD72tXIGYMee9oBOwGTe9l9uUgyd/2vBjc4rwiv1O
VU6tDKLuGzFN1j6T2B9M+pZWAio/FK+uBZnyJl+3nTVQG7TX38510kJuiw6bF677
g2ayQjLvJ/R0vRzPPg03ShqRvM9/4dJ2rLUBmTsFRUsGaG2edPUlQ6tE6UmuaF+i
1I1kNvJEl/zAdH0XVYN1asyYo71HCg0pcSwAwM/vWR5B5XUr8IKitNBueZf3zgTc
5lT1nVlFDrJrDtHcCmd6IfcthPcOXJtITE04cNqcyWfmHoW/LiylrxiSDyD8ORi4
iY1xWwugv/bD28nZeVb5oRnJVQWzcptfvLRoW5RK8ZdfGrU3v8zYqfJIhtrY40Cr
HeLVXvoxjBU8MIPfkqAjc+FO+wpsoBxN4x0JOFe7BdM7RsjosYEb/3iJ4xdBW+LM
4QoJ/fV85dFHihTbZSJ/4tgBxY/6n0pHM7/5bHMiiIDwO/nANm4hbaFtNM86sTuA
wy7Ng/TST43Z5/j0LEQLXe4PiVaEDPbydA01fd4t5mwLEo+yu8VWT3ZKY58mc/yU
QdN00NajdcQ7RkPzMzW91RLXIY+iRhnCrPIlI449ygTC37jKKjzk4E+wQgf5fgei
Iv5rSDyR/z//PnPO0R3ubY+UJUAg7BUJc5YOcsp3pjQOx72eqnfkcmij2DirbfSP
sbUl4/qhG9xzpwOyui9Xj9yfDIjK5vE7pKTNRxjKCRTL85f2R2RQhpoE6/Zhfmuj
7eMUtoqcaQZRGDWzWm3kq7xvXRy93m5j7vtX6NOlYSulHXSLjCTh1KzY0kDlWuGC
RLn8GnOXD6eL0yq/uLdI6LcXUQcVWIjEmrENnTssywa1BoUwMYp8AwHa4FUQlvHZ
XZuVUSqzZlmmzc1stgwFVLJKrvKsii3g3bgCqFnsnXyXFfKO7boC2w0rUekBPEMB
KOEl+JHXFcgZtJXJIyEzV8sMjalh7lhVeYXFOGKZQlA+AUm0Aqo9r+fsq411X8X8
lqYNCMSC9oet0i6PKxaiYqiJ6od8/Jg6mZefKhMOpE2m0t0meDQCnbX7g50Y/8Yp
SkHxyEXv4kFY2y6ig+vlbf5MRUDlRRB5TQ5sA6cegL/Ze9hTNuYok1+wIPYDp9a0
RYssniQRn1YYJUGHN8qFqHLGbO/FTpqrQ4eJgkJPSUTVnd55LqU7k6ZlmQagKSWv
NX2P/egMDIW6yYxV2PDCvSBPoBPhik6sDUXOPEK4ZrTarXVMOFa/tVs+WVZxb2gg
Ut1xXLZqhSuLEMknfAH1+VC1ZE7qtwOdz3qVNXtE6N3uz8hADxc1JAuBW3jB8Q0s
BvuBcHUwWrscSoxivioPQQinUzbpokoWvLTCKvUTW/SOLtR3EC/EtLzQLicVm57E
4YkmINLJr9TFFYNwbviELOZntT0/0d/p/VmgpPjeU9Upue/5mG869j1Lxjc3G7wS
DzIJfISrNy2/Po2lb9TetI+rPjDGZOqwezS1TFf41w3iakN+qL1e3FOieNAZDKv6
fo55dr6AT8pltgux+Lhs7l30erUG0bn+OK0Nh9BRe/Iwfzer8Qsqx2UudPRaeloc
Xodqw+NfKwKH9l6xDiGO69Z5rpH8Xeeaxrr6lyv5XkaeQ/TMKQ78PKUXfQKnKrTY
hi9RmE8tGAYSjPgJ/hC7jTIdWwpwbw/0NzAEvO/5S8Bi2Y1ymBAdXY34KrRRZ0OE
lxbfn0CLuseTQdn2attNamAp/lD/7NjG6VdJGRThbLIQ9AjnRHC+p8JZo/wEgrxe
wh38MrTuXprPydARXrm4cvYmHJ3UWNXCBfe9mQMV5T8IkttXgNN+F319Yc2HQmhx
jtZsGkulPRGUj8uwrn7NWxXkfscBC0sI+Sr9SujfQRP72BgUIqwWhzbBpP90CgKC
faq6E0sw5VnBQHk+sW+9sQ0o3B6aWClbcHzjIySvEwUSqEp/V7NxCJZzC3YRWk0J
BbdgGvJUDnx8niwr2rC8ykuKBINm01UVMXnHoDAy5IPh/aBpqlJrMu03LQN+o0CB
WKXb9xqEN2BP1FXsy7sRvkmj4yG1xhBhjUFnXsDLbR83KBt1B7KJ6dPCkdU6U/jy
36YhPHIgMNfSIq8O1BtV7MVlPQ15Y8R+xR1UF7G2Z/2so3THuw7ci+maZ10Tgn8q
APYSDH9lgnsPVhDtTzHCjtZSLaNx2DwzRMMYLDfndNXj5Cg4qk+esW/Oh1UmRhPS
eNDoVFpfFtdzyWMRCJldiACZsEUO+mmtrtkCRV+tNBb5fS6ER4QMXCOWtlmZWNfU
N8yRbsIAOAI94eXDY3BJbD1ZSGSvjyg2wqc0J5ROKiWsakbTDwsdV+WlabjkTpKe
Ou5SiQCFWkOmQgdSMdAj8597eec1NCPmdPLXdUR2+DmRhHHSmlMlQU6jW0KOLIPC
0DvjthsDWjdpItR4tnLjSZWv5JLpvRm6/FrbfB5aYV2N/18SDjFSQEOtOlFPRtGM
7tdeq4mMSFaTBkTKs0qCkiJLPj9y0d2/RGXoE8tIApGn1HE86RlMcr7CYf5NNkLQ
XEmHw1+SCnyaGhfd1CPADuw4db/xHJgeTE/4j7/L0KIoBBxVXZV4VGbMRcwSF1rV
0LV4On2sfmqVWIaL7UiEe39bkTiAQGRsYEiCYbFfUysCQF3XpQfKrRCfFzzazfzj
Ce8dJ8fZ/DoQFBSOdjd27Zg+vu+/ArT3RlaHQ3qTQ+XeCO4We0ekc4kvpSJjeLQM
vZFpR8V38yytHs4M0luUJS8LjmQ5/aHkOYmV4vNv2jlmoELBH148c6JS8gOYNkXd
/ZVYHBzZS6XQTkHO3t+AZMqdxS92sstVCCDOmTNfz7HwqE++kS7ERz6a6DdauFCI
gfzeQ7mlL1e+Z42a7IWRRoULC9V3kuaxXW3D7ittO4H14bCXFTp/5B7HPlypSkKH
kuf9fVv9j4cKInvjwN5q+pzo7qMnK2fYC8rNvYY55MVAd/WFYJTiAIKJjMWyMnCH
LJf79siFyiGppGg1rkEeMgebowZI6v3EF/vNqDOXZ1MTyiwFDCZ7198+lL2VA6Fm
Y0OTfltMBEUHgz4qTav5WMQGZnvR4cuxEX2yIM8lC7EFHFoCBopmMzi59tzjWjEP
EM+MZWsx4OEcUlqJ21W8Vyl9M+X/HcjODG+O7CGmKAhHhJq6PwihwQBP3piI1dwR
aroI95AKngRSbA2DddgohIjhRGEsOaiAPIqcnPSDUz0b87/SOGIj7BqSS9BgH7nF
jA4uVSLOnG4fhjNYMGH9MQp3gPLxDzQSDRrpUwCU87qRwhTesy1t2mmi1L3ZKCT0
WovMM4Tds7ed6XJxgnhhKfV3G1+b98n60WGzRKJ6pbhcNI0lL3GgeVQrlJirFXe3
kEw62nijEt1/6OlIymGAUkCA1u35TiqgSdynU+Xs0okRd5A+4gmRha2UwgpugoXt
HlGoIC7ND6v8DthLxJe6duEt7v7suDN/H14vBveiMYCZn5yFiYRuEEGptI+frhqW
JtDf+OAILrUXvWUtLSD7x6hDo3yA1NcZnelzBHbiWw9/p56sifh4G38SxOrpF1ZJ
NaKW+zvTnXUTTI4CJj6qd1pcnWj/bIRYg8KdZXybOsil6wS3xl9NWVmifGXW60cC
61CsHTaiKrBvKgZVdwvX1PQu3BMej1FwIq2z5SQRQCKW79BV7hGTCsQSTE1AxdDr
j89qd5RavIefg71NK4bHmMAZL1VQUYdtbP9wg8+UhWwyVs3BL/5qRc1wZ//1BfB2
ShkrohQ56Ua8YHq4CtD4RY/X8YBHyyGW8xIzj0bPHMSLdtweh9JAls8OIpYOuJLR
Z6ff1YobymrdMhtvOBMm9q66uqwy93KfXfw3sVcd3889NV89so40ecA3oZ300/TJ
Gcin9xqpVgSAuet1k0pHeK3RQrfsAYd2t5BBZrbT4BVUTyVRaCQ3BEQYA//EZt+T
vB2rf2RS3GERgxCVlmjQzqNyGnADZSNNrwrzCp48vHymw9xnCLp6Ry9Z8Pfq1gKU
hFDhc0rTuYqXr/VwRa3k7+sbkbn+0cN2+2mzq0vifUgCTg+DUHJ2BwztnB4aO5lW
ZcrlPtBFLhIjpQaCl1ybQuwE2cV9X6C5vs7W2aCO4xenYPxNoRVJVx0c3NxPpmRU
ThGhYlYXB48L2K8BFq1B9jmEKSkQzwL22Z9D9DRSobRFaRQ6LSAjIPq7RT/9oE5e
AwI0qABKGdPal9Oq2ofA86yKgTo2BlIzzGBs9JwuwPaGvnhWFH/4DpQquJsC45NU
U1y8uEVZqaBvb7iryX5Aas4OKi9NzYbfvSQAgll44uZqHdUTDZ9Qke6yt6cKX01S
QDM1Yjh9WeLklG9Blfr+yvnhIl5dL4+Aa8Kz9uS1Lq7ODIF+pjbKI5YD5WD+BoDI
TpQmPpPzrTCTI0BO7OD1xH2whZc17scLd/B6O2GU/rFBr+FtA6BJuNxBda1gWNip
q0ODWQzTKvRnVRwHTaVWrfbvMnjddOhr/ZGD84RLZoAC2jcR6Al3g2fDp3zLi6gO
XIZHqBEEmapC6SYAvIEYtJTHQKNQhQN67Sp7zgf58XRdoA5tRqPsrgFcDpIHrgKL
c7dM8tKQuUVM+rWSYnQ8nLy903lFugNuCcRRzqOxcoTpeJFkDmi8I1mpPzPjVDlT
qR1DBkeAb7uVJvT1dji4OY7CP53pSiHAaLrT1uJY0iKZiv1aVC67VGVgxhwW8j/W
a4AuWpfWuoYKtBtGOScOKpxG90Mmc1Y+2aufZCsRQYwwJJlWS/8ZacQLGm/s96tx
ZJkpxyG+N36t3YxlIeFLFrYOWTdkb0jQOiO6dwSxZMg2oYds+s0K8d/RITBmCgyW
gDmlxDWFqHTk1DEFOAsOAlRrrcGrWml8N5OQ3Ywh8s0eMwCK4C9AJjJMglxXVPY+
BgtRerDaSIrIz7eUz2C2x0I/BdvG7yRrIvPh0dSC0E2Sntb96DUphovaLm+dLWas
PuUaiV/FStpFLNu0Hd5ZCSCEqti0Qde4rZC0inoi/n5rPIC+JHHwxvhVIKuDh/wz
ZomoLFkRK1AkyLceVEHYnJ8+Q0nXDT9gj9IKl9gyf9IRNrTvRDUFEuuDSFxQpZ0t
3A1xmYAIAjrk1WJQyw294UKRmyUaaZejA+ZcwtuuE4Q8C0P3cpppEExI57WKGN/k
GC1yuxowX01hqZEoP34FE8xftLXlDqNTalGPaFjN3oCGEMO7g4zxvX0a/g//Ak9k
m2XdHPgFi99n+LX84YTKL14J6aPgzovEeRhVWjX85ekPnzmtI7kQrXBt1teixfQE
Tm1N8tijh/pq+dgYVWIZyzwaI3r6BLuQu5qc3SQ8mulqsSQXFtcrwP3U6K5QhVTi
/qxEN4CaOxeRdKJjTm4RpNZxfPcyFSC4qZdl58Bo0gJ/ox1gcxNIS4Y+ExhXxBLS
pFs23eUIIVwAG6Z8brFuIFjLLwJpSfMzecPmfrkwF0RGgBCfiIa7fuKNaqoRIlpp
FoSnJco4o0kqq7RnU8iL6SODu66+WyFH4ieWNTq3kOqgTh/sTAtrWgjrptj+RlAR
zfaTWpFF5/k1AsVsMeZybvpbg5fO/Q4lK/BiLovJK9Vyf+EapiikR18BMqO2nAd8
m+zfAF9x29JGUnXS3C7/Lq8ZZyayB75sDdraayw7v6KazAX3nXjOXWDNzhnWcE8E
i8UMSGdJyGTNbuBQgVvQ1R3VrEkRkYNVDfqszmZ5Y/Xw8Bw0veWmK6PjTEjKDM6J
tFmg3B4n2yaTfBECBtchWGpJcB8P3Fdv+lay7iUxa64sdFS48v4VGPxmBT58e29p
SLAbeeatB/I5WqKg64lxvTEiwY6dBxktRtSWuXZvg0gLxNjo/RZIe79CAT+bwsN2
aYrDzqQeB1jt0FGwhMDbPYAquWeRny4Y79hvX7uF0xZ17jU/SFWqF1FtUlaTJcHI
YrAk41weYryx0+PfVmvbdQHhHtnXvsqyvWXhz5FG2TAuOBJKZm713tjSv+G6pVcv
Aqr/2QPqkND4PcfM5Kjs6/BrosA9CvdcF8pVbb/Xy9uMNkq3JMFu2F/bjoqbUITv
Uk+IzA1W6+DNcASsK2mxa9FdY2Bfv6IBtPOGZPOQH7T/N7kv/JQGV9kT2BL8lueC
GZnveKvx/HU+tvKl/J9Xr6FkynBr8HcCoITtU1hmt93MXKGK8JLmupGg5k5Wn/9R
weHRL6NV9Iv+6qFZDTE+K3AG80sHYskjAUzLeYGNvenrrYJvBQaN+FuNrO31nOaX
Acn2AQd6w/KsBope2AFEXjnrz6WGMnxdZDBCnJMwD1Eu8hcvfdcWdDX1IyAr3JP4
j/nlmgsd5UZDxlCUpjkMYxP4DNqUnL7jJV3wuqUauZdZ4JWShCG4OXh4cpuAgLTQ
deDdsy7dj1q440KQ+ZVaP5gQ1b4aYOCwxLT9mV8LkHpQRS/MOTiIwkn57EJRYd7O
JUpNbUoqgOIqLjCDjhUzu6IcYZSHXkzpdUf0oJggCpcmkaJ58OE248Jl7/pB17rS
j0L0EMSuCF+mxz37W4pZ/zRI06WBNOQDVluhUGPLWUnzNGqU7QLfpgi5a4rdtNPo
w4AUt3CF69a+8wP7p4hW1q1JLWqDAo8SPqlO2IJkOMDT0ZGnzxee4HSeWE7zouuJ
/kU/ttvG59+JAltBSvYQH6NpHWFQq3yaI1eNmHDn2bQi0IiWESO3H2Nf1OIQ8FYz
xdltyJVTjbBP/g5M8OzVMI9sMMk2IFsMnLgafedkJcJlTSZ6V8443dNVj9DmvoMb
SyDUNX85yLYCc9WHkRAAyL0nW8BhIHfqQXnoILFWoJVXSlbAyBs6P8g7PZIftpUr
NYJx1Txw/+7J9vF7in03XZbiPJ9i3lvnaZ5t2t5ttMOLPaXbyzX9zuXjsSl1Iefz
1unvFQsvZlAA22lKnNgicMucdXfBSWE3NA8eLFj3BSWIucVGMYMeUFOv01gveEYh
RDZIZj1xKtowAn6UJ7m0gFdYb2tuhALb2p3u2BCor4qtb4wG6nYj/DQBQvtrNuzg
O9AgDER11Oxc+0CwGSWLBIZyH3fuOsF649uaEXk6bG9h14Zr4TxAHwfsuvamDqPL
xtdpStw3BQIRL4BIt7VRn8Qw8yS+banIuBA1IJFPNaV4QHiVpY+6nCziymCcc8Ca
ud5qh1AxVyMKtnpKAMIQK7Xc7+XBcJxel0aegDWz5eDDk9cE2vRMH1Wv66LF4lpo
fC/+59nFC+osiV0CNVG0gv/9xBmPy1G/I2s9rfUkTaipZSA1ID/i91ZgMtTJuMdv
5IOHebdXo2M0hXHxNJhspQ8eU/BaPKLQyv7/BkErRpVTxyQwfQFzQd89RG/wHRzk
HJr+aNRXUr17zDLcgaWnypHZ8iRCChHN/Vz7v+UjkBfKU07kpScogQ90zqQRzx0y
YgfW+Da5mG6b5VUYdmxz2u7i56U2glLZOZdOiklry0fqjyJ/u20NYj7zlmBOMGeC
md0yjOyfoYiMFNY8cePRz6flhxuTdc5Tp3KnuWtqvOqIFmg1VW4i2unkaVUJw/QC
JockKWl+TNeIcSlgJmS5b9j7vuzmnGpuBdrqwo7WESECaOwHFhFfdcX+1xYPEvG3
Kgp/A92qLw9u/acaA+4q7nkB3/aUVThdSY9vhGimgyNddekv+Yctkf/RY1lPwKcX
wRz7go0xdsPxHzlW2EopGb22KZClZEtharBBFUgiQ4AfFbMIxaHBQytgPSJiotLd
h9ctJUPNhTkAc7/QzpRCmB2rrpmpzszwkZDRoYFdedatwa9uY53tqoa1GjzZZ6fX
fX/FbbuXQN8JgsrXZ+vIzDKngoooANHKXEYs2POPBaMp6tZkMHmxwPKaJ5s6B9RM
o25/otpWMwO9XY0KWvbOIH8UtBlstJpn/Kqm1mJy196XgTac1QMxkVquNQ89HQ5i
wVhRjdDDDXXNraXu2+RNasrTBB2tRBUqospXzcJhJkrP/JvC55i7qWI2xfcwXuLU
IKGwMTZfCw5rlmXKwSYB4Wzej+eUUWjrPRp7mHufiy5NPZFcJRmnedTinndMKFJj
a7mx3y5gb7PlxnI8h20/ZjJA9GN+tSuIOEUFm+NhoOBSSypzppBkBpH9jGvBDoBl
LrUF04Q5RnH1wW/Wz11TNkNEFlNCVsLGAWDzklYU5Uk0uTtwL4NAvAq4nuNt7rhY
Are8Hbg5xbBRoMO8ze7zHGZw4NthbggVhX1ll2I3sdpKLBtKHPHl4sqCfBaCdTNx
GErnPa4xLEwgNZaz8/KqAVTqW6yu1tGNTBdYtnp2wuVhy316wpb0dX6aAKyLIJSa
P8fPf0G9D5iwUdhznX+cL6X2v0jh2wZzlh/Y+ZmqZ5165XKVmVbuntkq9GX4oV0Q
gooJo/fWhO0VAQ6UDJ1vHDOVAK+hQP36YR8a3YVLa5RWl2dOh0CTDVEO6+kmXLKL
HCVgAWoV0h0PIhQjgZgZX5DzDmJJn6wmQSnPT28o5GmFya2dl5p0bNZzhjvLGNPh
hen/HYWsueyaQQMubhzDSVw1xLl64tNbrfEsbxm0br/SdzoKpq74tcQxiznGXkdl
MtQDrYv64b1G7ZdX5V6X/N+olsbIxz1kbHJEQSDBiQu5N3dQkwTgG8U3OqPshW9Q
6erZ+0zXRJ7s+1GGe184zfNdspwuuA85BQ7vjJmh06GxUSRlKdnv8voGH9zV0gAI
i+AIatYtDpPvNAhNzKEHkvGYTs7CtGK6TxerCicGcKx5a3ayf0XPK/sbyYIi0cCA
VnAdDHn3j1yvjgcUQCkutF8H1F6x/dYbu481ndADafbRaF/mE69I6uKZYFiuBOfW
T+DsLoOiudCBQtuw6wcBPnH4+YLtNzd6XZctnEOqk7XSOd0XMeCbCUaubj0N8nII
SbT9wIlrIdqbSJ+p5R9Sm1OBw4PmdPsKclQlqv2Yy5X7rtyUX8vXPU7e4Ag2BpnX
L9JQfAeGpBjY3o0djN1ruJaZanfZBPqRymZDxu5Pey7qZtUZ7ZH9/R15b9/IQNY0
SEK2urwvNrf2G7BGCY4bCj0Ue6sEK2UETsNu/G71toOXG+P3MlR0aWOPFFEmtp0V
+8Pmcfa0T0SFLZs3Uq0Q3DOUwifq3F+ZtY6rmVGiCYws2gggU1LUmmYQJXFqVtyN
71c5UwY3/j6wB1ORPft3FTDSF9pyFsClKT1REZKN+3ehA59IsXsWHKG1CANLd6MQ
I2kWHUlQ6L3kvDJWSniFMGXLhZcyOG/Uvx/5SdmnLNpI20BD0MuInqtCk4i3w6nh
zhy1hTK/1Ft1aVTjy4Rrx4iRcN6sp4NYrzQ9pqkKwkvk9JortNIhfm5xTPWRPstC
GuKE89VRF9iuDizf+IPIK5PPvLKfMCruxSJWGBSf534Ry7jRSVQHmOubbpOP0Pjh
4eLZkzaQgQw2a7Wbxw5vyQ+p6KI2gNtHVWgozUEY4/es6Rq9m56YGCl0OMjcVEwo
A2gp6d4U60IXrclvCnMYsEoVIIhiceaRIr5/hPKBmPvTk6N+q/lh9UV6yzpZYBZo
RSGHiDacow/68DgfRs3zIwBu0rBcPc9jzpGuFbSsePqKod8/8fIy1PkZRrJTGuKE
jdyKFgVcE9F6N6pOKaGzXppnem249NigdfyWp4Rz7v2Bc4B3/GUF1bOjAEF94Zy8
c5GxiyizFS/qaQs1iS3Kf4sclmU254Ybn9y66+Ml266UIiU3bCxy5ygO69zD/+oS
aLa21gk3bkvb7gOCy/rY99EH1wchE0ld7IDzw25vuIO2ETcwNSxWmFo+8uONyWr7
jRKKU5CyniGiR2uklq+W3pFT+nhgIK6SthXGcNFV3/4+zejdlrTElwG3RhgvxzyK
xFUPE6raKk6l3CNOddWHaZOs++10iMvrsmvLWxJq3aJmkHEGQdIU9TSlZWto5BPW
qOaeieQZXcY7+MTufsbmBiRB3vwU3GCurFVOwDDTwR/LedOgxNNsSotNCLgwadD7
r+OKQgD1Q9QX0EMyIg4YyBQJAsydEM4cokHJN2qOv3FL99sFQJFETLc3B7h4h7L0
t7Odmfa3C/yj6JGKW9Js1eIMefof8YDpQNIveHB7R3/am3BcCj32QOS45AYxvZBq
PfLZEtD4sA/0tVWskA+zNT/tair0FZBpexOunnALVlNQwRPZkcS6sojM/X9tu5XK
8kCl6YMum4P6LpDufdcRQKttj4R2nU8jE/RY1WenZNYHpipLAMpkfsThRPvxuQdq
mvDi2TGs+idR1xYQKg8/9cQolgPSmo0+ZEXHbwrfTOO71EnBKTu6sgCaTxhdBtzR
uLTKv2M4tQFKKPmh2F+oInm/W6CMesUJ0V4jWi5ISpMgll24CnF+MkFy+J2wz2zE
BlR9YlREOfnkv3xej13Rye4X9lE5xAYMeqdixYH7PSpZHFOe8AVdeZuPCHBMqYvT
IqgSsSp4V8PClK7JTg6MMMdjy69zydwSw6tjOeOtPZ5/G9UlTOctSHcN9UVcHg2c
dKkRcJQWap0097d4EW0dmm8IEh2bcU7MLXGEnN/npz/dFMxWgI8gnF3Z/RQ0YUc4
5jBhvP/GFBk6WYBTmbuxFsikAbcxUwYOQpsrxuPel4laH3R7ns03fqstY9wx+TOK
LPfrhPX6OfDWkJnRis1LqAo5LGEkGvAyflpvBBgSEw9PxtC1ptnfGUP6OwfBgD0I
TWeuKE5HeSdZmcwRALjFG+HQq2fKVNyY6Qwcrp1+2fBnNH7TWk7BmnR3M82wRNN5
hqW699vYa4Xefzorh7fBAzDAeFZy1/j/vdXKOFSFlT07UXAPmjFSaexhEIxtAGJm
XGWDHFOrh0S+n2xQTQygRMweNwMAP4YpSWMfxbzoZdUrWyUFrxyNCQ1H8W9G4YvP
y1jiQQqPWFu+eyohHtWmw6m1zJhKKtteNz0I5vM4cPNEXsEgScN1JvIuUWs/hWsu
9bopsBAzd7cZF+O3jCGdamuoj+1ByQIM+xwwPb66+E9NbXgYEon6YCdYBFkK8gVM
3duoU00owuyoTDdlt6VaJ9MFzwOUpq3qNXY1qzdO2Kl12q0afyqAujfYa8Ld7dky
j14Xvmac0sILMHaxlh77WDUm7OP014qgVqMVfmCvP/dbv9GwRRggsMgN72WJFtkW
YN9QMxFGxdgiDxwrZ2NQobsFBskUvaXH/+OIR0lUuy0vrYCtQsrx3NfRUP8YPQrK
AMLw3CR1rGj94uR7oQIIDZdYDrlM+gswI2ajKx3Ok9KhQLyDXtd39mfa+6DYDstj
ZoXfia2qR1I6mn/fFfhWbbyOla5jk13HN+DFkMj723GCGHMdopPUlbYVbXaF1RST
NsMFTQLXuB9Tq67ySOs9ILhEY5KaXnlIuzte56KFmWmO99unu5I49blTgc0FsG8J
y4b019wsjYzqu9jRXnmawF/uClRtXzYwcM4t+ADQqNxSQLtPXGk+98nZTU9KTaor
SMh3qQc84uZAqIiRi/79Bc9adqqJZ074ZpaZP2+FkR7QAPhQGQ4KGsNx8bnNYc/b
xw+t45lvWO0BvQpVTgJ2GuosHD+VTndUbzx5fnQdwm2EwjkeqjBujP52VO/lbBRR
rCtIYGrOWoBUO4vGXjJm6z0ts9ZFrwKDZJIFQ+3IEU0ovR7BJZWekyoCTut+rUaA
7oFWubN81btymVPe5p3TvMFv390txcoe6XbBDdDoo0gmbTaomHn80VLsw9qSL7Q0
X8v6KtQLvB+z9rM1+iCUZyrJJ+tKzTO4IP2U0i6wcg8PyYdWlFmpkcItXunmsNE2
23Fo6Eh1oPXLs6Xpt/hu1CFvlprh6sQz6nqaEJK2uoULa/BSIY/2xbjMt2IEJjOP
iQcDqNkzFy8myDbGjEjRCvhnYQncdb5OpJtvhHwvGeBbWReoU5oCkaUhM2b/CRF/
8JohIW/4+mOp71IIXgNVIL8DNxIQ0pvylUCudhEs8bp6g0YPiejf/lnX7MoAV+VC
5kDlqJ5k6d4NVDx+oeZzISRwlQNxYbAqNTIyWEf9wi9C44ZWgbB2c4/+2eyySICi
2bG51TWcmUWo0TO/yrHZWojm/d+YawakhcHeqnD8LARGIyqgaO3MstkL0OxXii+m
c8UyKuTXfsVhRgB0vSGtseoUJ2Q8KHdY2Ntjd815QE1PUNsAqHkMMpe/kd/+c5Jw
0JzbHE6/bTc2udA45SQxQRae7uwpxIOzGkLwPYLIwKFfAV1Rs2VtXboyoDDjOanZ
S7zgqcny1n+LfawaGh/3i8uzog158Z0Rw1DpKZTmIZCQboSLS2jCz7RUZQAfee4X
vDTmx9BaFsVFKofpBcoZCv1ZxMvNZ0es/X/S6yXVghLL62Dc0+0lRfRX9v9YkjOl
/9nMKv30x2tTh05vdfFnfEVJ7bw9dEc72RsGfzeb+RG37hr7ND0lOHByptn91sct
3A3woXUIXvlOUUxxt+kAHUngX2rbQNO1pIie2jn+Glffek1n6+by9xkyEeoJgiUd
PDBmh8d6N3b7aTryjFcsgz6r1aBYHZ+TAMzUCWXk3yRg/bB4NQ8n+sL99HUL6V7o
pi5s0Gol1qzNfIJrOmp1yd0h6C0taG3RHpyb6kxU1xzYHVBd7snz1g+TERheGVSI
XMmRqptAxVj29nxaJIcB4edwI9QSLUiPpcD7Gob27AR3675CVLaduvhysHIobFbB
3w1qNHm9nAtQ9eY2w6j5iVLoqLN0XVIln2i0wqK+T0wBvuKiRmqhHAZYxs4Uo/OD
Usa1ypLC2Sh7yOrsic9yzYSo3rBs+v1srooAMcTGLskPFwDzhnTu+fIh0y0TMOui
`protect end_protected