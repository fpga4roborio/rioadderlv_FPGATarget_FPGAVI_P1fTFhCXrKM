`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
ddtXksX2+yylW5zu6QL2Lhnb2d1sD00763mmSITNX595NcHTEkwn0zB1Dry37fOW
FufOhVzEJp80NC5qZ/+F0Vk7Ik02dIR0elf3clrjeJRK85K4e3Hoo4xn7YbFUIms
l/8VZSb14+JVGURjfswrIyCUotIzlzVYZ6gzoZwDXIi5gQIBf/gI+KxNXPaKV+PQ
Ufys/12rjO6aI/pPlqSm0hCvftmBcnezN2hk1UeXgOIuKZnogjOsf0iJVX2aOOWE
6pD/psybjbnsNB6kH5uFTA5frkzIzkzl5d9+YDm9OyC+k84E83I/7/j+rk4L2dah
QJOvksSIzN867/4Qt8qYTQ==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="MvBXkzurAa5VTw+1JJ70nePUfoQXBvZOku/SMmg4TwQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
oRtzZL4VJ4iwysPsC8SXYCzXS8Fw2gtZTOskLcDV+1B9Nzn1zTyNtlo6lNICRmmK
ZRVu2BmCc2G+fmzynYlNTnSa7C0Cuel6FYpxCBlOuk3OF2tzAmLAuDyOH3Z1Yjzk
a0aHuoCdIRKv7BrZCdALt03JeUmXKPdOmIlkVGFl8yw=
`protect rights_digest_method = "sha256"
`protect end_toolblock="Jn9CQpRhJt4rnzZPRk+dOpzAubz7omckX1MrFd4p81o="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 21216 )
`protect data_block
gD6l00tciPUa6pDNTk/+t0OO0nC/UTtBwLB41d4inuAUA3i/ALrNyoJVcBnAmEQW
ptbcNp5fxEUJjnOxnedyZEuEBxWRieZFQnkRdF269oOF+Lta4I45UMMx7dZRCAtm
QRnwA+2biV/0mGF2lyI3v4miO9GvEY29D+z8nbCplGFtfpNqx4+ye4kKJ+syucAG
of5Tg4ET3DD5AcSGzXiRp2dZdku4Rw1WQY+n2nkQW4hp1L2pttwQAF0diz6ZYMhD
ltGg3t/nb6GVOEUU9bjPgPANlBIGHL2VIRJcsAZVlOrlFYRQsgrP5RDgeXUEdXvu
D+LYZicd12hgeu7UqucS7BvZDYjcFpU5t1KqiKTpfrVe4CxbqO6TIFVBIGkTcbJU
y27UbdiX25UB6sw6IR0s8ytGS1t1OPxu1VYIv+ktPJlImmxcZx14wzjzJ9lSM7VD
djDqFaAmyVxE/Eoynj6CKPRoLJFC9EQYnN0fQQDGYI9WFSvFPDxIjNSOKRS0rBv9
fi7HRb1YIOdCRFEgYKjXunGBJA7KD8sculmm46QqvDiUzrW2lBofiLoqBdGLlIRi
7J+p/7ixqMgd411a7jPjWmKGW5rBA5FP5dGcKVja+t53TFjH9a8FwXM3RLhORRgX
nJPmcCY4M+ROrqsNiYQ3c15gggtA1RL3kXPwsnnb35RI9T1Y9YUeLvlyOG7wkz0A
EpyiTuR5rK2I9pad1Ncxn70/KpjPj1jwnqo2RaQ6OXvoNORRySzor9LPWnP+ujPk
aKrIb4mG3uS3a3M1DQplTX37A6QG0mrN3BtrOQpLlmmbCnkOBqr8kplfO+XGgZ4n
XJ9r1+1uaH4+/adXr4KUpRjdhvl1bZ4TuqDDDtn5VGDAifpSTFflesxldXlVi4Lf
x/jAmrGJhZPAYcHu8jslj5Q3f1tbI5kWQEDsJ1hyyhidhX3DZIh4D3zXi3yUd9kJ
xSzV3M+f2SaPGVoD/6ioaasavrz13fT9wxYyQhzs6cZ7KZreN0mDNhVK9PPS2U/4
CA5dnePO0okO48ptw3+FFU8haM+jxnHbPKX9XYUt7plOq9v4wi25DVkBUJ/t3d4a
ORQ/KO5GxR7UifCRLfeGS2OsiDXWnyEo51IDO4fVI4Uu7pVxnXMfjBb9BOIXjEls
wTUGPwmjFFNxs3fwmtCeclAVWA0k9GEF7zax6DXqM1Ark4jDjAnrbdSU936d28Qj
0bju6C+0HALF1ZZgPIIaxCdX+b+gz0ZIVAHUBExm9H1M6LVP5OnqvvvZZKICeWrL
nAAYJul3j1DY+mANk+Yka9Pa33xPMoExPyj1D5IJKl3fG6T98rep2+q/Ayc/Qdh9
63E3/9oreMl9x1voTvrLxG0wg5P6xLnADeeBQa/2sMPBKGUpaj8sN6KJHY/dYi5b
vete3JpVQfbi3vCCzSmdzqpb0liH1uMsecEXxXvyg3eNTbvBeP6wBHK/WE1hgreJ
OqzXaXa7bU59MEL3CSBdqaDClDgy8cllGUcaOHXNCvmiS4MLJ4HDnBml22bLgI4k
H3BC9Yb6FLb8fJCNdh1TpaHOwAtj9+hXQD+rYfP3mX9CbVimNBvKCyLum8i3/k3f
QDSEzw5jW9YJcJ8MWdnQu+jrMsRtI9K2KhyEZdgcv4IRlV7AGzoEBIokt7wbqX7E
RdO/1fBoOrruZhGvKUGUJJnAjtFwObixSiTwVeSuNhd5iNspysYIgIkwAVc+sW26
hD7dElS6cYNEzSlLGkqIrOh1gyuJ2bAgqpRPxLXkUeM2e7k8y2I70s7djahLSOcr
IB3McLn10teUFbCD2DzLlaCDimlO1ms7StN9HO6YwpHNfekEjpnTC/0EJA0/b3x4
qDwXO3n/GlQru62FnNlAPzomyh65bvEz6xhuDF2LcxyvUdLW26RzM+e1FLQkFBHU
UL5F/c9cDLwZxpT7fXe1Cw7RVYeh4OizyWMume54golAdCYX5TcYz327h22w5gUb
lJ3BtcdbChQLau2YEcWt9ufhJESN1pvPFuWMm3gu+rI4px8awoeJZDvqIRndAO0M
s+SF1yRdrPw60OFpS5ws5lIjYN/XAReDThrKG/Zx0vXvBhhybrcLc/LNTLM+jUE0
EoxNRKEWrWpninvfniCCDL0OP8prIaxWR4JjeekHufCUvnAx61bSI8MB0h+8N/ls
04gga9LMFVa0IiTTSmPn2mnij4irpiLiNJIkLjQ77VDsQmd1SWSIcyRHFUTUfPtn
8ELCVq9E9kfIll5MXS13S3OX1UADqZpCcU7dMhK9yr9jf+BU+OtMu/o+KYnWr5b8
BlopMT+1FUfKqVAOJkXoTEhyID1Ek+oxNav/JFO81+T0JnGGdHegaKNc+g+K4NLD
L5HC+1/7qhi61g9O3nm/PbUGYAQsihidjyMeDRBpAKGyeb+OQB+AN+qEV0wwe00Q
+qpY0Z1JPutxN+anRRJHKrSzJlcJq9tNnxoAq7p8z/3CpFuaJ7KPtxPjGfBJEh9Z
Pjwatu8O0VZvycTFDbE+Me5isiOgLUBP8JCiEnZRTIhw66E2wKpyQLDP7Deldgdb
Wp02s99U0eqv6Zyb7vqdCU0Ha77TGcIpYWNzUffm0LiYamTZgD5JWRSR+ZBgxt1v
gNjmA54QGqnlnZA2OEbUY0GptQZAxsQG0vDJAJrCTqnc84kbs4VE50c688owgQON
c4xkGvHJxro/HxQOE6sQ0vB/CFjrBQFJZO3VRF1u2PVcZHnp36UQHG85c84gcxWT
tJ4nVHA9AbJtHMo6K5mjVn3HaXADfRGgSEKT0z26OCdcPvaROkZ4asyKn87WgRAv
NvyloeoVDagZpskBiLIP/MrNT/fnKzUImyAsBYgA8eQIrGrGfyTqWDw2T5BmkEUf
kvOHq0mX+4hDTcrG1yuvtnF5Lmf7kb2f4ni+xa2niTZ1KaPudJilfSZQ9S6eWtNU
e5w2JSaawu4AYi1cy8ifvBj24E7JSQ2z9gZki+HVoVDShCZtCTkYzxdkBYifQLcX
kLvbaZnfF+eRQBJ4qPwtNjUOVMbfzANd3TpqGDr1G4qXnGrjRts4+BElarC7etym
2b9O4/k+sxOPwci+r53cy/chFQhHqh5r0gRGy5ecXGjFRgDIJ6RpoKX/kcoF6txt
Rdri47xrl73w6bYIGPLlwnM4p13hXsWk6HrCvwT3y174u7jDD6MmyN3NV62lAvVh
M3WDeRgmX6kCh+Am8qMY8hHXNck2KRS0aBu9TevQLhlGEvg6NpsHQfldgcsMQhqL
sSNowkhALC1eBrrfwtHLQgDGRolrMv0dyRkkl9hUdP6ejmbXDlF4K+YYVrmA5mZA
40KGNuT+bInOdhzbeCek1dOIpKJ5dfja6g6rUU6jAsjmPFHXEgz/EQP7sxCljoiX
VGocUSHRyulWYduvbN4dPe1IRrKSZkCLHvIgfFQzgOux+wcyDXt8Ua7ec0BSEPHg
1YqqdgQX7Wp4bmz/wk7l7abU00EwQTEp7+aF5L+t2i/23yjBUAIx2zE0WX6fW4E+
E8i7/y90N+FrLCP+tWkUOfJFZ96eego/sHksRVR5OIgC8CTvfisSAlr51iGgYqf6
90DGqfxOFF/Vckpegs4xuAv8ewCjk1MqI+mGt6Drt7LWsANOtPQPCk6a77gLIIFA
SRH16nlQPNaX5/Hjl6aR+PRrKKM4foK/DrNijgwuUKPUJx2X6izKxDA8K7xKOnz2
iaKaaryo5ErH3uSsZqgYUapBmUk8/fiZqCzRTU1qSGrBgM+7uGafUeCGjxuSGCqe
AZ3kzPYkFRTKxNojEGgyq9hezUuUMECprxNDB4S/WlWRjoFQFzx5V4dKTLTf+DyU
f2e8M9rT4rKEpH5pWrMU1b6YLf+e0OQdH9ZFSJw6HRbsGbSqs85Z1GcJWI/Vwzgz
Jh1EqH3KHi80d1LmbgqFgGmyegW98iJTvMo1sTsKqgwZ2/Tl7BlFguXYOWiFWzeg
fscPJgO3B22NZx0U0DRY/5NCYBHkqKRqHI4VKeROehWQrCwGNMal6T9L8G363xd2
wT5DF2p8wWId+xdTvIHrOfPt/JDIIhdNG0/+WAjvgDEhU8botMJcplX9Ob7qqVkx
2RVmxrFWPrHaT1fCUMPu00iICm5RxtY1dopGCoFFvqXDeb3PdRzamhS4jxHJEqpv
redYK3d3nDa6bRbcnJFh0EyW1I+dKTXTm5l15QSEcFuX+VcAFfWi0H5RiOt4QmFH
fxkmAtnLhQidZRmtIjaMAw86QfhEPFn1irsXG54HTrAjEVpQBpjW83Cs9Hsufca1
6kcTEnkHCJpEDcLSaeDqmNttDpxLSmAAT95wJmzshDBJ+ocgfAvY0Oy/YP7uh1rt
kl/QjGeryUKuETAe85/V9kuMaBABP97MBNkUVXTqrLz6b45qLwhVmL2iw6W6yNUg
07Hz2YYvftw42QeMaUtqLKhHoC2yw6YqDhTvMiNi6KHkBzdDOmYcDgYavhWV3O+P
E1PZD1RSxY/KouknaG89J8KWBS5NKpPHFXeWuttJUaqh/jkUibLu0vyrlMvyf0CN
Mh01SPfcGUTepII4G76W3hAlFWfEjAwpX/v4xW9qA2MRuHwuNSxHLVnekkfgllzw
yXX4X59wbOR7FWisbANloqmVCKQ7hAcLq5TN3kZhlupRMvIOYfed1C0p75nIKyEE
UfZNgfnZtdcY+uvVN4WAAE0Lq148hAsHI3kJfZmAj5thKgvrfcJkYmNt+hCRAl34
CEFiv/cEG9G/oVmfd1svZEc9I7XMbGeCCzt+BIC6M3w4ylB5awqIPawsmXJxGABe
2GUOgrXlRggJaAvpaO+vkRLtf7ZCB/4PZHHJpw3NhumxvYxg2QstHQQ8TMfVrfkb
YxPVs/K98ro/8brTTWmHBOXP0X4qlM7nDSAaYztlivW7Szt6HPFzoNDhpiEBPBsx
1GOln3dGvIw1Xy3FyXpUVo5IU0mN//rFncG9ZFb14wcJrvLDk63/EfIU1+fi0pUl
RvI5iXi5hOUs3LRW8UmPDBukWpq7+UOflISYZPYjT73BxeOfgjg3I0d5PxVW8w0T
KCFTrqfCHlVeazx9Y1FGeSsaZCO2XzXpPsAfG6b0TBFGrikwuW8VDrb/mOqS1lZr
z3axQKJ35YHOVxGaUj/Z02/cNUMR1Ph2QOLOgSIAc8YhgyC274YvSACaS2vetVLi
0N680rgvmysIFUmyxsHJXRZUmMaKBPbOkB7D25nSHOqR/GUZb63SQBYjGmIH/HXp
0QkHp0a+Nc2QaJRZ5GXOll6mHe38SwfmxEnSW7mxJ9V/NaIDFvg9vmBlemjGzx8a
qxmKrhFd+9QouIeetKRBAopW5krOUjsTcrOMNXFRK7AMBKOewBBoMj4TCF8qi/rU
W6tscCsD0ThZelJanlMgAnbS0IOz72oW6LzTIgCXurNoHh3MWN5xZUX+b15vVRBQ
wvBaBhkMIPpj9yNKdhvCFLJtIkksgrEmM9PTgwg/Qixpg3CR3jB7al2qmCjVFigc
9mjSWVkW8NBZL1iDFQ8FZu3A8BoglvzkVeJRBS/BOA0R7OS9ASJPJb1dhEVTE6Hx
CXQoV3NvPHMsVE4YwB4vYF3MkDoyjtoSLXRXmSyUgUsipvF6wWVYv1iAl+qvT8FN
Dx95Ss+v7EW47SwIyQW/doqsLCGOvaL1Nnyts6W/dJpWYqTBmCPxg7hQnwq7Pl4d
R3hv409s8Dgk2ptB9n1V52PbnQRqr+9MlKyBmVPUbP45Drevzgwx+e7sbQY2umMi
I/KoKdcMdUS/NguF+v9/gdeYL+xrtvIY7afJQuEQEei1YHTyH6ORChxbyh9zfLPB
bAiMNTbpoDAwXNoG4d4It/TVFm4/xNmwcOaI9A717nbxcouto1IskQwUvn7cdw0n
8aHMsWNYMWIUBumY1oYcfbu3a4at64kl3ADkkPRrecmP0GIFoMJaJp77rQsuZ9+N
iJmFaY4W+uvIFLnpvVgx1jx9Fe1TEcxU7GiCCZKp4USIASsbfHbITL3jO+o0Zjd4
nPFWazisuS5Q6QTvSBMlWBYnhNYfjkW71tl5z4hqxILPw+XCobng/+6meMwq7vnl
uL4zh0hH9dI3l7ohTUHodM0y84mXo7sgvq2xszpLobO+QCIsnL6eGaOdxBtOUl3Q
fpNJSU8IQ/o2vMg8vgNHDM90SQ8ZeoeOZ/i1Ca4+cQRG8ohY3KUAHSIJ397wBdBx
DBknEBxyHa1c5v9VRbvwltlNJWu59GUVD/H25yesStrD2wJbJxk9UpkdiXHY6lgW
AEw2RMuKMzQpeMOy6kO9aIz+dYiFoNLSwNM1XraxDNsp8dm9TJdWRhuMMPpb/phL
AMR19BepcSURIwIVKutjJ8rnIcpFpq8koHO73HferDsxymdztYgqA9dvEDZ72gzC
BOm4lJHMPOFiqCOvDJyMRRYWJnW9ASuaRBtjMZG8rkV0y8sz0u1gSsVs7bzeJzyk
fBo/mHs6Hl0tYxy+tXm0TCcg4wNr0ZVkuVrKdsiprWF63kF2rr03d+RKM/gGJQwf
i9EJyWwjmm7ofeDjVOhJRbxBzdkeYmwpS8APy1c3kquuMrEh5n1k7kpPx749f8N5
nG7hX8s1SlM7dAyLKebS75xO9Sat0mMCFlXppDo/bfM4qqSQrB5gviWws9uzQEAN
wTpsOLg0KLikt/z2wN3Kw6iWOpc/7ullfxRhYgcYj5Njb8uBWt+vl/Umiygpj6HB
/C2XGliruVXhIgsnmD1N6PipDh1EzmIUTxYhB/cntBnqKCFH12YgIw2ERbODTD4U
C9Ou5rsP3flBhZhm2oeSREV5c4IO3UcxKOtjahLnlA8PH1+TJyt8Re+/JcYSk0WS
CSQJm2ouKu2gW5sMkniIO/fieuDPHTEUXQFC7/dzI76KHGZXMPz7bDiY7cVk6BJT
Q1T35+WHO5tzOU6KX+f/L2fT5vhXNdmTEPLeyOxNv4yxw9EacOews7eiyyaqFPcq
/Rt2M1f5U/sXuEP2AYICvLdYbazmgXNpSXxntM9jLAKekQBbAubXpyGuroIOmJuC
wfuF8vTlpquHm20nEXwQJbJUruLmqayBR6BtP8ewJCgB5m8i8voGwv1UGzGYJ9pa
782ba/jLO5IZO6irjfEGVlHTywKLP0GVbsOPVwBaCXyKpJbSjnW/qYH7tpV513wJ
A0dWhd06BkGW9ucBxjyBMyKziPlblxKM2M1Q/Vfl55spmT7NjCuXEy1aj+SiTn6A
opv+dtK0KJZolBh9kny1cnt9xHRSy5QkX+y2ux0mrjWQuMqRxfsTpRDAxAt8YxD+
5Ml0Hf52kwrcGwB3ZAA/6Q/uoSWc+EaIDClnLJta0036ECwJC7n6wjNuxvgN9QFF
CQWJ31m4Glrt6+QG0f/IWIRJfQPZPZFheHkJ42xw/ByKyMfLJh0kZ77ZcoR3z4lk
IPaZTDUtPHjxQit9CBnosh6xLzcFaRDqJsGBjRGy0YYU+4dEY7IyCFn5NKgEzAvo
fO3A3W+13xLiT16ibv07o6RPLPWqSyvt+8yEnbP2z7YTcRMiRkq6+Ak17j0nPIBY
eYKCDPCmR8I/3PRfr/UpyoooCuBNAswWYe7mXzjyodw75ki93vPU3E2ax10ghUxy
S7DVK0phsGqq5A8cDMhAmyysfqLvSemPTUp7dlha8Bt/YuP2DW57zGeyvh6va/L5
NNd9nN+w4/4cxiDUc8nQAJdMkdxn1EXAi8XzU48C0K+zzdWnf8yYegi+NQ9siVuo
awA1ATlnYwmb8s3FpRT58wykuVhRSvts3GGim6RYoWq5ph1ArlKo8Q0VHL+0Iif4
nDbrAY/tcdmIjPnpwlSy+a9o7RjbFLgAeUvFfMAzkAG9j+bVQNxLF2xHGjuZC1+8
iiOMftU3MTtWDt+L2g2o+nVWch8G6Is71ubMfbvxF0WgxsU9nMfEUPtBus9Bugy0
XUPMpd5xMP30ynmJue0WQjLPnaFw8QKJuoxcKbbRZ+InG++YC6AxWtzStDjWwmiT
uZpuhe1YvhNfIpzcgXLbX359iTG0mhsgMiNL30mn7vYyw4x2tqNmoibaFNptqOA9
fz9bHBdzDGlQe93cysn2KBGQPKw3v5Uy96apSxVPxeCDgFI8zcWMAvtJkTY7ocNY
pAaEBM5yMEwIogs6b6befQVhY58BmGBesbLJ9cbx6p5K0hRgW1rlNEKUeUXI3PI7
o1Gj0Fl2CSXidZEY2lpNSL7lCJuIMYmjdDOrKd68Qk8mKmhudqtbgN1kU7eJSEAI
+RPm8ww8hiB1NsWk9mSP0xCGzubQqyyWH24Ixc83XHAqsIm/0Brs7h8VpjbIhamY
2pIlrMoUt3T5ges+j+LIcyDmVfwXJl+cKBQSGEa35mlO3UO+/tK+Djmbr1KD3Poj
fk9q8w5XywXsziqZtjzpP77L+vRv8qxXQNsxdN5UgvMykT+4ie9hEeCYJOiJyab0
ClPI0WtAN4eGm3ihTA3+fNxSPVtoGUksUdehmXTWTuP063ATLXZEafDyCjgryd8w
fBjU/Hqjg/xummllGrw59XCTjdL+FzxFbg8hc+eYNgHbUhcDLK+whnu4G4q0tWF1
nCXXVd+6Y0BJ4AWEQW6F+9xMUI/DFXW2dA0PIVINeUdJ8RouVPKP1CENZdVJBfnV
zsKUkqFgb0USUtAbf//TDGbiCmhiE7BDsnBQnIs9ltbFJAzjsSqzAmgl0huQ53l9
6DqC7KpueA+3cXpjL+mcAk7sQDmFYJV8BOWOCmmZ188jxnAK27f5kTl/t0cJaqUh
oKcgWpobzZh+xFu8J5b1SMPX6SGokc09Kl745DrpeRFvgH2P7z1q4E25jcRqedTa
PaR8tTrqk4jdA/Q1WUFnDZnXjHPd5VUJXMh88dxRoFTKBbJ0BPoftHqACrJ5PJbd
NmlVekkWYJBUvMPEcRMpGbP8fBL4w1G6yAiROClUBaUF0blnI5Yce2Ddw9g7S1gD
yzmxfgugQijqx68hy3IsTX8g5dOiJaEH2MnNhtyKYAp8cw2+DIITvVjO0AOsRg5I
n3J+a1mmi33vdVN+j+nUuG0RSlhv2KEEj8u9O4ebUd1FOVv4tIqz7zkLyrYaECil
vbCsPNQYs4zON2Ippu1SUNGb44VtdE/tpMUYEW7ZwUsPInVzQ/tV+rgQPixGFKaH
bj7LiwXPH7WrzrZ8jyvOfJPIPPzIUe4j9B27j+xXJmsGFamijrBOOPoLNhbTiRgz
R7HGs4GY80GvcL+XnestGEw/kY+2NmNV9XtcQytTdLrPt7mQRnEmCDdbuW4x4DqN
jdpttS4hjiw5v0bE7mHuuvV34Dfn0t8iWHGc4yBR1KCios6p6QVUZR8hC0yntmJj
Q6XfwDeblBYilzcoEhFDq+8aZ6b5gGcvWqvWEQWFPrn9mIjU7QoTsyMet0Fif9Pk
cwxwj7CBICv/OvpgEqYShFn/iow37PtjBkMgWd8wD368rLQpTNlTjHv3qmpviDJs
H3YEkQea4oWYj2J8UJpfsqQy47exazhyofiLTB9EaAEEkxtAnIaZGh0ZrWzu/y75
QfJ8i/vShoLogYRLm0hmtTfz2k36Kel+98nsdYKG171wW0hOHLI67QymhwKV+tYn
gXYwH2EHqsapKM0exfJVoPbqzQUB4fERyLHkURQ+SKQvvqOasX5zXCF+JjT3rlKh
tliNuJt3RBRn186cMNX9Zp028BBXkwEGz4wucwuTph3XFOe+RvjFH34coiZDAKVr
VMf18G3gD2sZTdwmI4M7R6nKng/ECbJqqGggyrLMLkpj+O8nkRxcML2/HSoplZHM
d6fRy3ZU4M1U7qTEZFZXUmT59BJDhXj+Zog3RBfFDFkA4WxvjVEcvDddagTItUiX
6gEI1gVH9+3JuY7xQCTPv6qKO5ybIuvKmj/yRRKuXr3/JnVdAyzcORJIq03lB0WN
eTjKSji8ZXNn6MzVdnr5kXoDlREMeK8YyMmS5j/4wP9jcM7mwKe/0CZAtAT1uqAx
pnLtSCuqUUKKtBrke5t7sOxRddAcloJJRTYaldu8pW0MbdIbo01TwUidyLay/9MF
ADaYRofwgrNZAg0FfFLg8VgeFGmTSrf5B0D8JuFt8+DbTzyEoJS/1OM/T9qJAQsq
oYVJ9tvAvtZ21csqrkQvnjZ8OhVJvmOJDSb/Bz+4WN3LkRQfcOwBp5aGgo5oCDSR
GOLA3Zot4auH2DiQE2UNx6/rSp4Mqd9UzzxNtL0SdEinB5iN9uQgoJO/htj7xHct
2VKIiWQxQdfSEKjq3eI0YxO6FA0dhsxes423RYPqOanTfndwLuqK/M9Tfmrk5JM2
nebkyqPDkIs6vEs1CddMYhYtu3MuZuLsDGxYKvhs+lBDnsi65aDkLLuKpBAJHRXI
Ov7vZ2vFNmknYeDssLODhC0MX8UXOH8wUKnpHca8+JKJvtCKj4KUjtJHSHJG7Clm
b7cSCG8ehDhL0roYsMJDpt+tAc2+gdE/UoTTMTuSbyPhZjWHcIaQKjELF5urgBZF
BCRfXDHUEuAiF21ZVH4WrQwBjb+ycsSZq9MdfSGDzQdxqomxPu5sEcjjMpceShVV
Ratq/QgqHYd5AwwMRB0V4N2YygqJavjy01jZ5MduSy+0Ov+JppzbvGktqPxs7GIx
LaP/IDT06er6t5IboPq5me4iME1u+4PImLaeZpRoEpO45r4rcOGFptxHo0JiSwLx
nAam0GpEREfgGzwHaQGDe//UbkLKnhCLXQbsu9Gv3gERO7oAmuFUYGm3oKXu0jXZ
udK3fTQQ20vdCtNQHe34RaI22udqBkxRQGjeudEIu5zyizJKXx7coG4MVcMkaQ4b
ryGcNKsSiqhcrC6IDA2yZOoYQuIs+JruXRXczNT00R708NTdJ0KhHmSbRbvMrqlQ
DrHJ8WPmMDmNEKnhfkdY43VK3We5hI6EXFrhfGgzpGf3DMwApnMCt3a6Wcc/0vGH
WdePA0M5UXIY5tWQq0ZgJ50Vsyt9qhIVAxDvm8mcV4KwO7TYWoUH0OxuAYtdPw1k
+uPhTKYeu7Doab8heHXGHHDwvpfi0TCfg1EpZ8q5BRT94zvi9TZa5YwMLr/Zsrq1
fEKrT2mtVmHF1hT0+Mg7y2mjPCp3I4198mdDjes2sYkBawIydqxVWZvK+H2QQdNz
dM9sf00p8kFnopdMz1De8qb2+u12qgvw5gd9Rn/eY5icjTxJ0bdf6Qb1ckn78M5p
mxcWDvT49R8YxUgj7vHIHYcna28HBA4Txpy7tQPG6g+k6vJVBgCV33ROmALdbZfA
chQjONcVibgT5Qk3H9GqeinUVz/xn1Q2FvqxtC9TyYsPVbcj4atY7ZVABRsp0LEP
xSakrelP5YvOS9a2B9RinXEHMoy5PY6YXKO6ZdA4OSJuN9xY1Bu8OsMaW/Ob8yBL
tYDOIZXbMrVz99xR1U5nga3KUYS1HE2zyiqafcluw4GpHZeDkmApxCqLCv1HU+vV
fp6hHgnrhwisTK9aJTgL6D6+phn9Ke+GGmvArwHZI5eS5d/acGwNKHcilEMC44AQ
7j2BIbN57M4aBzAhWqh87WvA32fk+Acm0T9csYCQ3Wl8o7AwbhYkXpvVmXirBtkp
XpxeHTTZiM4kizKJDgP7t/rcvPwstu8oExDmoJlXH2pbvPIzQucY8ZKLVgRtFiHA
N3CbDn7JKbltQ1OX5XIok/3IEZzomDVFwtBlPq8m6UDlXWGagtMDwi/faaoy5LJz
Amaf1MHgpB0rQnKgNXn7cyFZi2DrVTeVZSOjamD2otvvFd+7YCcLdL3+TBr7CFY+
tWqokUOo2Wk41SWNI4yLvIAhDWkOFs9/Dn7p3j7jJHcWYZzskU3M1VuIIuztl1Jv
sdkujkRWUCj6KICLVzpJPlCxtN+sQJKO07RoTZCqg99OGZ5mjzxXuNzxQDmWtJ10
HMm1taGpxBCCYNDDw1LEyAFw8ybo66+BmN9EE2Q5wvNY45rZmpFxkz83IqRtRPdE
I487lvYDgOHhwWyVbQlTvSLBS84wY06sNVlybRghA7+jmdHNsXVsaYlzd/F73cM6
lyDUTos3cEkldyvqLpX14p9dnytCUekPlMz1iSGMw+gx6Vtqh59YLGXkUIX1XAdN
zZgfvsEI0KLeqGxW+qzkeibu7EwoPkv99RemOe86EGAU6DCqqjlTPM/j7Bjm6QtC
GOXAVqHeK33TlfHbpYlN/Hi7KHtoUXY9UoFP+FZMjP1eYSrBinroRT8weWEfKGiJ
pXctESOrAGZ5Y4nKRPypQt3zWbw2RxDdZu5l6QbAvqxZ13cWuTlRCjT8m/89yo4K
LZANS7p3Jdy2fErZ8kXO2DXTYf4NbKaOKlZSGbxTRYB4NlB7j0JEAEdy+tJ1fQ4h
YxMPj6FTF6+9o32xWmej6K2RDvLVaU07CAYkP8nDxWuwf/2n6UgKDDZ9ooMDUmp4
cnLNWsbt3gmGxlyyT7JCXa6t+bkhvclCS9sDpjhTeFOkAK03JB4AVVdxgmoh7PJS
e94e1MM4J8EiHMcOvPMUqgdzxRfJd2QuRW4W/8XLzA9m8/dM7QxUU9Hn++WZkXxQ
fmBrEU7DXsDa9kGl52J3CE9Iq7eW/wGsOUKsgWQuiPEAkgUfFfAsO/cxTJd3BHMQ
Lms590GZCCWJWurOtcggdxvzea/inWFzme1gVWU4kwVLGOjc19/4jTnkEeerh8hA
GKbMNe7SlJZ80ahaiD6+tGLm/rRyRBjAjBtIP65Mz26HLF4l8tdc0pNELVSd9QYj
/BICVZ1aQPUJzCgzW36/vUrnWGUpEuitFQ06hFB0Nxcx46tunqJ+h9WKwFcvqmdm
xnjZMh5N6O6hkfr8vyfERqF2Cf76y1W1kLwJuCDiwh+RFWmadtbxmeNOEO/JO2Ig
TWK1sQXblFrSpJ6ZrYcZRi4DipYxCRSJKd+PFavnlvvoAqxerxHRE0OfDRy7si8s
sY8zkMZORgsOXjWVJZBdxF5FmRRrPNoP4Ffh35j3hR0wNBe4thCvtiAujpnJjRZr
q//bl03d5pBnvcRpwbm1ExKVf8/aQX04hKxgXNX3evmb096Rl7BCy1wwhjVz9IVy
ipSPb8mbqGoMgOoQ+o44rWPzqmjOpybCvx19+1/zK5XEeLx5lOe5qnUurlNgI5cR
BmkXsEjN2OLUNyrpuIrC757UHFVKFB7tzM8cxRit3hqVVVl1obonmsiwnUSX7KBw
njmR7FdzX9Xf9TtFBjU3Epu3h7g/S5gUTboDntdhoye+sPI2iD+MT5mCuDSosuyc
HZ3dvF9IzNqWevFGJ7jec72sF9JhG3PNZkpOvLTt+VaxMCHpQt63elNguagUgBnw
cXNXKLBnaJVbpUWIlXSyEUMSKRz9gzdBDDeT1uFKKypWUgIwsu5udFTVBkNnNPT7
Np/LtTwQAeKscov1mfTwskpkoefCLbAVZOO3l5c73hlysLBfQ9fFaH/+d4MWMZ5/
/2DRP1eXK3HjTnLNsqFdNJDLVbQinmMglyVt0OyXEI3JRzgQZe9lAfpbcehXOALP
MmMk9FOQ8k4BweiIjDHHspNN89oxRmTiJRWlLi09dFU6AGsQvUrd5lVxz+8+46tc
WGwRV/G3O6iLGZWmca56m73P1s/Y3vIMf34qIF89/HGj3DJmX//2jqjY66N985oJ
qybdwcoy0aP0VqBUWzQcqi49EIW/IWko4tXh+C8cRUaHosDQRmOtcGRjNVi4AG7b
EbSQF/Wj+xJ6OJCnYhx2hbcifyBGsdYGHOSv78IiW4mz3VibJilg6nRtFAre9UMh
mIZZXU0g5DO5ZLOJ0y4TwSR3leNDaKN2yFmr+rWLRPN+R61Ht+PR8MQSzdGBm4+k
kAp20g3b4uJ9GJZtwC6ys7B1HoGYGiTUi2hlnTm/KwNexmvrKEdO3QsTuY5VwMxj
yjaTc/yJGDGTNQJ1/YWR3fBD/tbfvh9dkhjyv9ADhuKN9kp4ageUNMRFkXkn4brU
22yG79EB7I5YEjCFfDzcqzd7Ufh8/dGS6b6OyEGNQaUz66m3CEq1YWHyc4wQAq76
thrY3nZaNYVFRqM+GQaLh915apBJIlQdrDDi2h82TyIHmfzaagNAL9L8jjSCUWGu
efB0zR9eUtVLcNLC+6J9SfbQIPGs3oRwsUTid+mspHFMhwT7lCCepvycaLfe60Wl
7FhZMKB/6UjYQj699aGE3eRFGBPp64nAxSQexUVGnbWfblRqrHrQbQy/2BqyHV8w
ZFYYUAzp4vMcstp5N8XqUOfp8zHNFceLk0iQS28Bzf7UUZgMIPyLY/djIhQn9utF
mNHuxUUC9wt0cq9SNOMQZy/WUQWAQkyWdo82O8e9iE94HiY0lLSb53+MWMZyaKJI
BEVbLd2hCBCcziyIObG31RltbVN/18QUy7fd5wSMtT787ov7hqMaJkDuYjEudceB
gjiCe4uirZQf/lv8nf8n27Y66+hutUNnitkOt0x1Ce51cRKHMEjB6J+gQeW26cQO
Qa+jE/lyHlpP+eZRWlEkmopaBBQYNXKDzcc55sT+85uznxnDG9tYZy4thE+aTCfB
vG5jhLTvw/nokOQRDUxclcdPCJoxKKM303pqLOOmxR62Gj5waLxUchP0e6wDPhVb
NogeWiDHvgwB8hUflypjI1nbPZSghFt6uJlQ+339lm4UP9L1mnMTIjMBl9WPfaFC
b3TvSc2sBDIdO7NEY4g0Wj62qbdHPpTcOH7zZjSdemaIlH/Gzkkgm5A8Rn/Vbli4
6KY3CnZW4/OnxePLvd7nK+SRz2L7yQdj8W+nEsbqopIGprrchldRPouV8kyBD6BB
+MXyEkdaVt5DbvZFvAfP6/wfcvweCXttxCEuWSZ2dPWxcWXSuMmEEGYfsZ9oMRbT
yu8BXwUnq/jIgDWUKrZqQA103ZsRkMCb14yq4+u1K/0jRLW/ZAB+0urjaM2YLaby
B2T2mI/EBuiN75FNM6gu9vv0bcKkw8UYMzyWTOn/p27zaVqCbFHmBJ4AkSaty7MJ
zqNcSKwJ35BOUws5WHw174gZcJCculP9SrKKoSCnSnuB8Y56q64L0LDMSL3lMTij
FV7swop8drKwaH8ihWssHmGYopo+gv8qrz5jSRIDmLU22aRXl/w4ssmiVjv2Ajtx
nMVtWjQwvWO4BhpPdVWClAUH0ullFIVkUEW7vsPWmU1WR8ZSrCoFqyHUlrDj6og4
ApFh+PkLBz0YUwmEhUYZfH8h5R0IhgDrEucxjYCPaAtYQsufbwRTJHrRToOvMYGb
5X47NPxklZn34VDFY/6vR5Rf56omIb/tMbu/vKLcvOgYPxtQXevnaPuB8Z4QUJLX
C1ROqWagdik1/LMF5h4FeE8MioHfVKfvumD/gq0aczqIgnOXLX39eV3Tq16fQJsb
V/415W40zHXcaxJF8sG3ZjkwUWPW3nXYYRSUQlPsRKeDCmhNYQ1qhhxWcBPlRHZ3
h84VK0TqsL6ndArhtWfgrqmrxc3qOUIRa/yNMVifsHUTeaUFtotxHJnISXVsscoO
6iBe5Lpirdr2ZXxHM47xmeQv1883hTzsv3YBYiSht5OfdwQYfqwUVKXqEdf8e0r9
h1YfFD/x/c23rMZyR5/esTg/+ffiGBQ5a+OtVrEmeV3AL09SCMsvM/RaKCgsEOmk
eH8/qqaW7YBeyUgfCbthBo6Dhxai8awQKHQpULy/SzuQqFMiH/8GUITBOvCVDpKL
DgZ3/quoekpA/8M9AwlS+KjITjEFL2RHmn2en+AMnXmq5XHIBTF4b3sy+VHxGqK7
Sn7tbCnNeU5gMqjikrCvZSqPuuwNitauTSz4Kcarh9qOuZKDEDVqP0Fpew7D7+Ia
DugjHElRucj6pfigpy4wSeQ3WR5RdYz/iUTmZSp61lHOMa05UxAzBSJI4GrcNBWe
/RNeHpmMIJ7G1PeTdeEZSoWRv/YLPq+RhJL3G66oHpPVoQcU7mOd7gLgd8YyZhak
ye8RcaosfQmRYzjOU3kVjry4ril+0ADkd0PP1Gz2rALQKeNcD4rGabcogu41Ih73
31Ii8iHeRmONAnmNHgqGLHqnXyDYyEeZJGg8eV2XM4rk533op3Bb6vMkd+m774s7
auXYr5QVMde181hvZ7uaOpH7YOZqINP6QBVS7LZw+eMEnnKbXR667Q4XoeTEVBuW
GsYef9rqIyRzoNUI/FQhbjRYRgJmA50ZfC7ckekru6rOMqewLndwe0XXAmGJg9Il
8OjUGpaNVz/8/4uyWE57bpSuRc1OcNe4vbRhxvPMx2b9YK/HAT202tfimrG9AfNb
/lywZEivc1sRng/2DF7xt7FWZtIeW69jPCHyQbOc/C1cbEMpAQSDNV53De3nK/QG
hBs7PVUN4x9jGH31+qf7qHBKz11EQEfptfijZjKU29xxwXYgfKhGyts0j4nWUbiF
gFyDBU3uVgh8wL6/pSQaspgZWn0NA8ubiM/mQE5YTWtaE0HyFxtF9pdLtnMDm3b2
Kz1LI6Bsx2LS6phXrQu2dBls9pn+TEPMey3hJO+Rmnrpu/iRLDdySLxOjnn0SeEm
k7QLsnqoop2jFJtvCtQmypNaN0oSNn9NWhCrLJqaXvC3CT4yJzsnjOixA18Fz7ax
igjS03hs9cNR1HS/EW/a/Z95+mLh1sKU/2cTW+n/BqTPHoKH21cuV9zd2K0fy4TO
edVhA+RRrunL49fYuNs1ymflvB+MyMxGG/6Hcg4//jEgNSIz3uE79sVovSUCEgqS
vqEtSA/j2rMud9iuIte5VaS7UDC5E8vdnuLz7i+GSYuupHZhDBWiJrhTVn6XjBf4
K+g/lrTpQQec30qdb1AL63C+pgr1H4MtDk8BnIAJfAS5A+0M84PLV2p4uR/7jU0V
lkM9tCxt3Mz0dRGkkueNUrmiVO0VmSxCjF5HlsyDbqH7H5fYVPcwZsebCOBDtN2g
Dc72eH0XF5+0Y2BlbQHzpE7JdlYoaxXXkTwIJ1h+qMV5WVNoG9gg31HUn85aclAE
ZQG1FX+tOB5/33258dg5tQrt8RGyU8qGwIr4P8nyku+kzolT8Fxe+TdtlZ9bf7f1
b5XOazncafEjfntnZkIEMIIylKKYdFXpNznSmHGbnzyqTou5HaeYQOFfynMO2yT3
AigLT8Qn9dislX0cwpuHbIoxSAuEcyssobAP29iBHhxTgpMpgvu2qTSi9OhCwEAo
tmHZhVzygLRYnwikOuPCb/8NhBQ5W0CVSSG0lzF6eGtr6DtEZtxEwr/GDin8gVRM
B6nZ5yasDDD9iXIKcG5FOuGz6rhZL7STcEsl2ZyOdKSrfFQxFRD+TgZeZnfpXhvA
9Mn9tX7rD90EhVO0asQEc/hvckMqr+seU8zrNJ2CfkfjvKuEj9Ptv7B4vwWxlk5X
ckKO01wlbASV/1vfEItQETsPKXLC/Uw+fqn2YtZpj0+y33ZXYbH++p9qqqTpMGeB
X8VDlfixoIwhKeBG/daO3VxkbbTHw2aYMvFg989oOwd7V0PQ47SnDipb8DrLM6Si
8/UDTdiaaz3zEZ6T2kb48aPS1SsX+Nk7Ff3BQabn/a+3oqoQssFMOLjumGLmYvi4
s3O+vHBH8I303ASDth31bDQfxsrmjfJ75TaJg1aAXYMoCh7PNYnZKnb1MCB+es1j
Sk5BPEVuLDzRAplHuMc2I8uTKekHmleGhSY8DLSzva7nfOD1C7nrUgHfQKcGbLmW
jE+jerLEdj6YfmXEeYy8zm9zIQromjjuqSXIRJmt8qrMaR7kIjeIEgqci9MhPURP
gw/MyLamskX7oJKvLY0F61QBjr9ncKTkXYszRUMm05HWy1YHwQqfQXOZc4MvxDQZ
sak9ZXZ24l5d9pmIYCgrQmoyoFU6uGsIekJ5uZ9a8aGsCwFxEMxYmoz0sWEbQtVf
WSC6DB0IOTW3YRfkNLJWdE2oKQZAKJkXBivp9sTuYl16VNsJ7lX9+skvyMiAkCt1
uAFxD8I1OYY09A+AgnxtFoRicHXHbdPAhR72psWp/1dN1ID0MGB7r5d56CDjg/To
3v2H5+smNf/nlQS6cD1pAteWP2Miuhy+kxdwTkSC4JrQr0d+YMj1IIjYqxdzj+Dz
rDGcCzIB1HAD0qJyaVjvykpJ5HIjSFbuC6ZtoS0X/6No/ufATWngBHJoF5isBKpG
vVNCKZvY5gtnYSE5gboUMph7gs2OlC7tbxnqEGsAgcvfSP0dCbuY7SPuivdFGw8/
AZCozPUzSrFnGDdbShcbjWEOj4e1EhXAxfs7uOY8VSncpG7+RDwixzBuGqgMybC0
QS0R62E5PNzfa7Q+d8TXUWmIt2mTKVX7xqUK+MWV/0Drcgh+2IiYY0EQfIIuRHu8
A/yet/5igcMd+fu/vybNRs5LwJkFYunON9P95ennBF9e4uUVU46e/L1OfgBDNA2h
mzHnJUJ+zDTVAHy9Ckm8lyuIYXB7ADigyMkXVafcKCpHPGv5LfMlYZygRYjpoBda
4xbO52v23VQCZBtxtXTdKWJ7WXopBPEhhOe0/MSTS+tYa4/1+WBenhQcFMXX2ECL
IGQL45RbGiX+iM2AAHU5oIFYMtbabm8bJI8ijNPq7YeiZNXP4O3AFM4a6auCuVgR
lu2vDFZctC0ejjrjIInUHGeEAZxPDFRB1bNbW1ewUTBTIpFUjtRfcieoggNQJrsY
qreFh1sgf1t54Lh9NDB9vydtk9Lmgnl14r/Rpp+fwi9GwNn1Njrc5knoanz3cNPh
RnkfPIqA1IDZ91v7E6DGQEc2DoxZ5UkNKTjpnpbxA3olF7D5nBX6X9ZFH1BkinIO
ZUrW3vqYboKtstid66lpLDyzo1xaxUGn/58Yd2E6cJFoqhZO4+mS7LHqR4wxZO9V
MmLthuwrNXov8i8bkdf7PteRbig7x75IKBW3+795EheVsvYlmgjIys4SsnHhBWGq
0/X8eV3tnl/1D1PFSAG4bC6yhQhJFrPEMFuSIqB49nwIjB6zUVVFfyqwyQb0PLPS
bfOkdRkfwkHXvfO7Wk9794aMl+HaIYS0xAuEy8yr/1fuTPnYeqzbSrQZwJj+e2dY
vP6Mv2kG7ORHN1PKQNP8vyWAV2Ol5cqtAa+hi6CAsYnzjsTOhD7mu/Yu80HLI5dx
h6auEdAOhUFh5f6lijAnsV28B18LIufJSmmF9EGY1xa8s3pREwdAfaXClJIENqfH
r6ihPpG2KLlZNiliVylqsLKGy8WB9D7Owup8/dvhevbx3Ox9LJ1nR2/ggQJMieb2
oxh4DOmtyX6p/KUVX4a3W+Tu02rr5ZO2fm5eA/aXlDWYecygNzKuJo5/lU5zZS5H
C24GZnA5vYJvavxTAv5LzvUtO7HFbC5Y6wW7HwB4szzeSW+RGCDRO9VLdh5UIWdr
/ZLqldkdt3iyHA2PgIOVZal53wiRgQ5h5JojIcDUzaawgdKq/Msja9dZWP5PI6DT
fYJy0rHzAIG7zTd+c52gixlKeVcToRAPv1Nd4bZjPdQoi4+Xs93/uTsuvVYBr93t
SoVrFp0liCNdRAWLN+1hHOWwdXDohfNQv4L85Qq7epKoppN5LlvhCHZtI/akF5x+
ht2/l3fL9sjidr4w4OM4mBWS/Vm+XvrnYAQX8TzgcsHQ0PV/e1Rpj9eP3VGFk4cE
xsSW5iYpssWOG2zHoBsiz4XPBRYwSJmyw+vp26TKoEIFjjfz8jjoa9w5xikBii4G
N1rmb1geKWNEtVLrq8R3mq+BWhWDnULGptFSCHmp0H5Z2qxJloW1Iwqo4yljtPWo
9whziCvtZRsuQXz4WWszHpGyFKAQZYLRwylxt+dApB90vUt+WTy4m1Jtdvs+/ViB
IdDIUchMD7/TiSaMCKa7G0VBdhiKuN/83PI1EE1Ea1d/EwAyk6c238sFxhOcRZjE
iqN3sxXynC9i9E8m7wsA5qpRTqCcSHix+JkkOl1T+EFL1r/y7taOwiJujgcetZMl
efiDVnK7VRRgpTh/6AWh7QVsGJEHhMk971DR7QoOp2Jrmy8iL8pX7bAdFpoocJDD
oRSeQKNUN1yyKxyODt+aBS9NS3Ly0qf1ebNqlI4a4ZpUi1vwqBVdLZcdEa2/6sR6
rQhGmaHW+ARf3NwMZya+tXmqKGs25Hclei5XadFIhsS8kHpt/QdK+pgYvCPGPpa7
Fp8JE64ldklW6B4RF0Reb0pqLVMdhPa5TTgPaA8xlJPJdbQnbztPsPNdaEe16HXl
Ub8AFeeOcP0AXBv1eqKViSwqVpGzavi0eT/FlL6CpCQ36UKyl/AfrYx3aY4CqqqP
ZL98R08xippwSYptljpmV0bqeAl8/G0iJuroKYa8hVyl+X9FP/lWwBpj4N2XTZTj
zKx8SfLI5WTpp2TuLZWtH4sRM8EiNm2EyuLKrB4s0m2Bf2XJGlZgFiNagSGWEYwO
mg6YkLP0m8x0qhle+yMiR3mXKBagBM8FOlvXt3GPnWhaoG7fkgpzBzDAPCttM8pV
Be5augdMhGA12FJdL2HELJDytZnitjVB8vrtnJfejXfXNPJm3eoincueHMGtDsQq
NELvf59oP/asmC85qSraJWqz3hBY8wtPTaTtjO/0bynNXRnYn9IMxyMJbf0ddhlO
+nnaOkw38176+MdxZaCDzgEQCVX/1EbXJp30p7Ltet/9JWN0Qh6UIN4HRGnWqU4H
Hd6u4LusfkczzM/lj1nYGOfZnvtTl+Z0EE2gqOZ0pvg2EahkhEAhTHxGjel2+CR1
EtEiPJ4ibN7T18r1Sf1yPpISJnPxr3GmFt9vRGqBW0y7GbXLh/FxPPtEpu02yxKh
qZHy4B0r2TdH8VbE4bWWYa7AWGyWOx5nfyUQ5jMjAn3MlP1PYfWFLFh++aACdbPi
3gnaE4zDvYz75S6aSbzABd6XMAI4G1jDYlB6T2A/zVoiMfqvc+WwSl0F7dr9I6Tc
+qAka5CKe6j3rWaMKAuCRGkFw1e/d/6DDpc0b/OQ+c5M0NrYgKeTEz0CyjkbI58L
DA/tQo4crdG1ALC+GjY73vgDyPA57Gi8qfjZyblsbDu46baC2olEQyhHKKbZFZH0
QKmxINGrNbhd1E2aVMLX5W37rry/OPXb1LjhNOUIAeKNnBDkIiTORkNVru0C0J/p
hrNbDgU+NdSnr/+a4zmgTqUCHYVe9h3evcJzkCKZX2DBZBvReIreWP06OsZOvgFe
jEvxqtKBhZpMunaIsVRFDxminrYSd+RxEeFvcCvG8MxbGlu+9OH8KSqHhN7Tlckk
em30VGnKijB2pMbDuLx9q2EwfBV0vhtOowKaBy4lsPo9O3IVehvhdwdC81AlxpwW
M7DmTVWEHen72EVTeBl9mZwvEgloH+IcCfCABoR9+/K3Ou7BHjlMHKWcKi2h1AO2
c/RAUjgqzCRTC9m/1J1CuGomBY/zr3IEAbu8NCURZ65lvBi6kD01ZetRcBpjBSc+
8R03aGKsFbnNwz8jeOmPn9aqi2VThexk40h3ixgAoGEP7Q8v3w/73ce2WJwc6M4y
cUk1WE9AAP3UlqIKSyeP8t0m8Fej40c/CsYUJOkhdkQIRBsarU94W4xfocFSsKgV
+aEMMrNsLuIcUiEZNqYBSZRonAoDwNT03DwaqrnljZBiB3UhwYNo/LOZZBL0UslX
9kgN9LkLz+x3xQ0BXwrDgc6UDnVimtyk8v2nbZdrFUPRAnZ4nHlfwXq+2Xx0y2GM
R8Xvj8WJwpc8BE3wSbq3d/ew3MEBPONH47VD26GEJLirlpBJk3sO42SyAFLZMM3T
Wxu6O+LkawQl6wPluo9yhlxmLxUR1iFRaWIsCmhkxZ7R+2pRcIDp0gHPCPUKYX4Q
Y4D8NSySURsgi090tjSLLO9oYWMF97hKkjHz1tyvGCJx/5NYU5WinEdEoNEgZg7B
dfQ+2hIqP/FJFgdXZkrHNkvJ3RsCeauP1WfKHNoxKxNJ3mHMUKSrtyxemCeXvt9D
NOn6oLo43/Bwoh4RZ4EgYcKpYMrRtIUiJI7rMV+FUv8qluntDLGIQE/9IcROgSlz
T3mJ1ff0cuEPBquFyfRs8aKRCbY+Ag3Z+Lutr0y7nJuc1NcO9/Hs4Jzpa3lm/7SV
dYYNxUBLyQrkuLy/qNa/VieUxwwYFdN12W2z39t7axeoR2SzWBkZddBUZMVhOKOe
XRwN04xRlqyORAEkcd7EB/7ZHm6ZYlyTFQ2/qD4vzTVrMqvofVEj7xgq5wM9jr/D
A2NiZC1tDaQ7ZkgxeHj+fo82FxOayfL5idXSjlGJuRAepHrN4JPiabv0CGnPpnsF
9o8CxQlj5JASjLVKLPoHdn+UAIeix31Uyp3BpiQuE1XelB8vmILY6MOVPMAvFKgl
ZrP16+sdZ6UNbVGYAB59y6rDTDWJxrSDhfGD2NZz4XXV2cGIFfIDuskaOAcA2ZK6
7IbLCcDQAzSfDLkMmGCVmXnzAq/KS+Bgl1nLi3QG8u5l5SV4KhQ5pn7qXby6kLCb
MNgIE4wtoghQEpCjXVYjRwVQwSc8E0LHtFCvteeoHTlOEaAQiPsBdcYU6QuSbyUC
2d/oL7POh1bx1PmgSCoOoWVRve1CtA+4zvaL8FZ+udCUvZzZ1Di7YaqxqcoG5/xQ
LLwsY+B62vJhRi1u4slX0B3ORUvAtxtqZ2Yh4xlcOGs1Ws3m7C+qYMN7Jaxp1W2t
gj4f2oSO+9df6nH5opCQAfAYXQzr1ZTdo+OE+bLCcNC95eZIusBIvL0QdJXPSIeR
LVoK/zVqdj5xght23qHM26L8JWakHchcj1nSn3qUKxjuGu3UwvZYdsqcMoVyvYKK
bwLEfdjopvWYl1eVCdySYHOqGh8V9kk4750YhX6aBTH38sltR3dL/XqCaiNucY2r
y9rvZKE6ztxgJScn/cfmrb6dKtXKbjKNBvkOpYY++a7gUknu5m2Iai6kX6Qw5u2Z
imS55oGjFTsDrPSCy551MYYgCKGqnSIUtsiqRUiwJhcfWk14pkkbxM6JnP/NGCyD
I4/m5/UVRWqDuiZYjcUlowuEeMQnM04TS1mYb6BsbFdr9axOHfQk77mZfvicY0YN
i8yJd/c7TxpQmPOXtn1nuUpiQ1ieLbH7YFNk7LBJd+n9lfYojfJgGk0ii1HO/ucU
0RiojEAURnCdj6ck5qRcuNxA5xG5BAnvcabBduLBJ35BpyZDhsuwxLt+2DL3Rq9W
mJPYb3ubCqbWN1aXUHgTvtpz/qqtv4ERk99Tv663dykAenUxmDG+DpmoPyuFo0xo
s7+x+bF4BCfcdDlIUDgv634d++YxeLNNn7SLk5J2+Kzo1E0HabuLUaHWjXSsMcl+
fcsVfC1zkFAKz/GdRSA8LLyHtRkAsIoVDYcqmB8fA7XIOi4fwnSDbuH9DA4XZuBN
Fw7v+vwMVfCDyQjSSXwuHBGrrnLDXSNF4ShJ1Z798/c57FkN7iY1yhH0BdR0VjIY
AvK6SClfwoNtn4t6zgiLKW70Dk/SxFZ71qXOX8swHSc+joYKMlZUQsMnVRlNQKyR
i2heK+MORnjHtyKugSXu05meX2drWOinSAYw8ei695uGan+dODopPNgKEimcD0+d
cnAFJ0Fr4ymYqQ6+ltFmvsHjOlCRJnq6Tx00k0e6M9W8RgAlI1AH9MnuEeLf/RLD
01oQYvNjlE4r1tNgcQ4ydMk0cHwz073rFGAtQ57WWS0F4YdOtcHYB0eErbNia0OJ
iuyg59UreFC2+/ccIo5RtIpVqhew6txDKFHb72CSwxlm06qi+c47J63YEygOQfwS
mE5KvbZm4BZdXpxeY9IrfOqN+iMGRxFzZ4N0KWWn0YPvQN7jYmVuygiRZoZKweky
egpUvam8SfLfhnX2A4nFosd7ZBsbu3LaMfrOSt+flo64S9cKsngf2ECsY9JWq5m+
k2YKazmFkC8kMo+1iKIsWqAZUSpH5Xg0ERyHZplnYqJ68IFwf7aXYaBHAEpL98mo
ahS1gIqSSWostiUImIk3lz4194tsmNZtngb5Cv892qCz0OhuYUAifCseFzARokbW
s7lBJq8NhdGx+4dujsDm3ZzUa63f7vthvr3jKt8gK9q42B6a0p5nA9xGDIwM9lRd
sVSmrmd3Jtq1VtJVp9sUshuITk4nrqZ32O5b/0OzMxDOIr1HcFc+ypiTe9LIDSIk
rHLt/owpn9tMpycXKD3lypA9zgWVh2IHq6T1FXu/cm5o6MBQYNluhl/S0l/20zD8
wcTP1FDntk4RCtOaOSfrQd+jBLeS+Y2K+0RXov5lHv3JJtH6j2U+NA1+o3ueANqk
ZA58F6YhNdcdvZIuUd1ve7Dhq2NqjfldTf6nmaA4MWzqkpncBJhhA62dx8oIoURH
d98tcfpCW4KRvQzIx7aYBG/xf3UklVQy36Dk6go1qrIROe+rVW8vHR7houCLd7OR
HOY5PTgfxZBqpSuIWig7rTrKNJgN6BLoK7umxPtcblanoqom/JBKe10VoMItBU7W
GwrOQBeHUqNP3zFR/bMXW64gHUD91XjVRL/rDpMkEwp+hHY6Wo1tzfbUQSnP2uka
N36BtiIH5jJJDsgIyBlGfasEpyso5PR37x5cSzKF5CtbKxeu05Rkm5ut9U9+gLd+
3JUE9v3w8PBPzbs54IoLGOQYzOVUQAoFehtParI+jCEq3bKdhsnlSr5GeE7CqY0A
ET8plXzF0HDJM57NQDFIcqUUNGyGXau6F1IGu+hwBdn6OQ3UGod2ly1RTLMJ/ofF
Ih5rP0ATa1p6U2iFCwmYFDHlWq7FOpgrn5YekNFflRg/vfCPbIm4ej+2AiFAncQC
Pq1RvVTGxBxIgkL6oPGigtiP2iexoAtv1JbcWPvwYqMNplyqgCEUGlRCj+NZ2HNT
yfKrekPwB+DAMYuOBRM+CcdIMKcuDOWXoseca+UqjYePZuKYqKbZrHEskCotuvlD
3s0VGxBMr867H1Hmx6vf9B6v5B5DLAoUBMEE2AM1uhCvk/C7sSToXuq4apXsGpYj
qEZDZ1wzvcyeDc5oWizzqNXp+MT5hUDfLr1JeYDeLBUK9A2QV+Jmpbv4JkUkJJXa
8mgz9/t1S3iKlXApV1gtlBW1zpnW3nJn7StI+R4CVHsnuE3keBoVNWLnefKEN7LY
kSrBUrLVLkUX7XEb2WtEmFOxT/59GZigCRQHTZ6oS+tjPkiiV3hJqyCiqvKueTbq
5pGn9x4fr37CILpoHib+mm2N6gmtiBOqo4r/LH5bFz4qVZaPHgRJXc0vQlRTCxUD
K0o7X/l8e6+e34iCRSkc7f8XQTDgxfsAB92rwbGjIr7tIrHg/6/llkzSTX81O1bn
83rX3GqijYe78PSHbUF6h57LJwta4GnYLVJmVzoz06PJ9l04iZeH2/6ekxLClS9N
QGhEV+/Twp/nQmoo16T1ttztYIvStST5/qOaKVZKd22Uipv+xcxEnLw5WawtjdvV
7rDF6FvQxKpOlK1U4I6y2iW0LNZNRMgaa/pRZp8P4z6AE4P3XlylfVzWVbjPVpTE
SfUR/5ujn0+MuJqUBj212oWasWhlpe7AaW58mDNcpNZ8wfX8s2MrHe6e+kUZ8vZe
+5ImbtdYUSAJtLMFBKAz3Q/JVGLNHUZKREVhlaJ6u6e/VmdRudFAjmsrn0g25EJe
q2u6xsYv1Jk8FLH4Z/YCrQmjg2XNQ5uPgN9MXRrfpYcasUM2806KaskKaEpuFeTG
8zKRvzNURiHEIyjYc5/RlFn+adepU850FliuV99Bm6Pb8f6qkSQk8Sm9iuv888GZ
j7pclWc3k1dwpk7EWGZsKzCoZS6Q97dZtKE9ozhgEc8zjPhdLNHr07JpE5Ngj5xt
nxAsVnRRCvRmQSo3hzU+AZrrV2kY95hIXneRUuY+H1qK+HV9FWB6MAp8RH5lb4/6
oj/ME7SC1647IFuJB5EmhWo15fliGehb+uORveLYD6BmoneXzhLUMFB059Ov6HFF
Nc3yYsUBmlyZw1tHz85mVtQzOqxbr6yOFtMI+SCWogXJd+2ssl6QciBI7mg5p5WO
eKgaCpDP9h4rQJtRYdJYWYAfIFN8LhH4Sv4dKyj1AixW9kH/0n4UZY25sCfn3yE9
XlphjiwVq1arKagZWTye608dX2UlTt9xhT1Rj+0ysGwPU+3cImhWHkDDOgNjqywE
lf/PFVu30Cyt8c4rxDEbt4k7yFjTGi341U0vmV3JkbndNIUSSWybtZ6sWuNxJ7Y1
M/a4p6bGSBDCLDIjckp6PVIJ6LVw2jZqM8s3BX4m0JalZ0ux+W9acomhS2tCjsoq
7L1/pt1eY0M3A1/44XeMGpaJovcqXCBsW2DMOQvg42Ev3LPSGrIqTb6poGEa/skD
0XIxwEj6P9Pd5PQIFaXftAaWj3nOkxmYLIvPJZLoQy/KIHAWuAgJoppaGNsqlodu
gdMUrv51hv2uSNeZ5+VkohB7sNhfLz8rNtUTphNE8Y3KQ2XOzT33u3CgIgW5kJ8y
xhHhqwiEDsRIMVCmjnDarRfbE+kO0g9P/60fjr5OXJUObglAhV3pF0Sbues60Mpu
SsLVqgMc+f1ZIe5OrKeLSiBOSp0zvQWyXsIlkbOoFiTg4hBptLz9ciXn3H6XrF02
0wLmPGGhOglQh8/Ya77iA6WgqfGC+eXn7xFDOHwMy/h5BZut+IIoZXiEALyA85za
ITXKjVA/ODYVDZNIe6o/q/799O4aPau9qLdgUnquOof6QSKp/Ip1mYofCcJoHsKj
CTuANYq8bgu+SsNZ/uOLpD4evBXOImw4zuBqRfHMu2b2cbTZied9AEjWh+jvDaRN
VmqXhLO6zwx149qS1RpoPCMDJ0zafKH4wu7GBG0Q3dEO/9vtCbQbi4guZ7HFi1LF
Sq7fXW7ZOk17m5gabfziKeRdFs3QExRqKL2kRMAcVcJFtlN/j7I7HKCZIWuoaPPB
N+rixFbjbpdXc9R4hIGOecR4wOFBo2bQQ8gT4AeK4lMygiC0X2LrBEsI2OJ8ReR1
LRpnwJARtbUPpUzCHDWMDwJuQlMj6wdD2Q5tS+XSDWwd6gkBGdUmVmxX6nYHLwKv
wFlhaC/jzOf3Bu97NVTim1lGg2A4a4cQshS/j3aqUZwW3s091bsBmsWvpx028mbN
vCSYNkThoM7WZdMogcZNvKFK+VVn6wKxwqQ3D4rHXixfip8uBiWnUjJE2xw7APpK
mQHu5xR8+UmFtnafHHUhOompRozASVjiYFUhVZkDWpcluoUxgAoNOEwJBrGaf/AQ
NLAGA2rLgb1+inm8EzT5PAlfBnsuYR7O0svMi1iVuwmaUZwjRuchrA1wC9/x4+pc
Obcm8tuRsJwGBgWSnDV8s+3MzUN7PyxB1cO+X32ytC3n9O8QvutWDE8da3pzSG9I
J7NJomPymADGJqyZqSDI2x3K3DSy912o4dogAbEiQ2/4BDyndBLd8AdXlXP9rzkP
G8+WjkCN73Yo5DNS7quWZv/TKrht5hpy1IGmAXA8BKY3Jb6R16AxbsyLBxbjVupp
38kdrmBkMjeca+FOLsVsCkdkG9mqAn1pTnhuFGMGGG7hIRqd43CFmH5HAmli5JJh
J4z2OsRFaS6Odlei3lGmGoGJVGur/RyEcr8P9gKhYNQwHErRRmyc8yuefo2+Tcpa
X2P/CHTkMlIjXT07DxVzJ/gloU870O7i948tZ0HY+sg2NW07fAkj7IH4xIt/zlO5
hVS3HxnDLsEV6NPXyyKuxJEsFcpkxbLHBqhFBEbc7LxgT7CQskD2rscQH73eFh1f
hFYaQ4jHlq6xHUhS/qCUCJvJ5XjzZEyQjtLHnqMDgrB5bgGrGlxkSB32638QXpsm
ktm3iBLt8V6a6w2ocfj/xZS+yFqp1SwEwPjRGFPoco2M5U/I4YdrKJDPbr1eIKv3
28xLiwyUStHVfOwtywUzS5kQ6d57RAp3Tbb0FKZTFQrx7E4ilUyj4oYfRH0kvZ3J
5Y9Ep5evf0S9aAHwGk+riYCkyNdH2AQNpQ27++Umk6HxdwW7ITduk/cDVGmJ6NKs
YbIo3yimQDZqnNqpR6AAH6wjOoOeb7KltGxf0bdTmsacM4oKlcCTc/TVWItrVHsT
luPMdbEFOC/XF0Qvf3oW5LZrS1x4pxOVkniwGezUQrwxyiCZ8WqNlhk8SVIpF0AR
dDE0FMCOiTA7ehs3Rg1WFdjo9Q1J2zMcWTpePj3ocB/gbrXekbmekfJzoLX1h39x
PpQW8qPBB6u8cODZxt/r+losocwnaOkAmNxz/wdjWjNJ7g9WCcOKfvTFUuJ/fjcv
VJT9ubHv7cetQP0rTtPMtgMaEXv8uAZceqJc2IFPvZ2+qqi9wf4HkfJGcQn5wBg+
PZx3Po1ubDnWKGb7NdcdezcOqHYCbiNJFU3BrQAS3cTyGLLENysx+r9V3zTVohx3
`protect end_protected