`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
ddtXksX2+yylW5zu6QL2Lhnb2d1sD00763mmSITNX595NcHTEkwn0zB1Dry37fOW
FufOhVzEJp80NC5qZ/+F0Vk7Ik02dIR0elf3clrjeJRK85K4e3Hoo4xn7YbFUIms
l/8VZSb14+JVGURjfswrIyCUotIzlzVYZ6gzoZwDXIi5gQIBf/gI+KxNXPaKV+PQ
Ufys/12rjO6aI/pPlqSm0hCvftmBcnezN2hk1UeXgOIuKZnogjOsf0iJVX2aOOWE
6pD/psybjbnsNB6kH5uFTA5frkzIzkzl5d9+YDm9OyC+k84E83I/7/j+rk4L2dah
QJOvksSIzN867/4Qt8qYTQ==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="MvBXkzurAa5VTw+1JJ70nePUfoQXBvZOku/SMmg4TwQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
oRtzZL4VJ4iwysPsC8SXYCzXS8Fw2gtZTOskLcDV+1B9Nzn1zTyNtlo6lNICRmmK
ZRVu2BmCc2G+fmzynYlNTnSa7C0Cuel6FYpxCBlOuk3OF2tzAmLAuDyOH3Z1Yjzk
a0aHuoCdIRKv7BrZCdALt03JeUmXKPdOmIlkVGFl8yw=
`protect rights_digest_method = "sha256"
`protect end_toolblock="Jn9CQpRhJt4rnzZPRk+dOpzAubz7omckX1MrFd4p81o="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 23488 )
`protect data_block
gD6l00tciPUa6pDNTk/+t0OO0nC/UTtBwLB41d4inuAUA3i/ALrNyoJVcBnAmEQW
ptbcNp5fxEUJjnOxnedyZEuEBxWRieZFQnkRdF269oP8X9HpANA71fSaR15d88po
2nbXeH5hTVY2LTDfJzBhxVDxIq4B/zdeSi6JgIv7r4aYP8ucj6u5neBxJMf0oAXU
C2CJsXV4l5DzVLV9q3gl/ecKSLRsFxcuxhtGem39aQTA2+wArkQ8bfIk7gdEhnYL
C52qTIHANL+6Dls9Xj2dGs/PuWfEtgiXpDTxfN50OXs6W5rFY+irMFdFfLFxIy+/
AG6b3ut3qdwEeciMLbfsr+TqqNxNXTd929DLuH9+gBCtBOooMNnJqDn6NJi+Aq4o
tbDuDCN9KqpSlhh3gxPKKKwe+sB7oniuMSuEzX4d3zGcBuu5WEpqtAs7y08h0bi8
dtZxPXhQAv4Ia64bjtdDkLzFWmSQgi6/Z/9uh0HPljjXAW7v5UhfR+v4Dg4W2m03
NGV/4IyJHqlfTErE1Vu+wVD/Hr5QwVt2odTTTh7GMVme3nh5WtMcv+Or+rkLzHT/
I8+Bj+V70hDmbdGkTu6pD/Plc5bjmy9Vf4ZiG02vaOlb2BrbW4s9b7t8GTtP8ena
AjfE+Rj8JFjT/PNvSQcfygDL8KJyqbOLlIsEADB086MBqOD/1MjRO75I1OpFll0L
uvRnCQml99l0OSxcxn89Ah5M3xRB1kKaEA2soCkEXrYUZ53N8i6jzqeHtUJ6QiNo
uH56JXkrUAm7S3nJ8kqF7widbi/K/MBNAU2WhS3zabSA+eHo9JFCKi9iymEJSKJf
gULaRb9eaAdE3iStYHQuW/Ro0nfoBtHZU38rZdrN3qzjJf5o4DDPNVSCceg2dXnz
gaz7BnNIcdv4zO6e/XbjU2A3dQbzsnMAtiOcvHYBG4oyJZqzSx6KsyLvpEetPeFn
oDvASplhQbGkkXadO7MPk/hzK7gdQOYWVlb1FtqrlTIl2TX+vkLxkjnd0zLPnt5U
w5CmzZwLxS0mKrFxlTQo2Fv9D4TFI5A3enee1gQFJtpsTPtzp6YcOnijd8pwlbC5
FQgt+aHMXj9FQx+3xvxc96kNV032Ll74Z/JSzC2BV9p3ekzqoshlL7pBqVndd22/
SBm8mJ0Jmzwe7cLDM6Ae4g5oIAQJfaeyMORusTh1Rsi6VRCxTOcne8yPCQsUULWB
qVuys3DUir195wp0qrrPjZ5jpscEdXtRS7ord2MBbGBx+7mNRE1AzzTsOE6I+E6Q
mVYWFEVgdVR7Onk0zRgj985NCSyTbTKjdxikrjcxz2CSFzgAiTeETnhAQ58bAREx
eDWWlaWHU3b1Bbg4VQUBg3wjI9v3xVw5bjrlzAPEJyy2oyUC9NGtIAZgUmEdoS9a
/ng7L0wLb9oiRPCV/FEcYtELwysC/YZx6+T0SyCitS63265JTaALVQ3afE49q78X
yX3YDakZdwkDfSR5CUS2dyPmn53m7dx0cUuTIJIE2ntCrtyegPpNBeDag92MfXVK
DJ4+QBlsPlcKm2b1mwjCr4z9KOmpSVcVZi7/f2K8b6GqLBSGdna/yvFSJDvZq15O
+WRfb/bHig3+xMYwRduUCkEB3vN+pUbzPUgdoC9TZQgO+35OUaVIif3vQ2NAcvWA
1O0/5e1b1uRtFP7T4R2xvFKphfW63IPgDR8QapZjZN6SINcL2eycUfKo3cWmc2cW
CDnBS9/xM6Aq0sYYVq05J54L/zZbOtUU8Y2QngHd5L/A8HVn2kdRbFU+ToqMxlGd
lb0QCqJW6s4a0JhcOP6z16by8OMbeJ2rmgIMrtl5aAmqf5bA8+Z5eWxfZrbLnVjb
c6Lo2ob87kUt+zpaS/6seOzHcLNVbIncocgW9PyxnkHbB/3yyRFC65XujwRq9rgP
sesZuAA4lOUQGduLhnpHC0av1FjzVLZDu7s2QXmzGfC7iRECkqsg01MgDgqmQDn/
35j+kWzleZ6nHueo/I6fT5QYXUbaebhXcLc6Zs8cu2dxjMs/orgJPU+Jug5dz/a4
MpXDq7Dk5c2uFWfk3mS4lGhWmH9HexQt8NCszBa2Y/nYZHz6mzv5TtLwSfV0krbn
hYSyJgaSAUDOgYHpqbO+YGR1V21zWTnsgg7WqfPbG4rAVNAjQRv0WfClyQcv7Iqj
TR5ThlqbtTzeEL3/ecByYV3xymOb0Huk+5Q5h5LJmVbCbBDVSlmJE2878/u44vNv
mCz9y6gZeG9hBQzLHdIfSbE1iJmT9wW7PtEovj33VBry0LGUss6p/6rRsMDsNs1I
Hrgya0oi0XO+0VU7Bl/oV3XqUY44VEXie0QkH4lL31comTfVFIc3jiG2iqA3aBYT
SJlBaDPLf3g8sAS8WSZeMyBITmsv8cP4C8HU9MZTtEHdg6aWjjR2VqkjF+6gD+8U
oChPXT1osb9fTK8BhMlT0KKMwy45nU96Q1goVZQcy4EwW9qqMj6+f9e5BZXUXUF6
yOev6Gea+W+fPZpPwWujOfsOm7+RswXktoG5Yw68m3XO9c+DQ159WcEsR4Fj2fKI
UdoijuBkUeGZfpoRUcchf9UGMWBdh2UQBm1/s9TGlQifaSAJq/BJAsIYUjkByF/4
ksssTm/bUAR2udedzwskjZV0R4fXpkbOFu4SR55UUTj48NpLUVnFS9qqQmPz6Kzw
2l375luDs5ouKyiLZsGlnu93p6v3tE09+uUttwMAKh6nla52+ZW6+NEdJ9XFpB7v
VS2VseKbrpcM3id8UthtwXMs2K2JO3J4s17s8bPjMPbLs2hHiGCe92+5X6owg+il
IraspzHioDb2XSCLevMDXIVV/JlOE/XpCWYZ1WAT2L05AWh9hcImq47KFZ1um1xc
3hn40wJjBdPt0YkpK6qjZ5UA8rqTDnJILsZgY9sCrXovYPU0pwDMdozABOp2/h9y
hQk2uijt7ePyWqm14aa1XRH3iBciKbuZ0heKS2YUTEtlFwpFaP0iZD66uPM9Tv5Y
gcijD8h8l9qvnCN+qg95swzDU7YgDclh/FLo62dw3/iQEplbg6hXZqIpNyh7E1xc
d2v7asgK07TCcDd2x2wSnTTLF8GBd8VvF6V5ZpqxU33RgJAKKlmj5rdGa1ffRv3x
h24T8IY+FbUpF8Jp9lICOEWuhyXZBERr3qBDaX5bljzUu5okFDOCYnt0vGQDexGX
23n7/p+mrr0blbMasuCYbqtt/qcdAYtX+WGWxX7B+03ruMg9HTrlsz/H35LYRcS4
wIFjuVIg/MpwodZroJPpSi6o6aR+eX23BWaOe99r3LUj/W21tZ6Cclv3NzoJji7s
aX7IgeY0/KRVPe42eJKgmjIL5g0tHxwaE/g3YyjGX0iNr6RZZcp/YaLCIV4kLs++
YTj465pRveUR/dcb35UIlmsp3xL1sZHGpbSVfIq41FuKlsnQN0LJKWudECjv7co2
nGT7eHyZoZagTwMJs2+NpfZwxLRaK+J7Yo2WVWvSYGzeiMKhSxRhxMuwGyaVB0Hr
B4xKfaiJ9LumQDU0bBUMHrRMZJDUer5gv/nYxQN2xzaWFxrHe3oJ9QrMuZtTcZFv
J9ktjsH72D/LwIgL3BhQLZZ6qN2k/tHsOvXPUsKKxulHmVA6atJgV9Mt50KsjVLs
hIYsp/nNeUKDTQL03wLdRxIQsYM2IiTQM/be2brmrtdj9Qn+goiy6fRE3bxRuvWY
dqgnnm7uZAGYot0m6ocqm2Il5Vl7Wr9L04NsGQ1sM57HTXu7UPUzUv6jTsJaJZvc
zXXckSv/hV3ZiJWkz9BhzQ9Altv8Dfu3sK7ZoUU98FAU9Yg4e1h63CXyV4z35kmV
VEs43Nr06JqIU3sVpVCTP1qqcU0sRoirluoyIReNu4HTBLt6dCn/14MDy/4FPuE3
6PlFN8jdMnV29+DCrI9sl7Vb+gGJyWLTAqInxuafSeO0BhZ6GZUi8sGyqGybWmMr
sKyRp5lo7s8Cehhj+pSVjdXkppbx92tqErjsch6shpFlaVlF1IffOdyb3Jw79hEk
QbtIxuFtUMoU+nrSomqT4W3i5uhTt4FYhmUxAqlvOWwToPzlIIrlYkq72THHBKVF
ryZDenhqNumZTuDJf0pNXKfS1rxQoG45kSvQlNwYnrNTc5/P9OGNpI54RqLHIoQr
E7puZid4eycmfgEE66QgdneS8avnIniCKhzrpdVzo1XkRWM26EDWFQN8rdVpA8u7
Hnh6p5mu5uSYH/98/5vdNqUGWkj5V4uN7GQpB1OSHA/CXuIpkoLsaY+KqhRqnNqH
NkBlDlrC97uvpA0hi/NTWL14ACq2cxjMtsGl4g5g46Sd7sG5hG4aXAD9A6WbDDww
9sP9vVE8rxAUykp35VluMVHQOfWHYOx6XB+CTX5eg7ImZgyEd+rOwCLHdyVoIV4e
sna5rDpRP21VSBNVERgKkuPzVqCV6ibkkAZvAOlMLJ2YbHlcD/XWYchYr/W5EzGl
8yTMuoE3AKKJtNo1nuh9/FH/8i6cgXxrdiFHtQQwTjaoj/pVL7Sf8vBmyiC9kFHO
6ZR7JCb+LsZ918pLyLk8pCGDSUh9msEUy9nHWB6D3shtMvvW+x0BhU5q1t+iXLhE
oLM4/dYGLWisyltdSp9hwJZ4UEytFzD/Y4B7exkCtMZ235X6vXvJdOo/4HLFEUYw
4hlc323i+huZmTBCbiFp4DhjZMvhFA0rQocUw5Ymz9nXEZ8XCNJ/46+irc1T/1NB
DXHwHWjVX88Zjs4phDfJsYVold8y8L/apXWfZqCn/LBY1dgFkmYk8MoOswS13OPE
lkDnff4vkEBiHQgDN0bYfqcT6VHCp/mexmuzABw4ZMInBPxpz3Py/GMFzD644MvC
Wp2y2EPfHvKPSotqC/AxzffeplwGmyT2J3SyJQsiSyVqCogHqAiClvhqD0Fg6Zem
scOxt6TwHAmrz16J0mX0UDwYmXubL/bHYCKXl+2GubaE6UcP0bWz26PKJhzaoW6X
+hE/zM+7pbd83HU0VSs3wqEXq9brmWHk3eYfIG6e6I7+876SGGKIb9IX3ZVsHBFs
MFiZlZ4YuqfZqu1J4mBwjWhQ6OMAfTI6lit5yfUZ+wwPh6+ws1fEyJXXGqjR0vCr
9NSaqCmuzdAGa4ppeJ7ypK+lDkDHm4ofQ2aQky8uDvy/6XsVig4XaRzwJmQWXRgC
hiwM2ncsK8i6bwsZtkButORhPVYVMWPMPWvVDif18aRTCEYcxl2rNpjR1KvuEXzy
LUJNLXM5iOJdlLutcafAIDUA3eGr2x0lFcWVAnh2q9LG09E88RtXAau2pAhyLyEQ
oF/Tn31xQCziELAMwVgh0wlPrOYqttriKtmVtacy9opCiMwQCIgUCt7V/Uy+rN+6
+n3L4ftxhh8pik4MvXXNld2MeVAXHX/e8dh1xv3K5u70vsuKYiPz3C2+2JfYxP8B
yvsQwb3ZmIvclKuEOEL0uEVjk7LJGp5Z9pdILLwjKCb5DuhcHP7+Dn1/tA1M7R5a
fxWkv+PL9Ezf/vw4ZN7nFX1ceP9sa1XLAmTHiwk78oMr0OIS/7ZBjl6xC0D+1xe5
xNlhav3XnRWLHV6rl9FvADzXJ37sHfPiE4MR2sesn2Vby5cZfPj5NrQTZYpbXoLG
Vxu7qqJKw0ihbZwCRKvUskmDxzl0Zxcjm+SW16RJ3zq1sDprk0zJrj1dKu2frj9u
WlttWdzrId99Gn05+Ew6HoF024uF+WHMSkb0Cbn7mMzUzO+WXAQVxuFOXujG40lQ
vF9K75MiCLyUOwwC7d3G7OppUxAI7xO0pQChNPhJbEmbnRj22/UgK+MGILtjfkTb
M0DwJtZ5C9jMzPl5WbIPkL1kaUGs/HlziKihTu+hGygR4nhtZqPIUF4t1tF5pBTm
vF7AnarnVDjkFJpEogN9zztSqtbTHNVvWSbpIg5Sh1Ifbo2GQ8Yt4aeTGP+BQFfr
g1xYiUjgkzpKwPwOJFECwPED05RtqQB3hNXjLekQ5ji90y7/KrHz+NIAefRbtL7V
wG4AOVD3dlExs1ljYAN8jdvqWGjjVwK1EYgChfkThteZoDpgTtDg/8Xa8ThPTWBa
GVhitDnYx+S7FrscQNImf3why9ka+MXpWpJSx2Tc7lZQmFcd2cEUFBk+Fh2/m4c5
iROEkJGvZmbFZkyE7DZHe1rUxPG32FSqIaopblRw+Cc64XjhdZC7LxxTdSl9Qeby
u73gkO4yiDPjOnXGz055RTUg8iu3a5UQIo7VqomhC42Q6yQAutqVO2vEZjsAPt0c
stW44UJnsr2fCik1HSLbBr8rhqOuI6z7OaG26a3EFnaw/uGv/M7Pi/QdkfzwtuPQ
/Tk59TOp6UCsYKH7uF95cgtU6suq6CqhohymEUc5IU9DthBWar7P/zy9Wr96XJsd
uWkSRppMJtvhVhkDYBH9vsuB8LMYdt4qMpkCdBfW28/gKX5PgMdRriBA5wWPyXwc
69Paut9grlyBDMVsWOLy44Eo2D2xvIQzFAW+oxQSG9rL4aAr4SSJN7dZ6gQiKLKS
FfpPtUWj4i4bE4kopj/zJd214EGGY3WqHfjsDfPfcFJiYpiCILKtq6RCnMbUl9Ga
lOVojfTrINRCiCz6UzA0MYXdJ7A1xNv2ougfiuRsIvb03kjmyUV76+F+Af0MCqoR
UfbFuw8F+XdVE4AVm2yLo31/bp7S7uvzuYxeAILi7hFoE6K64XqUerCCB6+ZWIE8
RqAc3DzqwPtDYOYkLri/5+L847DSiMYeUo4qLlYUqaMrO/usOhWqZ7CS5vSFaDIz
PZpqJcgMB+TlG7Mm/AsyOCOlNT1wWtPlmJfuYq2twNP01lrG9J25imu8MtT6907a
QLKhxI/hNr3v8H8Z0JOMDKe3SLWOY4tkq241QhChUlP4Jpg5mnKL8r8dWTLl7ta8
aJwWR3MxIz4y1QCSYx6t6iyvhH5P1vKlO7hipZTpcYkEyAYs2lOtX+cowa4BNSLF
fRFboDyfT2uM9kSP3+TXAuD1dMsv90TMEZdeASm9Z4nWfOd5yK6UPvZu9O22cafz
qOp4X3tmaBzpd/APYR1d62PEYrGL4KO/PbSNND1g9mI+5AWhW1Ht07vlH05h9zE3
qTq0S2K2nbHuNlpq3/ta2gOZQkB+Uu3DrZPivQb2uKJhaFZE32fsbC7DxhNgqfhm
Tj3OVEW3rxYnXt3GuOeu/LHaOphlmINV7DIP79NDYZIrVYOrRATXooxyNXkSzkca
qcR1XD5yPP0vJHhXcrUZ9U+1GCVlDttzpTM25KFcELz9c1Mx9Zisom+hdtd2c6dd
PqjzSwIKh5vi+lBhgLdo+X7mpBvFK3OI+k90E2uAiq6csgpuSp6vbSbZeuypQvkE
4SOJcEFOzZ04v58zeIpI9SqzYdfm8UXD6WWoWafSVim5oMVSJcVHFm7HUvkbotPi
mU3ZphPieyYhgankq/fQuCXN4PG7Y2jBKSoGi8+zCNTInWd/6vCpaMg4R1mRHkfm
B+bY4jFKsZ11I8RN0RxELCIHWKRf5o8H39lqzi4BqeS+2/IW1fiitHFqw5Hajarb
dLO10UeIX1FXhT/V/M1P/Y0rshAl4HxfqkRNyfy2XNSz0n7qqBWrdE7qMoAxRj89
YnNshdQdNXDEys4DSUOLTeiVDc3SFfdFYCRzpVmSFToyIV2L+Jg9RBCdECVJt42S
W5CApyRIOM4wHYUVc8HC89vlGP86UnPSKhrOfu3xnalibVwxdQdx37NOUQi6vMr4
wArsB+fsFQFXg6wXty3G1ojlbodFlNFYfeDFnns1taqgGqHIUYSAYH+m7Il3Tq3R
nA6XGAGugvi+wllN+C9MXTqpyoJbYKcsFOdlohhSk0ssHAHr3Zt/4vr1/rpItYDn
bsfbwZyXYxeMGv0X2brM8o7ycNr0YtYwBoOt3TgFTz/aPLCRfHE3SobRHaibNLz1
tFtnT8Yn3Y39wOgo9ZOCtQGZLEUoN9PvqCIgIvpm5/kqnrxuvkAn1/9tvaOFz2aN
x/3YYm0O4GslKbaa/DBVQlMh+eoC3Rkttmzz5OOmyJ01rVS1KW7A3lSII4dWIHCh
9CO7pD45BkW4YqUYYAsCrONY9XUWf/Tc7YoomSbOr3uRAH76Gyz2TTXGAHlQx7Vb
KXeu8stdVHGgex8Fp/LDIrOO0U9CPbxNc7XObCXGOoqQLmjoJlJvhzxDQXY5p9lP
9r5wsZ6f9ZUICqmOiS948BDV8MeEVnzeAmbWhazVlizYxvWVQZcD/Phuzk3XqPTt
iTClyhYIPWy7XVNUNDgBhYTkxd6KIpKUuTiy696dLDhP2QlV1pOXUe5SNrm6Umv3
J/YS1XreJcQog5f2Bts4nFfbE+N5kFclmti2r2rcY1qhBxGrB5IUEYlUxnsJlXak
EAtHLHTplgwyjKMT5zGATz0xmc5biyxxyu8XggKbOp7RSTamWGMXBx6R4asMWjAu
q3PXb0xj5aKYTCv/T2Wou6Y3lFelgUr/I3yl6Q1/YPUckAsJMs2HsXSoR9YnGw6c
P1XRCCgZEEINgkVwBlqb+g6G5JIwwU65aZCVX9r2rvlInMLjkpdxhxJlOUGqcWfI
wPMKXVyPxGXLWfGMZJl0vBBgSyZxIoUf76r1pbqLHarurx04+NTqQZs2t1ynRPmY
ie1ubthEE0jmtpVGcD98SpPNiIwy9ZpcW36asjbFEndjs7mlCyE9tWvpAgTwtszC
akHlJKAeHgoiuwdiJTzUYDhDvsIv8LKYiQnK8JH5mTE5m+GT3Ga6Jv+GcMdxqsAU
2VxMpp/Fb7SPMF9XJk4ucaiy41nQ1XBXboT9DMq8sEhU7kYvFUv0CSJMaiUT6s8e
FtXq2KcSjsFMN2ScwAZ87SFo2yWiAWehPqdxW+m35yZ/Dh1W5He4Y7UXn6kq8r1w
TUcWAwf8P97lPH2RyjA8/IbmqMhZrul0aLYZl4fK0uc3i9p4iIg7U4LLLqpi4iis
5AoQ1UbfHkXjptuzrCQayQYTsUM4w9SMqmfSLYw+lTPBeNVvhrU1Q0J0EefSwziT
OxD1T8zqmDDX/8iDevmrs3m6jnFlhWV/nPKApO+vNAuPxjjj1bGRDwj/QHZANT61
9ezNo1a+0BiqFbYXglCPU3hP6poXD5qAuzt4VXLwbKIBPaJNMzgkopt9jXVRn62P
iJ3HjYdcb1yzrEKqYnT1oGrYK5rOe2eWM4Gs7bW8ooTGUw9smZtncY3/ID5L9G8o
egkzvPeV1aFf3EwUr0zw3n7TElpgANneE7F3xSga7icQasLJtTkLzKvQDDzI6m5Q
pr76+G5Zz5HVwL8lwOmfGL1ahIyKgSMUBHm4UKY0UGkodNwtwX5DG6VmWi1tiatx
cF3QzNpBRBxwXsTEyFsxF1Koj9dzKGc+JjE5A9DY4UQl8MHlbyLAjZ3HkhxX3Q0g
3JbNhIa8tq6E8hFDXUzNDi0kxgHwCC6YL1Yhygu1WKrEfPnAatt5tASISA9zpkyr
9UGAjbS6V96wGkz/vd0jr9GXm9JhBFNr72Z/LWEaDzIhUuaGLbo7dgD1tvDfb7Ar
Gu2jtLajTg6YdEhCT33U2HsrFQ+5PgRgy9MpiiKGK25QSHGBtKcRKtmvu7HeEZWp
qQmh3GRc34LfKUdblJ494FJ7BFFyfobzDwCslfUjUuKkorf4ss/7b9zLv3bGTBG8
Sd5QvBSjxR1LhxdAlS6XugmNMG3uoHweqkNWYmbhS4qXfJQeaWuuZhPWEAM1Vguh
oRupFLiZJzwnzvwuRqrZjULRd1NwZmDnB98b5phs8CjYwBV3paAYnxXZ1KW+SM+J
uYU6N7bA3ChpiCIKWSdZlQxurO2E+oEPfpm1fgN3OlZZFyidTyeQns49ad02WMho
2zPRP3izYBAxexur+uQanyGroBl19LhvULl4sQCCxFMBIwLvDcTIxfE6JbDdJ3Mi
XoM5YyyHTvyxZWUV1hFQSzz0+SxSdiyf7XAcf6auVdfiC58mfjAh6W1zhZ3YMuey
SX6sJonSTIlJkMysMguUS4fVpwyFWTgF2Ymc1YKnV6Jar2za2UnTiAEDaTCgeKyl
t/eEyDWEhcogvONTi24mankDNb+Qz2pU+X3Y1qDCoHMvmECuT2/A/bjV6CM696bC
dYlOudqZSsaIw96Vsogzspci+qglcwGSzX7vAUtjXpn9t74rawYWjKxbH788+lsf
hxGEpfS2LkLFtB7MFfq8dEIEHhzUru+DWy1aoK8vEZ/nqFgkPInKo2tANjoDYB2Z
ivmcRl71kpqM5tHhF7Bzd7i2Iz9hdsqdX4uD4J1oUiC+2EfEst2qnoFxOMyRojrw
4ooAxTSkn3icDHTu0LPb57O9rzEzE10WCJIzQoH0xBwS6y2rZ+KzUpW6olnoPwim
OlcQ9ZFS61QkL99K72JEec44rHLkmr8ylSQhsXdEaFmtcjLnK+zi7lNzu0ISCyze
HrroEfSxL2SF5v80MZHTVQNyoohSyUjEHABxnrCrtop6xw9kUj1sGrj9THGoV698
LhjB+NiBU+Qq2RQxXfXqsd2nr2Pe7NQX9o198++FxGlf/NBjWnDqKQnRgbY6E0wt
r3JEy3Pu4g48zYnt0QxenOGZESYGiXQNJII1p3XV5xupdA+yJv8a3UJSkPcquoPp
wC9Saoaw8lY0kC+FxMaRLG0qe0WoofJOBvn85MtVdbvjnUcvGzUnm9S6GZGGowDz
T8rS+6a+PcVBtfTEURaVOJP2eOjFBVRjOPzLxua02tc7rold3EVliR9A75ApFVJo
DuU5a+0T1q6/XuDBfP+KY/dqbuhFHnpEIUJo/OFNhn38/8rrvjTEc715O2e+BlH0
cecQNP86p5d9Wt+4qpeQTJPvexjMh5GqDDOscT7To+LdF9fQWbnZHctn2ueOF6He
dtAmHKcdTFq/kjeN7NASp6vXwZ57yog5Qr3dRWOxKfKRU6aUS2wpdu3D2hEV7wJO
8NUkCKedHe9AR6NVJDUt3mg0VkusP/xZ//DRZYHatkOfM6HhWwyDm8jNI3kTzD8w
dxRIwAU5WlGouY89HSeHn0yAVg2OYRZWJjbSsYkICaQD1Q+QZJFSDgz7zCGwwD8F
A01YAlqyVx3ah/TqJFfFcOTByx5Xpd5CEiGQHAQHxEMS5xP/03UiesMieksryc6W
o0RksfHmO8KwbWgfb7F1CiXdaGlyvOBrOCb3Js4IkHBYQr9FwJicSXaG6S9M08b7
H7clqdmZTW7myarsbf/AQNlb+cUeNAdMnG3EIwjWP1VvSEaNO2mWVv4Ye/ZF/4Va
zyD0bXVFqjTpiXXDJmxewD30aACUXME6SPw2yLd9+R7ZaTiznRvHFrSnG3dW/mST
skb9Spu0x49jju7bS3pqN1uG08GFjBrmGX0yzoFlm7/LJXVdpX2QUnpZMmGMM62C
uHC7clMwRLYa2A0buEC18RbsDWHrNB/SdsufluyQ1zcWFMSCN9CqCKZGlHS+5bun
An1z7Vch5gMf4Z1q3lpyFXwj0o9syLjQLudSFxO3dT4F4iuCZowTz7zTeW3Ohu+f
qwYLlgTkKMl8+9lmnxqQQoZLli3pWy01GGnNGOB0M4ylKhlF8tlYcl+M+ORwlMnc
AHIQx7R9ijOqdvHBZ/ZEYIav9s6FlBKOM2E/3WrUnhSa+MGZZkcWkqajSP35D2Ef
c6PGdW2V0thJHYib06jpgp9HIy1d8cFai20+qIrdGxeHVyzdeFT7uCVA6vJNHfIg
uFBrRZsgVuCU1Di6+rGGSmZAPX3lBVMG7hYH3Or7vy3mG5WeFsE83kwXnr5UBgou
VXT3xRCVTHZ27T9w/DdgI9LoW+d3CLQ6DUYYPsUkz5NdlPV99ZdcrG8ePR32dop7
vETPpw3XPkwiBRM8vXDAhFnc/4Y8kaNPSJGak1lRMdPZb+2S/I+dQUjKJ+SWXpbH
ysYLn+RJ5QIskH5Hsx3NLKuG1Oxj0N0Kpqvmktu1rt1ZISM1wonBxeec6RkTkQmq
+Ga/NgSy5wanjrNvXi9NXuqVRu3Gk6rsi+8Z5rxCylKHXhDXlhO5YWnZRccCQ0xO
it4OhNT6ZzJLj/rqOvL3GR0SYHeTCaezsawFS2Zk6mukv+WU3ZX08o9l98fXWzDs
IWYzAv+AkNJIrJiLkegEDggphf2vx96zIiR7ERgC6XStDdTtMUzh29zasoVdYPaj
oUKsMkrid0uqk7mhsTiZ9xDYe+NFaIUDQDDt3AkgFxEw4L0Rv6gJG/MMifayJIMM
xJnbxncUt0tHVLiHBg5xN35U1Ks31wU4QP2wqt7AanOnECtRqxmH7EuvP9hwaqnf
mrv/vBFEAW0rxn65gsCwGUjxLpK/Z07mBZd8GCT0835+Wpr8d52tY3381s2if4WX
rFwfw0PSB3LV7VJvBhps3SFS38w7h6j5didoFIGdRyT6OVUcbtWox9bTHKpTC2Lr
Yzrunt6zzP3ljsqBxPXhREQBpK+WjPdgngOQqARpluG16Ci3vjhOGap6AalxrMem
J5A8VZlVvfApgULjhdSf7YUw18mXYO3x1hBIQQTQhJm0FVooaDfW8K00ptIouilB
Op58NQ00UhmW3t6n86nYhxEqQmIRlzyT1GQkC2HorvFUWiBVWAgZ1oyd4uhQJ4u5
KRVRdPRontcX3CHB713T+aimlNYt3pwwteDdluz+7czlhQgNtidh2bWCvRO2/nQj
rFyS/ZZ3g0aw++TqhzJwWRDnMWsNcbBDAov14VkcDvHmUnVP9E8yTDt+hD2zk6tn
w1K2cht+vqqDsJSycfem+Bw4tt+Wa0NNTyhj3eZ7Y1T+UGpmM/hcRM0qotPbx8KT
4B7fXscyxNKy0NNJwOTX6rqF+zFx8W54BLA9/QAX/+UbPnS/5LxNaiwqi0uHI/HN
ZC+VRUFnSxniL89ElofZlSTsMcLMSicZ0YrRHdr77fFvwPDmjMGmmZdjLyfhBtgO
R5ndLwkA/CaU7T1kfgJDJh8oeXbxSdEZIEv1jH/lvwuqOi/dcp5ctOg6PcaaFYA0
vAHo9wBsh2QHZ1ehBbcRGpH5jOk3psd+MxyU8/TqH2Fwp2mattNjzyFSBrs1ndLE
UeaVy7aXHCzlNxNVakQ5t3TXDBDRCgViEr3jrdEFwD+5APExZu8vZdNCvSoQ+nAp
SCGnTNo8blGhjcEE5u/OdJrA73+Jma0eIErWXJRuXtfiZ8edOcZvkuvC1CC/tk71
vILqeMq4Dp0w+7OAxgKuLCo7Po0Oll3+bFDkVN6tCXX/xnZ4AJVXvZXcCoCZ3Eka
5hn2lAwCEmbYqTVXJAAjn9Dc5bo9aEO23lPaK0+FV+cPpq2aogY4x4Smm1cifwS7
DMeNEbMLkUIj/imYkI/3dMKqDsxvzKY6xbOXbOWRIEcZw1LOMK3YAHsehlFQ/XeO
psMHHsmPUygG+e7OCki7bwGwF1a9wHxtnNV9mOpemj68ncIxQ7KtkkHPHdSpNZWF
kVxX0hw5o6puhMoEkirhCOPNtbgT4s0NMIa9wPXyyh/hhPvgGeS1GIkobdXIWfUm
XhNYyx+b9vpbjAYUOz823AYlstdGkEkzmy5GC7WcU55+WskHRIJZLF0/6YU5qSrL
OI7EWlx8phKypZYLvouFs0eMPVYrGlBykAiNNaJYz+r5HBoA605vFF9Hb97fkcbJ
3uA9mAza+/X482nbJhbEKSnXbX3QzJ1X7HUr8IVtaa8soP2cKUs/h8ZsXuKPuiBV
6mYpRJ6yjRam1dxCCSMSDbaxoFWVJ0WJpO++OPka/KSVRH8NUvreunMNf5dt3pZR
lLIz+GFw//8vBVeIXR3Glf2awymcn90xktYmqMP00LMLv0jKBWDu29Y1rjPo8H4b
5y+NkESiLSMSJVERtpVyYhReyJJ9L9AK+ygEF6sgS0LnkfbHbQQYQU5WLAMjLuUd
IhBdh6P6umn2x2o7gjH7hA8ai3ZunHBzpxYgYJbX2oAi6Yjb0p5Mwaqd/roH7toP
+RxC248V+iu0tlAscT8aFTb3wSWYiDEPwzLBW0BEFkKqia5Ac/DrNOEA6w7jj58z
QkwFRS9Iac2LKJHcPiQCQ4MUFpRSayod2udCYp0k0aaskHkAHhzz3cN3yhbLYWYd
Fncl3ITGPHbfcIux/YK2QGqVCLGMER0i/Yygv34GwP5rvKA9eJHaHNZy/3K+ViTs
E+T8u1cILln5QJ9OTVaOSP2lYJbtuu+5moHcTuzIly2Zt+FNdshJnBKhFRhWsrFO
908UXuQTviiN6C8OcGgKfzyeMaLC1s4fet/VlG7Ne2fnlZHHgTd8kv1zqp8JZZUF
GMW83XonZ7RgmftIT0CiJ+g1F7EFcxy5WNGGpiGpaeXXG+1LE14Un9OF4knTLb0S
TTmFu1hoo51fAw67ElB3zKxVOaQ2GVEz9bZiYfLs0cjeXxSagaj+1vWDpI3B2KPW
u9UxGHzDdEU4YNbhfoaLRiXJZrXs0L3Ix3I+pzpB3ExLqb1MhBnpqWkXEFWPf24W
auvWz0vCEEMKlydIRe5esfDsCv9T1MvrKn8uedrvusHK3e8zoEDfbwlHB3y48LWL
5MSWk2zzBTF5cNRHX7fCkO85C3AOG4GpLZwiF7x7cIZgReCBDrCTKLf/waIsdOQV
VGnrRrQtwJiGpRRp4K0sscLp9eTby+vNOa0iLF5HBnwCxiQ2+4RlyaGS45UpRBNk
axvMFxM3dK4SI5y+bTxC1eeCyJQn0nQGrristQ0Wf3h9QFF8h10s80FPmUoc329Y
9ul+223AQPik60mUVQhwDXYobCnj0hoFuWaQzkVAyLnNsQhWSBPK+kQWdlKO93iR
5448PVzN1xNzKXGzgJDvffSP2IcNtjxVo9swoqpVdv6KAULeZ10O3KV0KzTWSad7
RlreLYBRFjWr9q8m16FjCiDStNXGVY+R+RTWhBfB4zb8evktHiJdWpwguA2F/8sG
Ldb4bI09IHGK33QW67sReEWmz31u+Ilfhq1gsly4Dzx2V1BDlYNePyXztwTFvJ2Z
ScisCYO65vGG1oP+jJQ2TmhleNuIaU7FWDBN47ycgEYtxHwAuHWeMjBdMUPok+QP
n22i2MFaqrrgaEXNf+rWAxozkYOOeCs5Ga81yejasRh6g8yDdO1YzUY6syyXYUNw
Au29FECrz06oOtlibTO3YyYfov2BUKX5e6JAYnqVwoBm3OYC70WLYxDp1Kws3hKh
IZSUxoxpqAGVYYqlPQSnTTPjX3x2S491Nc0Xymaug/eCk5pRSwFrwDbAJTf5pcJ0
S6v2W18DOZZnHkUWODbszsPLnv5XPJvuLnhaBF9vEtZJ7cd2AFuaZNvPA5/RVXv5
57W8O9dPUkeJuJspJCP2tbamRULcwCn1XFX2YuXcyX9AMh6TMvG8lB9j6xL4Osvu
ye4HWyB3tsnWbzq9FKnxrxWAHipwPKTqWv9hQw3NnN7O0zHks71p9XxC8ItO/daQ
z/sEHcoCOGXGGF98bS0p+RtCqwQ3y52gfOiCD5eh55Kss/W8+Z4agnj+mh2o48S3
FnbWttO9JECQSkMWdXlk1qN6KebQjT+BzLSh3cFVEXtk2BOhczc9WvFFAZF3nVze
NK36amI9Pfe2Wmqeta4q16dAmn5ii8Pa+RwQQxrMNmJma4u4E5a97hg+BeeorHAk
LFXkr6KbzpOjS4mzG4AyBGXVZMunS6igUBHDq9FuHnlDT8SpQNxMq+Sn3l+ONKNK
FGRI8ddzW9BY32dgTcozaxq0/UM2xNTmbJ4G4JY60Nd16Vw8LrB3B0dXi1KjLdsm
Wq+l2V6eUytbmkfh1x24qng6hwRJ0Z5fUk05ialWWwiK86u/IGtYpW0snyEMPpUF
pJDFT8SY18OK2QvxOWQyGVQKHGO3OVlcFRCOAbIWH8DvvxD81ymVOVUVwK/znUkt
jaZ6A5QmIBWeqtM0t8TLNab+SW1UeRl12rUGip20k4pPPoq7+Rgq9rRFs4qvC7nw
BrbxBPGCKjZxALERq1LdiDRZicDzEPLDAq+ukRilW9Fmt1jTcFvjmLm8Wjz1c/Nf
x2YwwGUbxUpvKlmkF1cx3+LmnkQU6YKrI9gXuJte68QSaJOW8GjJTJ4J13x16+Mk
lbmcXaXFSeUbeSDXGZDyrRdnqZeJVQriqDX9vl35lfIZa2Z+3riejOfSdA0iOt60
bW8o9To6tBbF327dZTPvSYj3l5BN9WwZu7Ci5I1hw/gDCg+L2eSMs/Jhaiq4iYfU
LR+2bMupdigpkinOwa8dagnJO3spBRxrbcoVM1u6i1XnRn234vt29vDDKQb6VqtX
TJ5pvbhRLUjEm91Fm83Re88p/XRQm+qtkbXaPQ9olS/H1anuOkv536quSpnLurBb
P4hyvKTlwBFYRjEZ8TZpIcFvmXz/0S0Y+Dv6+oZh7MiD3CCRkx7D6QnEUMfrJRgH
R6T8uQflTIZdQ4CNv7qWZakcW6Glfqqe+8F/huEcjgTg3eXvduOZIBd6qMtB3b0M
wvhY9gJTO85mQPM0JSK1h5lIaKrg9TAUhsW1w2XvnjCWkIIgfW7IGzWVd+VzO6c7
SBWRfBk6Il7w0xN7KDppUY2RFOnO46VpNAGBWsxqVFCBnoDz1Z+y8iFVKOsHEv6R
HmktbTEf/HLHtTU0ASD/f4UZ+6l65n0ANlImy4niG1ig5r+XsApOQXgI9XAslqIo
eFTtRvw3OJLR+bdAPS8aHoD3Tyr0DHunDzAvV4Brkkoe6MctHw349j5p4AQCSR4v
3Dak/XAbG2ETRuQexLeZITUVlXu9RjzqhtKnp5oRJjfvcri97lTNgIkLlQQ/MS7+
icRhEfZr1kmAGZj8+L3BRgx3zQgUwqQ2OP9Gh6e5JVpmNzoyzdl6FZ6f3I2bI8S3
yLwLdS7KAlF8IG/LOeAU1qLhwtPXjX3G6TEKmLSos2b8I2e2o6Z02iFXMEIcC6dE
IXg/8LrLNKeyTw9X0wgVrPUZwtvpGVmBG8vuF2OHs4fPunHS8Wh9GuaLbeF3Q9s4
X9OH/K2iXgEvIQflajUEr+bUooZIwDkN6qzTyyx0ednteRshZtlvc4HxXhP7LMcL
/In6m4NtMy7Y42Nhzf9LlLhTQxQGldUoUmi4vyslsqO7mvS9tnSsDFfLAg0AGtKP
Wm04JsMFyIa0lhanFpaOcWBGsYEW4fe/BfYbYil+cDCcq2Req3sVIu0uvS4C2Mzs
Hm2+L2pUn7xP7ZmC3ux0T6lbiXdJ0AzkFjqzb8xVUFTUq1Bqw6XCvfIv2I0DKhSi
v31wio24SgxZ4GxDI9FDJF2oJwSw3bde+NF8148sdKzjMxzAjQVbpV4lwVrzxzQ0
1iiFa/CId2C7F9Qm6WE0j3+3y+zT44gOWgVQoLpgFgF/B/1oI+x8FA0inokYi9G9
XWRWwNansVXdGNltzHLnxCipEJ1tFib4fumtQz+WhFq6MAf/N2upzZ7osAGF8xem
28P1IipVG9u00Ddff0EWqDVgw9sNl4j8C5Qlbj5oO4/hWtIbGjcYhz0zjMW2R+fu
2XQyWuKyBP3vtSRfxqJKQUPM3UmZo3LNo/n7fcz4Sx6NhnOHd9jroIPluDn8yHKv
Owc5bKV82sM2DpxYhc6yAvpHBUOMiHGAGLUWu/XD5TmsXzsZ4qoIl7Ihaq00wM68
fhBW61HUTxa5jLIaHVxr7guJ+Nu7NVRCdjSp7ST7o8rZYzLUodkCHL+IimZwEl0R
6i63VUVQjd4KEfHLM+oCfoH6m/oCzPXx0TRW00AhgJ+JTpFmflIUGgu3qhfqJ5m3
079AbnNUONfpVtKvp8pX0zah/B8SxCJIFxsvoR8+GQ2B5y6L2M5KOW/e6Q4boMAQ
y1Nf6jXBYrD9OfAgKht+eyXrDyQ51CfSmUiRt7Ofr4PkHGhIxeekgvNBGRIE7Oai
5FLxuHDqfNADZbTS0LeBkCfGmN5+Z0AwjH0WjcQtC2BjmXtx8lWLmtfRDJO9Yiv+
bBrrIYigRjEfGGx3iFAsdmwQPVBo2t9rpoQVv6r+uiBaxqhdnXflho1BIzutbJ2n
VrzZFSMFK9uj/r0wTwV19dyQ7f1/1U2PA5EllgU95CN+i8KgVbjmcn0z+9eCUZDJ
cQ0xtypqX/osAbripbOjfADRuyLMf5kPvQIK21eAFMI1t/9rFuO7qv5iQWrkX1P3
JUaVXdvq3TsEaa8EO31MO33MC86GWYyN5BrN2TkCG2P8uUzfLi6Re6DeP+rpRkQn
vfi97JsFY+Lb56jpMkCmefVdVOqFBUdw1P/4Hw1yU3OvAm9pe+Xi8WOXTg8MQD+f
kdUVxiqJ96VZy4rGFqB79DsgujukHz2G9qbT1zUR5rcjz+3SGGq9lS/t+vJvoowP
1HemtIbRDFW/b1yP2bfSaOEYqHMqLd6kvS4L3XerBqFa6MlJneu9oSZIG8JNZPVv
SRKp7b/pUW7/+u4ibdS+MDFjd+kkXdYm9eHR6/Ta8OSOZJeBBoAQbOW7cvp6DqNX
EguRMMgnevA9/Pjq5FnApIh5XEMpqSXKsAbXTRJ+QtYYvrolozjae7Yt7LqYdM9k
NmsdRqyWujKkxpe6m+kK10ci7jQfGkmOSKLfE6e88bjlOLXj11MxiUPcQ57fNMkF
sGgv5ybIcVILVcDdVkiQDauh+/lmNogC5dDRXG+CkT0msVEylbTWFktJvSBPjgox
jdlwfh2FGgvaXA4sfs8sQaPLUzpL5z/3O8WE665Hcyu0RAlDLNIwvWbhuHoA72aV
dfvZNmdlXSJL+5IalVr3euj2vXmHAfqR0AkuYlCMAsbUYxduKcHxXeWjIvDafYwr
69JHnWds+dOOXHp7cNOcCATI6mgjXq2ATiEWKqAgL1TPwfe/Xmug68FPZOfrnenN
YszB6h+egEfoSB8XD8nTvzVKvynqChmwr8eDv0vESgR+VLK2kRhcaIIA5YI84swY
2ZUaZMkrGXa1MFq1d/Rdk6IpKE8+KfW7S+nWqVwOuJzkRECK8D5NmTp3AUdPmBG2
3ppGgzp5raeIpRMYSWfiQt+NO6BfkxL8S7RUoUlOaqiAogRtefudqzsIIRaHJu5+
ag5DNjKQz93hupCDRxGYSPu3xmc9Gydq/FSpPM5KVxNLKoDZVhGqi5KtycnAI1Hb
yiEbtDRAwE1bbrxgjVX3XXAm4+WM1kSzwXAzoUghj7hL1Ra+LgPABmqCXbEB9Bgf
usg+ClRo9NIg9Jpc4ciFh3KJl4x4N9n1mRyLAZzLHnOTkNxBkxzlA2l6njQdRsbi
EGWolWIm1DS7TEXsmkKNkY2EgS2Wt3Hsjdg+PYLvnfMyksh5BKaoB1y5cdPhPNsi
9AqD5Ub6IOI9p7fxVNgepkRlwQMU4n0bLIdNKPt0uOEE8KXAiiitjuqI4WYmrJ8X
hJmhV5WYWG6Ti0q6QIPSSk6tEUlWSvZCH2M/R49jew6MSjbRoW7wrB2DpFzvWcB4
FsAEdV25dZOmGxiFvYQfHqCy5YxeN+EV78KvWVnJx21/I5TPfRfkKvPBjgTCqQTi
GLCDBGjrrhHtKn51SdiW4+OpKVcukH4mK4MuOW7rSzADS6SN8A8Xvt4N624RA2wN
vwWYyENeJlp4CGw9GVOr0g117HG14Q4DpZu8b17Bd2g8qKHrTH7DWyC8w4YYD55g
fWVk3IYSMUh3fwHHyiOmzUMzF8dLczhvRjYdqPfFq+Uz90OhJGycuRvBQD5bYsB6
C2dBzLBNZpJPqLeAueYF99kjgj43bTXZziGCZZPf+dUNG0BIv2iqmMCth2Vqf/rr
QLk703Oa6Lb+lRzXJhaVTjYdowu1ecAO7NJAbKb/G09DOnkYzQg7tLp3WMo75gvm
oyAns417mf4OeImIo54VwmLd28ew5AZWuMLKzalVOA61B0PWimzn1UyKlp2H+gRQ
qlmrpYKfcbgBlapxgLnipRXnJLlt/v5LAkg+tdEBPXfzKULM5q7G7Y+K+kxdYhCy
mbjpwUI3XGSOaD9wlBH6+mw9IqHEJTenkloYdReJ6sta0DLka/tJdfSvRZzDCHTY
4nJlFt/Kpj7mim174KQXKdTwlRYgKznSevNZXmVDXCYR2G5jwjP8+f7bopxyJuWQ
TMH8mtUpHoOUKRVdupi9ibXEpZDRchQD+mXqna2HOXdssU//WAAwMEVGitY6M5TK
/mGzwV+rQirwJzsbslnBVTVsN0TvK11a1bV/lnPLI6mgDc+wuqLU39UvNoyR2Dli
VZSlgKlg0uXzhz84EtOPZQVYjUhjsFtXWJJb9oReCS4g4pbvEd/wDr9rzWPBnWcL
h7A3DnNhQEMqZ7jbpP8mXWRzZ8YCQYzrKqZXprapJZ0W5jST2TWK3WQ7S6SVRrhS
1WWsh3XwQiP+9ov8/aCmLuTfcHTqoNIqcz3kQwg93gWDNy6VRpK+jLY2M3ERgBoC
+1Qiav2AAsutFGWk4F+xsIBDOtmpuzd+GfbCowKFMq3N4/ZJtMg/V74dD7JTWL1y
gRc2lCwTFrkJurMbzq7qHrQBGIm6C2nSouKzai8P6OxR6yKP5kRJCDBb/AVqEotx
KWW8oENdejFZp0dPrXB229bhadDS6xrZB+Bp1JrqvurNPm8Xw1rk/T7UwbONsb7c
FvBf7xTOXE5kn9u1Dlqx+wOHGe7qCXJlYqYgMAq/ic2f/F5exW6ifv6f4EeJklNH
YKrjAievI36wuTuFpOqhjc3TV+rTodiyW6XjSDDqz8xTI2l/o7FXZFhmV6MOpOtj
f4qyGGVgxGnwVo628TaW1GKoa2Zp/EPUHgISyYJ3Mz92Mh5sVHftycBsv56WSEei
0dsGbKhdBVTWNBLErzGT9O3BLleQQD8P5XhUcXnK2hKIAziASDxju3NHku4li0TV
kAD2N0rlxQ5yejTqS0PlDTnu4Llb/nq6VzB1+OCLkNdAM/iWuzJWLkofQQuvuHIt
ozQCC6T6Bh2wu6GJHb58zA3S7+ZBxwihdfqPfhfMZT+jHA1/SU6DCsn7J77EfTbq
iceu0NTLMNYgyWskfHDN63lsd+uadd97sBMEmm9pW0ZcjJ90JdQPCDs/v89aX1NM
bc1/biPXOWSQlvTbj454o9xv29NhAHk9Y0CZM9aQ0qy1k1MRbBzlc3uCAqQpG/ts
boGN7QdAwqlg3cJFdDbRM+dxgEeXA6bhH4cj/bKcb9Mv7vKuLtpdLayZ8EV60Wdc
zAAnOv84Ldh+GcLYHqo8bde3Np/6nXAVg7mtpFy+0k8Yj7knssrFun9EfSix8YKP
C/Kl3/sC1hVEkmQyrTGUruSuTBDC78P3XWqZFytKBvKBwaqoYzdwkiSTaMENKu78
l5MfKwSYHaXVXE/ghHKjXjdC78rwjLvglNKhgqIvA4911jMlAhHeNBOT3MPR+l8U
0nDDNuNTuSHmk/BBfUrQY9vAR4fM95rJIR4guG7qsVaUAF/zsDrvEj9HlfTOrvHM
U3uT/cR1FwykrmwVbgFpEI9iNAHwB+Eicqi+fx0GpfyAWIFPvFXigr4LB9j2pHzl
qFhCF6QvCQu0TEnhXR3qF7tyxbJArFEctDnpSwdQN0VERpxY2x4LYZ42sMkYs7WS
WiIOFUbflG7vzeIQYkPcAenrhCvX40QTf19GXzmk679hXgvuejHpTpk3jIOBr9fV
+8agvghmvp0wd5aum4NJkW+R1l4hoTx8UEBbvLtq/0k1/OUFM+bnf1qFeICF1H80
tFu5qDnS1zaMYXq40SA4OlibZKhhedHyxvkLXPGUwFKNrk0V0IQqtz/hR8Wf4yKQ
OtbjQZ/OylvNd14DyjC3ywitKCAlXz7hx3TsFQs77mj4xAdnWL0lXNjzdqGLsG7e
IjZoIYURj6Dk9MWxwQHT2C9jAMTznDxcV9SPkeqYfHvp0Cn0weQ81WH1Clkkr4za
MDHgbYeOEnFiDmQFZ+eKzxNBGdQZ10k3FqBmIt9dTwv+9LJPnlWnjRbSvCyf1Spl
Kl+bNNv9L/OyGxNQLaE5J1cbE7nmY6UXaGK9LVlSiJXLlpYMh5+jVai7gqHsnGQv
Gyu1z37ZIdA1qBa7huL6Unj/p9arFL0ZRg1IJOeDp5XZRC+c7EhdHNjKwGf2KNmv
4ishVpXljQYo41BBgjepWjTFt68wzFAoHL9RbtncseFhNnHZqPk1B5Albt+2KRY7
VmqY+P/uPiTpo9cjblR5oi1d3FqiVa28aJWesUgYAlni3Bz7h7aHtN3N5XdGGQXr
7An4L93ZXf4ShcxhD0wYFdSICIGOig2FSllVvpLI2q2+0HwBPHBzDQ+DndNcYQgy
ciUCIb97LNbPD7JoDweb9WZ94FT4muHFhXsXzFE4FCsb4qvB4zOjUpyYAzZJGB3D
pUQUuZrVM2V/HLCOkUyJy5x6jxs7E2E9pTIylZMNFcoLXSEz8gURaZQ6IDvk+fil
bPLgWZgYGfj+cXJDBHLnWVcVl2WzbZAejH/79cpvNHHVlsRVANIBYu39mexWJn2J
yIa6CPuOI3azltv8TuGNwr8hC3oCNWf7W8mUUjxAXl1/L1zHVmTNRmAWL87BCXXH
6hfTQ+spm6Lyw04Cgw3zKArCSGTZZcn9J+JrUuItAOmxlk27xuEQ7R8HSjFV+4q2
e+XxiSf1/R0HUmzwpXNM9FuUJt/UDmlfC3Ga6svrYaO+0P/gJq8ahupDiEudB5sd
IsNzhZugz5WHDQxNa9UmeuP8nKvHXZeLtHcr88FX5aimc4bl8YBOjCvYAtE7FOMG
JotEeW12l7q/3ZAtdA5Dtoqc8u5xG2+iJLXpM628G6bXrFvN98J6xS4t+G7yLq0R
JCK0aMOUOw2hNUu536WpCE+k49CBy/a5NJRf+ftaD/4Ia061KEzRIZGwG6Efohl2
kLutoJMWh5nmduf0OqHrBOHuxTKl0MyxEUYhugH0WuZQHJydJgGiuTXlDfJ5ngJj
hC+P2kAmkK1VOBI0+5A0atwFvLL1s+Z1GCsMQ17ugnKg99yI41I+WWRrE+shGcGI
QPJ9Ae0eo8JREVp48HJkzbpa5PMrVzub/Y8X/dY4xySNX6es9tPSvatgFWR0y4xo
JY2qj+NrBiKwevtt2RTyaoE6TXC+A6Omf+q3hFvjS6Ua4zrBpf0CBiQKfURe+13a
VNoOoXLH96xM+Gdg/47GwYZ/Ve2X5mrji43mTtWwRk5I8VbmoG85vNttaCmuvPrs
GHj3VaSl2CcIMLYR/Z+v2aPvx8uEw0tp4ywo6L7DEIDRHIcebTeS+LbzXG+CJ2dx
hvZhjbPBwlqDNCcT1Pj6DeRIPBLMJq8T5zU/hUkb79+bXZdYhmTccQZUd3yUaUFu
FrtwLgEgDSQ6hlaz/OceSQLmb7FJKg9OiX3Ku19m0HxVG2MvCXy5GjR3E1FUZnwL
0GMiUXlZegKN/+nUAhHOknFcqqY0YUnur/PnWI29DwWmEOxshhjdJfIXkdcx5NQV
gFIpjNXM2FsCWPyRu7KaTVWcr8p/Q90WAVJqh1MIDUHKKI0ml4PLkR8TskN9ZFKI
yGro9u2JYV6jVebkEEgt84AGko/J6vm1d1rhjPcmVnt+ixlZJCFNqez/IW1cs5s3
93neUMpBceKwQq5EQJALHG8VgyAjgjK6xKQOGBohtDppKfM0+ZEm36sOQmVoBUqU
2lx6HQnQZHYrU6WAPrrUZ6J23DQ2gr8tlQrcqfUPYqXQrBdco1H0U2UDGKhUiDEJ
muLUdhqYHaoZLMTPxZ6oj9I67j0xrs1H5rpWfvO7q9oj+kUppmIK5d8zLElZ2OXq
N7dAtjTMTJdx9oH+WAYcBxSjxhK65p6En1bfbmuNSCwI7JLYWrfQS0HqpXovUPPC
hLmsPBo7HEH51XIMm2gjqH20IJtSQ7yq76HtQ+Yq45KYRAmNtQ3cVzYt/OlErbTB
hJk3X+soxP60E1e1zakUCuRWTyqqeLMH3wj3SKazGs1dGTYUrAcgXPzmWdMFYQrt
VUeVhhjDQQoftFropD8l2CJ6xIoackYQ+h591xh3LA4yTpD3/vTlHjg21NPOGQgD
VDKOhj7esOyg8aesIaHNlOXMmZZcx+BPZ4LI+9Zt/TNQjBYPu5vljFAjsJrUBjX8
ZccjdXGnpZXLwPL0yA+NcnCzjzur2eR4hzHTmDdZG/jGjIY+3TKzUgplHNLdGZxl
kvjW/SU5jQ7DKVXs6si0ca7OpUZZNw49nxeGHqyhr3hu+k3fy/GMkHFORO4xRf/P
SDavfHZuc/izjfucknL2zu2e7vhZk/xOv6UUcr6gihSzlYIPZWRbbC6SAX+K8lDq
84fBSfnnzjC0L9uZiMV0nHCkykejDm1FsBpCn/dPK3bFJ/vM/vPYDT7BVmjL7m5T
ADI4eTzdIO7GVsaGlfQv8yMpl0BfZg2vddQbB+2goV7dLsmfcsuXOibSYmg8X2s1
2x+QZFozeF1hIJbUvUl4z9ZkaZN5AALB5R/xBOsb/9BMuOnyDLkTYca0TTs7ogPt
UbP5X9qTm2oYFQ/tjm6GaxEMFKB7xJO79/uiVAzjHgpf2uwuAkSMC/2gh3/iR/E/
a8m69FbKX0tMwsgoN/K+4/gXmm/AdgxsNKc5xZfzUJ/5vdqIG0KjQvv+U2jvNacf
Gd2rSYfifyhnqcxQBFcRTmuDjQFszddY9b+MbZTxan/j6AcZK3h8o4R5eK3r49Ek
Ncv9O1azo/FTezOtpF2qmx0sxcSLrlIdYAs8UdhwMNyRMa71I/c+P029WC29fzgL
asD+ohBTm53sVEZM1yOXtrTTCM0LAdO8TQQ+zCH877mdhldbr0bF4Dtxe7ZTdaYd
gilt3aqYd/l/zOIpZs+LP1ke2fuETB2maqetlWXnK2MOedyXgXqql2U9DpC8Itro
rkRjAHKSf9zO44YfHTW1AfNNhZh1acamWzs6CcY8lM3G6GgzcdAT0W7W/0qzcNTW
XcYKtpPbvwOJTt1/MiLU0HBA2iCFO7jFPXQhb85YhgtfkFpHHjDlQcA6cGRUYl/1
+oMxG6Li1+/F2c1lkrQNZ9dgFaP6Da64l3lqLHME6FMQvC0K47MSKVdJJw9DAaBG
9P03JG63iHQh4joUCSfNDoF4Z/3LN3wBFjXo0O9oOVF0MsSAIkqNS52C2xcKLXoG
CN+OdV/WutyemOFak3cqknBw9Dc57CRzHV7+G8RrhkEbtkUi8vv17NTpBi4phPVX
Kn4xnIpdNlIGAoJfXlbXsMUAKn3fXk73CNQDsLmpUE4arkmRuBBImjgrboH2Inst
yTdDdZbwRNubudXhsE5XGbgdDWyx+u2g5dfJaK42I7dlUTYD0FRsCPlvCqukc3a3
e9iPVaG+vTtXAsExJddrEdzmOBukWFTFlVoxmOK/OKIwFDesGD3SRssIISi6CCXe
WQHCcKlrWpkSx8WFDUgqU4Dps6kz7TGysopO4dmRralLFnt5WPuOrybegUDzrdPi
WDimawhCvk03bHF4GGqunpAsX4CPKRVYxFAF6b5VrjRaAVX6qZbbq4+qk/7kBzUz
U3fg8Ge92QU7JaTzMkCQbWLnyNKX/OtS+a+K2hmQ8wSKmP9TOm4touHnYMIoay4T
c46HtXGuWI8U9G0k6Yynta/QERwpr/Q2PcORaN2/g6C5EiBnJVDWD5VgFPz2UHf9
4Oan7OR28mb9vHVqS+ZMC786L2dD+vWxJZoFX42OwIpAzGdM0tSQMvj+zbmgrJRu
9hXxxXnaxmKFeh09yfni0mg4p8Cuc/gbJwIoNdHjTg8s1QgsVVe/SCiFczgn48Lv
g6unPUM/4FvGcighzmTxTHBoctcf8GwFB28m9Dqjvu0KtWFhB43U58KoWKJelJM8
BW/9ctL1DSbXBBAuPe5A1SndXdDSSFHYeff1QmQYBflFtIHZN9Cn2bR71KgRMNLF
WewzaM9vg60vGYKQdaX6zEuANgBrpEtMhi+zHKEodYCREforQHz8xDMh/Z13h3a0
CPfO3eMFJpIkG6Vwj1uqtR6hQ22JAdOIT0sZCRlFYOxW7q+3/MKD35CybPSTeUWW
6JTTNX6Hh1o0ARcBcED+RV5akGyA7MwFgpPnSQd6xpSIn9yfuqR4A1YNrviPbboU
2lKSKG1jC/NW7rLIE4oPxe3GZrZO35P6xb9csqC/umcI9Fp1/QJO32+7nht8BwZU
yOoFUegEZms99Sc/rM/6GRFzgOSjXDB7B8mfGkqe/u7sfK+KyQF5RZ7d6KW5sXOx
jB6Bs9jBoli+dL/Q5fAnIRvJ6nnkHXHca6sVyFC07dyb+qMVy4nXIxVTy1b/puuw
018dlUUeLAM6+Qk+BARnvxVQUbcBqSTA81TYfNZVv4d273+8SQ7sxIgWjTeNT73o
qwqjFe2IZErXYJmNmQBr4vUQLxaMWKZZ80M6Gwf14DdJ5t6jfGMRiMEoH0BlfOFk
oZ1WdMRZpdDF84fbLvtZ8KmXMzKFo0PQ2mcZlzJD910MwMi5abZ/rjfH22K7xwlJ
SQp/BqaWxzF1ByzXyyCQ6Wdh7GgHVUKWkW1+pJXBeipCEaJiCbKKRdlq4uJSTrJ4
P0YFEuqJGUUUr0n9UY92Hn1KJvscVPaMb+Bs1qU7LW2bM0fcPBK2mW2CnpAdkb4A
/gG4tyBGBNE9WpRA+/zkkYhwYHS1qsFNEL0uv4AA2h5rJ+nASL1UAOpVssYdSFSA
4iDk2qnBcbt9UP6n8kBfdNlC8N10tKVLzeN9a9Xfi17WoqJ4u8DUSipulePZxXho
dJNiv6J3xNP48ovZN/tN1NaW7RWVQIAwXStqbZhW/R70bU3rtLsMDDL7wmTsoiS5
4LNYexexBuAaFkF0WZvpcPBXwfDzBEJoB+nLuxVH4gdIQtY1D4Zq/nzgDeJQZAkA
GobKhZAG0ebRGNl8ck+nsikvHaMWbCjwbJzPZ9Jy4PUzqWry7bKAAfcNSQP2mq6j
neg+RWWq45HM00UniVyJjzkLOZE7lsxP5ZpcYZUiyrUvbJLY0DeCoHSUoWnlKOWe
GY/8KH2KcdTwr9U1FGn78A8zYDFP2MfztE/v89iJcIS1dHhCi6/w+ARHk7GnXMF0
J8knx1Jy0E2Y59ILNhEvHMznZIV8wEczVfhehghSWSEMWXZmYxOfB/mQGv/C8mns
Ci4T4O+fLCI4PYqD7TdLiUvagtgWVsEjLTiJFY2qJGAsccAj3jzCVygIS48WBeE5
RVno/bMD2zDNu54/QjU85dUZYfn8KjKfIeADnWgiwvxFjEaB3L4ArdMxhCuLsILN
x/ZSLRTpJUH0Wvfxxh90g/3S63pDUdPjlKdue4y6KGzmA5xQB9vTK/OV/RF2OSwY
GrtbuHIqzmoyVlmxVUiufWmoZNplp96N+4uOziJMN0VPP2N8t4U0vM6NdEuROJ6I
RZLRkLPeZaVK2vERxF6M0+YXvt+2na2Lrplq+6NpiWAZQsEv6p35JiFYanGQ1uVf
Uv8J8gBE0yhu5bX81rNQy9S06QsbxqoNkzOa3kLDH/okJlwBWR1UKq7Sb42ZV1wH
Sky5avZvJHquPaxjg+Q+0tT4BEkV0LjZ1KonbU6mRog48veiVLAjFNHSy8zPSWVs
xg3SZ9+Lffe55PZGANmW+rW1PZ30AEHCOC60G433BcZnjg97z5ydPg+kTL+fAp7R
SYS4y/pYN4OGUtPkTRXq01/+iOWD31kvs4Gcu7BAcT97EWBsLhDUtL+XSdDY5RuN
x+jdPjoiR0Dz9Lms1IqxTz+LbH3sYUc/MOlRFItGz2wWdbaM5lesrsEJ2TOjnaSD
mhuC+IYbaxi2mxXVkFt8sVMZRTM/KPiDnUwdcu9gbcZLhgCNIwSn4PIRqrfQTUna
VBO6tMuyuUxNHrivUPndBYE9R3X4g2hW4p8EXdvUc5s9jP6JVKEsEesBhNNk5Ikt
VbG9Y9FErIEp53oQiBYRg7Sqwlmt9AU4NeYHg1fOsET2xHikPqjumIez18rz9l39
wyLdzohfjAb69iXLnhl1wuAZcxEQc/GOXyoNiRMkgCcSbvzUjcsk2ou+xasVtkDs
PcGlxVo8DIDWm3KnMutx22fiYUkyg+h5VZm35Dhg0Xcdjs+1yJALEazjfS6WWPGH
XwXc0jAMNm2KYqoThmJlTlXwmFCw5Z0EpX13Ajh+WeH+pbK9eX8MQXodSbWEX749
OvIow6c4Au1JZG0hOVvYytCbebW73cOOnGwaFtYwZlny2S5ugoA3gqO5w8kKpRl4
rT2Bpcb4K1oFcs8FS9Mc/CM6Hg02oYloiCP/SfdKZGuHjD0hRtdkOz5BGOTogctE
OUvPIKuZvXyxvQ9XqgxeKrvDluRsfHVQax+uVR7ZbmIFESSB8P6mNhStTxUGjjA2
dg1CpiodO5S8YWW3451tI3kztzr10NxyfzFaXooQZBFDM9ZgIaoeCZJOlVmBwBVH
zClyYKj1NKMJF88m44/cB8cRJt29wb6a8ujllTN9RN+VzUfAcYZbYu8XoveDEWjH
xxWfaAVCTrdAc7xs/mWcXJs/ECQJxm7WElHLC0dYYaeGy6893BcJx8JVa+lP5hJn
/8CiqnJZxnsBIJRuRzM2KRMKTgjJGnlnSIYn1sP87uoyMa0l7qSHue+eawiX3wJn
ixyPo3gJtCvBL0oavezNeY3s4MgYpcOo/e4FJrz5iUn+owVWE626FNGcncA7VF6U
GmqjdgmdgmQOEe7ZW6dZPsNHWW4OVtX1u3siBenltvYyJc8iEYY4FPKn5F4dEPyp
KdVjdoBD62/eHj00SKMzlrXiGL5fSI/ZsRYhXEaTPcvIM/zEdELz5u566WUy2qyZ
gJPn7pYWToY3CLarjVeWzHawm4C90V5Fq16h07V7KZ9Z8Xnr+bHATztpNkusJvtX
w6SwiyHUjnZ159Vd7lrb+gHuVoRXMlOAGIH79/4X8kNQgDp2ySea2n21mhg/+2cz
9wFSZcADPLmcN6DqP6pAd6Xb67Amc77uIfqF4NpYxs3T+rOBw2qlSwibvz87Qknr
TzcaMyge9LboZuNJq1+BK4a3zttng2QK8bgm618lpPIjv1yEfOiF/NOAGciqc0VU
8stwTs1LFzbDqy1CPRCPrp2A5lnXJKpq+zD6tSfTfodLrWnlOsqS5fgHCcenBt15
fiSfEeTYNFKysDRLUygJJfH6BJMjIExRCJbnPJxXV7FDFySVjH0lVNt3h2yWUDlz
QVMwuqNRzpSnRE4d19TnFVj+OAbMSXomneMmDv3uaE4RDkOPZiJH9EGRMCrVfzY7
ysW8RTNES3LlBvfJAwEYDBUDbikVYfWtjnkXGeB9MRxFhz5NuIsz89le+kGAgAFE
jTDmZ61k+dL30HUhvIEUeAHJeSj1rpNU7bowAtS3a9Ax+I0BXmBiUnjozXKfM550
rbQH+GbxFATQSHfsjj4VqPF0U9PubKlQrhtvTqc9n9Q17/kWTppfyJCgy3sOYwxA
oFGwY+CtxnZphYl6PWbe+tROWxzDH1phxM+RBiwpVjRjEbRYf1UbYqII57E6U1kn
l2SQDOA/Cm9Vvq1z9Kc1PjHOKWqCN/2Zo3PsI1HGUk1r5g81QE953kwhd76lX+pq
gTj4pxI28GCgjBF8cuHhEZ2clusUY7s6Tr+5oJLBJ0wlD/sPHxaaOjIEbcxl71k3
yiRSwmRvdZUVdiqCkHYThOoEiDeqdFzpRdGKdd8iYh9JISiFyB9HeyVLnvN+VY23
0w34cGZ6hH6UJUrS1PFfTUEgUIiOhHsxRxwk9h0U4IXhz1ShyniMAkZwjgED4RCT
Vnq36ORCjJk15CJryRdsIsgsg5QrjMY3t44dpdQXhiqtzqAGaFKj1XZw3RsgNSLt
QmO7iYe6jPR7gU4KkSvF9GhCcQzUdH5BDXt/fn+MiPn69vCJHGVfceM1O0BDmWce
IryTfQQgp8GO1wIggB//7OU25bR3Rk7Jv3k/Wl/xRxnDtrNazSVy0gzkLNdRJuIV
Q1IuSHeflzXX089F3cL+Elld9uBUzWNRVE//xKWH2OJrFtr8H7Lak8MztyuAj3kS
UKCblKgBzqpNtNkhq3I1zR0zSyEI2DFgplsjNJJcM3zK0iOWMsRPUCwDheIGG5Tx
Nu0dcr8LE8WYBDLT2NtljaAWqFT1M6QGTKSK+xVEdqj/DMIAFGDBULLx9wiUye08
jsKnCMyuq5SpzGfk7SJKC/AajlNSr1QOxySc9SstufSFWelxCbEHgBopwnJmwZmX
6GVVKwTpGRfGMv9TM45GjtQMwEtz/S/hion0FlIe729+QacwStEQ9w7OnNI4fhu+
jVvvV3WbT8ReomUIoBqT8TflPdiKJydnlBHeNZbbewXfOv/whv7I+JjWnQvXwdwD
pHoltYmecKneEqKtWGWuD+MXpgexGZpftxabJWLRERYnsyd0gx8pbEC5B72SbtDe
5YiCJar7/x2s5VP5GhETnl0yo48tbaA3/regjwCoUQ3v5Jg/cxuDA9LZB7+5j2or
HtuwaGpHxDTa9NONAl56Yi0s84borinznqclPCk5SfmEkXx9pVy613dHAdJiSsXa
qteg2NHNilDdPaPhiMiB7ppjG3epHshvCjwTfHogU5gydw9NWPRM2ADZrs37CweD
zmZ/K+iinH0EAmG1kXLefZO62nFzT0zsvmcvHZgJcV2RFEOAquyRCGuzPpoy98PY
VwvsLSgtdBpWma5rnRlbwykx3TpTFegf/E5VMtTckDJR7vrjICKL9eKZByAhvZv+
3yTdZU1kEvbmon4WXNWLeWsbuP+Qg/GsqMhZt9X0XL9MrC7ZcJymmeZogLqYk/xN
tCPUXCjs9W8Dc2VIBnPYj1vFaqSaXET5toiG9rZT/7CkjnczNEOh2NrWY1uZgkX3
NW+/hhIbK4A2b9rJjVKOEu79vfPIVTq86+MHyUYIvkXOIG8/e7Pkjb5T2MAShoE9
uH1w3Apuc6fx/skI46wp2ShR0H1ANkzqA5yZcxz5CGq9LF9jnjO1YTXy4k/aD1JD
rxAbhyMhaRE2yz1GO/GVPG6PJDZkSWYFn7gDbx6V5yLkG9Lnjy9nZQwcNMwIIitY
ZH0lVnmTiYGLz+AFv/BdRou4LIQcbHJwG3/Alv+1wMr9iMl9UwB/GN40uclG950b
H6wObszFhqn7tSddDu/ev0taZezuomcDxsvWYT7ijf+7sEGKHE4ScRD1leaGCOtg
KP7gCKDoOeiVM/+Ao/JG7pfHkP6qBupwn4Y6TYF8yQmwprwAtacThoMOjjUfFXN3
xKfCIz7LDFzxei/Q0hXexpCRnLK0xApjK6euL2q1lz3Uz4/w9yndnfSC637mPzlG
Ojll1GgM8Soub5+GnMct8xX4rcMMQSoDsjdxKDyj2HnnelpEIgWmG/tHl9adf9wA
zHDnXQHmax/k/B9e9/wwmvkkFe/GgOFlghy8lf0XZWwYZnfpQEKueJH/LY2H5gnb
dSjae3U+JMfuKkl+JfNrEA==
`protect end_protected