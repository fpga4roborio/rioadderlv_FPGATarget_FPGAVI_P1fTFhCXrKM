`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
ddtXksX2+yylW5zu6QL2Lhnb2d1sD00763mmSITNX595NcHTEkwn0zB1Dry37fOW
FufOhVzEJp80NC5qZ/+F0Vk7Ik02dIR0elf3clrjeJRK85K4e3Hoo4xn7YbFUIms
l/8VZSb14+JVGURjfswrIyCUotIzlzVYZ6gzoZwDXIi5gQIBf/gI+KxNXPaKV+PQ
Ufys/12rjO6aI/pPlqSm0hCvftmBcnezN2hk1UeXgOIuKZnogjOsf0iJVX2aOOWE
6pD/psybjbnsNB6kH5uFTA5frkzIzkzl5d9+YDm9OyC+k84E83I/7/j+rk4L2dah
QJOvksSIzN867/4Qt8qYTQ==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="MvBXkzurAa5VTw+1JJ70nePUfoQXBvZOku/SMmg4TwQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
oRtzZL4VJ4iwysPsC8SXYCzXS8Fw2gtZTOskLcDV+1B9Nzn1zTyNtlo6lNICRmmK
ZRVu2BmCc2G+fmzynYlNTnSa7C0Cuel6FYpxCBlOuk3OF2tzAmLAuDyOH3Z1Yjzk
a0aHuoCdIRKv7BrZCdALt03JeUmXKPdOmIlkVGFl8yw=
`protect rights_digest_method = "sha256"
`protect end_toolblock="Jn9CQpRhJt4rnzZPRk+dOpzAubz7omckX1MrFd4p81o="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 2960 )
`protect data_block
gD6l00tciPUa6pDNTk/+t0OO0nC/UTtBwLB41d4inuAUA3i/ALrNyoJVcBnAmEQW
ptbcNp5fxEUJjnOxnedyZEuEBxWRieZFQnkRdF269oNdXhZKOXD5LJut3mwZv4mt
PbMUDKFUcZOSzsBM4xcEzbBaKx49imNUdxOlBgNNbhxd3tJV+vMpfT4RN4qEI3dF
7j0JoxLMQIVTqYtT1333mXjt+UyRR097USEB/hYaf5XB/J3B2copbqOqsJgH0ftS
oKl7od1uQtnNoZHOecC3NxZT8VNGe3Bu1FtkPCT/lPJCs+ZQ3ZlbHpoLYBUa7p8b
dkNcStJPyLuS+RpcmQFEJP0It7QTnOLAo+7RyVmImecPAVoHntm7vqrQVrJdEd6s
ClzDY1/DUwkHtexWGbUApMZvCdH6p9HtIfCagDznJsLP5X5LPFZ9mzgibhfm+gok
vHh5ZVOa17BlFRpyVdMG0tEAfm/kLOQSjghu4qiF65t0WwD/HQzJ6frE9l/+fFmb
P6nshAitiOqseTBpEbu4xhEfxBvT9w7ANade9LubCGCK8AJCUVBLBwXvr67CVpAr
VtpX/c7MJCssV3DWAXkI3bH8HRG2Go02zMQ4SYjlxCuXKeS2IzUad1PXAEbLtYLe
mUdOSqB7RTTkLdsZx2Dcl5KTxGHs1mqoVZRASCC1AByas1KVyGQ0u8c3Ma/RGVs+
VTn/gZbFlACquSBqLerdzTgQ1Xr1JnS40cebC+/X6KhtadqUtyq1BUEHcF8V0oBD
AdzrrWldAkpda1hsIOpQ0aJc232s0UVxA3ZEMcgHuJOhcFPT2SBdCrPx+hEoz7sx
WpGGl4qMH7cbzEde5cuQiHglC+usMhETGknYTlSdAz5GBFcV7EPQyBy6TAyZd6l4
sM02x3w5SclZsf8Ze6whSVK+I6IfOypzPMVt8TLcozXqjKZ+zEDzkE5s1Bb9B8TZ
d3VKcBidvCDRkXwMza9dGZO8JLpjrtI2SWMQ7pHAyD8CAKQ+1A4GRodDOGtcuoV+
1HaXb7wLUgNfKVb2w2kjLjwOJeeJ2BvYW/xNx8junegpMbozowRL6WGGhK5tCvoM
r0oNYESOj1npEadu8KdAvhmA2EhHz4+ZIFR/290K+0WCrTXC4noM04AvNtYC73zL
z/5PckuF7hTjuOuUI+NUw84UMBCCFzcRuVv9BMfzs4z5CGImzzj6Xi/2vnjIcoA4
Vd3tPVtACxEjloqsftLGKLHCITK7zO8Cvo0QfjpL9UCbumXnQ3qYT62VwbqmiRUN
KqMTrRW/6irrAiLhS09YANRu3RCchJOAv8U5RqxAsBzIbaCft8CeqVYCvdnOoQIe
wAnw4JKPDUfP0i2KNlsy4qml9PrTL1PriP/SWVb/M8bu/zi2UilPTmKnlF3KWn3w
uc8zLUgQyJsoueOSBnuZJYBmfjr7kbvO+k0FN9KCn6JANGFwZckTfw5KDTPgJKNZ
RbuFW/zVi58gWtemzJzkNYZaOszmBtxXnYn9poNex/dniZbj6nLjdMVnOGD9Nj2/
QDRsmAD1STtGzHBNtrFU9LsTrcC043WeVvLl96vwSYqB/DJzulU07QO2IOHj4mVs
XcdVqFwGig4/kBPlQjNmZOSHr3ZE8eTgQ/zZn3y06amDPJHYgiAPUOxylxtxqmfu
dVULV+OU1Paj3MI+7EkuyHID3Y3GquACZdWax2C/NuURjAKq7Rn1bpqku4Xis0CU
a+0OaM2SCpgZVIorda8L3gyB5Rfh1ftI2hCWpG24qUGSyKiNVJo9NcVGCQFMb/kl
+nmImHUu9QuYf34LKC7gybhY/3RSYhcOVAfekuVx1SyecWru7nCbv604b6QfdN5Z
qRoFajtwGj0Gbn18HFeb3HrPDctQHBwC+gaQ9zcCUFVXSFlWZIFUoLEfhS1INFxF
81Vts6VL45MsX6pJCcriJM/kUxA+2KD1tX6zl8WqiHSYAQ4QIzuUl2XOwwqlUBJm
1n36jT476kgYZa4wJtahtl9mdAO1YrwWpcTOP5sjsFcwsRA4a0CcdzGHHPSRxOKb
JktnBGggICnRyg7qjZwBY9izicMzwWeQ6W07ixHv10e7dgEUs42ioaoPwKwixF4I
joqOAdtJOBwa0a88tEl/9TcclXuHgFQ6fD1hrCf4KBECahvMzEnwD0Y61qvA/qTY
+4JQCVATaTZxRrfi8MuL11+BUS4sfUk9hyEH51HRFjaObVbWbHiz2e34HO/L0TSK
2efhE84+a5I/pxgdV3qR0flXlGCCIlYLrxsKUBDbTH2XZ2WhRprSQO/4vGj9W+Vi
A8HXOR4fu8PFc3uP1m0JvYiRrL2GThQcKBMWDpp2tB2vMYt5bgqK2aoB6hhbflP3
QKNleNEzIbg88BhyGYNbRXGJZmQqX7wNim2CRezrYQLYoxXKahXuaJMhmgRFzCcS
QgPogUOEjg50AyOwFXXDAR0Hldn4PTxaYChoNVA3D6UsImDifNdSukR7uxYNbEK/
iINx9NUmhSNXrvVVq1BduDbuLd5k9VDPNq30vKn5azVWxIZfXfkxTh9W1ThEH/+D
IryBXbhUVoQoMQSQZjvo/LfTszK47wEvBknTJU4pNAfUTXVJrRFuxE2VIEHkB7co
uQILbAz7+kLeR6e9qisGN9N5C9mBIP5jBuvS6E+NUN9ZmQzVNCQ+zUNNo9o0gAdp
/hoZ3Jp63N23SeNKEvbzn9jpS0OZvvBfSbHM+Ty10duKp2ftP7tqG2eppnbdsAd9
zRdquTIRod007bnQAASCvKgEls2YTQzfwCnxhK1yhZ5Jkvh8fb32ojCRmW/+iRl0
Xax3VSMHBkRohtxW5NZEQ3jzsIjy253YO6Ceze9ZEYA9kaEBaGahspHIRBj1G/JU
kAJhd/P5mD/G2zt+zfpslI7fEyGU650CbbTXGOSjbtq0nkiTwqLBAGJT1noc8Jxh
j3gevsrROunItWCEbkLoCoh2yVGuCIrW2G+cfwRW6HWDoRf5W5QOSqWsZRureRYn
Ju9BDjBQHIMZFO/FpQI00i8FVIbmw538wz+mAC54y2j/hXChVFpZylTTYubYDFGd
y9EiE0ckmr1ZKRJDvO4KbgGcSO+IpazO1c91qRbGEzjD5nE4AoGW1LB7VoYVPBHy
8nkmFnoWdlRDuKzbEAmeSha98YNO7yWllN/baBeMpqk6irBmcba24TbwEA0FTN8M
M9FbSCd4mPhEkEoyTf9tE2MZ6DXkseg9zuLUvHfih3827KajXwF4maMTMTjKwkTS
vDbQHqccHlhgAYGFHuwvRwRqfliJsSuopIU9gAylckpOdgiOmgIF7/hXWrf/KhsE
PmZuEoj8GtMjeKvMOAu5f3TeLFePyjItS0oyotttytvxK8X0iyRO7UGvsW8QGaBQ
Otk+Mxa5sme+GEqv0roaS2S/RNDraZ+MT76v0LvbeOtr3gLdNdtIbSm/1wYHfHUO
pdlTinS5WyzfZ0TGKSWmaZXxJOQ1EneS1vgc3V5zv/7tY6Lb++gQi4TFapDBZOix
cHtoWTjZr2bKj5Nk8Dsknu7bLhUGs0MVNWTRmOFphh2igRVCH740Go6PuL+2mae4
BBS+szq/qd8rc4vuQYvVH6mS+ZSiEXXJA5ExqfjNK8OZk0GjclRYhP4HQacSATZu
Vv7Oif9AJMVbZdHcgJ1gt9oCtVBYFBtXbpl1BKISxuiNm77iED2mAxTnUWlpvCx0
skZHu/c0py2vfNDzfilicEnlGQRngPuJXRf0haolq0ZUpCRAoR/VsnC2ULltdzk5
aLTs3IBW5Uqr2S/l4o/IEyB6qOzytzvpgsQShjGvz9cax6CqsoWWqIiaaJ2K+99f
kn5/MoAhjYtRSAeSA2RjLR/esJ2gFyAh1L1GK4uf1KRjJ9FlrWL8m+BcTdUL34Cn
u4yUQMmcO/RfI1F8jmgP3A9n13haRkbbumyomviyIQg=
`protect end_protected