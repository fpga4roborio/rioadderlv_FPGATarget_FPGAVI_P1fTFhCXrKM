`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
ddtXksX2+yylW5zu6QL2Lhnb2d1sD00763mmSITNX595NcHTEkwn0zB1Dry37fOW
FufOhVzEJp80NC5qZ/+F0Vk7Ik02dIR0elf3clrjeJRK85K4e3Hoo4xn7YbFUIms
l/8VZSb14+JVGURjfswrIyCUotIzlzVYZ6gzoZwDXIi5gQIBf/gI+KxNXPaKV+PQ
Ufys/12rjO6aI/pPlqSm0hCvftmBcnezN2hk1UeXgOIuKZnogjOsf0iJVX2aOOWE
6pD/psybjbnsNB6kH5uFTA5frkzIzkzl5d9+YDm9OyC+k84E83I/7/j+rk4L2dah
QJOvksSIzN867/4Qt8qYTQ==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="MvBXkzurAa5VTw+1JJ70nePUfoQXBvZOku/SMmg4TwQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
oRtzZL4VJ4iwysPsC8SXYCzXS8Fw2gtZTOskLcDV+1B9Nzn1zTyNtlo6lNICRmmK
ZRVu2BmCc2G+fmzynYlNTnSa7C0Cuel6FYpxCBlOuk3OF2tzAmLAuDyOH3Z1Yjzk
a0aHuoCdIRKv7BrZCdALt03JeUmXKPdOmIlkVGFl8yw=
`protect rights_digest_method = "sha256"
`protect end_toolblock="Jn9CQpRhJt4rnzZPRk+dOpzAubz7omckX1MrFd4p81o="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 25856 )
`protect data_block
gD6l00tciPUa6pDNTk/+t0OO0nC/UTtBwLB41d4inuAUA3i/ALrNyoJVcBnAmEQW
ptbcNp5fxEUJjnOxnedyZEuEBxWRieZFQnkRdF269oMa52/CXJtY8Ewm3j83LKVO
mgEZaR9lnBAZHSPygHOPR4WjYqr88v3XHoujjyETw30EHZEz40utiFX8H1Fz/owh
r8THFhQhcphg7i+wGxLCO4wbOOs/bTTj1QEFpY6GspxagjLnFbmDK52V+dwexian
+gtTXyUWTPCcSk/1brC6lmMoEfN6hRgRReZN9CdDm2gij6fJRDvr6VK/QhsKPJ96
zA57G7fjM7QL1AU8o3Tds2f/a6xgx0ABdlvT318ZGYcW30UskUEFTwso1AAs6mS8
Bs4QK0pLBOqu8dYcbPCCsCq6UhGDiwiVHeud68SZ67r2Aztx2yK+IU8AJsEpW/a+
gyn5P2lfgNERlPRTR1jUsW1xHNesw82isG5mr6+iYgwo83dIp7ntxSc07DEyfKW/
bmKQtFjwIBBIxfuvjomLh+fQN4Cz/ZhlCFVkFTrMkD1CADNC7RbNhlEwkqEh0VHE
TbF9QDWXnzkil7JCb9GOnwaOInAusKOdfOmP3KwcgQYwtqMlGhiasltnUVFtuQpM
3r4OxLuCt5tcmiD497zFyXXX2pwXKCKUyDWH4HWJmMIwu5Zj5LvhG+eQiIDm/b7y
92vo1oXL/a6/6PWIqIx45XvD9alPNseiBScttBKA2ngK/mpDBV4YQZ3YwbUl/dUG
70rIVUa+xR93Dz03qlUmIDoG1iy99VQwiULRpf1BLv3Q6maTMZs1rxUAv2x/BUWy
Ofk4Wi1JqhDUq7V0Ae5fsnDQTppMEDOuAhqeMgwj7xxqsvShVekdIJoBNwYleV8O
fKBneZ9iCnwOlLj6vGLMxqNDYMVTga7uEKa0GMVEBbmOAXyWDnZCMQHj6cTUBOe+
fIUMHZ1pL6nd5Q1tUgGYwKKu2xSxP9D87/HzURYtBER7ovynNmG+dggdNY5HbrpG
ONmzK8k0Kvj0T/nx9G99jm4YVgaD34SxFXxF1Q+FS4AP5RmVtpOqgC+Aw4p1jLc2
MskTrNPGYSfX+pUMjgqGR+5WBxRMRtQkM8z+700hSlQxrZqyxV3oKyrNov7M08MZ
2IByu0+jur64LupAvMNpx1vC89e54JMuPyqjndsySK8bxzZ8hZBywAZTkHAUAbh3
GPLgKpETp+YWDXugu/Z83Q6ds+L6VDMPJaNa9uk4dqHI/8vWEoCNUTI8NLWpdSD0
ygryHAVLaD80BuS6cp1fVM986u6kosXCaUXVBICnYv6qDtajunJnUTV/VgoIiY1P
BiCi6mGO0tfXZfU5rgJWWdda9QCnUam108E300I/45ghyKpycdtqXkgX0grEqFJd
cyvgsTIbms0QgL/65wXXowwEjvmpmNQ/V5aJRpgkTXj4ajXhN6hSVd5ZopRXlXqH
WR5vssr8x3ARLDMhfSJ8t3QW+jAsXndy3EmXuXjYWloNC+6+nM+NqoZ94XCnEaDp
oB4jrLYX/IQXYwvL4mapkjbrznKym1o85sADMZ9W/jmpwux2mVbSH61/yQ0XEh6l
j2K6A5F/a01L9XVfxasBFs5mDxD4cnGPTwjp3zK+GYfoEXKOsczPtl3+ZoMsbxvy
mjqut56S+XKleIESBRFKFQR0mEa43MnnjdpnJAd8ikLV1hRA2B+pu14DgiBqHf7h
LEMfjBE9dDseY0q1E9zTBdl+OcsZEYN+bYNR8wVBc1xbL8VXu/v6YZ2ZxnED5ENL
z8Q07y7RUATCUgBgmV+kLo7/GEHmIii0CvuIOyQk1HhPAwqnlX+sRyAaOH+KU21n
TwZy9fnF0J7GmoYHC4xweNMRWvAhed68BAIJ93VNEYMtK8xsBFtvocp2AHx3Gs10
r4whi141vpBDywtphhTGW/3yWgvgxtYzraboW5rOwatPQfxZXCdWF+0K4fHJJwfn
ECVZyJQb3kTJ6TNzWnceCBeloBDHeRkEkmLAM02BOth6iBdWSCuMP4BVr204zoeT
lBF1vvNHLHydBDmAfPDx1RBkadACr5fWpmUHs5FfktyhxfjbellsOEHAZSnymcGE
6UQDsrQdpJUAjPAUwBKYn4U3YpWgyY07cw53EWkLa70jEUIoNZnV576kmMZxr1sz
z/UU4AkHQbD0clKh1PPvWEpSQgrIsbQ0LDmalgIYVBNOAWdMdrd+NWfTe6RdEf28
TAfl49w7K9u3l5qXmkrxb7Ndx6eRLRq6BegVEnk2dsMpIFhNunWXChT2PH0P2p3l
qcpVA7gfozMERPfKEJd/rM3oMQoaLvLm8ibbg6dPPl7FdiDmWa0DS5oxyAHEAs3y
XXa9ZSoWkKhNPifZLLDDmgZYwKMbuZG/zudB4twGjTvNMXSHxna+aH/GuDolwbic
v0HuXYBiTv8Ek6ahZmFD694mQENNLUhssoQ3Hp26Ur/yMmKaCuM2/+1sQ+WRI5kd
6n+YuhDVyNve7454sI3xgmKkBmOfGNy38+JcPsx+bLPs0qZm17xgsMwbXrTrXFKP
vIuavtGnjZdW1D87wQicX1KzSOaemzYVosGQyHqjj0i6w6670Wk1U4IgYaM6DuaO
gz9jmzPjRKxYPy0Iu3MCNZN7+jp6vonXOyUplYRFHCdRw14qzItwIJiNlXa8vTKo
1QoZJSUGi8aIkkx2Xk9I1yDYZTQeGWuch2fX+FI45HKuTbU7diuOEarqrWBTqyNV
Aybt7FFvgj5V2psdHGLRQ81yPsVz9ycjJrHQNMSQxTleTlqyMO8qg8YhqsdYEY1r
2S0a0z6bqNg+HyBEoJn4mXjVTnDQlphi2lbAHfw4yhrdw/3PCqZtz5+hXFVcTRNH
D+qtaKD41WQFo6g7YlZLsZs7jOaHpr5rmsjwNnl4VDXQnTUTteVPEDA+A5fxnRa5
DW0OhCfvMWZv8So+1qjkaAdHPfPHq6tsb9AqUp0XyqaIvxf8wyTIqvsEAF2f/iep
f7tEwHaif8B7VGq4AogsfMkG+zZGXYUKoUQdpDXvOs24ti8JRQoxZaSaR87HO9yG
X20uDemVEDC/5wQSONhPkzKsdWKVVYUW8m4Hbm81eVkckxN3RL4ITIU7DhzzkIBu
JxlFAX4TzjA/Bh3j1h4weunwq8XwOWX9wCaxjMV07ku/lLFnBEaJc+K9xRsc7TFM
LYcGr0fwNDKnpMUST+B54CO/qQiuqAFgQTsdAAwbsxwK4zD08+7tp/lsPYgdcQ3M
hPeRAUUtYBAUBTk63n+Z6Qt3DrpY9RRtF7rLYwZQFC/dcrT2gwGs92TXpRWy+NoJ
UXF5bltMW2pbP48SfYN7O/YhxJcjB5WbxmUHyFbfI7m3W+p3Da23faNrL7Tb62mM
lISjJXHjzVM2axhJTTe6wYeL0DMJPBVe+5VwBg1NJz3k+tjzEkF5PhdzKhzvz2iE
9P4Lejrog2Y8ywVsTCEPzMOFh9jTbcjyDy6ax/lz/Pir4/BLrQikSmwJeKBE0Tmv
btnBu8823B18yCbMBJbt+4wrzepIZkEUhmOn4bh625oD4Ucbyyi4fbxT/crOsJLi
IGe2bhi8lMcQRnUuNkI8pAksH8diL3ZsB1m0yqEIQF0N2qUk5Mz3L3sYHCeHZWgb
VupYoT0LsGT15+SKwrkDj8uuK6InttVsAyFF055ukOLHp10VcmxOa3lrAEbLA4ra
vaWzC+8b+ak0+7zFoNvCo/XRnky+KRws7+4ZNMU/r3tY5jhP/qG4BZ/pKQi0zDou
DgJbSK8vkVP0ujcLjsdcF44/5xrNkSgTBXJAT1pb/3532v24akE0hfq3AuOwRB3P
+vvFh3jscSAPuWaJUOUZ2mfrTaI1JZkEIOHvPP8ZtxYG4gE1tYgw9vIcbJAT1p6C
adcJNviiJQhI8NAPBXcmNMdos8bCRAPBrOgbYrBiF9KCg7pmgdS9oYG+rNafXlU0
GjKR3HRh1wT/uqLWXmqYSQdHG9coFJc3e744r8ycmega/0HUd2kzrg1Nkwx2Dhox
tOkVH1JAEdE6J3GyEv9DUUQvhxJGXqzFp/avjBPbeB2pgRjEpWONkCwnbqEeyboH
tVOlVHBcKEcUL4da4oSwcFlE8flECCshSnNTad1Cf+9X3kOwgHGNMIMgO0pTGwor
QomgqefM7/o81I2KeLXe7R630pM5fcS3OaFD3jjaGsuwS8YfGDT1m5mxBj6EiIRb
E+0O1ttsWE4YoWVDZryWfIF8gXHI+UtZfBGpsR8SkLy9JjLxskbyMW0w93gkLKYT
/G3bYj8mcbxFB+rljj3To9QwHGXoa9n4BL6Om8+H6hgV1Yc9/rOuNKrJh4jd1djY
VquVV/2eEMZB7M3TT7YlHi7LDK8UCShEub3O5kduNqnzTayEyj88ce5G+K5si4lN
jAcMlhpug3yaJz5n9K502VawzjXNXoyhW2Qhtvs4qD4zQb0UKzc016lGD6SFsCbm
cuUtXXIuhkj2xl3PHsXi/lrvDSWSEhgNVic4RQHYggtrsgT1dC/NJ++vBxDEUs2t
TNYBUfBMX7nYVHWLRtAfSIsBWqJMvx4MTJgzKc8kZpje1xgbt09URs8CPSnOth5W
4BdWZx1wrnlS5sst8BfrtGtDa1CEtzjdfeGPYb6aqI+OcmSF2Lq4y39mEUFSCad9
gdfHz3tBoUKcxfidg9F/GTWl392tKs9xbVo0E1d+4ENuMYygLjczYVK4t9ktSj06
Q2T5Aa6d8nDZRV60uN0CmI+wmnJvCjfkmTO85p791my+p4eeF4h3bj9bpf6gM2Om
z+RsKbuz59q82MijSAaBNPRa226qBUrlgKQ8LfEtf/BSjDn3cUd1NVn9iZ82rHAE
oTlN3NbaxIhI9eK+prFjW+kAay9efSxFdBMlkA2RKR5pHYscpsBp18zz1T91i3hF
cds48ry7UkxkIxgTzAyOAYdHqfj0nxiTbGSpCct/Z40NkiobTMGuzYjwcY0Znqrv
URH9KVz8YDARQBwx3V8Z5k0DMiy/UmA8foX3XUWIpe32F9oDOrnpiMxAF9/UbN40
b7T9rF7bvvyrX/KanxB9wdBgfwwHSc/8auxGA9/bUB5XBp7jMyfauk4dSXlQYLRQ
D7eHmeImq9/vNP4N61u6BxyZPpYg75ieTgqSuwJc4aMulby5Myi07FK1bafHJ5gF
sO0ql2fUWrggQszFrqPr6RH8Zzk//yuBEwb/WUcNrRmLdiU/TCJJLMD1w6Pxeob5
C0bhf6JO8ePqr5E6iaaPL/dn6tXk9X82OCmo0a57B8yalXj7tFSIHjjaLnlsaTua
6pBC5FQ+JNwPNXvY05s+ry2TUjDA7RS3BFZTUQavsCRMs7njuH1nYn4RAnvbDVx5
8U7pO5kr8pGiJS3MwZYUSzqarVG7gMwWP903JlbNdrCIMpSRA2+tj0ZYVNrSRrqh
Ym9DiX4/ZoM6gVBwZ2Eo/7QKxf5D/LFQlrmqIugjwtzqmZtCEu8yW4onf07fUaQ2
gH4fHDO72tzkAMT9UNKzbTx6SJTWZL2w6eD1szYEwYHYoSjgFtsZDQPvwgNATKcb
S7FqrRHXBNZJE13ZDBfCHnXY7hHQqWMsSGQnR1MJBnzGZYXRGcX9WoG/SSd9FS/g
uQ+C0BF4jC6q1pQO5CeN7eJUeo+HyqD79P7jei4qQOm2mPUsPDzYEX78mJmLSDTi
yilNjxdPlYOxAJlUpZZEgxvdN7L6BoqCRovH+VALX28GoXiUtFjfpI+aFhgMtTaN
Ed80bWGuJcAt0v1ItBwba+RyyZrFL+ywjk5AAoLPfx4WdsJo1Y8WRYpI763FP2eN
mR8+G+lsQ1fCQuUoe8VFMBw5ru18v2TRUOY2gOxIg22ysG4xm85q9Hv+3/7vcHO7
VP4hkWn7tqDTgKODwENCqU3KkTr3GmhrsoS1GrADAOrpR1hlcwd+xBoal/PHa79n
uSh8dlPBI3Icof/K3OiYG3hZxDTNSVscevLAPvji4klCvrXyMWUsWacVDXj5l22s
h7L01xbKCFSAgpjqLJjw31nmhPqu449gI3U+z7d/ttxGHGZMJz4OccRh2tnXBRuD
kaxAFGOM23TzKBX9UbjG4+56rr7vbvAajCOrIuy49bmsNNefi4JTMvraB7BU5HZm
PD0GiwFf1wvXcGlXR1DTYUPWXZGOzXlPIr1WnptG/s0iHHz6HcJggrzXqTb5awgb
Fh/V1Ne23u2XImeng6gGTTlR1yw9+crGSGUyzsbcUkUTJCYbsbou8WkTvA186gVo
8Vy35e8jTnI3HJB0vyIsycyQHYyd6/CspN8jLSuT4jgOjn5IbOAHys2R0ZvMYQio
994cWdMcZESN6yZr89GlPR6t3NnO+A5P9nE4AtvQ4uHnY9UFdpQzcLHPCrNVia4e
gfBM2ppxRRJNVuENioHgt68+cfSeZigsvC5mmXgkjZVSjpmiNIIhrKpUhTcRF9oB
ANk1wOpl7b7mSvaNpNweAu+uoKO3qIT4EkMPtvsH0gt7fojhBNbwGQp1/BlH+j5c
3XjzLj2QcmAnHBZfbTZ/DmRrjnRvwRLUtEVou6q7MdwcmYWzOuCBW/+eg1e2mxcI
LA6mTARDVNI2rCWERz7CRIHzEMU2cWaVDHaU+8gyk4qxuwxbDmkm/NWWqhMaS0Nq
XB6t8IKxfEX9ZDB8g+6mLZfTmuPQQF5/Z+9DJY5b7R6/4QNCNV5A/oXci/wiwr2V
wFGjgnJxZ/Fpze2iNqJ/YbIodPyu8wtxbA0ee0LEku/Juso3aJy1ZjVKA+6vVifT
PBunGF3UitriO9aCARkX7slbPBLWBXq456Jy92I944Yy5W+c1wwA34ijnYw8hEzp
gl/Jnl73EfojL3K40uWk5P4Xo3SOACW7v6pGV9gLbR8qF9ZEsAcMzpbJKbGHFeut
WfzBdzv9sKBXITvlM4YDXDVCJAUPzt/mP+SRk+8YuGMPffuzKZqw081Iyik04DFy
b3aSVeorGaVFH/54adZ8zC6t0PbQzfHp7uGvjDI8R/ioqB04aSLraNAMc0sAQTqv
tkwdl5snG8NQczzWr63QTphSFbavij4toCqOmRfZOSwvDBPCimeVSlukUVn6wBUf
TnQy2Vd3tAKDSB3jwog4lN2FDxD+n/7IZnt54Rz310nffuRNCVJhMpOzyFGphMvZ
8j/7F2+g6b1+ZJmPoEIA6IVXIITcOJiPAbJYWIX1DRJpe7YN5uN4n4eUsS/Em48m
axu1kC3OcabMUMPzpOaT7/gRHAw45LU4N3kwT1Jd1KwbQnhxni+V1wpQopBBYzrd
ghNuysxDGrP5KWFJSMw2E25c8B3AgkE2d2cGUnyXUiP8sKDMAlFdLpMwIPmGLLvO
U5sA3mqmZY6qbs0I/V4IZfiWSZ1YU/K5OGBdwIkyodHCbxubr8oJdFDoXRMqPXvl
RNZTE63LJFPRpDciV7sqZcJtoJPvD3a/1oD2X1zy6eD/dbPvQF4XZJE2lwDq+pdH
yMJ4q+SW9YjeLpj41YA2SlduHWiczWQsEdYRlEg3zoWvLEGZlA/qRm4PBG9yiDf4
vMTqeCncb6o7n68XVJQW6n97HCexcmDB0MLSCGj33DePHCAMnU9+GuCBw1CZCC06
0SRj/kKzzVWzO3pFWZVTHxZEWaNMrcHRp6GQHsV5upN6W4cFTaFXJvAVBpYECN4d
Z7B6Fo6bAO/AzqYLRNgn7zhYa2ApHXghr+VgrF5H9pssZajV+Z1xjhRThE0Gwt9r
8Ns9N71dxPRKbpQ91QQiDB67ejER5hX5HtmZsmkc0Jzz/oiYLlonTigBNN5mHjJ5
AXQKDnlvqXu4RxNstrIli5Ir8xwPii1l5/nWigMXyhGBQTIH/s8/EtwbQO0gKGr2
cjpTPryN+g7LosyeLF9d0NTXZsIuw5TWoPR1rmU7oq2DbSyhmsWvLEVX6474fqhi
aeF0qoxi12/WVAtHEA+k1+I1BQ84m0Br8MttTQh/4Bqrw7APidQHV2QsJght01Ow
IcGuRIcHF1f9Rk2kSWoq0bz3m9tGPincfXD1obpLLWGW2mHVLo28/QJUlZQw0jfE
XSwDaN1t0hB/y0Ue3RZll3kU3QwsKgqv+eHTHXR60fbK/BZAhoMzonlPb8XcSiS8
2AZPMEe9m4oxH9HkHTtlXn7jSghVHoAg90+lNF9tHDvpBX3TGWsPTOPJ7tWJsKqO
qm5ym42WY852ARYyaavxAX09gYNkJ0IuWI7A37+kFJKkFtQty4ccAEjH2OmYCmaf
OPw+XP+xom2/0eQ9GU5UaoZKrppYnBLgLK/oJ95O3HZEZ77x6M0ZPbQCk0sVQ+Ai
/zntPAZDYwfHcynDeTAwKe7CZ/y/UKJr2Is0r7owtXb+q5wn9gbUD32wSglm/cgn
bnyORwek+YENX7tELcFDSn/Vi3Cve/rOvE8mgoPhE2FUY0xU6ulWHX8e5G1oPR1e
QOEHZg405WAhCuCNfAtE3tUHKiK/Xq1Cdgji8SryXxXQ37W1G07m3EeYkNfrc9C9
Q0185mCGxkjujlvhK3SeZcOMKgcAT4NpeVtn0WDQC5UQtIC0Z1Z7/jMEe4amKdUK
48I97ngTnYhMr65a4iAxAUA5MOlknQB7MYhOPdbaxdXrr1UYtI/fEbFNLpIMpM63
IJckVSr1TyFPAwZWpCpfBalu1Tnk/Bfzmgh58cSW4xe8ziPQND8UIyhswrpSUG7q
ldi+pajfqzzXg49Eo63qJFBdYNGWko2Y161Sd6RftpWFrHRishgyT0QAqTnReR86
mr1HH89rt+xDIJdq5062u9LI/h8OTvfg/4CRjV9494KIUVQE+s0+vFvxhfZcCrtA
F6wXlNPdON+RrkmOBogoqC7/rkIs5EbYVtgBbDC2C+EVfJ1baTFMIixPe/Q2mttF
xVEEhnQkmN9XyUCdAwqJC4sUe9QNipjmvOBIZANlS9DmtW7xKameaSeH7Dx4T7hD
JSrQjNVvLieakdTtEkMx+EUxWk34A+7Hw9B6Wih0vm5ZPCxSTLCeyLWBLtWhARGg
HnEfom0/Vq4qVU1cJvarJ45cTSTWSf5f1PQIKIW7fPLErPMk8pT+YQSzVqKU+WJR
2mcUgnKf/zYADfAIMZ34uiHZIt9rRlhfPcYracDyvmhY2J1xfcj4ffqAlf82QMuI
9IpTCxjixaCH02LnopclALUAaraHNe/2J38CEyOckWnfEi0Uv4rk7UplcPnDU0ex
QT08sd04aHUcuDEqIFqTTLXnnsp2RtwHjVJhB88wrh1hbA+87Ammn+JrGYxbfv2z
ByIL36F55tDcXA1cj0RQgJUBgjXN6fdWGcD/sy9XB682sqezTVeJ2T8HRdSdUwlk
V3P07otdEo+2IaCoIQgv8EW9cldZk6ce54dzXG2R8VdEanvkoL8rUg481kKOL99E
oizBwGUWv4F/CsLwm35EkTExVgkSjVaY76C9ArV0eNC/v2M61Rzda0f8B1myNBvt
rxuWY/teODXa3FMORLJ14r1zQxrs3w5vYJXUy8IdURcVpgOpDoVQRd4k1GgvW/8g
ga8I2ZrnUPFOFKZSfj9/14Dx7zeo+4mwPjBG5Kn2ffuFAWLo9liZ8uZPE/pK+HCN
xMpCSzU+l00b+5vjyGLUqoj0djWpXyr8wCb8cv7cwb0nnBpzl7qyHwk4KzuNaYrQ
TLmY+9/feK8lw27ETJShlE5RDrkdjm28GLO5LPwMkV7aFwYEkgZ0PaL5DCC0o8gb
EasCe4UFR+Tm9HDok4fh2ktyYwTr05L7WpOChSPLy/gocywVSBSkRcNxzDF6Mbw3
TvOc8UfaARLZYb2wtX54isMFgDxDmkD7SXbbfDCjEq1oJtNaGzdI0kskz6PQinld
mhb5MUET0sxtEWBFG8XIe2D9Lqo+tNDwwyR/lsOHeXchbVQ8gBqM8Y4rWoqsOhl0
PJI9ydhuoplQYOkWUCpted3436W6qJO22kNi/sZ1ChT6I1hWa0gHUKwSqx9vJtkU
FnWwAAaCyZ3MwzXR747wjSXgCjkrckZb0mA/CBFvkzPtpwiDf+1DehZsDYaazKsl
uhwLuPbr+6Ub3RRAhY5rj9lDRx1tSBgkEMkxyUmIixpM3jlSW6EO/fYFaHTQErSI
Bzr8ZUcCasyEtj44pGVeHD6QoXbiZAmQRTVKS4s/TLfdDc/Fdk+25NJkaKe8MhzX
1kVdO5F520V8yHL7ovo30gNJRIwcDb8j4q67y5TOL1qawmRS5ySBg58TqLIh7JtO
qUI33fp+ebsdoHNmd5mIxMj9cdSm/hKYY5napDiHAiEYueeX2j5wirmnMYc2OKkm
mtOp6EZS0dEgQWjprWBCLlSDUfPuLMDs+5QDdj4bnskGpQ5odEmU/YdkBzL9d0ZS
lpcj4R0gfW5vxg4hrf+TskUL+WR+IQug0ErjBLu+thLpx+9Pzsx+fQNwAAt2GEnC
6ARQssVs7GNsscU93beL1OX6Ph2PTMthRVyhn25MNO8KNcD71CdtIhkp39EV8aJ1
OryNEemqNmbu9lJGdOV8oYhVJ4nGO1k38lcEw9ZeyOLuH4nvB1ZDvFXhhWkoVYOF
JJOS2cx4O8DlxskBe4IiQP2Oa489Gqfi+eCiKFwtFCESTC0u3NU7OdXQjMefBtQJ
yBCIFh5601OW4xHBqKQq21CXgqjT59FSWIXvxDY2/r5a3EweqPy27T+Y9/nYHWd/
IhLkc5B11wkLtXMJvVnOFHnvoyOpfX7lzdjeKfZZnF4o+5G7QWdUsyBNQtG3JI1R
gba5xw9gGWLelWDgae5OcwEVVWjS1p60bi55qPfLIueZLIp8BVVZAqgvFU0Sb0rC
BEeS6jDmTmY24msYaa8d5s95BvzKkS/+M6BZmksr+akpBm1UAcGUfHQMv2LOw9Fk
K1P2InbKzW4DHkT0hPSCLoIZqVLvShjRZLtgBBEvZ8diQwMXTai6C3dATMxRwLHn
DIVNFGvPMtQhEacnzGlww1OA4SROH0y0kuYmUsvSGUpToEzv3KAmj4+1gALCdOUN
wRYJYq9kPVAD/iOxiPbB8ooKtBXtoMaLDcz4Hpr4D0kY45E1gqwaLtZmRIAP6Sfy
FC9DxeYqfTy9Ao9Mx09GiwCcNejHCs5CqWVhkAs8bhTQ+zWRpxYkMNRgN/vOb6Qo
i0zEI0D114E841Iex4zRjJAnTZk8S7LzCcHlb/Hkn5To8qRPbQjzumi0+gA+E30j
jBt8i3cOmm7oAhA6K/fayDKPqQeafo2BbCLppTdnpXpttOXltYzwgNBVcObftKkf
Nl1OkTeIgi5TilH0CKFD6sYucIufbw3vIUGUfgIYL0C0PzZ4NPOvrX65cPKqFTqi
U1Kfu3l0kynTRTw2BIJ+Z+UCt51Aj++urNdcM6Mrb8rp9FmoSYkHkgMutcigaUlk
ZAldoDa2XB1pCdarkU45idqsPC/JdM7R3Vd0Usv0S7i+Vdx0xgI8r3SCaK/t976C
kKC/rlyma9fhOdgrkcaVQ6Y5M9BcZ2pSFZlYt5+ebqAt3HuLq8XovVkrZWz48kO1
ZonbhNCWaap1PjXm4ck0ttsNtdaOJ0m/5EowR+8A68LLKhVFOU9SBhrhg+hZvRe6
J9pOj/dkxEe/pGtefu28jVQwKwSZLry1XCPCHJ0mB/EIUrJUlYRq0ywhY6fCymND
LLAr3mgXdLTA179QZulhoONCStBJlgaYPK0/bb8wjmBDZ/p67UdvXjDLbzqSETC0
eRbPFQLYGk5Oh0i8WwcI/J1uvNRPdbNFgV/313af3WiGvyX+HIiAuxgRdZRg09Pa
Y6lJDjq3uGoNPzABwZyoHcsbuwD1WIZw4RngkIHteH3qeG9+cmn1A6oQ37YVjAmG
AitAAppJNoVvTxqZPYBPjQZYy4LjNUMd00ALqgIOynGdtCwEBTeeMMgbAY11T11F
B5RZNM5PX7speZ0Mk7hRCQEIDEvubkSJynJK9y1uL30Extc9sxVRKXhLlha1ShVD
JBpJkN+PLmVKsCdOkAPDpnsdxebi7x6bw8qR+NL20PMO13IUOQEkkk/pz1Q2r++m
jxhrCwLpEO7Y8d3onXHoA8Z8IZW2oWLWwBkcAV4Ro+fyygWOTOVngurayB3wCFJj
neTX+5DFWyud4DimWVKKXOgjoACCMfRsSjwQCR6Wkp0E97AhLqz4elQeE01Rqmu3
eSrELB2shQwK4/lJ5xTkQaStTl+xdTNcttwu79ahe418nlULiEULg/xRhvjoDeJu
fuC5rbUKHZ6IpSkFmhQyy5rTBfBBu8GRzlSVHwCVUxXhm8ua+DnlkpNrB24AwHFz
R1pLbVB4NWxgQlL+clT6ldWcaP1fXWgOozbgKyyTQcRZmu9JdMKfCuP6DpIMdukv
UwQLU+h+F6CTWGkur4G8aCZIGf6kkjf7/7MCdaEOoGVDy1rUs49B29ujHKF+VkAY
QzgrAP5xvQVmGKDDodtYsmaTqpBu3+8GpVtrF9rzv1WJCPM418bdSc6payGAoUSV
RppOn4W/d0YD5ups0l13L4wh16zOFBdPlcVSU6yZ+J6w7YSlqGf5plknBQzbpIuF
gtt4NsE5RQccrTRR0/n2JdT8t0anrCFnrgxh/+WjMUZ6x+4tYAXwaO4jHLFMahJm
w3+TmxPkpVikQmP/HdkABYEMYOc0OE1xCKtaSRGjahB612I0xx469lPGmlLKE2fs
Y+5QQnFFx3WixnalrI/BKGeIDAhiLWXS6s/1FtahwySLrrNnMUL4zH9VY/87NQEt
DTJJwqKkafnbtYp4R66DLXEY9jNBkdsiFrPSC6KPb8uaidSFr6gsavcacyUPDJNp
Yl9mpwEkMW0MvhwVdRuky0rh1NawLUUEsngwDIOd6Wpu6JD0qfA0orHW47WnS9GL
+LInDkcyMDauWAVYIii23yT/d7DzeP2mPyKcb4RPnCzMaQ2aZE9OvNQTG0U7X69d
C+ckNSne3pp2SqywdKcevv7G4lLAvfQrZZVdVhLZT3H5hZkVzZh0M00U3rwnpcWu
tqXawlJgtgu6EvmvlXrS1KMTRDzo5WFN6qeVyFQdJLn6eJVQush4CBWNC2csOCYY
TRKnCzsdQV1ZtiQnogZmOJNWe85GoJda+Qh5cs6Vaa8Q2+dLGJxqQNZ3fu5Na4Hn
Tf8uOqzhGDztsZFIq5xRtx+pfvnZH5dejYZIwX0lR/veRTf6tGomJZfUkrv1McDH
zshCvhVFKs6cAS9KN3rnddfBpdePuIF5fKIAKDu7yiuBjXEJFOT/6VxoHiCJoNbP
3Yl/tFyC+UMd/Ti9VYE2TXqKcvAqGPj+j4PQJKJ8u2Q7spWQl3vtIFdT48aO/Snz
0+aRXR1wDq68FFASWbIOeRXlE5Eg1xK0iJ1O2BGCrq/fv9qc4M5azr+I45olHgSk
UHNY6lS1IOl9o7W1Q10gu3lSIObZJRZyxYk8h1/XrTTxhfVfZ459rfcZQFn+9lYO
5yAZswAS5QLgfjwRqanfRVwb64doyYi11JldGxIoF5zsnYbQpOmQhmBgptBfajMx
rv36g+G/ME8y8RLZyCkU7Y8PyvHlK9AO1vzTi5Baur4kofMKVeplsDFM1fARYK4a
MMDs/tFW+bs1xQvo+8nmIvoOuus4Ym4Ap12UrdlI8kw40VsAYaxhJlbUAPZRLgrY
388q+pTTE4bAfv/qfGl5N5iO8V+dorapR8JwHlyEApkXQUq0l+qSa2u6z2nebMoO
UhxTjp/xlwUxF61dtVEvieFGKY1pA1fHLbaxGEyjHUXMpBJ3YrLEC3sLCqp0+74a
wzpKYOiPt7BRWCeS7GHCEeoTzcZ8Ncejyj/DaUJpwuzXueuddNq4o3f0VuxaxNG/
gpdMhuqZhwuVPLswBl7WEBNIccMv0WmScIwOP6wgS1e/8FMYPeaxiDmKNLAKHRvo
AwydDJ+TJUIWwb1c5+jHsSMtfGZCIjFiFoB99UoOiPgeO9VnKHbuenqzLht/jUSq
DEFAQtE2DBrmP4XL/hBzcY7vhPXKuQZyQ/eqSngttv0fPp28a3ZncBG2TjxRMRdz
iR4cJ1QnbGmDo0IJfEK7RKorbCgc10wQRcOzYrZnb/UukF7/rsu6SIGrT2albQe8
ZAQhC9VDTixS4256YCOeNo3pD1w2bwoN1hhCPqtJCrgh3/2R+qzFg8baXNBVfmZQ
7B5M5DYEBxwZatLuHyv/tdWa/UsU+ye0UC22jORVmoHEwmIk9opOMfwcKu0x5S4y
6Zq1TUIV/ha32Q2sUQpLyk8CmfkEBDNJwxUbH+0NBh47Y/obZUyJplBpED+JjlEH
l9nc0o6tHYN/WTEeSKbKWMIMoSv24P2tg05MXMkfUI2EEZLWeOv5RNWykdF+i3UF
BlZ3UojZFoN2eM8KYqGhX29mFcsn0lh1JD7SRjLhcZWFqmMV5eGSnKADKaUky9AB
6Mt/0nWcGF94vRNogyLbaOFiCJJM0CaTTJgNLRBCyUJG4wJcB5Y+seZt8sCSJxN6
Fx9l7WZi9Wt9iBjs5NFvVZ5FrNSfMQVskq6DgUFWOhtpJ5kK4jblwjw69hkDJtHG
fIVqAZdQf9tL4vvvEMaEoHe7rTuHckgOTYtbMerA3QoTX4Hudhw2C1jB9V8uvUnm
xplmtDb8pFuCMqQ3vy9HG4SVBgIZttnuXUmL/1LO+E5VZJ0XS97qHp38EbKtkdFa
o0F58Es/Y1nwoCV3t+Fl/w8ihgBZT02Jp7kO5foKy6GxAHAsDVNBN+I+Zji3IvhZ
4ZvVMRZ2zvRpm1/wjgHGkziLYs87NANcLFENpKIt+BQEITjCl1phYjlVhgI6Dmvr
mzU41CD0mKyb83KLC0iNzqPEbxRjohHuT8+tItp2gb+jCfx5/P+im0Ra1cs1snD4
HXJ65svJSZYrRdfPGOtxe83y1In3JyD1S8XavBxRrtEJb57nqHFzXh3+0vIkufpf
vXJfzpsaqukZrMCGJin9pB3WEolf72ZwpTjoO0V7EbkcUw6ujoV1KH7Z9qoqtCHT
4p0a+1EjQHYZHWI6Fkx9NYuRrS9/AEgnzgUrdVw5kxwkQvQI7lLgnlK1OExpUjQQ
c1NzHvVY27fhOkLbDl3a3YwUx7RuYPxY8Ics1Nz43uuB9EwYtiQLP+YgO8oNyRZx
Vz0jBCMBHr/6qHHJ10uY66l4mSZfBWlAqUvenhmp4UvEoIwKZsPFs2Rn5mypLaLq
Fm+Q890cuiBcEIt00rH+zoRZcoHZHbqqwaREuZ8x7W3G5D4fga45YJGUL2VycYbs
fxEakH9jJdi3LzGHcNebFTOUs/9iBw23ur1sJiz1VNxe22TIMqHERPjPypkFSFCi
lGgvYCxe7PrzojEMx+ncBGujFLn56tODLyz5QK2XFo1OfjlzqUQA9Pq1Va/tZkEN
/R39h3/roiGjz3NmOVzXS8gHnaA5bX8kD3ojDF2TQs4gtrB4RQaggM6gT36ajJgT
5SC2D9AcRbFFZcRsuHDRaSNIyqVHkw3dfYtaoOb/ZStEc5DmAOLhQTE9BrsXdIXt
o/6RM3goQ8HYvvVn18e+w9G9TNYBr+VpELp9X7XMIM6/ig6uVXtcRNuWO+DpI7HK
eJs7IzEnBv7lTbhlNxAtBEYIK3bb3UHCZs9BzE0ka0ATCp/G8n35fEv++OSxBJTy
fcqHwnhXWR4/CLfvIUuVRsdybGcMnzTRv6zt9QbdBB2jZHZ2KfRrKr4hNOp0xn4h
jtamf2+ghlf6BNGOrPbqq5p27Ve1xrNXMbE9TrlAqD2X53obqMXSCBWnXNIhvPo7
5doaJmyu/rluEB71Lg0L7sGJv4++QI6umAvNLK3P2Ii/OAWN2CnP/A4RByNuLEdC
qCtk/FhChqbdHS2s+xTdo08i2pt4wf1epMeiixOvIUs5GzmlRDAXIB2sh7uH0eHU
99R3YcsGs7Zf8yVD/0TLz9xK+FGeNSyPbm4MTI4AWyDLabTELO/BEVxHA5XuJMLx
L5xhruFwy352KkxVIa77VA5ZQaMrVh+d+p6xitVqldoHD1x7q8753jIOLUx6YNqW
0HBXJl5Qaw4hqFS4R7uoA+FMq1AkRzBftWNgf8nOgrf9OKHl4sm4VK8xCkbcrqS/
TQsSRy+TYNLLdypYJRJCe270n5S+daQP65I2d6lvPp91ZB9vLaXJtU30cP1B6JJ1
pP4fvrXwOwRrLkxqmdb20Jy13G19U6R8Oa86LZF/8XQrIjwx3G46dKuZLUldmxIF
iNAtaL/dr+ewJB9J7eLzjq6Qnj04T8iHPdvmBQokyHro8HX35elgqTGZICySK5Wn
00/P3v5NybzEsTrNeRwrxlLee7S0zb3wNW6xyqzcc0Gxahc6O9v+LU8iQgmOWp3T
6ZQU3pm2rWexKCLP4i36EvIu3fs6B9jQFAEcnsDB5sfI1WWEf4YaTO/5ao4r0xjp
pjoC3UDb+D+VcrMqUaDSbaGPIqWPCKgVbDIVsg6OhfhbKqHk2Nr0o3voY/zL9ht4
kQPYTxHQInyCDr9YQ5NAJi6HTn8pKmpRndKGd6Msp6/Kp3ai4UTQYQrlacV5kHEO
oOxD8CsaSzrUV+mjw0lY2qBNt9r/HXZjCO/q2NXb2dVGJMqSVjsDME+0FnfcIYBP
xva6Po0XAbjm0tY6dBaAw7xQk44n7kDdjEK3dFvVlDrwQfeNavX2ZeW5zkAjFrTD
8G/DGq5CduRDKyy8fVP5z+dNaOwXc7tOZp9jZZGpq5HqvxS4OTWeoJZms0Vs+/7b
XhymVU+wVxBd8pDsOi8Q+Rq85czw93BggDv0/ULGJAPYR8OwQrvONz5u0VzWRyTZ
EPvsoedu9KGhjX11/x9mNj8l+bGhHCP+++Gemht90GWaNliEBU+X3EaUT+DfmIVj
ZTyW9QxXXfb1tT107pNI3+cIf2hsp4lczvrHcGp905a2Ek55zYGIc7/zKLtQnkvL
+pSOD+my3uZEdj68itBKSZPwpScO9SIMu5w1tSKZYm+Uh64fsMgJauX91fCTeAjg
AG2sDn85FFhtXv9NL6CYM2y9OYItb7so3C2qlYUKjp4RJzNeKrF56dzmLMHao+UE
qNly+ckMzuJFO1Dz6E4o1zZa25e9EG4CeLYyWd+lw2uQdrlZCsr5gvomWD5a6CZN
wR0uA4iR/addQj0KqOKA/01cnJhQHS4gl937Utx3jAm2cM8il+YczL2JjGjIKIXY
NLNofzpzM9PWTdfhSon9VZ/JMTC1yhx9zayrjlF3WB5Ul9AkNOJz8lFVNUBzyTm9
euyidW6l2zrORQnIMaYhH+Sov8Fd0PSdPT0tnDQNbj3fbaQFOwVf/vJdfXonSJHt
uHFZ/+qA+K46jeX2A5dUnX4YZQVXt4KJD6yUCwuX99KHt3htktqKVUNzluD8RHe5
JGexLdvbUJX8fvGZHM3GqqMog58maQU6xMV0Z30fVFmlqFa8pQv5iSw2N5tdXVec
gCq+BahEoiWQNNxYESs6Wb0tfr+hoduy0myuiXS56432jV5zmtGjaUGAs01mzye1
o9KBaAFW4NN6zmIqmJ8+s2tMvV4fF7TlHeqBnk8YWDgBQjjklrwYJZbtN+JR8W7x
AzsRpy3vP36Pqx65CELx4rNLprIyAXxsvqHevDZLHntVod3wsUIrIBtM8Tw/OpTZ
wtehWG/hZAd5IEgCdJn7b4jYxwAqRKXqx6r7yvrW2DAgO0ie3C7R2AscQqQ4Tp6h
3lmsKuDfICpX5RumeZybwSV3/DDHaVFk45INYXHgbEtZG5NEvYxcwu6n///HKUce
T7rPXnHQcms21GDF1BT5keLiqLwEmuHyKp1pE6Q+40OHBSiraqy69M99ZTjLogGp
CXU2CN5F2zvB9OXp8OYK7qh+y8YV7mTaGrMi0pgfe4ns6b6nNvsH8/fkl6itSCuZ
MJE7GX+GBswJJj3uZi+wT+NkBtLt1f7AHb395yL0uQYMk2T82bC7zRRu63MPm2OE
i5cDwnEBbJYFbZmzNQHy8F7dBWXdm1YEWj+dVlfuRi+PFh3rDk0PVS3hbU9HOtV3
o9uRjGB99HYAbzaT/FXLDsrQCstvdiTfAFEMlbhicUnyL0ZPN8sqYVVTMPVJD/8/
1iLTLd4kH/Y03t6CTpVP52uNbXdGys0pY05rzJHhteN8s+PBxgzUb/rZm16OpG+2
ojEwI7G1Yly8FPB7ECkp87iub97GplH2D6oYPhIXk9r01UfejFLkNZ6J6R9dgQin
gVbrReBXo/ohp+RGsJACnLfrFzGkWiX5IhqYn0SNb0tCSNeUrUFtP12vJbwOKeAx
Rmwoi/iK6Di2RQBrVw9bnac4BKpyc+OQarvHqojDnsq+WycNhM0KoUnkbVhPHe5H
YOZQ+TyTOzhbI7pwltRBEdYCL5TpARSDwa2NgG6q/5duRwoQZJ0aZrNqsiHpCFs3
/qMLwTI2WeQb2bBoMLdcxxh+8tB007wN0IN/rloN2yn3CdZ4ACdqdbrhtZGljFlK
atmmHcSwO6oBEt7eKXEfDVpFxyiMjb89TDRRbBrs1ertFbHSHfsq25ElepvE6wqB
gesDbT6DWaTQCFEf1zd9AGf9+XiEEwHCiQ8d2rJge9OXIJiv3oiDuu2GiiO56FV1
v0VHophxaYx4dQf7lC9kqkp19x6/2JRikj2wRSYkNArifyqznX4rp+6Eg+k/lDtY
HLbKSS/IyQfORbM8wziSk3dKbyVvWMUZayFP8Ew7Rh6afy2kIBGJNGYPbO6Zic4q
Qmo5ws1I022peqegO+KIcM9fQJUmfjPCV/YIZvyEpnr+PTDZwrXV1b/7JK/hPRqi
KLEgC3IucxJ/U/2OshffJSJBpsrzcXnFKhkPPN6UDLv8UmjHho+PUkqLqsFQ2i2z
1j1dH4snkizhd76rBZAPjFYS2UXhLP97l7hTrq9Y/VVGjlzOkPcC7razMI1gzt9L
hNdwpxTeDah80kIVg9oePfk9+vLiiva1wP1kJNF18Xh8co18pWSCUHo8mLwXsfEm
pu2kZoAiFBBoPcvD1vjDITVMY7Q6I+W5EVs/rHGktmPRhUTNufHV4EyMtYp4d/7n
FTf9lknoMiaRcGtful5NYyBglB5/6jYdRrdRaynyeze2a4yJXptbcjhzaACt4XlT
qZayCNpmiJRprLr5uXQwwh6zB+jaEFxaP2uWqy1NyiK1r0zXk/JLEM0fdcjJ3Fso
UVT2pUz6xa44UQirP9J6sa/UEebOF7HhDbx1YsLqkkUS3x07bmEaNVXv9rOusw0/
XfCm26AEEDB2rPsgDE2WNQPpAAD2XNwyeaW4CfIwfsvO5o8KXEEMVCP2o4n6irvW
2n4RO+eRIFnw+HhMmql0FRVSG1bPASVLgPvxIR+SyqEw/AgSMcOzeeGXs/zH0Z1h
/9jqkPfiG7DXVmRoB8FlbMYmwdr0zqlwfebZ+a4jdv1kPlMhpLwsfLMyGOnaUDy7
8hh9EUZn5y2hEsa2sjUgx0V5r7t4E7YaifzxkBNC3n9byJXi578KfhrVHoI6/Ozc
zZOVLO5rh0FOy6I5eH13yHD371HuP7E4H/HGJf8Hzgrbv0p5S66R2MJwBsPvL5pC
d2hxr7USy8WDnpg2mjJaCaoVZKU4e9Sw5zWgtwmynnt6fZiAEH8ipkl0GtmNZ70x
wNEm+HYepqWMRGIkBG+IP8Wh7sj0obfgrrILVlES4h6d7l//gS8H86yrGgltvCtT
85xGxcz7PUfmR1Eu9cljGoNwNX0I50pQh5oCENUFfW+CSHf1xX+0gGxsLCkpdilF
s5pB1bDXHsghExWjVkPRIqeEaf1ec5rwVd7uMmco295sYGGnALVCsDPzBdVMM6vw
VN+sd9p6/A8asWefu1AjAaJkDdCXGMn3ggXBJBxstF0XgvyVs50/3tPiTyHjoaC9
Emznpx7hB79uCy/4KGIftC7dKcJ8CTpdfiDo98WphYNPwDcBH7D4AQ19Xw0JZ7O0
L0SyOza64FtxsDjdRqUzaXawpjH3XbHc2IrkynaSTxg8JRpmwxUkwas71CXZL+Fi
RzZSyZ5QEaAYV1GazVsaHzYptcXU0rIq91ZraZJSnOKxWdIIVX7r18AffKnq/q3j
l7iJkAc4NcZRSvTXYO0HLQfdDX+9l9/P8CNSojqey5zKuyeg1HcM7POSc7iPRmLj
HhWo7AFlQh/bbbq26tf7GRC+xSz9Jyb54CIgZn8SZL56Fh3fVM1h6y+5yExUr0Wg
le5e0R58ULvz54/nij/daGXI+TOkSniHA58oSUUq01kQf28tjV96XmpNGoMu8kr+
tc9E8T4cy+FdRUfALOm5NrCjNszZmOjgSnYWc7lIlQHGgIv9sg5m98KtMZUE7l+s
AcLjPGF7iZeLYIhIJt550eylmjV9e/oHmcATVzYwf1/soewvB0thEItAUAEeChU6
R9C45Sc86jpz58Fcrh9HyTzbqdFDUi2zuz1XJ+meIusMbrJCrIuab76Nfa+2rQFw
su30uEdFa3BQCvQ1npgz5BE4zEcPGhK8WV8Vd+uiB15QfbezsP9DD3/+Jn0xhleX
3PsEG2S/F78Fqu3AjRw9xLrEEljSEmDKhBkkfnNP9W2kE0z1YLjVrR2Wfj8AJe2f
k1hHhR+DB2HTBNXjnDSwEPT1hHsKXwx4UP5XqHcsZGQ7VgQKbwhmtA1BJyS8iTtC
B9Y0O0AMbGaZoNRDcYl0n7mG++NZEPDhv4/QzMc6r1628JNw2vBSAgtRks49EOtp
p0Mrpbm1XxSs/y8VuBUvDH4hyscUw/xl7rkca9zCbwVhrtsygQvYjaL4SUFgkckA
Clx/XASp7/Tx+bTxIdZH81N9yo9bLuQXLarXLAIcVIYJsZfYuBDR5g+97HfAFzm5
hUVirX/c+BQxWjlFQNWRrUlWtzIWFjPEjSqtMQOP3kOthT84kU4xNs6GPlWSDeS7
2vB5E5Myg2s8bvVzO57GYLsajgX8pksJGSdTK52DRMNmx0pdzKxbWDOAHyU0Bicm
hmFOiWP2XFaOsgYb4vhzrajXwg2FVOXp8nyf2LZn5u1BXd2lv9yS1QOcCQbBCp69
aB3cn/orpK1uf8BcdZ+CVTud2jNhxsLt1EK+qMJQduYEYblfuEp/tV0ZHGT3DlDr
wOYKS0NYkeytWykCOgn1yMpeGdLxdH6BwsUE23igm+MXPXoNbf/khwO8jLOIa3dF
Ptuspie9qi6LQcLehwbiOHTNkfx7PWkeHBQvKvXScbawEFUtXg/21o8CKXwkabCF
3CDN70F1eVNGYFs5PpMsmkx42DaoDKSL6Mp1dOdK87v7/ftHGddXGSRLVrqGusgT
uOj9RFifEBGgqt9n2yloueywK7A0WciUqP6Ggd5JEr3MONRWFwSukKvkVJjkPrJV
TQ+a/ItgOBGz4eAGQPGoNGnQw/LrAM2MtCU6emfrJlDVgfNKV31K49D+fw6yYE7q
nKbFrjKgumhl9FvQCUEGmAtayQ1dlQ6iLnw0fo9zKlTZd6SwpeSVS7BR9m19U1gn
nJH8gxtMR/w8TXg++gmpCKdEFgameCT28KV8+YD9LrvGCi4tCO6+0eyrFVvZAQeM
0PgjtDyvsgkAMyfwYCFtTLL5dt4TYYxrJjkSjG4mjqH8cgyZMSLkLLDTVzOO2fMl
ERBDa8utNjVmSeZVvRIkNPPMEYSEupCH7QcXBJbKjEYdqjL/4tPuifXDDjddvnNT
1WdxrpNo+g1YghNnl/bAbD7m/LU0LLfaQBuFPaZ/5J7p8dOnaGkxx7lvv6+fe/yh
xR+y8Nt64chSjsD+l6NjWJbwTMIXziLMLq9i810hUIl8IJRN/IegfTTg6a9ziAHr
aGw0pd7Gv4Bn4jNYkHMu7SlYZYPoca6mNbK0wajQ1/AFiPmWdASebrQudu9yVreI
jB8rrCS16rOem6+YFREC4lQAgxRRXVInUUhXVkg3wMX2LXqp5fxxhEUVoYhqvTnX
V3mBrYhEkSI8GqeG8EYhxQa9Vd8di+lr65mJdO2PvfE6HcE8TxifgVIQdwqbb1Vc
YDlHGrx1uT97KdGbEDaTnxRmjAhdSD5aB/Orqxr4F/L+LcCcY25yLQ/ttw1NZ+c9
uBM5a7Jphp10eQuD9LQ8Z+ysaNfqE+gieXlWxl7uzLihvVT3ZloUPnxgc8A8klGR
wAJE/f+j48dnxU0EHSBL9TRm9BzQodu32RNot00GGpiMIWqL+hi8RXC3OJsI0qHH
AQbz4yj60Mgoxcs2JmG0Xrwm95gWi55blc5wEJObxf6KQK9XVCZ2v+2MyMy4LU3T
DvDdJ3/GQLWM6snH00KdLY2IMj8825JgFTfeG5NSmUVOxH5ZOp69FasSSHjoHxsP
q92gD3lyAPVidvyaBwKYYl9ksLrKnf6guwpaVQ2TSTarcfEKCJk0VohTdUWAI3Y2
/sDi29V+utQjfvOohIz0Hxh8HGLblIT/TG2gVOVIvKnABL303h5ip6VcjuuF026t
cYxMQ8IgV3OyR9YnqDEwSRepI44Fq7nI1nq8PA9OvScZf+3ypw1tU2EBNql2YGtM
tmp2R/NAlS1QECIyYL5hUUaNks5Kw7YdxY99fYTernAbZLuS79RQRt5/L7bRnSpw
m0WjH9yeyuw4Zhj+f+iV9w8sWerviqV+JmCjh5tE6Qn8G5BDLs6sxwlPPkqrlizl
jLDAph6Og6NO8YP6VGwG9aXHdm3CImkPmXm7q4jK28982C4hrTUj5I1LsfnMDtQ2
G0WGTHMhOTiJrsaApXfOuI3d7p4ZCvUxQA60f297RtWvyrQqzXfMUw9VkhA7dtyh
7VdlsWlIZecHXsnJdEijMeyZaYCFwdDsizpHW2PJOqOOzDIUlhNIXTWt+4OHEN2J
Ie0Dt68L8Ds6CxA7y5r3wTcxCjecPQaJR/4MgG7xbKEGpE/GBYbB/qOUYOkoTTlc
h72k2UvMaOBlhNe+3y55UE+Ddhs3+9qf4FV12vuCfZrvH/OVBbpKZPSgFFxKTqgb
T2uZPN8pUMunB4nHd65RHAX8a1t9sY+vZgCrqipXVMOBd0LmkKa3T2rPL4lgAYKy
H6TBCR4BIjS68HQwDNMw9xCkwxUkXsKNUNGn8RRVURhUeOCRRm5F10MTiUv0ISm9
kaacZCthTTcav2EwUXqSTWbRroyaVRR0HG0bjaW9ovUusxLlL44gFOffsoS9e6hU
QiSWO/Hl0TQM0nyYasxg7t9jVbrGQ7ZkP5Q6gMruD0e3HLkSs0Q+77WH6fjP+v1m
2+IJ3tmsVwyyFfLKSCx8HE5/KHN04U7y8ldWZ/uwTQyTre8GJuerTiIf98YCjccP
9unJEJ8oeFsHHK8iUPhg06ZedqRv2z5KjY2g0IPxrQ9FBB4lkYrnPs+WhdUaicE/
JQ4GpjRhjRuSzfDayh85LjFg0fn/B5CJogFmdET4G/TJlnoRwFdl1uBlnTQR9hJd
U214w1/0ukB7+snlC8xlUjo9iYOgshSU59unUumNoUeMk+mZWb5O2nZ3DLUaX0zX
BXNpDi4pZdfWWFvKfeivJCj4a50HiuPk3pGQablTOTPN0k5+YX06ofmnG1XVDbhT
qM2vcVyV/iPhFWn2iObq9JviDNw5/jlRDMeToU2lYfZFRMnkNbYMgVXGSjmjHkgw
ja/q1iWwJ6wJmiQJwrXlaPLhEyn9MqgQGJqLvaLlVFZn4JpXiXXnC6qqdm+MT6h7
RiWhzJ1oMoGXUJAVh+UGLZeE0KzIPrj5v/UAgQfer8xREfEEjJmTopmu4O3BVI5w
UOXxO4mSETF7Ibg4dn39lJtBPipu0CiN7HtxJYRqkojhvWU2XgfntBhIewynvC5U
zSbrQB11hA9XWZi2La0h/UjJ6CirRDLqKetxR5NanXhLpzm7O2fIEpbL33eKoiZ7
AQAiFTHdpB5FO/mQJcjSVEDehaXYQHBJXb4v+yrqNObGyLFecaaCPQaKo2BikyrS
ADkiuZpxjy1vEFqTtRwOOvsEjNBJYBjq3duAqPKrgKrTIEPktxqhLhWOfwFaycRF
K1Sev8UOhRYanCP5mxgnsSc8TlVkneagcueTqHIcxD61aVnWVOK2hy1Ay36oCof9
CJsbCeEucs3j+wIGkwRBdB4B862c/0k8lcDABrhhhvHhkZc3Ev2IwvsYfya7ylnN
xXj/QvK6oFty8NTcHZVdAPAgj53xwfThMWeDvHYSUWKYjy86r68T8vLgxCzsS+oc
b+kzzVxdT65QlnpjJjfxw3qT4OtdA+TQgfXn1Dehxr6hipz9mZWlixtN0q2UcLWk
boTJKv5Yno8aW0dn7LfFXfFsUa0KVGQzEURTb0TKgkmrYyRWvCt29vv8T77W2265
9Zki2MelkY/hTRonb2wneyyTPlyHX3IplAoJApLEhZcFnwurGvRQR4JLfvPQCmu0
FnoG+fGPuQaZRPc2ziQ4qNGTLP4LkgpxIekwNUSWghkF+b4MzdsjupW5OSNhsUDh
UT8vGdKHec57vl7EqfMzqFzkWoM1Stp8IC1yBKAAs7Z0oF/fru5VZAdlHdLsRuWX
iPaspTujjLHGxpwiawSLuFCr9znYz6z7k1bU41klYoLKoQkrlwJ7A4ZBo0TJT8kc
ldYVuBA7gMPujr1A+6GeB4EvbMYp5d/M12ChhxTOqhvRkQdF642QCvJBKjWhaHAB
EoWzDfvMrjnrMmiRlOwAjiM/fHSmwZkdPoMtq232erOwzBBKAHRa8zUp1YRstu0p
+BhPRJghmqnDztl3lyiqvn/m41jYiMEVfHrRK8U6RAPb5z1lFKcvLjBGYOjBMDU4
wSGOItxuZTqzx08X4IaFMEhlE0FpQWtm0KoQXvAbkl4p4XRFnMDCZXIBczROId9n
ahKuw66srJ/nY6KNS7d0uoVe5J0o4vtBQxkKSRBd7NbXfV9yQ2SW+cPpYYTywL8R
mdXwo8H4pTOzGozX+NyqasaPkkXjI1TGAG09LF9CKy0+fW1w0L2a2foPOoV77vKb
/fMnRIsGTxXAWMsRz/Ivti4w1oRmO4Oxhh74tYviUjdHzfQN7H4f4prqjryoUaPX
Yyc31vMeFonbXxO6kXelpnHLA850lY/15ifpc4H/fgZQ5bNyFOuP0ijMGSjQzxKF
b/uz/r2InmJxWPeUCmqxRVE32Tw3+PYxalx670yBfoho7YMrc8gs79GNMSwev4J7
iXfWwk6Ry8xqM3zk0DX9muix7bLpRwOt/wwMLuLS3dPa4PBOZcduYvAIJN8aEseC
VY/6LT5vuj2lnrnBkOoQfBIByxoY18MUruEYNlLjGTlbRc6CDU0KVnNqb5+KhazI
VNrg4AYgtxSRnf8gJ2q5q1LiuuxBg3vnsM15OySndvUmkiBXHCniawXMVo/9yXXW
EXWHEo1GIfgNdPuxzpKvHgwgNpn97+v7qBxp6ZJhQ0fsN7wf/w+FZy4U4crXox23
4ACds4S4UPbFrRFndnx/wRmMA+a6SB6QLyYHPlZbAEx9th715fBGPwfpFIx/3MAi
gq+ybZoQ2AYcJalqXm2Had4idsejRrOkD3ghR638nyBA7w3RXtlVeHXYOxhJDUCX
SdKVttVuOpp3O3Rk3omQFsi42K6WErn9alSh2qP3gqnaY9lWNpJX2VPalNoZsFlw
NUOIXc4yLmSvWbqvUV5FgmelLIVosxZzNXHGpiGtwjo1O0YnRLoBshXZCeV/v06W
d5kdw2y7ZWCxeSBT9QFWPejUoXqRKK1D9YQ/VGzlPzOptJffAz6Z56JKlDF55Uwx
R2PVZsyL4CLzAizWC/7EYojmn0ZtozMj0xGlsdr6WINWHLLDtBm6Rq0N7tE2sr9b
mCCUlbgYB2ft0Mhb9OktYT/oiAtm9zW7wzdl5SnzA9T5koBVJ4PWYPaAysa+9hBA
WDJvdhO1LPZA65e0lk7gmsxb1PEJvqfotps1QnfUeNdCbphbD1PbJX/WA0ALQAFC
y+k2zZGk98ig6TA8HGcfp6uONKzrjOH0S1qyZCmC+dnTH64h+YR+GORPDG4ukvA7
Rf55qbKYM+dPvnExESAjNCf0Bb9VJgRzXWgFU+zEXZwZeH+2t0BNCKY/2x97hHc4
ytsi6bXFkR6SK624SqjBAitrMLF2tXLsqbPSS9idW0LotiZzFDBfRTbGmRzgu/9v
Kfmln0x41fcemHy8xVnpDu6LeJfO49iUjTmHK+ejH9kVJsIiHHlh37XuE2sdd8TF
qJYz+vzxzkLCZpgwlO3YWcI3D2LsOWnkLIj56x1e8Z3Q/oa3IbYqlcPieLebYUi5
Fihs2CRTfPFdfq64T0YD3d3bMeHSTA95LJZcy/eQY2O3m7+s5U/tWRe4QUdL/m0b
CMT/52GcePTFTKHn3749lVgJ5evOksyEYQB7ZnuE4lo8EnycC7+euoELwIOrSdCU
r/f1IHCU2rdeOFDD8t7Ddxu2y7MNqWcLSsXMUDF3QfiNvZjxzNyue9ll+4X8PTrp
AKRkgux2iuE9Q7XCdAAmfR4z2NHRm6PCWd/fN7r/81fMD8hUS6+mJ2Lbeq6w/Aaz
3RA+mPzQAhJeR6KEPraGpqLbz9HtLD0KBtdMxJPn2Qg8qS92lYwX/6hZRyuEdHNE
BnHrWad0EUngAvcq44yeZ6+gJhhtZDSTJ+AYBnPNiUJ9xDMNp1CmVu/pe5xh6TaL
u3PD0N/obm9qSvmJ12w0lbofWxAQfcbUz47Olj1GMOW0sJ04cg1Z0n5cflWIXAO1
LB0Oh86IUmBETR7IUqNsABDltcmbphwF8gi0tUjoMKU5MGFBgiBeghy+bK5lLPOf
A1ggyZrqHCor9CUG15aGU5J7QeVhHlFIgOzNLRsEtu9dkueHUjMWGZvToUgnzsjf
Ce5qfMLJo7amLdklOUkKb4CvszbV8TNOC+Ati2g5Id8Xb3I1I7dxodYvmRo8IHM3
Ep9+tFzmkEfUVwlrVaJDpq/LpRZ6MnEAElskqKeudwdNrEmfJhsvIZmdk8pjSTK6
7pIkzkhVFeqq+8LcijylYevCMlL3J6Nv/boETtFy6zUq08zwjlKnBOE4BQ/dJZmX
IXNKvi9BBvnvTEfxEaFWydLMn6aoBwiDpmoA2A8MlrTxlcIffmWVvE6UTExnx1X5
rFelD7bqaFEf88dRTVNwUvnfScbR0/40b8vW3dJSlaKDR9EqrOOBnhAayVZAEqRf
JxeMcGlxaAZjE6b78g7QwdrsJYS/hS58rhd9P2k8ZXv52ILgmWkA/n24zfIAp45G
Nk8BQCkFV2kiNxZv8jCR+sSpsUKm22+Cplk1MSSjDqxRO1rSnMjlnLoF9YSZQeCg
e22z3VjRe7C+JsrK9cWJQU6iUkXnBL7ui6QCF3eICzZjOhKOcrnK5UI7iZgMU/QP
uYh4h4R1iLpDuB1Lsnxlo34x4CtAQCrpao8s4KadYYKwpQaAxXpSUCGO1q44owmS
ZyPT5mcrZHV/LqvwI9YlMpX/vzhS9OuSYKRcZHcIin/a6FC80URrt2yDE7Wsdnos
G3x/A5aj5cdOlLDmwaihB7iFYoim/QheT58UZ+I2uq8Uv0YXMh+3X5RqBcKWCfbF
vdZlACVTLZHEM18Wxz5NncOtK80zQ1dnb5I1ua/LjPLtmrpN/JTUdDwmxzH2ftDI
CxkA6L6A5IqFgMgWNp/wvBogGHKKNrYAeF0ka7667TEsuEnsJg+S8RYwJsnqNGgB
H+C9QHLf+SHEnbemKOh+3eSmb5shWlgXKql5FwyJCHH28s4cUs9hNF5qtXMUw1U5
18fo+AJJVYazxjZff+SGNF7PzatUbBaySoatB/nSjRXEBnZKP8GV7PXoZhjR21OO
U1KAsJSizsQkQqjDgnkb9ba16p5QFzotXDvQ3kjfT7956aHsKZj10c1C+l+JukU8
VSbbEdYXSi0aMfFbF1toAXi6LQ+VTLCnoQAsoFZ0GnSrI5dqlN9oZMEEy+1YbCN7
zYZEQxVJAWJHQWN48cpTKuYNzzSabdNN7vCjgUyI+Dsa4VXoSbq8DVqzcz3ZgDON
27j2iw3GVEy5seMlWYDEk1OYVUz2xj2t/43QZ+v3lZmVIrYhg6ODS4iKCTz+wAjv
prBEPlkJ+Ql777G4osNhYml9vykHMmPrEuvXSyRfrQLG0wO7DDWD2kzPdPzcRotQ
xSRRYpTtPC7UapqbCt9Vn5TqacOTmo6uW+xReCPZ1c3/tnv4gmBB+JbEcqjil4R/
lcScsPOk3N+Cksub2xtCVhENrG/G3V+Na5GkXBUWPwk/YsKEcU/6dpWvsaYR4Ygm
vFIZ9hABTNfdM7bfJ7TtNOVdCxs8eHoyXNaof+iRO286D0BQbHMxV4GEO0amLvSQ
HfeqPTXQTl7cMlA/dBUckEBENRVhnW8X9pgovrNFWvJ0O83cX+S7SPsKZoJGI0FG
eYsvRDUH9ijR6rXOU76Uo6yYH8jFVMHF+lZNtTPyY5hNek4Sp17Kvp4DE+opVaGr
kIkk+0gH+T5a7oGwuYQx5Gh3iBRSJcNmUTnCaQZN3xKfmoBznrQV6ofU7Cd0JPw6
Se1pJfvj9qdepxcUi9zwH6FH14ZdVIF8fAL9cHIa7tPkU7OkwHt0JIrEkcL30zd5
AKrhiYwjX3RgOVEVGp0J/meFVc6iPUANsxUsLayy9WIVsFiP7WotdMyafr2smT5b
mmq85j+tATucPXwCN7TiHhz2M/KUTLK5blt8O8CvlNCgAoSWTl9yGlRiBY44Oqr5
7G9OUTzCn3qV0esXR5EJXWZQZzTeRC5ZNDEWXbTs15moQquP2xgHAdf2OfUHCgfd
1TNuau+fjmD5nClW7C0IZJuR1lsK9z5d1IRcNDGHsV/+fxObT1DeJatWLJKVz2KD
4IgoAWCwwDM8+dDC7jkhHMTW4x6v6hYjdHmDGxz0aJMqj01QXJiZDJAfQCAmyXrp
R6GFNmethDCfekgz+dyz0zyTVhQbQ1OE781QbRNqbiaSJXT2oI2VKdKTmeE4AXlV
yC3qPMm9WMiKk/K0RmgEjSRJKG3YKxVm0Zn+TGmLbS5JjpFk+3aJzhHO+dkwDlVB
hJm7PnKPUzT2eua1CGOrL2XkfGFW4vMx8N/2C/+as6ju3W4JP7xAN8oghPpatmO2
fNOBPQphmFvnSGSy6t5RVPUfU4Mg2K7wf1zfGFOOObHmQHQBnL8sfch2WYxMAhOX
96FH6IiUtbOqqszxt08enxa2G27E7o2RxIAWA0Env7fhHcHzC4gq17ROBF2ZkX9p
vN+UUffeqCSmE7JUQplsWnGdLNDo3aqYqN5nU2dD+OHIEwsUf+WApp1NdJuAPbgL
OPYvUkJ7zb4DejmZcbJ9Lb9OMQ8qydnOzS4Uhe7sPYAS++XysgrzU/C1ba1L3wBD
bkwscekkDW1EunqMbNIEM9R2OB1lDM+c2yHAMMzItQa6G5ttNHfBVJ8d5JfBdYOI
EpMgDpCpklfm47SsvCjWWsPmztmqDJFS5aod6dR4g/7ouYT4z+jJuGosanLQHHwK
oyeFjXLTiJfMxY1FsLaN/Glg3xNGvV94ZA0aSznn7oY9/71sFFLBeBGhezAN9zIH
dROQGMgzHuw+lrFXkW0gDlboYX4YRMv0ViSf0v050C4GCAR9tHTh66SNxgSh1FHy
+zGZTmVrwSpL1aBJThzqle2wIa3kboN8pRsd7S0kcOFHQnsBkBItNlrJefSelj/u
DnFrOg4AeZekEkPGsO1xQ7ZI5EmePUUz0l1HtpbxZ2G3ANUsiMSYP+5TTp+BPiNZ
8KGsjCBvsqnzF12qWH3vmuPnWNoRdlX7Q0uLhrZUC6fypGaCDF8tnd+9zfKZDSDh
LfRb7Y4TVUgKY97geGKe4BBVN2NTjd7F4a5M5PxKjnaHTpzQsXHohAUdZNl+f1Lb
SBLhQHAIAsYHhCSVyXu1Cxnx56TFuaIMoJX/Z10L44PI7fOC4eetmSjdEZX3MNVp
BYONM8VeAs86LzhmBfgzJL4xGe+vYMs+al99xZnt4mjfKvHAdUWzvx80Ok38Fj9Y
7J04FlNmE/7wCW9JLvVnQ4W3LpIWRbhw+LhJp8DAXmEIoZASBbOPImTExy2maEHZ
zKlHghLlFZ9nA6al2DjYQ2+3ZYXX1iYSuYq2AfWwqnZu/tZhwzVOIqOIC19d6UhI
2TQo1n077MCAhDk7lK8dKxU75xrN7mnFHAD5iW/l6jgszxkjYJI91engXU9ToDdy
CMWgTRXQm/a54R09SBtQMMl0CwCkQIcbz0kx5sauMWWvNlhaTWqm07zie6rUPLeQ
q2OC8jcD0/26ZxytjE5lt1HKhJsUxTE2bm/Sf109Pimdpz1NEwh8hPf1vLSWcfX/
CneT0EUFBNyKn8TiYDh/Q2Q4nYG3qb4C6kwfIklNT7WVmD5tTcuLkGl2gIilHXNn
Y8+O89mXUgUdojT/NtY45l+B4Q33a2WgSjW31kyKD+FvTl5Yr2cQ4pNrlKehPB9q
jo2yAO9goSIFp22SbtSDR5lRnbwr1jyxP87a3zm8Uz0Ot64RwGP7AfytsptbcYEw
3JcwgWRLnA/KgdDLSVS97f/HpJBKPHLQ0sVXDUhfKSNkJFVOfuGED6yhm6h0PtR0
ZSy/bdGO9WxeXK8RpUJA9IO29Chm8UlMIkXtn8AJSxY+Ou91CLAh/hlayLQYEfXE
Yi/dKWFKNHgeiANv0VQeDh3Mpc0+aZt8DxxRNadcuyDRpwEltslG+mI1o0Lr3f2q
ispzhq2eL/tafogU91wYsXiul/pXJXN2Kzre0H5hbR0LCXCvuFYbSFIoHDfnWGae
JyY2ZAKSyfXOHhkdA7S8JRJi5TYKWB5uybABmi6KnYTkZujsFvr8D31jJiZlkFEt
q+mlO+xyI2O3iWthcCyzhj5VJAq6/u3Do1inGGpIp9kekgLne15RcxFPk8M6P2nP
oBJSssEQlJ5MUwI/o30pcZpsirdprrcAMx3WgCG7aAPUCtXCVPeZ5l/nBHjOlx7c
NvInmsESWhvnuGdQCxbILQ2ABqRdzgUZCf/EpQ7n+cgEp1wX48HbWw9Q8Rdtrz2I
1OgOSecM7xX5suHizUQbNb5UrleSU99tWAPsBtk9/4IKoXPVfQXwtoBbXbzqeR5v
KekLrnjLJV+xgTxmNcGdUWsLUiFrrD15WAZtnNWtLBsyf27nAa/jo69Hv/aE0e0S
FyaOFcGBsIahAm98ZzbUskbEDpdWmMeKkqrdDCB825a9OHv8OHJSFkxnMtC1VL/B
JVVsM35A/X0aQ/EBix78cPXrAuRFSWogJ/T7E0v31wD+4vLPQcBcOftSz20vTt7m
HHloTTX+fUX32iwttVm1CeG6o7VculgoQauVigvr2y5miD2xpqh0mTtK2CUHF4jU
XCyKSl/v3c1vvi4LaWMdcoR5mFAXJF2gWshVhqRGGAbKvWVPmXkf6wH9hrLDSYui
Cm/Sh9YuH782FxfsqSCnfAvjpk9vQSce/6z+v+5lRGZC7XAYprTkyNNz3FhDgIpt
8qZrocEi9RV0Zcv3hMrrs9hMKzKAYYc3kxX6v/BlzV6YFSw9RiGl3HUh/SEbD6yf
5aVHfFHtqK+REqFLtaEXUG60r9n7UERNo1ttLWnHuMRdlkp5EiE7cSLkOVHQN/5x
eJ12DNHeUf5X1FdAPz0aC+Eh5jUn0WgrNaq1XROaAKMptsGfL7PZIctWth3Bqbf8
oKpnqIV8WgxGPPLPQM/TMhomSviuJYnmQ7Faablgsg2wnTHbcgkM9OTRuqgHhxsd
oh7ZpvkpIL2X30nRqI3q1ZO7V1SuXDWZCJo7st84sTZw9uWtKkeTHpNEU1GjFwJV
6QG1vA3MK/KvwhBkcn1A/7s3+pZSxKY4m0UJ12mY00DCRjS0CItmYXuhXXnP3WYf
9kRJ7ObteVhEIvG8pvC0NMJznDCaK5u0Ho0TR0hbJ2euNjtotkWVxlh/v/wT58qb
7jkbDPJ8QRzbolqWC43gE3grqle5O06MFJOT3/Y67iHUfKPlRDojwrAJWDvmV25U
oQVUDFYzvy/UBYk42d0S1KSzHLtIvL2KU9/FByBsuvu79+7aJGllFknTsmw+CUFS
pXfP6LbT/oBuSk/fs5FPjjZ/RjQCuvoo0Sw0G8s843ODhNsLwef0gytvzAdHGd6+
wRwqW+JEBPoi99luBLFqpEGUuQ0RM5gKTuXDaCRQ6cwSjIU9vDOxaSlns/DpilSa
6CL2GhcO/z8TIKmcyBC5OyadU0vVGU82BjbFnSLXb9Q1I+Jy4nwLmvU0RdceFQVG
I9HV743yvOkL5vZEwUjlmwovj3OTzn4nNlS+3OIdSwwDKyhj0OYLd/xSr2v+gI1/
PyemwUk9O5kggaCskdpWfV/EdkAu+xoqjhsfEihfrUuC6x39no1eIsQzz25Gm8dR
DNT4LirMVLYGOiy6W4kUgai2JhZq91+71Lptn7nf5EuGEKj4r3uhRN60QFsLwwgc
MZVFs6kDVtSkrflEXpqvZSsp0P5naObAbRS7P5JMomwYUVUlKHHATcoyY478yW/x
y93VM/a6VG7crIiP1KoODXQ1W+N5vpMdmnJo+hkPMgcdMrv4hLcQFcOj9sQ/0Y2y
2Yx3fuIeLJB9NA+5NOwvX8/cGaCz6Dj1FmeaKVyNhu2Pg0pjVw4ADp/RXu2j/aox
ObatKdnBHpT+EpmnFOi3eg0a5eQoeiBlwcFlo4gOXEkBukusFNpSplOg5F9UtDwy
k6MLssbI7CCnVVUqn2n8tD/D3hmPytTVmngl82AfP4g7954uwbhAFsCzsVzeg/Kn
X7R9f2u3d5LbvZfa0PCkmep+gerJ4cufxb3FBBpcBzXlS4HhU9ACOhRo170Bgidq
pKpPoPa4fSWuCj84bFD1oHNAwarfNU1SPYhxd+ZcAq91oxUob5znXmIhJYqgwTdC
mg8yUoEAOy1CwpodfLxzU7FLBx7E450zBP0i65+BEJeUAYvGNkAk+uJRXnZHz36q
Ew4txiMmnTEiTMZIZ6VgW0YfYBeGMNK8QeQ7KSBEH7tpbVoha5Ag0aZgmOE74i/+
vk6IyfExisV4rMM5mES6lqnJVrKYxWAWevKch8LX7wf8QrwvbWwREdLxERK0coqO
L4lDcM1GZbkupI5htFpaktFt5w//iOuYFQvFcBtggFVV/T2Dj/iVu+YKGO0tH4bW
lBAIKVN5SSt9KjiJFT3i0KMzYn5w+MqmtKYwPEqZbajTHBUr7Hsv+sgW1hw31W/e
nWliCwbITl2ixNFFkHXnkKBIn9O+Wnl47HCDY2zcON1AF7zDhypnvSque5jc6eQg
NojTczfKObyjJKYuVSC0XPNaVto3oC+UMDmWYmflFouYWYFXNbJdsqZRp+jAaE79
z8a+uX3Toi+93KQOk7F6mnRxDlUommaBvZufQz9uE6oU1mwbutrYf4wFlv6hJg7y
h9flL5tRAMgoBppqKT7W55tSxsuh2cTCCw+E0pVf3RcktUlGBVYPxMvcsTRAWKz2
T99LhBfbGLbqlxvy0Uhi4koeSbR2K8cijFtEErrPkRDO7dFXLwfPPtI41bebnplR
Ypiq+kZ7SKWQ8fK0gN2T/IOwObWYeM/qsCxBYgS5JMTvd4VNOy49cV+LkRWqIO/A
mUUmmIpkzz/H/1QKzdgIfRNPMJRC3YRl3XdzmqpEI34Wu2GeZHAJTgqiTKvkJ46U
T4O+7ORbIMS/IhrqDdGp4WThiGv1EcbLSfkOl6cu1FAFYAgXRswn07pCigN3VPeW
93DnDajycvGWWkeRWr/2+DirQy47gQhZ3MALrbdBVvV59hj2V/feA4OL08BGjv39
1WGrwXrPN3BySHhTcKv3rDuxcQak6m9DSMDxRtPzqrysCs7gXU1aGw/LeuB7pk0J
FGwsamr6wr0M6Ls2yjkOwmIL+Lixb7VhxVRhzu+7U+db7bafT4YFVLpv+HnRYYfF
xTnrS/xEa2LiDW0ZN4/AnZdTJ4twpbgA7Ri8DTd0PODxnLKVAGf7xodkvlWBRvB9
fbZhCTuAdJ5uhBTFsp/8jBfbXEcjt8j0YeFGHZzNEyc0iV5lxjIbpFM+Nl95qK0+
PiPP4DNAtW2pnObka4UJEmlIgmVCg+BNPXTEaX+jr1qfYjZ8q/Plmi3ky9h/jG8r
4eB2rSFwkY54TpDhH0N9B1TtlQUO9/yJs9siFB4//M5ZsbxBSNLSbKM5oyeUxG72
+SJ+O8OwMNduxL35ZUfqXudNmzfw7VJLNjBFhwucdQRGiYBFFVT/kSQ1O8DEAmrJ
zgWsYMjdR8YI3aSO+jb5G/0nLdiMKsMZkdDfi39bQ4w8vzjWauh6Lg71WZ4lG1hw
YZoxgcibCLIaIu+QcLPGTA1WirZs7KaQjcRaJE3VyOfOTT6pw1xxM9cI+ZlBYk05
9oaNU8YsMNKNyTY2f/Nwl0Sz3bH3fhcQ+J+Y1DYwIVAqZ70RoWx+aNBMWqUmhP7w
3O6kBhBxOXvp81XVXiVTX2DHL2BJ+2R9qou74C+i1Z2UocFenHt3booSUJ14dPOs
mgt63NyHgD9gu3mKgBCeH3BPATJh6DW9kHHZqeqaE4Q2TR+PqEk5BQYk0L6WFChz
LYg5etrw6SzXdmHZ4fy3NKDn4UhCap+M54OpTfArizs=
`protect end_protected