`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
ddtXksX2+yylW5zu6QL2Lhnb2d1sD00763mmSITNX595NcHTEkwn0zB1Dry37fOW
FufOhVzEJp80NC5qZ/+F0Vk7Ik02dIR0elf3clrjeJRK85K4e3Hoo4xn7YbFUIms
l/8VZSb14+JVGURjfswrIyCUotIzlzVYZ6gzoZwDXIi5gQIBf/gI+KxNXPaKV+PQ
Ufys/12rjO6aI/pPlqSm0hCvftmBcnezN2hk1UeXgOIuKZnogjOsf0iJVX2aOOWE
6pD/psybjbnsNB6kH5uFTA5frkzIzkzl5d9+YDm9OyC+k84E83I/7/j+rk4L2dah
QJOvksSIzN867/4Qt8qYTQ==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="MvBXkzurAa5VTw+1JJ70nePUfoQXBvZOku/SMmg4TwQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
oRtzZL4VJ4iwysPsC8SXYCzXS8Fw2gtZTOskLcDV+1B9Nzn1zTyNtlo6lNICRmmK
ZRVu2BmCc2G+fmzynYlNTnSa7C0Cuel6FYpxCBlOuk3OF2tzAmLAuDyOH3Z1Yjzk
a0aHuoCdIRKv7BrZCdALt03JeUmXKPdOmIlkVGFl8yw=
`protect rights_digest_method = "sha256"
`protect end_toolblock="Jn9CQpRhJt4rnzZPRk+dOpzAubz7omckX1MrFd4p81o="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 1776 )
`protect data_block
gD6l00tciPUa6pDNTk/+t0OO0nC/UTtBwLB41d4inuAUA3i/ALrNyoJVcBnAmEQW
ptbcNp5fxEUJjnOxnedyZEuEBxWRieZFQnkRdF269oPUJ/21X2FZrbGiwDbqSKJe
+fTHhuakj4tg2oTDlDGFm9LCgXEzcosrnAtSk3vSmgIR9fwwlnyULKcU+eMNerly
l43R7srAmHPudxMqPzMisPbMLo527xQmZ0Cp9iBBA1b/IBG0ezMOsrVa0pAhKvHo
bgjJHTDgzvrtOSaLU0snUTAcCm8uMzQzL9+v6mdNxPDERrOyo+XX6mcLkpci0QDD
X3hUytKBGxv3YIc6s1dCimAzv8KUfHjXEa7GcVfWqucraePEjC8ihumjeH2JycYm
qiKatFRKl3vAFQeaIQlOejzgavApf48d2Ue5QNHd0TDiSQUk0c6tY3yB8IM1z+gU
rNeLsukQBFyw/R1cKwBQ4HzSh6usXwQyR39xoEMmvMQKl+DHLJdjtyrVq9pMc1L8
lDxRW9fTGGpys9MVJmCHXSvyBs6w3ixXH52fuI6QvEPZLZecQJPtJ+Iv8O1bZ2t1
t3JXzo+aDAF7WQPoEdpeS3ia5VUVH6MhkE9+icUJ2hDvkTmDosnOtGxAZ3VPNQ5i
zNxsULQPK/2NzpKEWiQgxwEh0+fEntcaYpVWGSd9X97bp2xyO4LMpk+1SNNmZT6j
a3B3O9r8OIzeSVLAvzcvMlAUZamnuNnYRBQp6VXj53arh0Q7ss0TUj0T3Kj9jBNq
eLq0eoWkb6vDMTC8VWEwtqvSVjFl6x/0aOMyKaUHkQlWfiMwbLby9IQDOgs7Yvmt
T8bpNYDGOpd3R+tAodZ+S3AsCnCFky+MEUSBN/1iSZSSvjINVmeVtHpAoPvvkEki
R/G6jI3XtkSdH/hyMKE7s1xAaP3FqgUZFzE65iV2oqYWYuFDI0cZKGxm1QvZ+5ax
k4d4sVH9cpBtrTogmQzPWyJ/jdjX3Zei31wJ0+cB9PzmtAuPTRYcmuCibrlDg4j8
NnnsOMHM4nvEKsek9/aonzYCJBgzcZuQs25MuKUQJB7de7Vt3ezr0NadHFjHS91z
2z23nnXKlZAzLS//xPTCCDXfQn6a49wvfTrkiFfEoPA2KDJgYc4ydBbPc4qCfg9E
aB9fGpIEhlUQWfwc0MhwJAJu7kFD4We7Nm2JiOrhf46oZZSQiXQCPY1ewTfsbStK
mDCvbHLl6RmzilJibamUe61GYFdvkUPBy3dhdicwE69LcvQOjLC6D4cziNfwGpiy
9nRXQlbGBnQkCMBoyoHAHNNI/JzABL5VHdTQfJffZgkPZVpg8ixtxccLn8OECOSx
2LR+rROW7TUqG2XxRYAiDxXsVMHfS9DP/YRryjE6ojNgKqV3KcHDRCq+WKEHiAX8
GUWBUTJPsv/V5jwCUuGiNr1p4ZaoxuXPQCLOKRbfzR+NzAdTFsUsEuE+POQgVkZU
QE9wiEfE4uTwoF7g9w1YbmQd34Z/mMEbeBg440wcSdLv4OHYDiPDPtJ94yTTqlZ0
vSg+V+4Lc/U6RZrYRwwE+KbqE2odT+MKYmzGGlojOsmRSuT7XUL2LAL/hX8pTmEM
yvzBJoNSC5c57h7MyjtXSTLVceJgJKmGR91H4gzJlIPTsEkptj6y6Ug5fjhZKf5l
wVJnELqrbwdkIrguyPUk8rDydXtM9bxuiUslRik6c98vk8o4fPiWnEreNj3c5phB
78moL2NW0KVAdiWwP1nMIG4PWN9NACft/J5bAVgpBJ2mKXLnauOOV/1mFgLZRNWi
o7K4tyG/UfPerEEM5jy7LXetjH61KnbNA8Ed46umv+V5JrBhV4Lhm1FdZ8SB5UoQ
qD1t17xIvuqul0U5qt7igU5zIKIxgZv6Tej/TjiLrkcMKvvFc8AwUntDqImK5zjI
kbwwZiusub7Jao3C6yxo8aVG64BwgCT3BacySkbk5LO1Dmq/N2CRrxIPPRJUUSzv
Fa/EwQIY2643ZK1HSyz7NsXaaEMYAdmCFWIt5sugs6e89+QLgl0ymukG08eQ3Xnl
f5OxOUBcWC5gQIGJYg69YltP2B5NPBctsMl1leET2Ha0VeCMgfTsFNy5hdV1w8k8
nJ/w/GPPWAC1/ZiYQz3usVEmz1WddufWCIinEjSB8psP2zF8iLy6R/ZEgYOsStbM
tD+8lGmhQ3dGwwL+Osuolwvs07SyfQ+GanAtveMzzhKMPlpzBiWr+9kL5gtiUnCq
IYxu8szCrySWekPF/c2tzbqGVfgAnxsDB0fWON1ak04NMrztYSaeRU7J1VdoFGhT
XgmffmInMwglE5eZ0KNbLpFOpZ1z3ju/NwW/R3ejYi/CHVF8f/MN+VwtT7dgq0ZS
`protect end_protected