`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
ddtXksX2+yylW5zu6QL2Lhnb2d1sD00763mmSITNX595NcHTEkwn0zB1Dry37fOW
FufOhVzEJp80NC5qZ/+F0Vk7Ik02dIR0elf3clrjeJRK85K4e3Hoo4xn7YbFUIms
l/8VZSb14+JVGURjfswrIyCUotIzlzVYZ6gzoZwDXIi5gQIBf/gI+KxNXPaKV+PQ
Ufys/12rjO6aI/pPlqSm0hCvftmBcnezN2hk1UeXgOIuKZnogjOsf0iJVX2aOOWE
6pD/psybjbnsNB6kH5uFTA5frkzIzkzl5d9+YDm9OyC+k84E83I/7/j+rk4L2dah
QJOvksSIzN867/4Qt8qYTQ==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="MvBXkzurAa5VTw+1JJ70nePUfoQXBvZOku/SMmg4TwQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
oRtzZL4VJ4iwysPsC8SXYCzXS8Fw2gtZTOskLcDV+1B9Nzn1zTyNtlo6lNICRmmK
ZRVu2BmCc2G+fmzynYlNTnSa7C0Cuel6FYpxCBlOuk3OF2tzAmLAuDyOH3Z1Yjzk
a0aHuoCdIRKv7BrZCdALt03JeUmXKPdOmIlkVGFl8yw=
`protect rights_digest_method = "sha256"
`protect end_toolblock="Jn9CQpRhJt4rnzZPRk+dOpzAubz7omckX1MrFd4p81o="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 2848 )
`protect data_block
gD6l00tciPUa6pDNTk/+t0OO0nC/UTtBwLB41d4inuAUA3i/ALrNyoJVcBnAmEQW
ptbcNp5fxEUJjnOxnedyZEuEBxWRieZFQnkRdF269oPBR20CDplsG7fa/LzC8Sc4
RjVMErUqYTfKDyphoeUqwS91+6S2WcNpCjk26FbdR1jVtP93l2cfCYT2mznXk+jI
pzMI10B204+B0IBFjbRXu+QKtzxhIhaqwBedUcVUV33lCLZY57eJ3199si6Ue1D/
v8J2tUM2gTmETv/omz0WwFCrtmgivPmyjFkiDgGQhKdH0M29AKnfyvsqysyuLdyj
GnHOGkQnVaZViwUWgNK6QqPSOmdhKaIazCBYGJo6/FCTw/CKFRMSMz6NCMpX/v8o
k63VQgf3TO1QFFiQh1X6wNLcwUu74G3xpMBey8SHo9/V+HgPDvCwviY2Qt8ueNcL
u6839jKf3E9SbfQbngs+DYCDXISMQ7U3hhfpENQIweAlKH34kYTNNb81+HfqieHK
D4MrTtnG5QhLhsf8ErCz/97pQ/ivxOVjx3quBmaoz8uovDbZWmfawlPJBo/tECGT
X+GVRN4WQPKLird/y7U+CH2r0cZ+Btn1+SUCFoufhPwqpHnfYuwM/5lHB2kSoo44
A7DxXcEiXMZHWsQPMWHZp90G6/ECSPXFRz9uyu4Nf4bebuqLJviwA3rfUS8QsaTx
b7iM3ZXOCICVAmV/BGzVJrMAVxCa5yMgwt4/qAjTYGtPcNpr9jYXP9aQI5tb55Or
famH3YA1rYObe+oj11IPw6WNe4GtcUC8SZglXv8fvl/eB2hBkXaizlzHzci96kso
gqV+H5OVk7IUoFo4+j/yZAzJXE+fcCCzCBKpjuhLMe0ysIfUi68N48siplZfUe6T
8nOSE0wfnbK6TPMvHzVqjXjRLLZ6mRr4++hMhgG1E/QKRAvE1vLJN+w+8fxxyzYH
SNVXXpkiso5qrjOSc8S5HaSPPVTf+WSsDC7a5BPy04BmjC+G80mrI2kKFbUHYFkp
eGiAsvYlM/zr7ROyBnbSjV/oFoCWYhT890henbhUCCupnfHobxe1XpOnyvrTz4b0
K63lph4I4t74cQKuk0TKIlvxARSbIKST2fYMnsifd0bsL7HOSjDTcA5NbkN49n27
rWG2s0qYfwRlCdiWxW3cLSHCskiZhYEJnzrLsE+ytUw9sJwCP45nrFkdR8uC03Vj
ku7t+s5AFIjW4MNE/2Fxue8qN+0SRXk9vb5R9j6V5PV371WOEM6rM7CBwnlMunyQ
lqDgANOL4c8505qyM1QlAzqW9hCBM63rJNMrMXjnPIWMxW3IndAW4klG5cD/Gkhv
sZsiGJh1qm59XEiERdbM7sMrW3BCbAbibk3dlH6r+MbIOnszCkGANjalsJXtAQ+s
WNVlavmCIuNNcNmfW1CihcvrMyy5C/eK7qkeOaQfjDampB1t4h/192LhW/Zh4/k5
29fRPtrD5whUGuKkB/iPivvSV0PYnSF4oRbadItGFd9FYqAD9b655mYbf3gqEGU9
tvRWUDI75QQ2gPgx6ZuGzv9rvZxSLaTIHSQoszULqbuKdCKyH8mZeIsWQQfepmEL
tLFPxxStYez66IB6+uyZzDDVE4brx9QH4OhzJub6o/uEB9WrkczXNpqufgDKrED6
GFBt16TneaDwXOdU7CmI2pGorvxux+iGk1rWzcw0CgajUEdtNYQDyTDWdLxAR8yo
rxD0Zp7MUmva356JGesPT8pKngRZhyx+lTxUtwcAf8jZc1P1AJzrHmu74bYzgIN7
NaLLVbwAYRNuRap+ImQ5ZPAlf3xbzIE/mTftPCJQ66DvKqk0zbcSpAE4HTlf+bvE
HzYd9WyP3gzOFQr1GoSRwFkWV22otTHFCkRGCF8D52oA1qzo6ihZctS3R8Ldfg4n
mRBOBwHz4K4AzOcTJMUuaBKj3GZ6DvNyuJZOeiDtGL89n316RnNzAaAlJDUUY3i+
nPP53+oFfGAKpd9LNq5nQhjjULL5EMsM3/u6tQLZLgXPURxJE9JYioZaFRKNLr1A
OXPNVgHygOHBGpJSlANDitbKK+g91mOyi74baKgjl576iiX+kOjAHtv8nZ6PInT+
v7CZw2k3/BxYhZmx4H+s1ejGHdEv+uWjxd/9vdvK6QoA2CoJOHnB6N0Z2iuFtxTW
5qdNYWKFg/W1hy4V1sDe+jmgV5q200bqX6hEg02DGTypF3y+hc5BJBZ72Q8v+1mR
uaGPaJTy4s/8xqivgfLIRBrY5xg5R5+taIb+musZIxUEjZ5hkY6M8Wo/63g9E2zS
MrnOgeplNuu3G2+3iDByqz2H7QBThTsw0UBZEb1rGc8RttA6LZtNhflkwN+qwnMs
XybyxjLyifhpatXkYBzsbNGWlSbQSyqpWejtEJz/QjmqyQMl90wgqWTF06ZUpM1h
VTNn73MfkGcZ7CK0JzvH8FXih9mb7C+Zyokh0qkxKfJEmH8fv+k9hwVLxToazVq0
Rg8b0OTYbdXGMUKM5i5AI0RngsYFDvT1ERBeM6+1QEV9yYHYpayCrGaSM/o+CZrv
U6IztZ5aBoDK7qc4D6E2Id9p0HqxL/9p3U8V9sqn+ANac8Li87ew2MrUYwintuta
83N4RrqO6d3eYcc5WLZm2Uo9QW+3XRO0QZGcYPysYfJQ4bJiLuydpNj6K6RAQhmG
62fmdHyr9ZXzAm4gFRcbmx/82UKjjrbM72EJm7ZGybyE0fh0FD75yE9VObjzCTBg
xUITGd8LsZCuFdJztCyt2ZIW0yfqiL/WmBIW9rSv/ohfyKfDAu/VY0l5wl2xNLMf
Gw4MqO3ZbW3Omb8xE+Zm3djordC5+WHSfYhWGd+OpEIq1/0+zAVtz41Vu2ScNyS2
2ch5Xtqq7IweKS0Y+XwqlgaFmsG7nLmjbY7PI0bNS5y3BczOMmPCwOguuNAcYkEJ
9QcOtnMi/blDj2c053xw2zPzOGPrgVxBcGpybhTzer7MPUCK1ALpQkWnaYSEIfSr
5ZXhcNDdAbzLWjJe/qHqTe6PIRwC9jE91o8xIF5oiloSdHnekGuhMUmvDCvdJ9iQ
mM98xH3TUyXMMkuuLD/N3i+ouwXtat37JRqJor5FqjlgWcEg6yRIvWP7mOToQKG4
FCui8gHnvWKtTCKcFS3E6C7xZbZnvp63yF7HkWzqiIaUJCvca5VmhpPpHNnzPF+o
7W7DJnZ1WE23ul1V4KW3y53CcCVHintAfzD7DabVN/YjiKDw/o/+f361BCiXEttI
j7aX4wvmfwp9KNLFHc8jR94tnFprUZpjJ6aVhblJcomYNm4eeR9hiw83RmYyXO9C
WE+PjR4LCMlHWf4LwWg6ojsWQ80SfDd5QVRx4J5UqqedaTXJTxk3BkwqC/wUrXGw
sF7bJEJltP8zVX72zPYo95tx8g4YdeaNkW6tJH9qdGXjq8WW4mAAlQj6jvyYl7O4
I0v+lZoBdCQXUkE9lZ9vgvGSZjhn6HZFMu2YcrajPB/T43LZMuV/UEkymnKaQiNz
xEJ3qPimydadHPnl0zyuNCNCgs63PNTnObHo32Br7luaOvoWakAvdppLNG25ohdZ
3csVnjj9pKFXdRXYwGkZx33Qlc4AT+/eo9M0qcs1H12cx+GNtAmAeJv80odxP54W
+pSS0kI7uq+4i6ZAOUZR9RLgZYq3UN22t/I/QR10hJOU7Y/UrKm7YzJd4d9XI7ZQ
EmE/fjq49UrTLRB2T/0xkIh5WNzCvOSNbTrtStzW0Iea6w5E/pUAdP9c3Kqrak7m
jkeoyj6xcujLy/8coZIxqQ==
`protect end_protected