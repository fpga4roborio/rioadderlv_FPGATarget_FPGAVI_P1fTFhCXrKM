`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
ddtXksX2+yylW5zu6QL2Lhnb2d1sD00763mmSITNX595NcHTEkwn0zB1Dry37fOW
FufOhVzEJp80NC5qZ/+F0Vk7Ik02dIR0elf3clrjeJRK85K4e3Hoo4xn7YbFUIms
l/8VZSb14+JVGURjfswrIyCUotIzlzVYZ6gzoZwDXIi5gQIBf/gI+KxNXPaKV+PQ
Ufys/12rjO6aI/pPlqSm0hCvftmBcnezN2hk1UeXgOIuKZnogjOsf0iJVX2aOOWE
6pD/psybjbnsNB6kH5uFTA5frkzIzkzl5d9+YDm9OyC+k84E83I/7/j+rk4L2dah
QJOvksSIzN867/4Qt8qYTQ==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="MvBXkzurAa5VTw+1JJ70nePUfoQXBvZOku/SMmg4TwQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
oRtzZL4VJ4iwysPsC8SXYCzXS8Fw2gtZTOskLcDV+1B9Nzn1zTyNtlo6lNICRmmK
ZRVu2BmCc2G+fmzynYlNTnSa7C0Cuel6FYpxCBlOuk3OF2tzAmLAuDyOH3Z1Yjzk
a0aHuoCdIRKv7BrZCdALt03JeUmXKPdOmIlkVGFl8yw=
`protect rights_digest_method = "sha256"
`protect end_toolblock="Jn9CQpRhJt4rnzZPRk+dOpzAubz7omckX1MrFd4p81o="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 3536 )
`protect data_block
gD6l00tciPUa6pDNTk/+t0OO0nC/UTtBwLB41d4inuAUA3i/ALrNyoJVcBnAmEQW
ptbcNp5fxEUJjnOxnedyZEuEBxWRieZFQnkRdF269oMBorCW1CTe3kJYEo1SA+EK
suevAsRAF/oTUS5+76Ce2BM7pQRVtwmbQUu4PQ5KLRt/LsZTYCYDyJ8Ag0Pyekty
uIYvqwnQOx7LX+JvwKI5zauFUQYBqMvqmGjKzDxDIFR2aIQHadFHbCss6Ckvpvau
J2HPiPmYvxPblknWtXoN+GsD8dQ67hCFXFmqTabrWt3EYwrlFs2WKhz86cgZJCst
MxY/GQ0zS8aP3h0FJUpLrPBkaHW9t/6kTitRqO+nlKnf0xDa9Z26RNoQmtsjDfL0
KE30zGjqH1QR3arhMy5LPS70FSDCoZQ8TctdtXu9fZnzLC7zdxcYn9TyDvmh1jdY
k8CFUcJKYiAoOYhgwpWHXJV1TykEBvT8zXfyzUnCaIMs1m2K6CpdatRoRm8zbWCu
2F7GmhjVdKbmzl0FF9DsxWF6IgQnE6YAz0bIG3L1k9sBt4g2sq0I1dd9V0rbC9nv
1j83ePGP/obZX6jeXWWLNU3X5ayggJxABt8IfeNvMwttto40d/9eMu6FCdCdM8qS
zb3zHYukWqgjmCH4GKbCXmO4NzxxB8gXgX6mFRC56vuqRC8G0yjhKrQwp0/SApGu
eNED+hkraHGdDOaFMlGSTcT2NUuX9oUfS7iHZ3dRiE8sjVkFl5QtbrMmCU8Vkxbl
KGGfFRFIo8r8GEie3KJp9fzEHtk6ldwS6dhH5ucp4SBZ6PBAksjEJeaM+Yi0lCMY
j7ueeg0NKvWjnKw29dEbXehHfdeyB9V95qSnGDZ6rZnTSaH6jalEFt/Q/NadnS+k
3BN8kWzuWp6H5TjzoXU8DsVzTz7AR5f2gJT8osoWP3UnFIW+q4ANHMrcsfc7VABn
WkRjBTmQuOlSsswTHds/T9/5StPmq+51KuzvL3oU1piXDIVQHrM4sGt5LQHXBND4
Lmj58P1PVZkMlg/6Y+KcsLQbevNylZIRlq2Fg1wBMJ+fdDLMQds4LUGEyxPg4Ebi
zTWR55Cs9NHOzyP/Ts2hs08MOUsjohSpDVIbfim9EU67ERCANnjfsVVYtFLYnolw
71/4H+hCrBm/depZuIfGzX5EWCaxPpreMOn2wzCJpaTHLTCA0fCVWE8kaizMpAZL
hcXueAm41j01llvQZ+AAGB1xiasOUn+X/E8cq0kvTs8FYeFxUKNf5/yx1uzvvCwS
YX45MuuAOGl8U/oVzzGtXF52S/IbISqS1n/pY/7IfEXozMJ/34YsW9svQtZT33rc
nYAEFNTs7l3gonsmWzoNpLl3NNHLPEeSw43F8x1wvI+RZFvfIE3cg1s5+0xCjtK3
Jaahn/INVt5d9OYJBfBzETemu0ZO5tvvwwCKUa70wpwgjzqCaLTlRJYCPXjnLQtp
Lg/Tke+yhtu1uGLY2saVWgvGhe+pEcvL0TqKBxYiVni6Ysqf1IubquAhbS7yJhp5
YjBORERJD8LZ1xPGj6guXorc/CDMAEOAL8vCuzU6lQn+AXViI0Aw9pjamPOOqGwN
8VOQ7j9i0n/Y+iWGtwwopv+AyZjgjpThCSN7Dzd09ogajCriUn9VZDDMV0tJtHp3
8c2OtQlMLbM/nw4midXstnfPG/x0OfDyDwbc9JPeTdzTVOvJzhLGGDpuf7z8X1/V
xA4+4aqug/DRgMawagishKMYgfVHSyJAPnPAjt6rlShy7JzVCKtKx7TzGLZvsa9K
zPbO3Eb+/rabYYeMOLhFg0DIi4B/TyeaVypb9eOh5maCrse2h/5aBL+3SoVs/JFp
YfvhD9iIB4ia3PE4AmiI5rSpF68feiFNhZyjadFOAifDCKYCXmj1jqRYSLQp6Qmo
okzVjJCy3xVWkY3BQD7kRDne5oWecS0e2RjYyZMkw0/Po5fosluitWOpL1rooab8
l75/oQwFdAs2z1CavbC9Q2ImbBa/IbY/oyXnIhUOdlOK3OdS7JcEU1s5dZBO/WLL
MFgZcDwvAffc5h1ZvJOM1/Ps3GyX8ym0NlTt3I3PeWvXJ39WYV2+/KsHHGllMMJS
atRZaE0ipigxMFEVwR3pHeiQd60cEpy9QaeqvIverDD6JwfstEoeIPll1O0XRml0
cTwoPajjg8u9/+UZ+2sq4f/fXw3/VCx/WDq1NjOJ5m6DUUyv6/cCZ9TYS22VwuH3
bb3pQRi49QfSnYEM+zEEORuCsGO5NPF5uaBIYTvFC1cQui2EW071TQJaGCV+3F1A
SOzsbnhyuIa23HH9FEx9D0i1IlsY7FIaosUxMvnm2oVc/WCt7Zkhkk3RByGsj1lP
vuakdedGmalbUP/jPyS95qTyOG3bwhCS3WA390bZxGNjW4vcDP4eNtypXIWE4F/W
BN6z3in4mbJjFmTaxj5RBAP8L54yBA2N5W9wRDfaEbzVXFfS/mQDOj4O9WBqiQKT
9NgZwRrstn5D4rknut5j7LHYsMQ8RkWwU3kSUM4KofwhgF+ymiSXqAyeDSYU8RC2
/++fLOcLF30LLxJFa7P73JRuRwEX0EjbPIwVvDOSMtLlG4UhlKGglClUHWQFQK1c
dB5FRHSxw+lKbq5vRrmElzkg6DvpREmOB/2m3yFUYr3SKY1bXJEvgE3Tm7TBgnjr
bf0YAfF3vgnRZn6vfy/2se9VbB633hf/nPE1fECYEXhmf3kW1MJ053z4yDLUP1LD
nHiezYek0nhdMbcFj9ophTa7uLIMKwruZ1hoYDdVd+kQrdNKzKyvKf9+7OTIOZ/W
ssyd9Flwn0rFr4v5SHwJzwkU0YPDh4n4eVbvvYhfrvF49kaPH2ZtPgI80aZtGpPe
PYZJOP6Oe0KTgXy9Wmf1UaCiGIlkc5AQY/YkmB4ncpCDpoWOr0zs7L9zsAtdTM61
ucdOTW+SQ+7DG+QZAxJ8qseUgOCWjbR6BgxeoRVhH5ECqTYTDVoxw4AFQEbUHPqp
+cifSpGDKhENSRW9MIE5NELwZZQ8MpUVAdLPjBPrNv1XbrLQoMHMQvpUKQxUZpts
cIpdJe0lTurl9W0pSkH4rqS2DXJy1kbfD/LjLChQ9Dnv0f9XmCJHM7Mwu5M6qpRQ
f3qL0z0jhtspPfLHPLOQok4exjv9YutHLX1zWK0Y0YxolcXbjzPBgmbDrTNepZUb
4m2DuPoUCG/RaaU3mnqU1nQ7kQLORj5Qkdqz+CrrTzUZVCs/BvN9fgvpuTtwWC61
5Nfy7iOR21udsxk0pKyecGxi4duO0nPddIMEY9UaFlPkS0b34MCbQforENpMcgZu
QPjxP5NYjXa85hChDZz2C21d4COtLkA5kWjNiRiH8d8I1q0cAf2NoKF+UeI/onps
6Cde24LQL4TSAYTXOEGnqUVTip3w5lSu1tNLDltEeiRyOSej9m7/g7KKrd2fCjY+
9mvuKDk7GHK/3U1zaK/HBqnAP9Gve116YVPfHOVU9z2+sF5rrd/MjXWiKOW67JGv
sgRa6fhvvuRdslH8Sp6hPmyN1rRjtSfIng242n7ztYj0ijVdT1tfSghmNBizvh7t
tW+lEl6wMJEqErHF/IB5UMbEDtxPCXZjUw1mv5S7/qhhDh5PKSYldtU1D0JqEhSd
VEe8bNdeIrphqHq1cSaoHtkHI+OOUfQ5R3Y0qkX8uPMCYwj7rZJP3qqu+Kfmi3FJ
2zQz6VA9p3abm5B8CsZG1YCAmqJq0Dm4zDJIhtU7T525268MkhF4QFR9WDxGO3i8
8KJ54+Fnajq5xWa5qMhFKBoClc0Bi/yZMH8LQs/K/kCweRfMgNNTk9FFIFm1Dpv0
/Q27VZ3y1mKrzUUtBMZdKH824zXeSieufh1iTMUqAmUQksOXAZHxZz/bVGcz9/xt
Ey0Sisq0nv/sdJJW3lwfCdTzczUGd3YJ3SEwQmhMFVMid98tXVDU3a06IGoAJdty
qGOFzuDioMbVGbIgOSGwys0vQJZaj/pqMVYS0SaYwoCLRkW3ZrwVGjnauHg98vJk
+mO7Fz9gUpvOS0A4e7Kqgy8lHBAePgxaZsV6CKrd4xdZhiZEILeUTOMo2GXu0+1Q
g2CTpWqUQbPjGTF6qMH7lsHNJAD0p0RJNUG8YYgnoZob3G73FdnrKGINtjpT9Uvg
cudWhimIc9oVr6VmcvyEOruO4bm2QMi4WQsn1wSMh30SCxfrgqekXvF/cjdxBxus
Xd3K7C+8EAULIYcuRLJIkIKFa1CRGtcRJu2Izfy/RzZA3YBBSGArDLppeMddL7Uw
JANQ+hhEyzgIEDiYzFojXNe0+/yMBqU/KEiafIBCdq1SX9jOACjLiUlKI/f4z73Z
05cQi9QxYdwBBxpsGvt1v6+mjHScVlnm8WJUJEP0MVk44zv88w28Rlknqi5TBU+x
iesnSm8/B0vcRr06bgPGAwY//zWnDkaShYH0IUravsYG7SDPN+7zNf2/PnElMSXl
dxBjSw/rzg9gSz9SvSJNGQ2ZhTMih3AHd9b0WsZd8Vqc3EAM+FP+cwB0ZypJWkfz
rZ2HlHSO8GAvOCZL6u8fDJUSWkSa8xA7BE36MYPqn/z6TI2FT3uyqEZXwxWiMg/T
GHvONhAolaot2GbzmNv1e7zauHB3ZJv/cYZKEeJGqvr9ubUhFNyjkw2ooQOm/x8n
Qq78jgcN3GxKpIZYtSZLESpnrHQVaCTuOd+cv6SkC9g=
`protect end_protected