`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
ddtXksX2+yylW5zu6QL2Lhnb2d1sD00763mmSITNX595NcHTEkwn0zB1Dry37fOW
FufOhVzEJp80NC5qZ/+F0Vk7Ik02dIR0elf3clrjeJRK85K4e3Hoo4xn7YbFUIms
l/8VZSb14+JVGURjfswrIyCUotIzlzVYZ6gzoZwDXIi5gQIBf/gI+KxNXPaKV+PQ
Ufys/12rjO6aI/pPlqSm0hCvftmBcnezN2hk1UeXgOIuKZnogjOsf0iJVX2aOOWE
6pD/psybjbnsNB6kH5uFTA5frkzIzkzl5d9+YDm9OyC+k84E83I/7/j+rk4L2dah
QJOvksSIzN867/4Qt8qYTQ==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="MvBXkzurAa5VTw+1JJ70nePUfoQXBvZOku/SMmg4TwQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
oRtzZL4VJ4iwysPsC8SXYCzXS8Fw2gtZTOskLcDV+1B9Nzn1zTyNtlo6lNICRmmK
ZRVu2BmCc2G+fmzynYlNTnSa7C0Cuel6FYpxCBlOuk3OF2tzAmLAuDyOH3Z1Yjzk
a0aHuoCdIRKv7BrZCdALt03JeUmXKPdOmIlkVGFl8yw=
`protect rights_digest_method = "sha256"
`protect end_toolblock="Jn9CQpRhJt4rnzZPRk+dOpzAubz7omckX1MrFd4p81o="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 15008 )
`protect data_block
gD6l00tciPUa6pDNTk/+t0OO0nC/UTtBwLB41d4inuAUA3i/ALrNyoJVcBnAmEQW
ptbcNp5fxEUJjnOxnedyZEuEBxWRieZFQnkRdF269oNiNwOtjqEgrTRkUo4Fd6k8
0DnWOq48K0AcsIOEhn7psV40+6Q2C/P+OJMx6hQZkZnnEXbgD90md2twB70Xo2XD
K4iD8+FpHg68UgUB9hS0aWA+TSwKZTmI6PbePkGf6l67mPCbwo57emeyaonojj9h
LMsLnxygZz/yJoTH4ze7I9pxjWQCXWsnaxzJsxupUpLTmdsIjgYHixdRHHRwRdlB
d546jcnvBlYpxAZXfpgayNcKu0C9/KglZ+t0A2E13xHsO28yS7Xv765BQai2+OrR
HQ5ZDbwLqtI9pY64RbN6QGPsr4/rBZH9Ptj/eM1t0OIDsAIdikFmrLibbjTjzF7n
SBemItuOEHzm3eD6c7g1HdCt7npN3+p9Nn5zwclDWabHHLwsfY7lOCx8chgi/Np2
eBgjqygIdgTbv9sXhyqre8N8cKz8QWmRIpkNBpzUD3yuvgcBE39i4sT1P27QJ/S0
M9EhLI5M0qzWluUJeRb/4KxWujqSpwd3l5GREA8Rm7BK8SLj+qxxQdDYlQB18aSJ
O17yJfH+0m9vX5YIxr4ojYTaKGXN5L1wnC/BnHh7SGwnQPDD5vZ5UT8WWveuKw8g
kypNV+u8abG3kt3Y3dBIZWBVj1LMjYzUPnmW8Bs2K1Rq5MSnL7Ur0JJvIgamBoZS
U3kSzd1lJ2xvW8FQ1LCfcZzsMrXnHUCL7ip2DXLvPie4PfGMhGa0+gxqmRVt/OfO
XBzpHZh5P+jKqRxS3LedC19kQ/RvDCMonH5IziLbSpLIxxAfkcB1LZBOTI18b0rz
nY7Y4kcSueHM4DWkhDoMewoc7mcNyrmaPLwfJ3j1f01yRj6K0S+whOg9yvdM5c9N
euY6JPMnhN6yVWHGCKl9Gh5xkd6RDNVpFtWnseJbUbwnxontTO/htqca/N8U1c8i
RRaMFl52zjKfSjfR6zVkMNHsyuy5Ru1AtQ65V8elHkbQdH4dTEEOtHI4PP9Se6zr
PYBxUZCoXxILcvGb0XujH/QNSR8ErSAArWFWlXFy93UsDJCHE7ZmZ0vS1ncGEJp0
J3AiJiTgHvug0kkPPQ0aAAFgSjKnxH780tfuhriPdxNUaKFlQgBa40cFmb2mOg3j
XFqdslwph2ee7j8ZLX5FlcgOxaXPyGMHKcFjG0kotITRwyl3rTJGDi6yMtEl76IC
GHyByzfVmDhfzMkysSEs0MFX9nUM/MttREn4Ykwl4M9ZM+V1noFFYCerRXMUcjLE
F7aZI6f/GI//q7PcpCH36ASJZaP3x8QfGMd/U7HigaBylMGvhsZJHmAPpdbE3vH5
K8ZBMCuGjRvmzK2mYvlkiYT/0GewkuIFVCKYto1UaFpymjtTY2pikp3UXv2fAIwP
T+/pNIUhAdffdKs3+xANqCsyWFg8czuuPU19/woIA63jS4EvCLCstpQxUc6Lor6f
dhfObvRwh9r9RK2YH8myFdfDVfNr+B1Hc9mVWsEolVQBv3bo9sZ701Ldrmogwr5v
nKdrIp1/1qbsqUI6ErhfZGu2IGAMcyRKoFdo6RZMHE0S7aMJw6BJMz6OfLiEvtDz
egnhZ89RNVugYhTWYmWh1IdX2e2oGitgOR9u8L5M4ecIlWD9jzzLjRVXNWc9fWwY
UjxVw3w5+mkU472Mmj2c1xSB54NorGIzfddLQh+sl9CWu/YYuMfftNmyMZ95hjpP
0pZ9qVDgWoIMlPBfTvDkI+QopeX6brhMHn1jPPF4Ki33ekCmIT71QM8kl+xH1FZs
xHC7UgQE7oGdg/BxMe5xNo6g3v8FsKRfvw4XU7155rSSvycZHzRY52yJfMrT3ZKP
mrweg4ebWX6F/Jv8YMr9EM9+W0FIQ5L+g6GQCS+jfrU8wB0Uo3RxNX/HVCNWH4ys
Fgwb0Y4RF3wIiT7prDpsvrULfB3tlNIUsV0MCFCfi669KsdztJ6qjl7Hvx4tWc+H
nPW9VeWLIbAakOB0DACJk5l+IJBwP5dgKI6hGrCajaOpjbpJhSnBfRYarBUXK5Jq
00TUJBmwtvFz5bmS+bXVciM9cOjYkNJ0IIotfDaHhKJ3QKApp1XV3KzxZlD0wtvf
iEJI0T+1v6bRgMc8cEUlCQ4emF7BAypCT20bj8K+4WQIaThDtNpGMmLccHYCfYkd
jKITET4KGCbUZkyTipQXC819+7X/p6nph15yn66OQ+vgxplYTKaZOut5tJiY8zBG
yOz5d/NCJTEX36XsBictLImzjW5ON/+HNfVnCOKTBuSq18WuN3dOqDXkUKGDG5SR
O0ukNZlNN0suEDLmtWILNK+zh/mRKUcPNSqXxMpCsNHduuhPnlfC6Z8Yrv9hbICH
nIp7tMv/geocOSU//li8N+By6EwD1lBQZbNsqkYL18ztRxIbguHHO3i2sfsXKNYZ
y1FEEbAGsEOCqZhMOIga1qhx+/zMAvxFlXkuYYU0nqioFyZqo/reYPfgCIZNQxVx
YLwngrReQ99eVpssKxrURIBhvNzWl02m2UVCvCfkIOR70YPm9OYCy5c0JDEe1WwV
oYZuEHgtzv79PaZYUBnggCpRpnC323JLJhpmm2QmupI+rBVozFQG0+G57Hu1xKpF
XdomK2rtN/BruUJP3ATd8rjWIjCGhPHjieqF2OAaUMcyDssuRTLLP0++Gs7xNoaK
G0n/lDrCbZIrRT6wxxIYcgas95bB0NvmxNH6Wv/m1VSo4VNzST/P3xo6LuwTRhzR
vmDTc0/chV3VQtNgg6mshsPnpQLZvNsJtzcDPygjPv6zHBaCfgJ19FaVNAJ0lw38
tjPq1Xalyk6uaP3wtkd4HgDGmAGWWbwr4Y/tAr4oRR0jOtWzGGVW6l8mz+izzAq3
zWC3FJxBwEQryh7KJIn2ciPKzc6qPmoOpocUtTlGf4kBK7lqhBlou4H80UIFnuMh
XMmYmgTUwx9NdryEWPLKTDj0wv1htw2088vjsBGCuGQm4JFNiXX6TTNaAzRDPzec
A6k6Q8t5u6TnaRTB6qsYJvltGcLd2S+x0GETtJMkbbCh1YNmJ0eFE1W0+QuNtF3x
pd3tm046Q5qR8MEQP0F26NLIEm5SGE13lxs57Zg3RIVMKsONpguL2oWhnmuYCr2x
hFs1Nf0rKKcuvEcEMlmZgM/Gz9K3gQekysdUxawo0OPFw0RH6b5z2vfQNAyVMbkk
3W5jDyJBuEsJJNxnh13nYL7mA1PdFxIutXpBAvM5qjlTA7vm2f7yikIIUBXSSfho
VFpQWaOz7h6Oeul2uQ1s/eyBCCtze4+Zuc9p9MQe39qHtB1WWzYBkrFNs1cgD3V2
ZgAJOablcJHIaMCXchxtgID/yWg4ZtmhFsPeGcK34q6ts2sKiOmC/AqhaXyDncLn
ALGip1Hwl2hyKEcQ/sWkYClKj1JahtA9Bp4U3j3lxtr/BpKAhcd1VL5tkDraHlKY
7rjdTqOCMsAdkgmDanxF3YF/fC5bCGJmvxxRMT989wPJVkJs3d8LWzjtn7f80ZO8
CA9eRl7Yq5lzIN05yLkcBmMhal7ItCl8sPzYj1MJ34SOXIeQttc/5R2OkFnCP+q2
BhlGMLUmgJJ5Ob3JDGh+sXTmGbQvZduzElE4Lm5E/DHJNQf6Cmao3MP2l2F0nSy3
5XEFVtRdFRI/vY06XrkLH++v/5x/g9TBJk5UhP2h7KZzEvVFbEAMMLUax5ys8RxA
JTGOgxOiRPL8v76HLMWRfjtHskqUaA3z2mLY486pV46CTtG/4+entzcl0o2Ve7jO
SwIuuDjw/kxFEQtclQeNPV/Rbj5eCVw08a7O8eg/xMp2ueUT5QREDaq2j0M3yPj+
kLpJdqunwjmj10GZ64HPvLaPydCVEMNuiv0Il0IPS6M7ZdhAdQ4almh+f5yULik2
6TiMGzYJsmaFCuTuiH0p+vGcvaZeM/G8auBrTSKGOMJtUE9i1TAot207N/tKkfmb
BL041yuFACvh67QpKS7c+kGRqLC7c+69IMuycgcxflYXAQD4qmW/TeV60ij83I1f
Wa95c/DfuNBFFd1EneRfUZuEYStRZYbtTerGCxFrTZPa7hQ2NaJ7mNZjMU+zK25F
MZv1IC54wfgE/AnrE4mFlZ/vvoYgQQ70szn+O5uPkQu2oGugXOuL2Uf8qNkFcvj1
qttNR6Yhtn9Jb2FZQ9vK9Och/8wx8fLGL/lue2HCF4wI1cdrpA69GTK6sy23hq+R
rKBqrs0aTn3YJyVqTygP/A3o7CK7SEudH1h//zvaxpFbkOJ326mV859ZoxSabLvD
pWSZhkJt0fzpoezWqguDuRzW1EmVjaUJ2y6JBk5s7BipDMeSm5IpYqT8NASXHoht
24fzHpaiUH/QZ1PfZN/FodiD5W9O1f0D6XJsqMl+9gksstwc+MdjpCv1c6c5YciR
h3x4i75FSB1yoGXfPiVkFuhv/ng+Smy7mk5jpqjUJr0CzoNxy0soUluNxrptkYyv
e36N4LejXjkAHfu5QXCHqp4/fvm/XQxYpgyIWTnp/IAc/0BG294pZ3VfhOl+iJwn
rrmLvUPf4thr/szqU1/5mTxwDn/ukgbyU5tLjhcfj/LcE1mYgR27v0LJdgiPe5Tg
XuPtAilwt3WZVOal38TjrFMr0ljKwUBKj6LIx6MnMdCAM0bggkzxdzVULyev/oRs
3QurRiSSIdkEJzfAuxezAID5qQlAL5tFFHJH4KW3jD8nPd9T4mXkUdE2oVjluSUu
IvPJxqPjRgO8cDWEzfMtioHM6BMUY0aOYCVOgjS32G05ixqj8DOpdsLD9JG7UcTE
QJ1epAYf/4Yv/NHAGZ8XgM9kZHq7Yn9bsEdmPqmncCwiWyo4LeYX+briAYwLJky5
nAzoi5U4RycQwSYF2Hzbc35iXc5TFGXv5k73/WAgxXuq66Y0VU5g/hdMlFYORl8+
8sKPFxgUROqxXWu72Y/jmkg36UOAJET9kl1edmG6Acleu9EKSejdCg0iiD79eBBm
0Q9mMUVPcNgFBkUveh4UIqLIiTQDd4XKq7JdmSLa0WRpgQDfFcCnbix3egIsWzdz
+o1t3g4M7flY+/qn7RsG5pij981Foa2YEh4c+MYQhUvoj5AG+//IpmWlvUv0miEw
+tc1+g3u/bsQ9w8t4E03GtGTHq2F0foxvcUPvNDn91TmYUgJqy9cnZ98Ly4Wi3RC
O3Fkts9W6VDCxsUKlYuXUpNPYj59ShVDLCf6gfO5OGSOE/nRBcQ/pF6/6ay27lv/
RQk8po8HvOeWcawJJui/iZtfZvtCWuIYIv5ZGuKIy/7CFjAL/NR0bGmu0GxE/Gwx
fjfDk0tUcf4Gmt2kflKCGD3MI1+SPW5AF+XVdH2aCKQxNwmyr958OTQd+wgljbqm
FF9ELbjbt9u8mrvfBUEQTX4dYpgpTxseLekU06CuF7vVFK+YdegDiCL0aqEupqDD
YVDDarazTTabiU+827IHwfvHSFkJuI+i9lRAZyFaWN9YufsNT6oKvnBUUcEhKyrM
LMpNvgduqseJOwMzU6zv6LvDa3eMiLBCfYPOuWYbX2A1TZYYWpiY9TU1M4hDwmN5
4r9JB4qiG07Yjq1e7cIU3QlCkyXhrpix82GjPYqLxG4Vd92DIsUQnYqrDwPT+2bN
qXwb+sfgU5eKfDGODpo5j6ik65iygDXmTjU/G55/+e1J64hMTy11wV+TV1sVDkt1
ARSAFihwvGcxMDVa0QZV/3tR6pJDlW8wbZYPuKKqlgo7Q5dYBu3VOL0Y5G08hm61
ZXdrIT/aP67X25zV3R/7XfqoZv7+dcUDKkewsymzPb2Ll/YyLPclU992HEJWla2V
7n41RVx4/nbAB1/ZIiqZ23R+sjCh92EFReirPtujK3bALRjUTjFku+njsRYc5hdT
/VtEdKT65n2mmxQi0oq5UIZRedu3+C+k6l6Ky9wFJK2t1FGdnClTe1UjJIl7IlSi
E4f22NZd09S1lNuus4w82cJgbsOnaHs0ZSk6BZjX/Je2hx73HCbbrD9eCl6faAuC
jwz94SYwa34OctTyl/RqOo0zxyo9dINiaUIUY26QgiBTaihEaa61p9gurmUyMRYM
8mKBRXYEkxlQIMS3zWQBgL/9oVcgENqB2k4iKBES2pjefiyx2ZvJ7lr+30VsFf7Y
qxlnoo9qqO9es3irnfNM+cN0+AeyKY6Cg+vFjHCN7x3a8z1J9B9EiU3SfIx14Pm6
L9LX/bppjPf4npvyRiRU+YtregVf6y4ybDedP/HRJvqhbvkOZr0D2/JUuB6KlZ+8
PNg7v6oWAMGGwxMsPaLTZ06CVON35zaTR3wprS8s3zLI/Atj5AulBMnL/bsLUmAt
dCOEJEhaVJh69r3nY2dkYW6pzEEJaKULfXvXBO31hPYGCfqlcRVb2/xRLYs2Po3x
G8CNjdaEjAZ3f25NKrSXNLpdHibneUPpEG0RTJZJUXSt8haCaZz9GHTfbYvo85KJ
zofHhTqgD/GCmRci1BvDNN9wsQvgbbFlY4La4I8ZiZ+SYAnhmXAEIrK3B1r2iXIN
vwEL9/oT+iFzeYYQGqAPPem3+lmgXSBxFNbS0RFsqqViUgla4QvSTKA69rtCwMDP
I8+Ewhv/z3vClrxgkEeuEiJWYWHo3ar2UVuODbDvpdAIlTTPsjykGLI2LAw12vNJ
4vGQhRamIdGXm5kudfwi9igrErtryxKxDruLKFehCaz/tPVADM+ivyQ7FU8efMxd
MN6f6wyZSrwxEFNUnSwLhN4tkEVmT1chmrsZgANXkEGuu4EZawIiUve9oKlGHIke
JjuvhKCzRUBEQXschJrY5JgIg9YtAxMAqY4LOV/UYorN4puRfswn6niOEZQpkPIU
1aWRHdjJOTcD2Hh3V0Q8tyL3IOpZa1mHTrRLKBMGUBsgtUt0FHyDf1mPhZN1l8gl
vJ/CiK3jXhnYqwa6dTfW5iQ0AxRYzl+xQCOSoeDlI57T26SXL4inoS3hHI+nbw7E
P0mtCMcLwm3PTWCRzOnewPuOhTpdkC5rY3gLAspHqdDckl1xjO3eMt7lvJI5gLdc
Ku0jEAlE5LkaFvFNzpBvoz2UlJPcUnJpIssutUx9X3IPo5EEnjKq7qONBpBckKhh
oGxE+haC6ywzkJ+tCT5H8x65Tq1eHvXAGeMnEsVBv85B7/EhX7oRm0bVH/+UMXgo
lcxrxnqRsjUGkcZkcOSs7P2XlbDQzLOGp9jfUGIvnajPZxtdS9GjLNimtj5yfyD6
Uvth4Kiduu0Pt5O8Ybxlc1bBF3L0iIVB9xc1DozA6pbKQqjz0l8DCcHHD+xVCVFj
pzl3lzPOmy1fusvfJ2eOQtAzYh6wv888BGzGbHSCmrN0OPXMn+NS/zlmfSdHgvEL
5ubaNpGj9dY/eb8q2jnKe3PMiTnwrzFcUCBv9Q9QlI0nSj+WKv1yaD8STMva0Ebj
gLgerK82TwCwWjx2c2hm7zLiUD2HFtlInL2Hj6LNGNCGw4xDD6GQvnvxJ1lulIg+
p+fhfOMzxd+GkFr6XC1DCmGy+TfFx6JWmCm7LX+NS8roUisIP3mwgVfDglKfQjH+
vKKMiCFHZDEyPQlVGHZMFWUMRbInoSCeHVa5aWB+I+dCWBgXDd5VCXIN/akYzDL/
KomvE41pzmHlUjvIU2kCQ+YFbQKFDTDZ0jLtnylGgQZHKnR6qtUlmV3yObDvx1fN
OOOqiKeaJAQcOEcGsDnH4Y96radBmYGxfvDM8rsNmXdlxfgmfjkry3F/21JOZI+5
1f/MXz/Sfxe0EMxJhVpBTPhF7aeZKdjemZHAEJT+OeBkbG2PkcvcMK306uhyAAh1
wLdA0BPR5wX5dLzGGCk1Fm4xaLLxPdHKzXO7fHXgdsHP9P4un63jhJjR1hRHfi3e
ZogHR/ojNM0jTqjsVyKCNIcmyKne8US5orvHd5f7cq6rlwmlle0453f6Sf9zAX3P
wD4oOSnTaQ57zZLJx7eZOJuLtM8xobIgp28bJx2ijrF/yAFhe3IuoOQqBClxqVDS
eWfHzbQQhJZ0eD03F8l9A5BjwkHf6geZhmE/cuZPbuivvW9xeA//0+hmwQJbfLST
4T9aAQEfYoQEljeve7N90pN/qr9dgJ/teVUwHSRdc93kVX4bCYXdLKw6b5rnfO+W
a7PvGR5NOGbvEAKRoAkxL6D8gzS9JnbuVCAHySFJe/P5M1HpGtOYlUDu9XFRyizL
DwIaTMlFLnIhNQ5pcSJelys6hkZnlskeQco6E05qXGfbo7k4KRCe6IYIYxRd3Joj
D6dwQxUifRAA2JpV21dBVIcAUGAqlzTjMbEjg1Jvi8kxLBsWlaAVdUzPMGm0JYPl
Fb82fW80UyAopYCVqPUv0UKiUvhtHwiussnum1JSnnMDpPuUv831RmSbJjUU/+b4
7lzbWOrnKNfuwX99xvNnzMNkQbtWiWdWwAFgE+CAF7Bhhf3s6Jyq3iufqaKJIxY4
NwobjdCR/Z3ihAiAbdWh9DWVnbWundKvmnPy0TMRB4cja8VV09AK1bZWuEJZRzaX
LeyJlCRLYEC+0qumZUUf8GKXIKZp0ZUjKVroNuOIASEvIBFwhPOtZ4oUmbJhraZ+
wKiroelHpTsm3I9/352pXMQpYI2uH8srDqNujFcwMFnHyJo1RSNoOHC8VSX/X0jL
NFp6LC1G5YkE06W7SsHmVVeI9rb/kuLPqIrk0RDjFKeN7p3zmpEGUj/D6+WnQXnM
Z2365XA6AS+AhtJunnXNFsG4jJnKdAELuNyUCvl/EDGsnJ3h6YWa7pHl6FaD31wx
vXcpWYzZzvOZjQP5P5WyThGJ2K8GyB0ccdRFjHEnkL8Xz3s42cd0Gzoo5atrp3ZS
dywtNUAxyMja2lHmdFkgRpSqS4muDDpd8B1ci7jsr7zJqFxekvVXntAYtpxArz+r
PnFsvb4GCMSwQl4+5Z9K/KW7adse8qxWiGIBG5Xyk3HfecVdy3QAE8O/BC9K9pcb
qUpwNhTCTrTpW90vNjei6WD8FxCpJ2ntipZmlWwC/bXnaUKlLTOQ9bk/foqHoM6B
NMxW9Eq4sPJB9G9ofhrQLLYB7qQO9L5fvtK9UKkC/6wd5EdhPi1TTIMe/GqcvPzB
TL43/o89VTnXRltscF/+l3kPV5qUOulmgxe65SdaRwVgOeTknTFp91ECpnNmfl2y
YePCl7/HIs9av7pdptGNU8wFoDcetfHUYNvo9y+lJLxVxabefDCW6aBfxvoebLf3
X1pw+dH/1dta3Abh/MirP6SqYkic7PrmbAcBWzlkSfFE9XSnr/+XQ607ME+C898K
KtNQly/hzkXEkv3VS9iru4PvQb2gW2mHIwdqRFWj7UytzEf2lOV4tamGNmBtKD71
HJEqUwAJrj+R9gpqfLFct4WxfT+gcgyX8cdsSuBoVBsL20v5fyJuEG99s4hOLN5P
y5AaEECwpVz/OLNbEKOwcFc+sy8k9xOkF8UvQeQgn0RXE9MFLPGZmzEOwUjtLSru
/KUxYIjNtYvF19vT/kWH7Hp73N2jv6Ct1QnhiU8q7Rk0tG6iY357soX57cBiICLc
orx8JKNhiqx+gmzPvyzYTaos79FGGXHpyeEvjb8VxEUTNIfmh1NBcu5h9mpmwmT4
1sueCOKBZgBoXBrJ8Ew12d4vxShH3jOZOX6HYvY7U1LZmXM6ZUKYbnDNoO/AewZu
JsVHa7pWljptUEbsGaKRZlY/bIgA/LQ6WH/UoLjuvcWKNu2C32ByKxU5uALjR3Xq
zW2lUXTHZMXHo0pX9Qb64Lkr9SP6ALPunZYPFZDxwC1tU7Dci/Kcue64iJJ5IgGo
6OAZRMhlalJykANriOgMC70vpJ9ONjieD5Pt8iKnPyjkGxqj/Ger2kg0OAM04XJb
UuttebknXmPxFtqLcepzDcDyssG1GxNeGQzIKads1K3u5avAVb6ekriwYJrCdH8F
nGZo57bMDQRmREeqYDT0hY13PlgliK1KvuZ8JCXpvefHoxIY/7cLE6rVD+JZlEzf
xmk7PFI4mx0h0E99IfZEac3ZFHpK9oYZRXJWLpSsJe9ihOtYMNWCDDGJJbLKP0W2
r2tX5VQFl45x97hyAIWu927iG3rW1Z6Veouq65Sr3gpJRV1uitdQ8cwySSsdy2PO
B0s40C0EZ19L3UR9HhPJPnB7mAbEU5gXPJAoBizTx4ICbcIdNJq1DWUxCnOcaf9X
7sCCoBYEHX2tSHV2TOvB8XYyDx5Ye1XSmu1f/ZFv+vvJIBI61xnrT0vwW/eVYsHG
dlYi+SyVMviZlV9p9Z0wQHaERi0hJ7lCI3AFVMMZZjVVIQgrBNIrQvEGmNjNp0Ic
fEmSg5HI5SRVEoWirQklMs9TTOOythbQQi5YdSfAgKRqgvow0gnEvkQlvX6/PDHT
iyVezMoy5H9tbdpgajqIeffUVP3nE+DM30+hUp7w0cIBCGc2FRfbbc4wOTh/mJHn
BaPCi3m2XZnTYBcyufQ5kpbXhhC8p0IO7NTriZbsRNcHHlsHSRKNuGdOFaZ9z+7B
iSnKboYcWbiNQgAVVIbg8b6naKPE/7kxpj/igcPHmmDS0f3nMyLRGpOUisKH1a5D
8Nwb2r8uvFJFAK88mDE1Ho5vR61yIzEvbi+tc5O1cDh1kdiepyJBEkvNcv6f0rI9
WFCtBgK8Ug7KwzKhmvlUZo/pNWHmCulM/FyW7i1swLW7GBJgx34FsSbseOUMoin1
vo2Sf+ks+O0/z7aEy5AlV0YYHJT2GV5KFLayjTr/GWkW0ZZFtcZa2JHd8NT20MEc
0x5FZa+51YUg3Cr/yVT6nU8tYjucZV7JqWpKzuPD3rycuHpQNb1AwomUjfZ3hTci
HEZAlE/oqATjgRYe1xHp4Por0iSpg6128Qw23WmmBhwP3ZMRlBrX8L1jdhUFU6qk
yEJiNs/q00/zmeial8a7MWKK8ouQ9Wrc4VEdBefOEHl8gvKy/R6U+Umzyh2xd3cq
mv30990HdvK1LqjSjHYHThTswBX1wp/ilOqFBrNHkdu9eXz2+muRuSanD5TaTGrt
J67k8Osyn/UCLVp5P96bvLVKc4DXgqHXtWRV3lsQX1OcHUzh4TnSyCjUAnoh1pYN
GxP4TqYzx0egtwTt3YznnyfTuhAxfL2/3SrKuPDYFE5S7zJFoFScqesADP18cR1X
UonKSAIALYwosnGITHZS4rRucADqJvJXsenZuR3F4Th1fG/5FzpwFF7bocYpavDD
RBVhkx9GZpEYxFlPxKFT7BCd/3FMOAnmWyG5QTdCk2JwCjPNy7kaaFbUy5huSCAy
MSCp6a8+qGLXMT5YMOZ0sTKoRgBp36Fvzbh2SexNYqxMmKbSrTJp1Xp6yexRZ5xB
aZ/GoEbzYlfby1q0+rruMg9L0NyNV7zonx7UbfihqFdTbDXPaeTmDQKr+dyOK/S+
bIYJtu32AI2sZ1zUQark5hyjCJ5pvrsz9PlLAMLeD3arbHFswIBpVUiqfxBhAZ7T
FI2z/QQ4rOJ6037Hbq7TGTBTch2O/hYlWaIW9lvrKc/753KQTGWgYdcElHQgyItQ
bo+YOjxSUCIbWGK/rFGkkm6G4FJ9wpOwJFlPYFLObhfi8Yd6r5HpXw1QQUAdG25p
GFlKWtQo13JEnDQKoiMXTsf12+ZgCWcd+mD/FGOwnOTevi67gPKlL3sW7Hux87gS
n3Ss+t3kpMskC8AlLfvnw8Rec6cEr/yzSBJtANRGqwVs8CbQZ1cAcSVtFMd7W6ra
Hi3yio8GkV0XAfBYAJdKK89eK+Fi0H6B/S+f1v7ey9FlPOp4PLJ/pk26By7cdm5U
qlx0Ws0ObUUbSQ2vNF0HTGVrW/HpsfaskCwO4CaRxmRFLCoqV+PL/g7u9f7xYSeu
ffZJ8+c8uB9RARU4qXxAJoixU4yk//Mi2P9PoeCvkWnaTPnENcXLg31L6XPGroY/
pQh+dq1DOZrkRvfsKowMnwA3cW1QIWbZSvHBoKTrbK2v7nKefh7ZD/P5dmW0ap9l
Nw7kTTN+r4ct//aZE5U3ie3+eE39aVV6L/tK8tDPNEiSUPymC8M2dpKcildT8GlJ
uJIMd8SXsKC1RRjvcwjdbuPo6kNfbRsdcqYJh9n+s3CoRjLwLVAidJH+g/mLh9Sk
Fg/R7btjvuE0kKGDN6mcUEJS9Is7ZoFvTugp4EWkT6eBwNzhlNscUKUp9rYgPMgj
RQBvhSWX1f+e6WVhIkA/EBfXLp435zsvNuNp06oSOsqmkp77vQ6PRXfIvVmNhudO
vyteJUTp73WvqJm4OSKrRBe4X0mZ+x3qjhEja2Xab57F6272oY8EzDC+IN9g9XFM
dwhoy6JdH4rdJ8cZhmISuNJTkxzRaqFSxOr1geCwae5vuX6AUT1nGpgV0fWUS66Q
10BxgDZ6yBmVv0DgQFVcHrKPzC0GBoj5YXEFBMXZjebzrXMRd/mi6Q52RP9L2vK+
K8tydTmAG97dswM8T4Yu6wTBHs+EwSYVHNMVfj7W7cBGOXnHwF3emu+vl/K9xJYV
eV2nhN7vwl08ZkhQolaFnBrQyF+OSx/oagYFKxN0H5ADEkti5Klo3yMYqgGhUxJx
Fc3ucEriCo54qxOwQ/YlTTyDb93AjWenGT2/ymxjZIKlOMD+v/52eZjlK/W5u61a
dcTY/8oZ3YNq1vjb+E+bYYYH2uUqxflzts09nI9CsYBXfwgU8Aj0NYZQxLNxXZgf
bJaXuhodtA9h+Kv677gq7lEAPxOsIvzxOU1+Zz+amPnARy2S8fqaCSK68Jr3gJIS
4p0QIvQlbWto2o2rC14rfmf943/m+jEBAYSKeTb2AVgPZkueKJ26bY7JSPpTUbeG
WLdJ+j337WBRXZz55+GrXq8jQnGzQdcAleFssNtm5iqhjEJzV+g8qwzopantk+6X
Axf1txLb94TjJk5yTXRN8dKCeRg82Haps+ErcvlJXbnwx5RPiFOqkJljVbe0dtFZ
9QGBZvPUsQ/ubbg4/083VZP3N3xkH00RXZ+LCSYhMCm747j513dv97BLe5FurMkh
heFto2bDcv8K7H3V5xYPniBdMMgxaeGPPdi420qEWElxr6rvFqYo5SpfOC1SHUYC
0er6B0P7v/mcfj+jwTv/7xqknHXriUrn2j4ayf+xchsG+KwCE0mHHtHBaHqgZOkw
rJNRznxN2bsxPhx/BZFlFgeWOSd7mbLocUlpD5y4tOEPIxAf1Fd67slQQNjXXVCf
KS0PZp/8SU5HL1l7AjltGLl2DV2S0HAkgH9/qd+k5/iCzww7aQp8uj6Rt4gHIOb0
DC+XDekt1JE46ZnZ8gJg1iRhKhHUQOsy1mXUxSrVwYUIGNYzykwnJlF+FMoSZH84
y8CfvHjzhuIeKXOirGU444hV1wTfRhHSQV8TnHSScb+BeONEadQdaEdcm3+U5hHO
Rm4m56ddMYRQ1vAorD9E6YKseBmPKpa/Bojw6HASEKaHYGCvxsM/+Mn42TjLHt8Z
CsFf022ines5gZF2vaamX0jWA2bst3AvGpkafzE6gwS53BbkzDedW1C6szS83oeH
dsnJD4e8YOAUnPZJxwvYj2gW0kKh8h32KWqFztL+B3jAs3EPTb6iB6pInFka57lW
ZaQ474HaWi563o62OTfpsJ8aVIcDXpmNDZQmow9qDruOtwz1TJ0yG9XpXtpjXiEt
qKm7+Z7ZE5tLDfdilgviqOh58uKpTmEpZvD4+CKws9yoepfNddrxZzXP4hymNJmG
8lYKt/k8wcGgY+n1NRCBib0nIx1LnTXLxeuHSp4pTYZLyicwQYkOJHgnoL462Fzl
e/HhmiErDvDu8DlUSJAFK6NaAye3mRCtelqsYdTKWCbEXcD4SoFs4GDugQBGqhzJ
ViC02pIF0JU9jVjNr/ck08T9w2sVJ50M3ZlZHB3rgT02KIbCFP2UD9zAhHZfP3jS
Kiv4QngtB+3HUH/v3L+lYBSCTCSYlPCXie3BU4HR5dkkrEdzjatsVABrUEOjx/TZ
7SNJm9aFEYibLzypMSmTM9bYdQmys+9mBSVDU262gAWDXZfVnEzAkxnD73/baGuJ
jsZGi0G/7taQavV62xcfg8F+a3DsY/EjO+lkItRqwe/Xqz7l2m9krdQsdjJuzibg
qi9TAA/lh3GnqQm7hIrqbh1We3VlI9s42I2GEaHXgm4rpbJ9a/ZPCa1H4r5tcz5E
tM3f6m9NzquKRmneFrw6BA3chLD9/+N3NDZ5Rjsb6U2224AIcvz+CUshoD0JEzrN
TcU9WCfe19DNxNpd3XNmjlDnBg0digWeyhfyPdDSXpTiaEYLNF9dXZI0Crb5u0Qb
UaPPZ+8PgtWb6YQynL52wRPkzt+XreWdR2rhfhu7zA4frZ5L1/H3PzyshnLJoUel
1QuHxVRc20VTYfJgwPmD2h/bxyPT9wBl//aslysViVeJVal1I2YbPSSXLBVly5AG
udzvz7jYwlFXR4RhKETnk3qoiZpYh7fxlBm2/KHZkK7hUJPbRftRRvd43NZVUO/E
lvnFXYj0tanich92uZB2AXto/k7oC2F90iz0fVdB5YmyK6jECsGmzjJD1sBSCTgb
TD74U6TEeMBJVGHHfVIYBGyVyZwK9LaglfYLNGNC5uccb2o2JT3h9OGuhtmMUOsj
kFhkZktgc9MnEHURM35GpMpNn2RobgUwxM4czfx+I47n9oHZS43mIKMobcl69Xjh
KDCmDOy1w2VFq3nkExtN0cADEmbkoRaRf2HSUB0DMUjiYmLoluoSKmj0MS8f2t82
SrXP+zIwRdIqP/OvZ6g/cAlIt2IsPNQcmOXIko8wMFZke/MTcwOxTccYChY9xsKF
CRcw2aJgFlAX9HddCa//CWI28OPp11IAtfeykH6RZeCqvrDudvMB9hlGaI30NMiP
NKTLTTqmRIgBlHimfOqVrrpZFtC0RbLetphd/3RNHXT4O4gE8FuU0Bb8SxvyDvZS
hop0KowiDgppNUFyqRnFkjKMzP069v5vRB5EVOH8WktkHowfGCtGLDczgK0v5nPh
NwwY+BmdaOR6go5e5XUmjgmAB5pViVNaXJpY4sXziTDs08p5/Xp72WXkWD85vTfT
oXRDFU1TKkfuxsKRewYyPxTqnWxRIDGgvyruqjp1VoLvDCr94AkhLDujgd3DBwUl
nmhOjIFaIr5IF2mgcE0WyrSUf86b40S+b+Qg5lMhMwnFR81sECM4w6inhEKOcehN
Noux/eOU0ZuKrsFqWwvh0uj7kiRWu+U6pWY/0dDoAd2KPc5tjkKnbbdp++hKzcS9
h7jeR6JLpBJ5VOO/ji5t5D1ZjU7GqPCtOvKKE7xn56bJNgLJIgbCekc/A2R+/PR8
6vOOcjDFqnm+p2a42ie+AOgl+bkJfn0xQR8cHrMEOhKWZGle7ItPFrI4lQ5dJDFB
fgYMRJbXu3kMBNLOSjHYoK6QHVQALHohHbfVNIeMXG+KXlnBephDfyz87SH6PPdL
4FqN5qMd5cjAeQ7+BfObrOkZlQYoqUqWaVgQI4ria6KRkLk3AEY2jRsgPWen6Bul
IEGYJYC+KAaHKxBBIherRUStCTiqY6hBKaVZe8urOXbmBsgUh5Dc9JmwfasIi7ky
tfIWjyXnmjRuHMWiE5AmzJhPf6K73gmkMSb2OPwyRjBwz8NXmqwi/ye591FXRlDu
6E0HuKXSz0vvP3bDoeo+QPJrxr34otYCdTR10SzqSJFqO3NMm6qgJd0XVfp5UY+u
3l4jkDp8CdzxPYZmtgMycwbU0e/dpKvWal5IR3SRwBUTHrxikaNFJfMNpYxCeHCb
xPNw90DjNIHeKRGCM+Uoveyum2+JizpNP3WH40fWwHNFAtXL4kPkb3VuDtGkgtO0
LTW7dLJEImHra1SU8r4ADNvT8WR2hrbC71PSBMQimvr1dF/V0fdpyqLEjDdJ1wgS
HqQ95EYqH9qb9p8GsOrRO0XBDDm8yjlKHZNCIE7w/tedO8iGHXXOr1MQR71qqQle
LpN+M5V43HEHi1B+hqmdYL+s1tQbXJWk7mxxiEYr/9T7gTwnv9mHF5hIGpQ6j2Vk
DA7rxTNGmYaoW/R3d0kMYIotadx1/zMrLnTiUaHiROUmrPvLQpK029Yv9n0Sj/cn
A3omeFYT5C8+ZQs4CNHbN10bUSfUdYJ+UhJFzMcP/DjQSR9h0+J+VgeA+5xD7+iN
1y+ufhqI/HgY/1uStCYigoiJxYrqg2ewqo9EoGak5zgAYEw4arV46YFgjqT5TGSu
gT6SN2byRXLWJpOfGc8SR22jdx41vK32clmWMaTLPYsZKiCFFygImtEp5KRFMdje
3iemiEJggQPYAjtnyTsHsa0b3e/c12J3XIMrLhhy78HpAJhnOg1wO60+my/rg+Or
+A2DVf/Qk7A/3pb7XXCOtIb9e9IVSLhs7ZXYHIN/oBmgTt/C22Kfqv5OXPmJH8l3
pbyycTcn06QQIhOYjz2RKPwydSHxIglSISTt+mBLjLJs2YxgQ+QW+9h3Sy6lgipk
IeEdKdwOzNMewEH7mauxsop5Hpu51uN1w/80mw1Fi0rX3tHcfh6hermiOpx4USjj
Y52DIuAmXpAWjVmjws1dUA/PSYlXE1J5gy+r3pElwJy1JQ0Wh5k14+B/A/0tJ4Pm
1XNPycCrc2ie3zMsUj539vcDbSUF2qN8YZvO7MEAV/WNl7elfvxXD5pHubOW4QMM
l1sNOjDnHJ4Znpec9ft6AF92fWpuMVRqXEuelemK5vGA7VqqfiMopuAMlWmaBvLd
gYyGlN8eUXs5kt43bdO2L0lJTgNp0kYbRp4O7gPehIIuhpcPCT+tkPmG7fV5HPm5
Lq7ZfN413mXe487rnS+2TTJDXe7dsaw20MjknFxfJ0kGq2p5hWnHV/zzV42gotSd
DGB2EiTZjVS2gIsD2qpzj7ZcOZIGu2/2l0WcYlTiLsc62RUXCtVpNWOIyGbu2JLR
1DRE6zmD9/0F67QrJ3Xn3V/tiNEhyk+QkWXeJLJUk32xSMQsG66FjIWgoDosK08v
+OyBagdiwwrATsbbbdgUf7Z9PcHo+JsL1FphVGH87suaqyApciDBy3aAshc61wvo
yvLaTncpRh+GsM6bE9Hjx2rsznSlZXIkeQ5Fn/iVSTQiM/K5FMNnFKmgP3oDhM1F
6DPyuHjwnni2EuTj16Z5enGn3dNSqI79oZw3QDNsEEYEaF4ZaoD/4FjdTvD1xNpa
MJamiYSRCJNkaVPk6DWOk9fwZhqWCx9YqVazuZijmMHW1GdvXC/dKYC5a+RMiTJX
teZlGDhGRXKUpmBybaHa1UCPzraPdq+HvAkqaEoyTqM3CEnIyhaPeL6vuvRDNds3
PLL1CsSpdi3r+i9nTRNDL9dFSeaXxVkY3aeh6wtfCptyAS1QCJnrTJ/72tR7LU5c
lAaIvGpnJ1E1GfJJmSW/ZQG6SHApLP/DgJYBn53C3a9PoIgtjYSTZ343TfKg2P2W
0bzX4hWk/xXlb/EqodtPd9uArDVj1hB6U20SE9GU3Vye45tGPHGjdg5Max/h97Li
Lrw7ey9atDdpudoHqQjLQVKde8eiTKxZqPfnPJRAj5RxEnL0Uoqqebpkrb7nbY5q
pWDdtBMUxibnGqB4hsMgvtKsmUMqnu+N7ewdvWBJEKGDmXg0WgRAdmE66ZTR0fDx
RQZaop8CgU+RGDr9roTvT1rFzmx07ncjD9sYBUVzRTtyXLOf3nubSn/a6/VqTzMF
nu27sibcE8ZwDg7TMC/IqHsR0DHF/Bc2b3Lrxt0DXi+KsB2EL22gQyfz091+GPur
w+atbi6pQIvvE7xnYgajGsZScl468saHa7U0V+yhdnzDeuFfSdPiC+Q9xc/g0x0F
R45hODtYdOPYPoD1XMFsWxSByjzIxdSXDanbbdon0vxPbY8G/thkdsuYj1KEkExM
8EUl0qQLoRjpgexVTD7qEG2whKXmajjWxRsyI9IRUjYmiIQP9Wx/3HCRzuE+W0oY
ilgfKOnp5TSHWfrJDDfMfbqn6jU1BPy0p+/m/p/0a/pQIR8UUPbXTKfa1fK9s/my
mPYU/Moq/G5Xau8VBrBSu5ZjKzZwZWwoKb4gIo9/g5+RRh3ESxBhjnVFJ0HT3hyn
0JvGnoMaweJ53IG2GMT7YpqPC4vdAhEM9bZfu6LoGSbcXxVM8E0WiE16ifVAvD4c
z86byMx/Wh5630bkxhChqc/KHlI0/7gN4j5MyGiBMWYR4qMYmvYEeIh46Xwk/QF7
E0EprtxsZyxCKai8THUWEAf+kYE6wfKwrOe9rLzxjAgom7RvZ4EtYonj6PxLFHoE
z/JH2BCgRY/2JPAyzYAbw52Q3V5ChGWY6RlyIsDDJwLBAUZJV8ftSTCKMVbPh306
ej1iaSgjRbtdCRAzG32k0eNCM06fFC4wOwsTQXHavrB4vvjyoOA4+p2zRMRDZLPx
mZgI+/u8kRc+swLOHW5UA4i7ilH9o69CAi2gC2OzSau+8B2Xe+cdWDETskzO+OBt
82vX/G4AyRIDkqK4jWHKY86SAjjiab7XwFxFWmv1la4yC7I6yD8kZb1tnZmnnWM2
p36xe6CZF2wpEAQAJJNyGN3ou8vB0Ehpe77lFJ2Ns7UFVU1KrDqaZEVIIH4eQU23
+TWR2MLyasHv00eHMIxOpwqF3QFGSE7yykT6jxP8vbTzA2kFRn5CUEoyXMgu9ZZU
vwTIo+4zwRzolBuQIXLrsyG1luA29ojal7KinxWWO9F9tpqX2RDpTtsSkwsZjDrZ
GyVODdMNK8eqESgqHbMcw40hvQR+Zcj5fqnJygGuRpJNWJBfyJnB8nXvrbI6fdr0
2U1g7WaaHFHnJeXwwxoJue0hbG9nuoF/pveUkYoEDcsl/qIf1hiBLREZDlcU+Il4
E33rpI/WLFK/fOHz9ZXHOyhZ75wrr4To51MJtube5AJlCEVMWEKzZgL3+Mf1M27j
uHBAqncAkDdgLOUdfPP5MeK2kbWbERotmZFxJo41OJNh/zli5XAdnNmUDf/0qVBR
rsjmzZZiHJ/9+vTg6FdStNwlwQNb2aXi/1CO/pgkcZqBRckSF3Hu3b8A9XW5jmC+
YK1vQWH0cnu85Zd4lBhYTQJ2fXEx+/IIsaC2n0WH4bebbAnLhz7S9iczKfb8tFjB
U6pord9FLJEjvh70fryzaCqpM0b2sepUI7ZaC5ge6hlzhX57KqAaB1bHFi/Tvdog
7BXK2u38q3pwNoLPlC/TbEV47lHfgdx+EKWzeRVfkVRC70PYRCIReayGwidiuhGL
j6R/yVZKxXeN+YC+6SYT79xjxsU1lDupWSzlZ1kLALX2rnxGm1nb0rZBVujmz3yw
Yp1GAYU9HKwD5JKfzFIc1HN2U8JS8laOUtHf+ub/F+c6qLmsleptqchW1Gkzwhdg
ha1YwPuJlzDY97izFjnHlGOhTHIt2+GHMhok67bEURaytEyLmdEfOHmJIGhSafWA
xlz/fZRNh0kUQNO+otke8eKqW2iGTZL+kxqURKk6E9RRDFYhMOdBD2e2WQ+rPR4N
VSxJPckswOBNve+7ZE1zpdL4ixbWA9pquO4Xnm7wirRibF7qcRMa+Depyj7OMFwg
nrAuOH0IxQWPBL3sK/m0NGIdF2ECAsIsUp8NRUfSrb366VtVYs58isQCkHklb9Bw
79ioQ1jNEdPpzpfVQrsCpXvZFzytZW51JjX1o8xFlEIydj+7wXwy3KugHbgLYHtI
zJW+ZouyKtjApqWss90JdbbRCNheDG/5AclqsWK/ZYMgQ0oFgX+2ynrLlhzLIIs8
iN4g9pEhr1s6CTWNgOFkkkuN7qaGWU0jtjSq3wjR2fZlQfSP3+9L91dJUFEjp/K1
Ro67CuhtzK6eoAkuppvwRsu5/uudgR6IK13xKrjTsZOG/vbmfqZ+LFHpsNcZpS3L
P9vuddbnBTeRY0kF+hgehVR+XvaWebjH3eiGY0O1Zsu+HEqfo0/GbAry3Pv+JV5Z
LKQthoOwdHr4EWCGpfoHqZdhhEH5BYf3s7LGRWwoSqU=
`protect end_protected