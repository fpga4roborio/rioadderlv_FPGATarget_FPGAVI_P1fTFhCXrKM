`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
ddtXksX2+yylW5zu6QL2Lhnb2d1sD00763mmSITNX595NcHTEkwn0zB1Dry37fOW
FufOhVzEJp80NC5qZ/+F0Vk7Ik02dIR0elf3clrjeJRK85K4e3Hoo4xn7YbFUIms
l/8VZSb14+JVGURjfswrIyCUotIzlzVYZ6gzoZwDXIi5gQIBf/gI+KxNXPaKV+PQ
Ufys/12rjO6aI/pPlqSm0hCvftmBcnezN2hk1UeXgOIuKZnogjOsf0iJVX2aOOWE
6pD/psybjbnsNB6kH5uFTA5frkzIzkzl5d9+YDm9OyC+k84E83I/7/j+rk4L2dah
QJOvksSIzN867/4Qt8qYTQ==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="MvBXkzurAa5VTw+1JJ70nePUfoQXBvZOku/SMmg4TwQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
oRtzZL4VJ4iwysPsC8SXYCzXS8Fw2gtZTOskLcDV+1B9Nzn1zTyNtlo6lNICRmmK
ZRVu2BmCc2G+fmzynYlNTnSa7C0Cuel6FYpxCBlOuk3OF2tzAmLAuDyOH3Z1Yjzk
a0aHuoCdIRKv7BrZCdALt03JeUmXKPdOmIlkVGFl8yw=
`protect rights_digest_method = "sha256"
`protect end_toolblock="Jn9CQpRhJt4rnzZPRk+dOpzAubz7omckX1MrFd4p81o="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 44624 )
`protect data_block
gD6l00tciPUa6pDNTk/+t0OO0nC/UTtBwLB41d4inuAUA3i/ALrNyoJVcBnAmEQW
ptbcNp5fxEUJjnOxnedyZEuEBxWRieZFQnkRdF269oOOkmPZ3uxk3yK/vcY/Ez/H
Bftm+rXuwAHd70XI55AcUQ3VGqKJGI8ZRLsP04Y9mWecy0v4t2MHg/1aA5caXfU4
41VU2mbAAKr9Eb1Ry8EEaWhvNcuVBxAiceqPflyZMOicTyNAVquReW6dDyCI6zjB
IrwHw0TE1hCxe3xk/KHBPzJ3SmBaV9NyGUJUbcAkXRzpRX3a3TleCIYT/34rBhQq
VCd5FoeavHqoGMJXVvhHuumCUg6BgdraffpkQ6sKRaf3su0zp2h0QCs/lDGee2Aq
Cse/tltMTGI3kbtjxuNvhpx7vxEqwa2vkrpN6oXMzMM3ZIAhByP+nrveR3OCRCrb
/30h7FC4OwRoZGNAbICqfMt5EVyxQcxWvCv1upvqYqKjjPiVP3DUzjbbu0jpNqnQ
+Ct2Y5n8gPfmjuv4asEr6cLzHvxBCgawEoqiFy8dbsqVdNojhDEFe54ct3eg6fSh
PqFzIyXCXySoryEgcNurFf/a+zO6xBYfajLj4yEz4JGQSb76wQn3HgzfhquSsLkW
WbYFiEtNtL7EtD1S7QyaA4OsszaDw6M617WGtbuDmVvgIpP3TknYI0/A+z6Tx66h
wPPtauNA77A7RBKgSc9SBXh++VAejOa90N+JQ2JyeciXdzQ3zijpQbLEwMHnaLqs
huXYCyhpqimvBU8fK+DL0qDrVEKwPCjM3Exq5WSopoby52iaxo/CDzBJITxVsDPB
/UgeoIksxfWrkwFEfGMN935tXujAWBMm5vyhEYDnXlSidKmCJ8jvDkTVNgPnnlr+
OW++JYnGt/RDIZp1silSbmPzzZubqV65oaTo6fw6WAdG/QnIQBlRsugayaRGc+Wu
I5G7fQULh3cORV+iMH4WJ9UrpwnRfuR6jgdGMoXAm1DMgrZltBnbjR/fARAtY5lU
sOyuZ9H36CpOEbpol3LUzGn6AzGfmmq2LLkDOJHvC+T2MQb7IypF6Bt8fh6jdgAZ
3nZkMa/0mNWVjdWwOrAnI5Z7nblzdE643doayH8xdER6nlIWK3nl1waEdbQtZMLg
vkeB2j2icgG5bP7aE8rDi61+sglkydcR5PoXBLZSK4BX6mq1IREfKMJN1M8lh45o
dGWEYlAutF02oX8MEmW4iO6F6O+8u3UR4IS1XQX5HyQQXkD44/VsuorjCkIP77m0
JctLALAsXy3qfMntUpQZd5Zp01cbXqm3lbC5fPs6S/kUlY7F+5dEB9/FFqs6hBoP
gxwomu9VityKc93MyHxiA53MaijOKKxs9yKjeHHKpNwlRCSliO/FOFN8fCmxVlpf
qucDxAJjgz59gA/cljNsI3vV4UZMjJSqhDGqvQScIBejMsPOe9hCXUNwZnin46Ud
3dqDR9K+J2V1tEaV4B89EPDcRkCdI4p5zsb9xaJm90rK5D4E2Nc5J7lUxn13hGDp
yr2IkRqaLxrny/e6mwuiIpfP7Q24upwLc6nYLtGfrkAWSSf/xQXeemt8d7wB+0nI
C3ijKbzXOPPNj4q7GPAQ87bTle19rgrvoZPUhr/FdTSHyhIy5oGFGusWDr/yvtdH
VeH6SoE2w1i/dk4l9z0PgmDvt6aUg4Jn/cNFmScrNx9fMehZ9Pq8/eb6LWMq9yUr
JE8Iqqzw+8+PB0NiuNmWaqOEaHPKNy2AO4LPptklTU8GNrRfB00lF60gGILuEIlL
8IKA6N10KHuyhdgHd2baXv7FU/tE4RxA/P4nuI3xI+mFnehZmUR+Xweskm6qKdfe
WcVLcTrHGgPgvh0DOgWcZpSZLd4UMBrjW98YsGoGubRep3iDKYrOySytRwiZIsZl
2pFyIDPiM3xeIlAp1mu2bPDVDWK9uGix4vlsYwO6fYbAOfRD08wyToHTax8gUkvS
puadY0XhmiUDmrmGAxC2UJlQatqsiJoz9p2u7oA2Hb7QEfi/t6e0qWXcpaR6ka55
c+m7qMBI1GJMQwxMMTcZT5l9LnxR/3qqA3WEIwnybNIMXj+VEdLYnR7SGmlNsPGl
MCdOZBKTrPMdI8LfPHoPozgbVIcwr38DfOCSGyki5yvUKSmMkCyT3XaATSbp5oyH
70KHBwHyFYBc9/7poj1mwClEVQXvl+xA6SWN5ufnj1sKxauUSMq/g0x4b3W6fBIB
oIPixxVtaNrAP5gakg6Cx/JbAwwYSf4QWNa1ezPisfFGyfburIy8tETCXM8Qu4Kh
MlxPFBxY58jsl0OlLQpiIy6fLTWOw7eQqtkYZnUFucBkAM56gwVBnvmuOATbDqCh
MET3n0h7DbQd7pRJH/i6MUNsscc6Jbfsw7ORtKaN4q4r5PVgOR103ZQjvPdJ61v2
+x47JAU/9TSyFB0MHjNTh1WdsGo/9Tb0eaGhsdw5n6KWlDQotBCDX4kbYz32vX4g
m8P/qjS8gqU1GkRQktFBQgW8i/AI+wUb5nj5R0sJbgKt7eoVzD1L4tpolrTstTg1
EZdj+FUSYc6cZ5RXKrrvIEA73lQwPRk6jkSQArxP6Yac4NFhGhisRd5fuoy3Mbc0
GpSOU/C3DkQIHb3t07hpSKSQK+rLw7shJmnWPo1TdqOZMAUpfGIisK8r2dv4nzXw
2z4bmeq6h9lybabFuTcq3hoZHqcMfDd4x2dIEdFCKGLHl5uTZloT/1WAGVKy0Vs4
osekD6h2r4kPgffqFvdKhprsFbwKTsPRNnw/MS0x2lYA8Aby8KHEwO09j8oOHcLo
L2e4Z6373qBf7B0qTWhuqLTXng01GWBAwPN6/9Cvy9YvRB2+n/u5aR0N567WmlVc
F8CEjhn49aM9B6RwiNm+DmrtfO53xTq1e7ZIoEWq7EIFsObr/LUgL6kI5p0AWYo9
cAbykfZ7bVgd6dmeUyY7oSfuIC2fXmgp6f/Iwl/zXWEs8IbFsF5QcAw+3PeDto7E
CgbNNF3lP6hNnrqga18pjGuf28tx8oVJYC9HHLr6hn1XHioVEgIgb7iYZfoAXcT8
GcAcptmGFwarNyP2W9cpEzt7pHZ4eqH+2jfv5hHMsXup6yIdUFAiAOHOqrtXPCc6
6kOjEvjAzz9ox6Jt8XdDc+KjGpuV5OGWacOhMg8Q/ZHgdPzBB9kTkmHfvj4rl6xa
l0UB5FAU/uVOPILd9694QXzLFlv4aOd0ACYAvuIvucKx30vpUemLfSFNas0UJp4q
vSsk0SMKfdEEVKcSbdlihQEcdPIOfPQ3m5PvCMsiMoVPtXjM9zbttZKq7qWwSTb3
dPYM+i1eDPy5LtRhCYMnF80oUnSuC+5sdLMxOu+VVtOGzTYuv8RM0nPDz02b2wB4
WDJ8v4uvlGFueu5NJyQcJ1ODZqYXVhOlH8sEVN2pKJ2Y1a/D9ueMGCIkfAS+A9tR
glSvpRU5uWahZ8xvexdat154bzVzMRd41SPsvyTU2ElluFZ2RGqCy4TXQ6VBjH8z
GeipyoeQ/Io/2uWpFJ/uHsN58u2BbuQLW7VuqTXOrPCvYyZr6VOpZGy/NwfHpSjD
f5TZQ2Nm6pQgw2zqQzASCDAzgfmM2ret2V2lGpVHS3/tzATj1IJwvuBYeyMxHU4l
Wy2BEHFSx9OEtS5LEGEirGjw39CZ6KSHZWIRWAdu4eU9/qHVt3YHCBj3vgyLFiYH
T/puSh0m+tidnx8uF2zH1FU/xQ6+b5SmvkPMBxxlKYWxzXdsvTurknoGfl0DtVjp
JRG5o73zYpE7FPL2XSAuSrf8mp2B+y0ktF5z6hREayWI8YzqCbz25FC2v8x73Wwt
LCbBzR2V94rCCwwuzVFLUwtu2gWx9pbysCWD4XfoECHDJEgPZihR8k0kwf3btuLS
/IOmXPzrLUj08AHGhTlqpW7RiCzerrtFPCf/A6gZZOqtQfJo64gRVKXXc05FYCBa
/KOCSm/Qloo9lDEX1YpD3XIXBBoprQ1/M64tqWC9/L9VOvnOTjy5EXDH0V3KifO0
kH6R0S8EyC+XY7pq5blCBHXBkdWL1hOannvZLpWiaOktJY1bvxX6yvgG9foDRJfR
zRKr1aqJG6ssLJCzSwVgS5ibgxmDLdlF3RYqN7AdUl4oXGAxQ1369xDrRsEow/4c
H8ipiKDYw7/8m2DdIGA26mnVmx8FceRFWJx9hEf2D0BHD/dAum8mOWXFpKCRkhrm
UvPDZtZeRdAGxT4IE6J73rIbDghrbDiKxMviz26/izNzzv+62vvEpdUeMoe7kvrH
690ogo6umZU1o3NMtk8gtjXdzCpBmMqoKvAPaJ0CmpTSxtyZz6noVnfTtnPtgtqx
LpzZgG5lrXnttRtGE4/T4dhMGw3Ti1fFIfeWcAeLxLkgpmCGRDLLHNFn/xNumg1N
ZrAGVOWTrvF+qaurlqwE7pjjM3lxR2JPcoIQVogOrAWQVA4ceAlsTXdziKcr28Tn
Nf7oT7+tUCsvt9GhlGT/q8cvTB6VzPDBrUuL4/96fOmNzc0n1fHCxFamK9RjVRqD
lf21Kd6JLCrfSLLLUh5jOsGMuMnAii9WO0rCnGggaoh4st0Nmk9Rd1i3SBmYLLKe
MKd24QNZzYEs5FTiOmD0GZiLPD23dVmSqcY6iJlQCshY/SwuVfai7DPz8hBt3sHB
CmpwjiI2C2wY8/AzIo4YjUmr4BaEHu3ChpZ3ij7viuI25ddLCQyzdaTaJDvXQLgv
SQE2yBunQntzWe7mX0j3V/4SCtlOXSsGMbmFe3mWuf5owxOMumzkjALB6VvRkCWf
/5+hmcop7OT3V3EkbJZwnbRc32KGYKdK9nP/XdPIzo0J7lVwhkkGS/H65Ms+Xzea
louH4ktNk5KkR7L4kdszAlVBi5AzXFRBssS813/K4k3kambCyRSqxprt5nF0jEBf
tcQiOAHCC5civdsanP3yPq5EW2GV9Nio8sk398tknX4OA0Y1P6w6Lby6JbJEA4hV
IxO/5IdMKVma8ghlRbg59cjXzF08HRzeknxIPUpyHd+JlUg4OhasVtCirHwge6hG
7T2MSlYMf6GjGNEG7v+VKfWhFi1yANg3XLYSpOzrBdVMfkwfD4dtBewhWaPvRZqd
DqTSWXXX1AVeVMhr0n87pyO9BOS5rIRY9gwM+UsPStBh0txgBQpFw1L7nUFWAdsk
O4vao9z+dm6woW3JY69e3rMsJJ8fZh0wElAjmtT28l+Hn8ludfS7z/TG1m+SaeYA
OCMwra7YXpzRhWyglno2wysjDupLpj34aZ7ua+aly/tOPqjPTGTcqxgSw3IQgYK6
3mHFMkA4lqYQYmJqsMhmQ1fRGMEiu1oQ60XniYhhVIvijJeFGI1E+thaQ7y/wPMx
M51qpUFALJu+M20wYlpkE2UIqqty05YivtCdtJkiMFlI1KfOgot2N+CZzXPRTgMP
73H7SeiDPRq1KAuk2f50xstAZbG8ABC7m4uyHSTtbFSww09UaP7sjAVTL9Akmjds
UDpCpQsF8pEKXQ0nmnosxEVb+TGV92aGgT4X0/m+oLKENwHHXyipCoK8rlzsDQp3
9U3wWDsVBHyMdO+VWnDXWzz+0bJ4EfmsppvOdLHg+hg5vp5AUPm01dd2tqfO1Ngg
x1iJ8AChUh0okranksON8BlQuU4HVSl3L3k9il8yL15f8kgpRcGMlAXbWxf6gl3d
6JAGJiet8X6vO0QuWuOzFMRY8o7ZKRa42l9nO/IN6wjZYrmuOSDlUXoaDX7WtAuL
9MmOHnmb9ni0M4mZXsa8enLQw+lbIc8RWZegkVwlRYoKBVRmMkzmP9E6Q7Wf5S9z
PRs8t/bgotsDijU9pZjJrGtcvHVtRg0s9UV8WRwpdQO9KI2JReTy2f4mIVl/LuEo
ZxdwoQY+axXphl5vQTskYbB1IrjmWkRtHsExuRMVXPZmPq5yLKPPAzEMwsWJAqRj
FraXTAXpAtm5rTnEYCIfhnvtrUEpj96IaUtx0ntSMtzbaRx0XRRtmRpCw6IhvrOS
Cnlpt2smQ2yXl7rZ9VIAZlqMRMNYPZhhfmyYIbqT69BMv2aqugf4o7D/E0/OX61B
+DDxcDgDWfhyIpKLBsf0L4BUVgSLjQIpxOH/rDJiUZSuYbb3Pzhu1n6jyx8CsbmK
edcpXqbOXxRgXJ8BvOGx9dMI4RedS7qmJanesuIu8oToLM5EtKnUOqcp7LlNwXuD
e8oe3hwEY7fPyz+avzr1H7bpR0IhMGLRS785pY3UofNspQpmMhhogM0GSKHllyW9
Tq0cjvG8UrFl82saPv+xKobtKo3YTpf5p+sBSBhl3yISyOzMz7rWxTGKoKq8duR3
MgrO6Pfw16mL4ydxyACW7kDoMpZpI7dUbh3fgGwu1B51aI350VpBAStteOdhwdhm
MK5rF1X3cHSXvZ4lBbbb4W6L4g3P/T+zTgnu8jejM1I00lE8geiVwEMnVX0I0qTg
7nT8RvAcClhXpzHV+EuNkdT2GCsD6mAt4cfYhNckzg+2n9EZuBD1GTU5yzhSa/Se
VBqQvxCxceG5BxpHDX/DXaLUIBXxdwGoqWEj4l8EOXW2WYpBWducIueZaIfY613Q
Wg6qSmnu2ubuyJrAf7KaE/17xM8c+DOGAodNFAl1LQdmUVKdpwge0O3DtUBEuCbG
liX9pLQ03cHoDClgdaobovg/voNK0iI1sQNsDXs5bh9hGuRO0peNgTkBMUUTo0u5
50tUD5PJ2/AkhZhZ2hiyEa5JgmuCMBHq9OMH/MDOaGKu7CMwA4Zd/ebuYeZwLYhn
B7BlXCOmpDdHNfasP9KfC1W+txM5CrP1EaEzx6qzLFbtUtt27RFl6RTMCm/iYdLY
f0FXjpYPIy8o6F1VR4C2I4hfMmWqoBzwb49EnKaqAINovuvigoVPXchVbcoZXI06
79rY7k1NNa3XDRJ25PBgSWmeqGYOt4se94Gl03/O5DwSmeuwbpSiI8C+emkmH4w4
jahoXEPASK2K2tPQm+PsMbZ6tIZA5mpGOk8MPQ/tYUQ8BOSxRXyPc5UkSP6tffSL
BN3f+MGyyirEmiZt17use8LsOEBR0rxPlTTcNy/gGscUYAj4CC2wZmo7LQdAhr1q
dR6vB4jGhP+UYJk9QVLrwScl+xCL5cul2E9xFJne8ByHj18DDdOUidHZWlzICb5H
zNFsSaO1bElVSRVLwo0TbF31ZrIyRu8BzhxOr8uNa/35a0B5kn3dHwRKZO9ru9Gv
MoyVDU4pmkUzAtx5suQO4pmwjBsOXmUTokEs6BJzwTgLxwVX4TtE39Tl/s6poyY3
h4QXdknZG1R+XpdXT2rOWKC7cjrl6hntdH5nFajo8OX3AtlkMarPAFbu5WpjYMMN
C2zYWGtS4Xdrza6nCc2s89i7NaeBn63E6kmWFsNYQRvu6pKZWPot9SPCukgZke1x
NIU1Tslo4kt9HGedxwY9dF3/lquHkTgP1LAzcj96relZt8zc8T2YXIZ0Jb/apFXL
dqciEwRyxM748fU85ziuZJLCczOxJhdRnAsIZG+Q0gZDCmIKRMfiULUMmyLBiTrR
RsdHvMIW72E1FnAdtywQV6rHwic58DEOxQcxfCZMo0yS/3R0fILoPNiN3mb7eAZN
UJkYGbHRQ8EH1glvsgk2ZFlnuGlzCmLeSOyKSBmBiGdxFXN35hPb4LakozDdTMEZ
q1RRa3+GThri0OvCkLten6x2cMPIaHiDAIdepdmILsguR9JaAk5tWRFUvDUDYiDZ
6uIXFpNPGSKOJ9MkwPdIpe5tf/7fw1elTFMYnRo4eWqdeHHkg6bm4n/+Z17C6OeJ
CCTMGD0LkP6AKL953UJgihEYhdHIYq3i29Kq3E7dveIPveWfZ9bBrw0CLKI6vwrI
BuOdT5CpBw0iazX2xCnRLS5XbqkPFL/u91robyq6VzRSwI4JkzD/2Z+v1Ofq8cAl
Zbcw0IfumRZjr1/Gpy0i4lv5JsgKvywKaMB2gBlm01N48Hm2CeIN928heuFcOrJF
6844yI5Zxtmu7gOu4zePniDo0RbR9gpybSePuW3YflbHjZEu8fNnMnipFI/H+9eR
bOI0zOflhbuMMSEuKTBq9/HjvdhnpqYDk0c/bNvAp1xz6wkaDzSwNU0918/4cQKZ
RMZlF0yuc7CpDLETMBo7qHFwdFkbSUyaP1Qs7uYcwEixkFIzJKwJh63u5UG0cQcu
yNo/fInOXipGR+IRgR8edjVcnCs61SOMPfMz5oQ4wtsKI+AYA5AbuOuQCu2xHA1e
d4Ccqh/brNa0pkVQ7onfDAAmARZfh2lXKtfVFnfagVmxvyxaUe08ConQDtJxWWyD
Mf0xAyh90xPG1melG3JxsbKsBPUeu7yLlt+lhE24axKhT/jFJQH+7BoqnhgTdJ7o
65vURvYN/Fog7bz9AoUknT/KKLvj32nVVFND/lfae1jOzJqEFoSN4cmd98QedGMd
fViqtQ4q2ziOzVQZzKNp2Lecuy14uEGiw0Vf7VdrXsrXGhGsWLub7UUVbVQ7Zp1K
VYuUjF95zR+vf9EPteOB6amEFh+4sIHlKIwWrSK10qXTmV2lrBp+oXP6rRcN+jYt
rRZn5dHrqcFxBwk5tlnMKUIVFrUhbg2KpOAk1xC60JHjJB32lZXoq+sCt6CoVIea
Dr/o3k7nKRMoFHq+NldQINFTYccGdD6JGaRyKbonbubjjfbUIRupdk3kqV3ZnX3I
/sgYOG0ev4rXYlbDnu37cxLR/9vmJvyUuPYpyzvLs0ZHBAQProvP12YjMWHfeGUM
yVVXzGo5hZMy8ZxfAnzpjXdgkJjMMh0Ud9/Vpm41wqxv7l9qI+cWRFaJ/Ush+U48
NXahm7PKNVKzqrKhBqTUibQT/WRtmYjdtvDypzudFJJ+I82GLW3ZYrrxKjHm7HNB
bHE8RuoHka0l3djafkgJIlBgT5+aO5MOOvS76JiqVEt3zjrm80y+JZMc58zbdQAb
5Z6NYOb+6XXm9jma5AWbr4TjYDFgAOCXx9gb9heU/FJOddGR33zMjm/0Fus+9X/i
tFgBmKdW2sfYzu3QsJErHPL+i6N5Enhkka6Vr3oOXI5Qh2Li73AGnJ7B2yL2U4QF
P3MnBWWjDlHCK69h6vAbUDnvtWxUe4ciYM4hMAkRM8UETyYCF0hSQW/tgzvDJ44L
f+oRiAWOMXDLo+BphsvjWepL0NynlJKwQRYkgAqMnoorPnPi6teuvvWaTRT4RWaQ
kdiKMGWK6aILS3gBEuG2afRZDHw5FtIbh//WcgPJlrJTiajx1VnnqmXduLIhcGzg
1JgVX6/P0JCu7sc1WJe9z9f8ScgiiOfJIS8Ou2ZDM/PaYPZqIgBb9/sRd3whVymv
VdprH4EtW+XSshEhyykOLfgnGafZT1oP6mxx4g7QUz55yJ5LTLaZy6+jB98WjNym
H041FkA1OiYLlxSdB2GK1BDGhDPe8u6Rzl3ZkrR8en74sWbW8Xj3MTt42BU2D/b7
VbbPIUb3SKc0HU2aLV2qeMX338X/dVCDjFMBKLxkV4PpkiLAJyQMn2iyaF/wAMQs
k60yTT8sd1ad0I24PmrV9mgtMhxh9rUdGb4qUjy2NRzN1VwQpDMv33Ku5c3nQm/I
p3Ik5isOd6p61SYZvhhFcC/rI5YUzOk9+xTMDNmqfsU2AQfETRPYvaMEu8r/HO42
Ngi/UBr3wergq6i9aIVHHLP64mIdvZ9vSY2+C9UyKPyuy3+0XQj/WxTQ0oVi+E3D
OP54zFnpGCq2bJpRgNPmDd1aGd1G2PsKDZi4fvsCKub093t2I8dLLG6hoSsjLaY+
RPJLxsXctNgaDaEJItn5EAG5eYcfhcTEAzw/HVRTxSxx2fnuqYNCkz90onVjCchK
uhalW5e0XfyBn7GOAtKPbhnZy3UzqIau+xdjJJM+I/9sY9DpeeKGSF2m8uXKLcFN
MaoqbANKUivFoxk9GIWom3lpMmsMgPamayJfkwO+YBYDaT8CcXcVl4fDUCLPdoR2
NhX0m89ENieWXbMmlGVVsESG3SrifoUm/70mjIqZZwRI3+vavghc4D4gVFV/Ywgy
iRuN/eadtC5ubGGXcp9f/FwbdnvyyRv/Sk0at+xPTfQG4mgWfqRxgpd2pgB05bc1
zphmJczMnZ4cTaclB0OkCpNDZCMsj9Mm6hwCP9SfuCfgGXtc+q5YDTWHXab/udQS
cb30UMPuyw+4JeJiP874/d01OUOs+AaT0EQGf6LSbD9ZSGkjpwdUsrP77URzvn/E
GeD0K2FJ2m/QhDjPj8ZFN+fXzRpczORLoucbNp1g2otVuKjc2B5nuibNsB+1XleX
iqKE9YH/fZjRhFgYhkBBmXmaW/7cNBorXncxf2oOQ44WXtwgwe9esiH2KOoFeP9F
4OEdccmXstzAhsZAQj4HgVXAJiC5mXo8TgeBh+Fq4FgrmPWzpuboLYysvBJqcjdJ
9HheHlOh2fi3+JF5Qp34w5Iaq4hQU5a53egBII8go5dolNNC8Mh+SuskLgs9tEFg
f/nWsxd8csSj0r75ToyvyBq2SgPQUP8mXQ2C83u5vk9TqLXQbkAWPiy5sl4ToAUw
w4fkc2pMSZm0MzGQ2RIV/baRO4rcAh3MRXdTcRmpz2dCQqHWt3V7sde0noe8e3ku
+yWVz9+sKneAp1m6AZJjhRdurCGQFegv7r0J/GygnB1eByeV0GPWOX4jU2ptX/P9
1lCELMl2ZIFK0Z75VkhNKhy7a55OIvFAEinER9qhhVR/5w0FvgdeaKxtQMpze6m2
ZdYRSbFL03EDgsqRewk5Sga/ra6qt3hSVTFCfKNqCRGZ8G1I0W2epMgHVXj9fL6p
kzgZpxvvwx/JDe/QAmoiibKP6VSoAgud6ybmP/lzyFlIETybyKq5WMcYPVkaxhzu
PSR1dKY7fGPZfjAaQTaZ6wa5aLd6f6+55hes8oPp09lq+UD/cgB1y99jAGcwFMv5
solMHMbrMVukwpFXMKEbubfL876pzuJkfubBfl+PJcuU+Df4+GMAlOzDt0Xb/gte
t60s0O4dicZxuRB12XPY5KalKGxSp0a8aDne11QdqiEyAw7wqKxQtMHwDMbHDXYm
ftAIr9i7EExRSE0BKDhiDluo+HvuhWOrgrW4fQL06LrK+1O1c7OnQSPIPcpV5OpT
YfqtSVNaPJrgD1dv0WsIvzc46Kxlpu8yDr41WRinKvjNVRYZuHEzFB8FFyrYaOTu
LHk1xNkI49brcwcp6bgJuqLh9w10Jtl+U1gJPc2+ql1l9Sstih9/c7pK+ton60QE
E+DwonY1c1RtYtWGHRkNPe4M5nH7mLs2iQFBNiz82KYMSzts2y+kQgRY2wyNa9JH
75VFTDyrnjR+wGxZtCu2h4mYVadkFJybbMZ5ByIYsANgt2nVTlbRAolId69ivOUk
X8qvEo4EF7fZ0NhU3uz/YbAXoxplyfIhqSuG0cl1Lta+k97gi2YQkqSQ+QuvyvJS
voYr50gbIsKNcQkvYGdPzBpoKUNLD4pUj4hJIEhlk4+QjLpQjxshkwDoBBQ3Oq5I
u8j54u5MUTCb91P7IOnhzEY0l/IkQk/qWijhZLsvcy4oOcFnx8QBpQSO2yDL2/UD
Og0RGjx1PSv6HSXSkqmVsR3u8746kNJKQcbUaI62beHmlt375ZPNq5wrWTURJkh6
nXnqWl7CotLhh6rQ1yVQKBP9R/P6DhNap73TT5/od3RvK6BWHu0a7qVgnXNfES6P
/uBiJsHE/84btYbU2PhdwvVAiy5EPew0/cilh5JBYtF46JQXbjiJnOfLQxc5aZMN
P9Ew5kE8ZpGCmXNKzkiTdjdclsnnkR1QTuEN3lH9B5Jav03FnCIDMpLx9pHKFUzV
DBGuZLw8+7sffLAVwkIpSaQFqYtJjFuRGhOBiz4mLUbMyaGFPlArKQTWEsATSeks
1KOFQDVmfsItP7li7MXCAVqXVfFEkQrX0cA+puDqdDVqRduxxYpH2KnyuibOG2WA
Wyrkjsp38Rwk1SzZfnjfM9jOpdt2ZfaIuozF60QQef0ij+AQFvTrFynYpXC5CtfV
euLKWS4+qWvTVk5ZlxKRhNfBTE/w6NF9w6BNjWBvaOmkrTCwjm/Bp0+0zajInSBq
8OFEh7wJVisem/ehzqbQCiwGuVvLsQuZIsCV68t5ny3SIVknvGBZlXI1eQzvG53Z
LzVmfZrzhZIeC5t0Yj59ov4ge94HYpv12IG4RkSLt6omALdjIP0xs6hbD9Oi+PrK
DxHpJ9Mr/hCoNnpyWOWWcZin916PZPXCj4ppYnb5Tj3fed0gGgR8ry8lwRfVlzdb
/8DZX+RdeXHC4xHr+nW8kPLz7b0DGfTGJw+EPl044FK95wOVXkPFuryrJ9knyIv1
6Z66O3FHkbjx7rGZK7ooO26gxfLZbRpx39t2J15GK4qbWqWAne8q6pLSnvq0EOnR
1+ZJh6k8tN3yiGc44EfyRu16EjJ7Cd1u8x+Qe9/zufrpobuYMkZ9xpgvM0C2tirI
bvmqTdgI4Haw6vcDxrEtb7wsTF0pTPRCCqC7DAWJAQ5f2IjzB5CzMbWgwgImQ7V0
CC9KG1BSyOOHMdbXs76Hkg8mrd3TPM+MmE7UrRSoltOO8NrrjXs4EaBtC2ILxXcE
R10lDyBqbcOWSxtbj10NsJfEUMbPbCb3H0Ucasy//+7DorV1veZdcnQrYT59SwcP
94qLYOjzn7E7V32iyem8JQEWS6L0zLMSn/fjATZ3wn1FMuCmR0YFVa0TltIn6NhQ
QLfb1pwb4oekwfJ+8aEw2BqQilfRgeHCd1jQMhOzT7zOO5FoGUGAWO/xNQo8etvS
dCV+3CqPRAvNZYCu0EDNsEadntMSMsOZA4ChBt9jbAh+tGknqxnNoRNP53w3CCOG
fuLG6KqSqOIRcZ8RZmfZ8PWB3pCOYFQ4WkqHKDD9OiNKZGgbGU/RNbz5QgPOKKRC
+lmkjR/Xl5U+rm1+bQasNgFEqd7pXvC4hwM66ifxvoPWK66MnWyFOpNWT0fQb0dH
Pz6Ps0CCK+StJGlKX6+73T61IMX2fBeNq445gGV7D0eGx041931po4t3nlPyHJJI
Vv9GuU0NY8GCqOhtKnhyZBvAAsNp7B8K6FpY4nLVuEf10M/Mze8VdYqdbtn9IhBt
jfuL1D1NlS21gri+Iy3WA0QJOccoUijrRM6Kq7xB+Ri/H43SCxE0iq/Kc5limBQD
P+AKG64bQdcghq7afcBe99tmJvLpEaqgOTgBXXozxV4H+fX8V7X93nemW4oRIBNN
csxC6zgd+XxhJuek3zi9WH88d7WEsOq2VujIb4685A5wRBJCP2nzfVUxOJ2Tjiiq
6PfpBu4podgZu7/+ScMNno7itPXGSVNpu6SyDIHLf4WA/wjwdPTwYWivp1nXAwUN
EYYV7kquq3PQSGjQKI3YfOuVghVkYhdtLZZ2WznUK2UoOLq/5DlqfFenhMVrjXXR
4SbHnaNaJ7JlfdCX/vdu2voWV1XHi8KthH7EYTjou71aklSrSmf7yfGKa6bfg2oA
5P/DhYvsF/fJEkJnHKX3NQyiL+d/60zsM2dYYTizQUyOzL2cEZ4JPy0b+O2qgYVV
yHXdmaSyD1HQmnWuWniVKzNZ//IH+CyIqFT42aUrZ2uprLQ94XDpMnVKaVVQbF3G
6Urn3yjaDglk2Oxlw0d06zpjkIkR/wGP3KJQFXHj+z8sWExcsvm7qB76g59qC1FX
DwzjLWc6pIgXBg30RG0lorE6BFFJg7P6EpaMNhT0op3CUrOQ70J3tNW8Y+V1QBKn
t5l5oRuu6JpLnJMbw2ZBBTrtkoXBHkUQ5KnQwPyKuNKgdQ6KQshHi14jxO5XXiPg
AM0/0zFHeyFRI8CNBqVa/yCo18sjC/YT2833owPdnCsMdgXEoc/FI9SscJKRctQ7
bLe0jTUqTDUqfsTDPRkZuYc+NQA34lD9IlGndh4jSxpvZzJcJEtAaYd/FS/0NSyR
vsMxMovOsuspXzGVMACfasjd2vt0ZIGSroPWkxeHve/JKVqCv2NLY1oYhEM++Em7
bX0hhaZSd/7FubiBZNZrSMhkK+LLiDUn1JNWatvMgnG2RkuOL1JM2jj7eaQjvS+K
CijUZGEiN2wxsIsACYK4W3Pwqm8Or/ah698fqagLQt18/SGyELxRPXVKcqPJK9Nz
9fmtRUwBL31CFGo7+jc4I3B1LF+H9FR7+psiN9TcieKtv8sYxFAnSMOWr9LlJY8l
rMZq92bSbPHYg1z4tVAPCU/GQX/hZdfJLDaKdfcroc3DnG+Kz6fhCYnSaFDl0XS0
eWF9u9bsMLE72lo4f4PUza2GwTX5bNOSMDxYD+CGnb+v0ORgkSh/aHXBbRnpFYpw
g7iAs7eniqm9hhFbmapqUYAO5DnYfW369cMqaQaSaTt+nNZtbdAtFRKTBIJFLJ2O
6xhtflmKRIVH7MD7uyXR6IqR5ml/mwoqD0IAvBZ0IcWeJycMIuX3s8aat42HVdAe
qEYP3ZI6w+sn8VS/eMpsp2naALc5z64G7R/rXBkUOG8cYBVgCAatXXW7DbQYppoH
yUPLqMcXQ+7gj82RH1cEN6pdD2G15XHLfAVZy8wRgPWyDoLBUbEX5wGjuyWTMPfO
xM/hoN/FOaQIJ1BE6ql52gXm9Y+Oo/CMEU8r9jzbnZq4b19UEhiwFkhTeN+jQJbY
2hIQvfchqWW/+bxmf8u3tTN0t8XcUPxBdwzElub/SQ0dQV/5o3rlMV5IRDzQm2ar
SDG60ES91ViSAThLSOOONcsC9mPF3/dcy9xi9wGjTjBrqnxxxNyq2HvwusVKc8P9
h6a/hDlq2gEQKANVhiGDD1MNGgYVCu7hsvHqinMQrhg0Wvcn2X10Vh0P244kys59
fqhVhP49EzgPVO1YaSQ35mhbuGeSF8CQQ1VaYO5RWNM+8BkO1pq2oBM//zswBNv+
9wF5diaS4L2tnrwHPwMmdbXvn+EC/WqXobgb1aVc/SaoMCJ7+j+GXbh/RDrOWTEb
cIENQoLnJRHJLMQOV1DG+FSzHLzaYPmpz1vpXT/WSCyI12y2ZL3ZmMvdlio3D+1l
I7k0IfJs7fIS7tfkTvObdLYSTo4aNkPbbXQimhKKU0q6xjbUrmWIf2PlLjAcToMs
O18zZVpq6/Q7NeD7Sy58rfDcY1+yWorusKqNQhjVgbRX2PRtDXC7KOG2xYQQWeVk
x5Agq7jNuhfg3cE2ogpBsR+xoa7CWJBYw0rZGDeYE4nVimdxQ0W7rdcAMevSIrZA
JzDVZza3vQ+MCthqiCM+3uz2EnGE8W3TJKimPgWVmMl8N8hff7MvRw/bVGe3NsLS
9Cqry85wWPzCIuwVe8LIv2m+tK9DUzJsilzlRMmZN+elhsmaAZk8h+1DijdSxQQW
yqRRT4LfIPzQCZa2NOQctP8R709PgA5L/UFzmaPbV8o9v1A5XUwoM3okZJS8R62K
x8FGdyg0nsBh1kfuZ+pVBkBtMVo1FuH2KYecD7rGykT4DFwsjZkcdF4J8XHeua41
79w2gNcqHhCdq842XlyR8mT8bQHKCOOjpmkVEOcYp7EtnxEkZ+kMPWTiYLgZQub8
RfCBmch1FGDLKOTfsVYtK2Oj84qrcIAYXxhq2UyqcPtKUFCaXsIxshuAZXe49spa
O+WpK9Gl/XQz5ZkADjzlzSD9N8+mS/CtMsuOU+3GDThriCwzZ+hVe3QADU5hyLG5
o6YT6xhoZKAKXtEQdl8uDUrhFdKXNv3z60eal2dU8oU5H3laY7XV9bn3M+3rfnkL
AA1rW3SYl+cDiOLwnIWAkf3Y/LVuRzRrHUgHAWPRCTOPA41Fv7ZApaNVWVVf428v
lmGZ4g+gCE+2ycpsOdtztxe+IWJsgwxVpyOy1NWhBJ7QqfFlOlX4iMJLGPocdHmU
CtBKGovnKUb9UEAdt2NftGvIZOEparfsm7UhIFIVvyM5D8p0OqhcWYwiDpbF9FRo
c3pCKzbHGFmpfeGbblf90CCeqdLxS/6RGPF3DX9na4Xjnkq7yzRS5uP+kproXHSR
khkl2D2x4Zxebwg5qliugK/SzOiRJiU1Xp5rdxtbgzhCLmvSIWMADJWsyoQhJMk9
xLiCZHRr//dBi/esDdgC4ut6/6oSjaREpV2wT2t5fNW/I3zspmNeR3AJJjea37xL
m87Hbip06qdPk9QCWcN+Negd6z6JplPMfRMxF8fo0XQpOOYM8lTu7nLJhvsOSGy3
5NCa1QGu8Rze8ifp+ARIIsGeb/VrY3t1lJ7r+tG3UH+TBIwIQkk5jFKuMS3ZKJ5c
FJXrx+nBLGlC3V/T7Fm5KbxFnfe506nsKJe0La6LV0f0xf8asw4/F7acGUXz+xaT
boD/Y9Q/N4BDodU+nb9EsV5cCaGstNfenShqdhdcy648vvM1lVY5+fbc5c2HWSl+
Jw98vC3KkdF+fTPmk6LblJ/855I44haRVDCoRqKGDAqroluUlMuJX/ht6DN8xc7Y
+1/EBnDZRmuXt3BP16Dbc3hKmf5BYBYKWDtWRQxpkFByiNhsh2a2yuB+52GibxlL
IukbTieUORK/MiTlVNMOvJ/ZRmIAGiJUmfjYIMJYJVfVCrYVQlPFkM8AwQmu8Miv
/x8khg4vWWmaSB+qo0O2l14JYxvgngE0lzi3F2F+MbPycPFiRe20iRj9PsEIsgTa
V/u7Btyqf02u9RpSrW1HLcSfOy2pdQjn/vrA2JaCQOfahHOgDYtZk4BgagrRii3z
iUszPm+GdEZ2W9Q3gSQfN8JdbEgNnKWgSrt4LDaCIOZR4TyFyGtMZT2FI8LPnYFj
/Xl+H9bIWFPncYLV1BWZrbfAblHsYR77eJtRXyGNeqmlCE30VFkwn/uCXk79vFgM
yd3ODzVkv8fb1Of7nmL0NupPf2Rc2dPfM/RoHVM8ftp1qsFF48XEmJWfPCS/B/cg
QnYToDfBs8H7A1uVtCZp8nLx3FrV89dfJp5NkI0Msn7yLtReCGF1IDfd40o0ObjX
f0LydJ0k4jAmqnR3OwLB1vwamKdB7hjXPt+9N/OuvVn9mNMCWqUa4tjGuZqFxvnB
QEbn6y4sm7VHc/lWV7RdjKY0N34BwIWAVJt88CXHV06k1z7xKyu43QINWHmL53pX
fVMvK44KHJYkOLadTudNLFJ+kwrdV3RI7UG9JBIOU8N2aOWlkwB3g4ToKjYNvC46
WrIoVmIeKVEhjifTNTupvVEqvcbY2ImNm/dgt4FRIhfbDYbjDBmRrMY9ND1Yufvk
So2l42+BM6Z0qT2ubDnfwlY+FJFq5D4wvkpLe/CJlF7Ic3J0Vhc8gisMCm9eYxFq
/pnGUGxEZeQvI6CI3ZpJZquoA7ngFpMZ+Y38ieR0nOVNZDbjbzD4aH8EevS0/oyD
HZtaYuDsIXSbhsxsoqolnsZ1ZBTqP4WQkmy77D+eK2hInerhXRFWKIMsYgkGutBO
c3nmcZVRfdD7PQ7QxHEfFtpAqXRZUgYRltv6AHDa5gS6qhaj0M+gzsROKHORbVO6
ZOhsx/PfPz8xGvWNcteHZTjC3er6JrIYIqQHZlRPMspxLtzmoWsgYEGCPedPk4iu
vJNawIk+WBoc7oQwNnkixxf8fMIhvZl3TBG3EnipLIKqkmC55N0QBdwVCa/mpv/k
aXwT5UwHJSxem+KZ2n998dj0rGEhgnF/X6ZoyJLuiAPsNXqxAYezgEYe+5v7R3ij
y8+i0z+aeZKFCIY9g4CN9f8KzJgJhiMbkEDlyAMoXFCFTSf3EmumKp1A8tFXr9oh
5jfwNGQdZB4IaVc+zDBAJZ6y9SYLVYEgOf9u/IUT2Co0WTJP7UEnEcm/9zrDTZZP
7kgivMC76amucOCsnGGSYkcEuxwaW1dBLIJMFZVAasTUlFnvdTbH6XXQUA34Ylif
BhfMx31uIKit/7xQFZ6DQvoGQagIJXxoEeZIPnUmKqHNnyk2fJ8dMgW6puM3kUUx
VR4dlsgk0XNVnqQGLBRXjXyMH3SQy7W1qTCygWmjo+2sSaCTgOnr2uLk3KrRn/Pj
uneDR+tYCC9ROwyzw8BlFlDpE32U3eUun0aXDDi2IWkacP5yyqrxNQNy3nWm6pSb
bCJFkxRT21lv888cGK2zM61uUmwqF0kVDKSYSNVxBH+3+ooT7HaCUeoXM9VLdzb1
SxCVH8lBgTN19Ui5vESCLLliYH4aBDjD9AzVB9OI8l4JuXWdkNm0O7MKPFDv5oK6
4lpZlfEO4ND6AT8iyY7iwgbh6SDyI8f92Wlj94CmGUHuzqSYulrFgHv8bIMizaJW
6+2NgAqmvO1+ZIoiGYNQ1P7nrpIU4D0akNvx87b1vJcpYLTpBHsEIU0P5BeyF6Zi
pdG38jdQrVzcRZonjmAIxEAiRYNPSjXIqIDLc2GqV59nGTRQgfD3KgjA1u5Se0UQ
zR+weQ+RQhoHXDSwEvd3XFuMxFjCAqb54M4RbXgpi0Bx1b7gM6K6U+2i8yiaTkTU
To+Wera9Gc71kycHnqN2hzt7nR6KniGI87h4y8if27IPO8zWjxYOGmBrNJVguQwo
/Lsx5fAKe44h4dQQTQ1FhXMqQI8B6nOcyO2R9ylqnCPgnvtVgOWHRJb7zRMH5oFz
yOjuxh/uWZosiTBNnjWrzr+LpNPWHSwqwUe0aYnDNTRrdDNsLT79phlJT93m431c
OFDETc521IrG78TtEoj2kKJUiOBQS9+Au3wV4kfoZmoPhW6vYSKWYrhvCCitXuml
xAW6aVJwCTmNsHYEZ9WnG7Athl9vtHgbXgo7PoS7fA/RIw5nmxuBsopRObpNDQht
dNsu0i9a4Snw8mvO90yujJTxe07KxfUvVQoxjGnoVrjRXk3YO2bsZLAxDqBppeWa
mf+IKmRiknPSLB7G0MrK0RRrJlXpTPHJ5Dwndz9uJtKees5MDBhiyPsIqTOzz0Qk
T/u+UnA9qqBBDVmBykBQ/0xAmAFVFxcUIHcY5smlr7YF15l8vB8nUs1ndrq+ZD3U
jM7wrHzAWXkadQm8Ic5+5dRPJ/DAj7PfuTfnNWFgOH/EQkRGh/LFnGjImKVSK2eY
rnj7N8By5uTtLDKIDpIjINGCbY3BhmwMWpwwzw8CYfSmNUIAHDetSvLktBigR/vu
zlXUpzL0npx/G+7qo2TQ+ZbaGCQp97Y+p/MjRoslgsynGEuZP8AmrsSCqe1Eui0f
42toF+6CKLEmwxbC4r7A5UfAElvG1DklQhoerPdFojPRO7WGxyaJTCXAw8blcCie
v12w7JBuSL2TxObIltR8FdnPk9+XS50LsuTIMt8hisk71j8G9FOd1h21dspTPN6c
fJXzkiN99GXvSILvWhl9KGr1tfImywnYRAWIF7aWXli/PILyWDwKGOxl9cFRRYGh
I6Xr9K9c+1pUM7vXmTNSQ4K9Y2GfsqyH7x4fgBr0A0VfsdOW1gXltqBTXwghiC9f
xPaMB1vA1CwemkHOxqNl8favjFMHupRwlmBkvb0HoTmoujE2Cy7IgNdwf5ThUUr7
ZOaqu1Ej+pvxXUrYFZBqGnsveJaLRv+u9PHjjN7qcwdtXh3hzJ3U+dA1XLb+NY2A
j1sOo3XtbRo5I7gDgXq/uaLUfKIhaul/po13uvH1cSJJi53J9dMq5oRW1HCM1KSc
13gbgr+VoBlXqIoWjjqOpCL6VDay/hudXklg+kCwcSZA8CX4t2psQb5j7xTOzbyI
fqjiscJNaDCLslIG3DLDvwO3WqEMseK+FNAc24ZguYljB5KWRKzCh9wVr6VVYFt2
oxVJ1f30XQmRwEWhyZPCgVYXkdwgg0LTzOyxf27mSqT2W2WO93W2DOe9VezTjLG4
lmoMMEbs1KMUOq+HSURCN918ZFOpo8PnFD1Wfsgn3egPdA5tcRivijckIEBrgZwN
UZy69gjebmF8knRsnKzmYMUeEDykNtAFJV1PAX5tD6rnLYuM72GZfOFxTPDSjAl2
hqNXq7gJ7s1BHR16Uvakgtr71i4EdmZ5NHKeG7bhYQmlVioBpj/cox8jFUoyJtFY
sF6vCAdsw5pQ/gGcrmi6EiTFGs7TQ4z9lEuC6Wpj+gQciWtMlVoUVu0C70/LgMiL
JBpMOtorrhPDI1lW7tVuBzfhbZVAbd06IOoUOMGbYi/2dG1rLZ07AWu9Cjpt5o9V
FRC6hZaB19uIC8ImFRC2YMrgO2uYHbLVWbL7JsbaxsAi/71ylt/TaUq8vk5ObRJj
lGxIXkiWwp0b4M528gjRZou5uy9aDa9n0jsCOLwTQ2AYjOyVNr7v/ElFqWm2SLji
ZNhR/udWoC6XgP6eA5oZCjATt29Je/Aay5+XtR3ZJmZINMYCO5jjMRGSoRKdmKRl
kekvURb/q3lLEMbWU3DXVyaHl/fMp+6pg0HHHqUIUaKT/COdKaJ1e65mYctukhvz
Mb85sVzY5Hrmr6fX7utPZuwZyd0qHXQYXImZ69q3blRvCxm101dbRIg5ux5gDjTW
AuWCHs4kDtyS604b3oDaiQUmVcCmbys6/2NjdlTQaH1dfA6iQsT4JnE4w7JAzAm+
mtKEHLdWDjRj8VJr8oqes0o2tj7xEMKbGuYCqfvDRnW0ZrJhobpDx1BpWwk0iaye
c8FQrqAfa5/yvCVdQnlJPNzyKeWI9zGolp33eoYhsM//hALCipxhkaouJSKFv9dz
kfaOsErwYBB+5vhHZLVRoYoXHa+eaPTpjS0tmCV3NUgQCMmQlxkK88tNn24YBJaj
fTmb63mx0JjBagzyS/pDJrjteE3Oh1VPlVAS3nW0BYVd+7ia9y7HjFPlZqviC1e3
LO8wPV3S2jXGs9QVGTNCFPkQzL0kJWK0CiSm4FuzuUKG8apnT+U/ArD29XmKNj33
jOWwMb5toxIFst4IjmtPRIDnC5cN6XaEOvzwdqstazrBbJUlyoGPomn0lHu4nptc
pLCCI/vZC4BemxlYRhFShqoIlqIABeUpTYww0L28TaomMqWjJs2oCAA+l8vJ3Uk+
AbSuLv7Dkl8TbUbeN4p5wjbRP7f9rzvpWfSf+O3Tigz4/7lMF4QW7L4XVJiulyzp
AbcGmQ/ZpFvAf+VTUEGNSN3ZAATAIwCBXDAj+7cv9ZG4cJS6PLe2nZYUMU4+7/Wl
XiYJ6e/5QU2c/rqXtHGOYqHmKCA3Otpw0CNKbA0urbJzuZPg7dPWQ2PVJ9wnV1uU
feuWns3lstdTc8JVDoecuJoj2u3ONvQjbhBmNUHthxNnTVyYgpZBb7WZQVKNB4HT
pk2I4lqogYTpynulMIQMJPqsYH1AtdhQhoUrJjMM4pxjHn9BCocEfhMnpnoivcQA
XXI7X2/NM05rSvq89pr64rgn9SaEyrTDSaz+NWJKJKyKysH4GvA5vfAeBssTy6qs
D+YTnj5BQ7f/GeC3d1pqHvZx0LjjHK0Pofc4oFOvnuVE4vdnTjVf9M41rpHILvfR
2FFh5w3jiTqlJdLWTRWvgjtwwovMFMYEHFBil2kjx3SpUajTwFC8VSPhM/ZZjtKr
lYDkHxGaSfJOIyYSeY/k8nheJxJbax7GiIiL9z2mwFz8NlNEMCCt9RqdMb4g1ntL
tOmkh7aPrXLOns6j/TOhlB3vfAPi4uFO9ZC3XntazmuqT5ICEadkxeJP+Bp//vdh
6rNZ8A2hjwVfgJGkESreOk0+yl8+kUeG5UAiKb5wGNZkbZl8ECQdwvrBy9Wf3G2h
xrbOxqVllOPbZji7Lcqts9tZTwekIBXPipAZhd/PCBXpvT/KUi58hPAaetBmeaoy
OnGXdD0J6oigywLFB3wrRfFw9hZXETcKo90RYdkeBQ0n7IzfrndJk9CKHfwUcGID
I9tLpWrtoZxvIkXUwFUNuHBD6sMx1Q3Edx0ZnsxAeXBNqAnFeDfVaZnGQXw5C8Vy
7t3VVobtUFUMogX+ewgHLtQSjIUZaY6a2fqkEvfLl6o7fz41yToTimbXcHW9hYZ9
plwS3MMxpqc/nyt0gCaUSZrHMqnR1NY8E1SPb8DmTDmoPNEU0R3ntIsoRwzgQI0s
4UJ3T+AldZkYPotlJGvAViXs1y4DFCyb6VyHC5XuuikqzqwBCukHtsqblQwYXlHc
dCgSuVb+KnbQ3iWIOwTH0GiJhzuWbTus6hyts1FRbAyXlS9P+C76gGgXrNRa473f
MsPdLvkTsB38LR1Vfss1Lcu+OK/yr6lK276XU41TzDlW8vJt7Z7UdBIewI+4N/Cx
w4NYJcVEMIW0zacxhni+k5qsU/OojaSh+tMliYENfTr/UgfzJ6mPurxU75dahD9P
hDQ2Xl8uTAfrtwNw7+y3VBM52lW371WwGbI/pUum4hbWVwPnCtKrERRyZgVvK6Nb
8+laqhDNAk88tGLBmyPE1Nbh9qHmP/CJ5+QLKa5xxsN3K5T1gSyn0aLkd1CTMkxc
6eR36uL0X93g+2qAW2mmVXO9mzPlbhszYCScBzgoTDoQkv4vSnX9i4Zti6iWKALn
if1hmvnpAd6vAusgbe5E3dlhp4DgNbRhoJZez9PFvnqjBBFVK4TiPhE/pAjxobtc
Y7fJFAUejqAOb0VegRLotexf4f8h97FQvo00CNJmD6UY561XUCFhob7zyTgtk7eB
3TNuPWyoL05PqqIYG3vm3VzA401pUWwb2coSpT10a/xt2eTgKCuWFYujTdE+9vjG
zvBf0uDdPXR6BC+0aCIHXs8mAuJX0boWFiKjtNcjSt8Y5S76RC006t0kdXug53Z1
rESkjPsgiCqLbq88maPn1s8jOtRoO2edgZbnEkJiYqps8EmVStF2PFnylcSRqbQi
zeFWMltltAixcJvjb18PST41Bc5/DzNKv0Fb13HQwYExUWigcCuWAQrmeQULuRhR
r/zwS0ohYzK5fJFKCm0Ujv+T4rNdSHwMKGeLofo/lUq8IYQrnxtQoPaM8lp5dW76
Lc/hM4Ifrdzt2FsXhRQ23lxKXHABbfCNosuQSThGmDzpgiwWkIMBvuuhQ1rkSHAl
s/j9gAJXDhvMGWMhHn6iMJZRqjQxtIJ3f7JSCAWzQ33Qp6r7wjCPuyKFivZcRyLH
ygGVqrNmyITC+toLQ6P4W+eIBO9sVvlFofVjl4LTf3fSuIFQ86G7+6DTNBh3Z3nb
1PZGwYrd79TF6oQdU11II+SGP3BQIGO8rL/UN0M9eymXLnw7fDDZQJ4CJ8/i5ZdX
YKPE3eo8uaCGvSy61coivWhLCjN00VE3Svw7LAO9fEisjCm2blknjJ/PabCx0YP9
SUM14Ktnp+aHcOXEELbyWPCQ+pZ648R0G1vJCU6Psy1Ockatn4JegX9bZGzeOKQf
3GuheTcGO+roTwk5ouSgAlFvlGZMDaLI3iqOT1LrJ6dzcpZQ9t2MgV7/BEbYmRqU
Do5bqZHaGxzb1j4DvBj+jigz3GePUROAcqjh17XWXjq2udjGRlykxUbjGYxpKmln
IN560lIOozUiVugzmIZZ3sUurFqMCAr0gBI+nROG5WPcuSYO//mKe/hOMtH+MeNX
dtrWptVWoWSg+UxMjXEnqcvUHL0MTMyCYmuaAr5yO5AYyjxD+WqIB+8N0FYVrtBh
4za1StvvoJLWJnvfxQVhqN5FzhwY+Yuhyjf2VsQNZeq8h2YoLRczIQfQpwm2K8rl
PNLBir7dm19IEeSokLDoDfY2nJK5bFz0ZtplmAgkNGRvisWJbksZauLiY6E4hhX3
I0Q+e+BdvE6mDQqJtEIdgqY4XSSTWlPPeSJWDCO4Br08WbeGk3wCWxtc/yILWZ8q
wudrD/eHzhM7xw+nDZtKjFfjKMH3zwD5rOxstO0PsbkiiQEHkLPOoP8GTOkebtR9
Bq4H6iVxYNpb6Hrbn8yqTgwjVS55rD+F+RSWeGy0yV6KF0q7kf/XyrzQ8GiNdoIU
C6rOw8s3zWKMJqBiXLAcaBQnGE3AbobGjjWdX5USfw5/LuGF/wcG+EC6H+Tz9OFw
S5pY1nXL3M8hPxCFHRxMWfwd2mabgDNYQDPQZdzNZ+LCYKAHhoZWCbnzS7+v64GH
GDwUSJPP+4q5qxun0BZrRgKlp21t+A0TM586Ube4LdoWtxrs0yMtnaEYABVZq5Zf
3pMuUcUw06wjhYw7zbdAtalT4wFJ5tQsKZbdumiEbenzoXppwT5eZQDofIoAM/5s
hEmATQAkUcUBKmQm0QR1JOBh4Rt6jCDKVNzZ2yyl4OmWBRPtZmX+UMBr+eR7dn9u
gHgn22ZJIki+0NkzmoiSBloomeAeB+qF9yKa//tLLqpOIaMfEoBVD4VeNAGBsgae
HQJW+/WaZRtfnCPWxzIwuWnxxb5lWX3lAKSvPtcDb+imYZP4E9qoHmsWpNrEasj/
OP90VC5AvabSU6buImSU9cF0mUqJz1mPmGFOHrYNqYHe4MAfJui0aTDu0WS10Js9
O2JmDgjFmSR+hvFghr2wbtyjPZBtwYCdG/Xk1OXW9k1UUPw0p9KYyofIkyaxPS6o
qQJwwp3NzDNpwnf3OczJEkbeh/H7Yr8imnAEVlkM5wA05SggGG0QmcOi6o6W4qmW
i239hOyht3gOsfOWQE9Bt2PaxsdhGGPjvNBlu5gBQVja8nGbk49Gkui/31qbBQCp
kuADQDttdRRw4eNnf/g2Z7uywwMD9O8jzcfupF6bzO+6LxfpSl7YgyvEqLWvBB8L
EA4uz/X8/x96V1sHsqGJoV9tNyOGEznuQCN11irhviBzgGzqq7hOMqkFupYuNal7
zd1QIINUrNaicsgbNgJkAWxueRsh0uD8daQOkuZ0yeDLYEYfZqHIPvFexHpnJaTJ
rRwO/TGoPO8/SUgPWdHlprh98P8RuuSSy9OiMA2xYpa9JtiQLE1NegcLbWDGyZU/
InvhLI2kzRxN/PC+AqINskjb4qY8zpMdeNi20WFNI6ACJiLZdN9K3H46lxif02Rm
Nd5moFal9T0vWWC37ULNvZIILQaKc84GFDv7R6codoqtHN2k3m8BMhKuUffIT+vh
ORJkcBYyfBu5zpCUuEE7hnp0xM4EkIIbUZgujtkEsokXM+QnA7/gYd5reJj6FxM3
SpeQjXW64RurJEgSsFddKMnAytpXx5g3tSdwcRp4xt4coqkNHrjtxEOXIB9AUp0K
BomPHOIBb/A6tpU6hjlrLBDq4T01vZdRdPC8OwkgALXBubDROBlBMJ0sQUmvHMms
DVWqEWut8luB1gfv9wvZbWzRv3wYlvCw7s6AvYTBnqb8HBIsCIk846e1Z0BCJnev
h3rUQJYBMWRP6yQqlvUul9ckR2FSX5MzjTYCSxCff9WnEPob20XrJNyFnzv+XrGv
x/WVWAICiA3bsevQvtPliKQKsUOOefdqYULY4YK3Q/L8Cl7zpmSsj0WMicTQ3/Z1
x1L5dJvV9BmU4cdPS9Mj874TLr2oSrsIz9dZLNRY6xvsSmV2Mj0KfyIPK4MwUxUz
diQgQlEmdeNvjqk5trm4lCF7XNxsf+4q2SDd00IRO/3loOXg1YFz2x2cxnS4VVia
DYV+dI6YvldZ4RwJSZmsBc19+QKhMv7dPyI/wyUQThcQv2sykorETy8sQcploEwO
B4Apqyga/uOfnzVzbGBYTBih/JQQbC5f2cTF+x3aPb/kJV4Q2SRCmA9DOq3Z1EY5
gMm3TAt2hvmCTWFKC+cXfn0ifd9YrtZ3lbeyG/Bwrw3rPYRPD0tT/sn4z14nux3l
b5zyfagZiIS9w/6dLi6fzhwijDH9jQLC1+YrQlP2+zsYW+qBsLTkgae1n/1c1PTc
ClIpjk+/lNMewOoP3gW/SE6vWZaGlA+MyVzhOxlnxeOndceM71wDe0kbpHDWbSCq
ygzfe7myAKHW1HNEtwW26lEZF/57St2g27NnG1nbEagAJ/sCiWlX1BX9tuvHgbxM
qC5Eb/+zci1dUNOnDyJmbgZFufpE2G9avz4rAzthVL//1I/BbHV7C4gE27WdBnVj
BaaREgx379K+JSNIofTFZ6+De1DgMQ9Ys0T9gAHW1BXx07YanH5QEiHhNmaTSoab
jUk92K4v1pfRru70KEsnvEsMYWjWK10Ge9Irfd+kBuCZSQ5uuO4n/z+ti9cge2ab
ytKGwjWLujtNAPW/4CB56WGBvx16v4lXk4mqZKuDMuEScmaI4IyzKC8mCdTot45b
j/T1eN+9UbqvEdiF62BlHIF56q7dMxDopSNDznIrvZGtExBfPf0eeydAaHYXSxuN
vYypEQRqMVjDsS9Qcx4xs+qTCRishPddJekarmvIAtOucI9w8cDb8mEdCvRPX0Yp
mfwmYFWNbrHqSzEcyebEE1OM77xqMoi4cNj6Y8ucSKdl0z/MxrjAcnIMO+khVHpN
dK+b1uDWjj4yUGtw7olsDcbL0PzpyMyXUUbYAQ4FupSQ0k9Xej3sMGvJ0vTDfN7O
DKH7Zi/QJKIbr2Bv80zkl/cldOTh+lA5ULvXSq2Wb9Ds0RVwX9FtkbKioFYWZU9o
GdE03q5yaX7kdUYStM/K2fTyP9dvVufq3kJm2oul5+GactL84IU82u8JsCIyiq3e
hQ9TZigkgwV17vcKCbXV0ub8cyzxJFIu2T8EGxC9WwDLVjfjaa/e7r/64FJ6fMS2
oww2Qp+AOY2pANJLd0Iaa0EuZRw55RtFCls7IwlC/ZF3QWXpsfm+piGbgMCAMdtz
+G29OvWyZ8THF0Sh1yp6czPWtr6czINqcrhMKDoiYGpE9egLr445ckAyJvvmo2r2
/GpdOuLADZ+TLq5nUagljTksZNUR77TijS300BzNCmB38kw6KFVs5GYv2lN3Nhzq
GWwUsQyp+f2O2zgd4XKJWS9DeHXjaAhIq6cRMyIGgziIupd6889I/MwoiKiR0rs/
u32TWD/Wssq5nDbcapAuX/xW+hYqnTD6Pf4y/jQkY6qd6ptwYKesFIv4rYiu6CVq
6ro3ip5GPSEuaOWvsSD9l7a3Bfy0Waij48WWkj18/PcU75EpPeirxeqr4Spza//r
+9ShO7cav3BddMYurU7QaJj8QNnhcpJDRhCYg9ADa3zbvg9fuIqAIbQri5Bdjk+n
f9Pks+xUhYsRTEh2X6Qbz9hz4iXqGI55DOLfMsldPRsQBau0wswXaZihBdwmDDBs
hUP7SHHWIbji/iMJB0bP+6ZJPprAr696TQBN+MLyW++ztU6ze4RRlNO5XO+IEQmT
DSvsQNRXaabRwDsVBUbmqCAtD1zH88v/Q4NGenFAee/TvdW+EF8y9Tmdczto/o0Z
wwkcI3NLQ4eKY6hKBUzbW+eJY2clfvVcc05vPnnIhN/U2DqT6Ife38OEMuZotivX
54X1pLZaqj1nPoTSR/gR/UeazToTTKe3ZqPIEWMbjPmpF+ygCyB0h2i9LRGi29Oe
mj2d4YbH8U6MGLDuTgW6CsUm8XdH9ikEltShmaInCwTem5MpvdgcAoXWu0sIlLjI
pDEb1FKqOBwi87rCjvWLM4lYXLqhJwvqiFCBWUEh9i6O7yeibqE8QQuEZ67ksmOW
n0EF0zx369iosXmaTpcWQ7/ausUF0shneQFMyo7LfMsVgXBK+1YDwxHsb8ZDSJT7
q3Zs9YGZrL6nENS3aCDDou9ZQGEZyUBfzZQedhsnMMWo2yDObMauAT/WkUBgfJtH
+bXoTF5CLBv6gRYJkmUmRNN6DnUqkVP4c4n/xeMWJJJMnzciV/rkl8LHj6iDtKoh
stYbBE8uXg4TXZjmdXLDkvKt0W/G/qNxinjD/1rGRnfWSiBm1gHhp7jc3dQrchFL
ppsmeytkOna7ijXa+UWHRQoKo1YUGd+nJuup7n9+zN1ZapyAACcK6gyih9RxN6G9
Eu3tOn0z+ZkrlVy1qydIxiKQxTAiyvbyEl7l2PpO1qDQ5h9E1d6ntoNHivKvIzIu
BsuKthO2paUlQBoQqrxMImxfhZi4dUo8xbHMrEl/SQ2giYw+9N5/m73CsBIyPqrq
DF9LzlHFAP+ToG1imUnYqHn+Z0BNb5FjcVoZpOJQMdntvm4QD/+zOVvOr2heYaaz
2oVTGWY5SpgK9qrIbARrLGOnihpzCSqJ1nM7D6i4H/0H6flYhnyJSBvzGET/czLH
HOgQ7/JrUm6gF7dIO3wgUDTYFWdG5zsaOmJtx9byHIK8fumKEGEqPDKpIgVH9Sv8
4BMcekxM/QhvPc54u8Tg/XraDlDC5IJvMxVFObhg2Yz0oogKhwp7s6N2ZpafVFNw
XAtbQHYEFUQQ1R444Or3Zpo1VFa0AkRDuHm5xZ2uHs6xZTH3JWiujQnuMHk16cmn
ODByiUtpr3Ft51L/dXp8zWujk+twG0C0reKEOfW3NXkiSQzVbAVbUsMjZhjzWIzf
aj89/dKbw04cNdkgWhm8YcT4D0FB63D/LHzMljHQ7hW9N5a3WiSACaCg+ohbSYnp
fg2bxonkknpnA0nOPkz0pDVa3jsN/7YrN4r3M0zypPdrds3XeHFHIqL1VHmbDLMp
UM3UI58FcJSDiy9kzF2rj/q8DeKFRL/seE1zjNrtspCTREXWJE100aEcw1tC7WiL
ebiZe/f8JV893q0GzzqwYuGs0rEKqQw960TP73g8I/FWiof3tAZr/e2mgxfORMYW
KTR4kXUUACnNZVtFhPXz6552yz0FO1sSU2AIpoZ1d/I9ZlFMzSJ528aXF/AtWhGX
ok04g5W9067BX9CLn+ovLh3NdMNzhMKYEFl2K66OOvRvodrQUtUUasJsKaJrnRmN
RL9947uA1F8JbOAcY+YtCN62veboI20lEvZnu//AkgdOGFVXUgGmTjRW2qy08czX
29BOj5GfBH5QUFmFmcVOhWLjm111fZSY0o+Srt+hF5DznQtzv6hniJcxTESREGE8
aEcYj4C0ST+pJrMd0ds2QIazWABTvrqcCPhsZiOipW+ptu/Bedkmir/GEqp0HeXS
y69EcCreyIdJIWCTMAOQ5xbJglXizQgT3SwRpDdoG5QDm5RnFWtn1Q1eBuO0BWFv
QRNAAp+LHjuZrowF2uPoEop/ydPfrM5ZNEM+0y5PyM0s03EmmZfbOZugYXjj1Xa0
1yuZqL1MgItJHyWr6ojtm7rimamQbcBgVzvY5COdVxV9chm+fA8xX+uaMOcMJcHN
+JSB3liFFNeMtalYBmAcuKSCIt8c/59jkNxCuXxtuu5gYFgLX1RGOoLcNKG6KkVW
zR5KXQQhqRo/L1z/6zGhuG3o/nsPl81LKh3lKevxDdLiZJ7iMwwoRf9bUnPX6OIY
Mm/9Y+t+oXSTZBEziO/xfwbDs2XUGZ/V+G8rwtEjBibZJrbEYrmxpfEiXEDdOY5s
uWCtyyCJu2UklVJpfqn0025W7AuC7JJpuWOIvuc/56QcZGofchgQsc9z3OsNKRZB
pc56eciH4QRESyWLjKGEUOBwhHTNoeSitmO4X1g6zH3qiRo4iAEK7GI3ADjgHBA0
SlZXSghwWsQlirdbFYIcOeL8v0xmgnYsqRO60d9PUTOs57bs/Zpvf6eKIrwoVGOF
oxR9WESQLF9UkWaBcYCVasBA32DXO0WULZylbXL0GTYl296sTzRh4ge2NNlSiYET
S367Lg9bvPTmCXjf+vMlX9UZxTDlR7VM1nFYrHR4si5tbWqgm0/XIgPxy7xaU+ik
jGcN1r+PwyDsyzhy2UXw1/aVBBEOhVEJBFAcwP2KW/WlsNCbT1RISgccWrKfjZjj
hKlkIEh2rXmuAhgOuJRRJ3q0LghpwY1160nGXoX1Kn1Lq9QFMRQndLOsye9cBpFA
EfU9xQymYx4y/04b/hMmGAlrPu/koZ06ImadHhK82+BHs4FnkU1R+TRT6k0e21cd
3w2DcL3PNkJHQcGu78JaLFkhCLlZvOeNlK0xwn3hRxqblrWfBZ7xGBOoocxIOr8B
RHXV47/oyeqKIEA+00PVxkvm+PcT+Q6iP+y/Rl5rvv+ZRwXnetZlML76Nwlw+E+A
AtsKSHZA9OJckeTErqVQF/XdAatzpJt5J/wTm5ffbmBMECAbeEfLFBW06UXiFOmv
WDLKU7Utfu8ovIQDVjq5cxonEtd3YrIW1pr0v4FXhNSakAi79JdWfaz0/LHRe9uB
1cfDDOYMWKlomASvBMnZEF9nFIMWT1TPRAoVsrLz7nAUBQ57DWBhXZsddLDMkwGa
zaWpNyZ0SYO/P83HrHCkNtn49jLEybUbFv7OunLf6vdeOYeytRw59Z3NBpA1O1XY
Afrmq6SSn03IiakMkfk2v94jfRENSo9A2+awK5jEmyBp0OohEaJpCxcw0ULtyfWH
yxIDlpj2NKA71zaHz2r9w5EgJIrS2ctJm6K68/f9a5AEQewC8N9Qgrf9ZZA7C6+h
WTY1B7Prz2FUzqggc7H4UpI0fP8QIQftTwfzOuJ/5ic1AvV0vPripJVjrNtkfNl2
k6MF7pg+mR+alMIl4blx/KQW1/i8/MsI32SmM9TchPFlHpQujK+35/8LKI3JlaLw
m3OKqdOwUWKmhpyQ9x9FWVko9rN2K4dCexECfM5wOOCUWAQtZuEd9xhFKeyQ83/n
Rub0ehTCrZZrcWyQzvHgzuyMEDfpIchuqoOEyZc5Ku6ZZha4WMYF8UBG36m5uZw4
1ltgW0mk5dGLMDcr+1AT+46ADdc8zJpTkonYG6KAAAoQ1V7fRMp/2Yl+nv2f/yZf
3D72Hj9wGXMVflWpKUmg71E1QHJSF5L8t/ahh35/yKJE6TQVKezX6SgFLcvXyH4f
eUggJDYRtHGkWcmDOdfTeSNitnh3HAJuDXt0xtkxrmMJQ2ux8A1kfP4MwrIg3XPH
oIfTAbl0fFf2x0Tk/nEd/Ys4n3aojUAlmsbDwo9kPi5DuTsLztRHv3uTLVzI52I3
dJ60C9uv7Bc+oZEepHQbkQe7t9+WWVDgvgZkkWqXvgOTsqSR1pD2kMIeIDs+ISxj
ERsjv1ZuAxh/WEl6zLZfm4cE18/3XiHomHMNB9f9LLfs1rZiKuZVQnSeRochz7iy
j+MrdNeZRe/Qr6H+7hLxLFbT0/OMsmcjoVyGCKanbZpexNcdIYHcOx+ZUEvgKjlD
+Sd5i/YO/+pBubfWBwUJ0DXtfp+gH84W8XB57rykRKk6AeVgXRJoqCX8yQoHBFih
VTQNopRfsMdCuj2kIg4HPNmLrBot9r9jeDBZnuHvneLQnk8TTPZ7sCskj8UYriWX
p2V1LaQ7PTNgeyiO5QMQejLbwHI2dOGWiJNVv8fNIQOLxqIe1R5/hsAhal2yC0An
BRfvmOQ4de+0FPrps2T2mr4HoqedrQl/cLXGGNE0ba/chO1Z8lZAJzitCrtqIiAh
w7UFsq8n7rNOnA54mpcv0wiDmKJnDjeZJr71bQXh0j+tJiLct5VlrBKCUOhGit1t
3EEsIy8gk2x8Vr1LhU6xZ8L4Kuv4iub2CD16XlRJQoaP+Qb5dkn7/VD4ZBZAEYGE
bv90W3mDTVmqes8AULalszLILQ0ylU8ZCLruU1P1dIvOKlBihdvKlNMTydRb2QPF
1N1u+aPhDcvf8TIK44Hj4fR20Bbba9I2OaEJxbbExRiRG6Phgb70C7SSGKmWMSOu
FEjmEl3aCe2G3VcmeQBjdQOpsgdB5QSI2Cv22trqtx3qoumcIjZg8Q3oICGVTxOR
uZy8sPdWcc/7AJLUuwls4umtFtufO8YXkmAVMH9kJ0J6I1DZ2VznEWkvGF05Hnj7
naKPm0w0h/LURU9qaN93gG/x17ZOVDUtMGCdDC/mirKUyEeoDhhj6a59EzPdiiLY
lR2+4Ha34gURJeDhonr3tROqZZmM6qZiVRgk+kirHBW+Bbnqmf97wux73Fyw6itj
mZDAdi62+1T6QVSGpWD+VPUThF5N+ZF0v4/bbYzoNIhV64p+G8mgGf75PcCZlsJX
c4iQ9MNPLzZZtjOtaF37XpKHR638EcXpD1dL53OgElOse+roKAZKNT0+lMWidASR
o97R2tfPenVPh7lefL0af9B5xAcVcAi2a8miGOKPBjEMUGNrmn9iyW4xtbag+5gH
KF9JnQ28MxLZnJni+u9FTKZTg2Nzl6aI89mM6znr1jCg8RMx7pjJO392h0nhDHid
es+hm3RsD4Ep+Jg0oTYGnp1AYTWA62KayXzvL2r6Dv3PrJWRy1eKpPZmXcg/2DJJ
XYQg8woiu58LhO34TS9z9TanAjqxiJL7rPHhatajitY8JDk3nRn/4SfIGA7ITOTc
HgJXZF48qkfeLwr95ths6EB14HSQQOKHzpJOo3we2XD6spqti7NJLyF/USeCqfOi
Iemikj6BdPkIcakawfNf6Jn/cBFgXnuxrfdGbme3fBWzGvIC2JbfOjfeTapLiAIW
ROCMx6Bt1s/oaz0tqKcaKOm3hY9iNLaihcfKXFobPzdx0s0189KqD1hgcmQ0K4BC
+3kxjtca2eGh2tDUbzuMdDa1kPOvpuCCUD/C9G2mfZGh1ETWSgwgDg5PBWgVypVD
v47sk6XrpQMhLCoj/PsJuM3ObZpk0PHFJOzZjYEQs0pS/a/jJxdKzgnsqqIGOQzo
BD5wysEVhIcN4iGL7n1WOceWWxvRJ78fMDxgv+uyrRMgupH/A3MuhK+0WBvbi/UB
k01sm/f4+NLjcXhQreR/9HxMaOfYc5TpbPq+uUX306K+BTSFkhYy+XDHuFbBX6bt
kGuLM1UzsCRs6KNJTDnkCWXzIPBPg8FMH0TyzzKQI/z97Mq3DfV90OJlj9Iv+4XI
uRaTawVXAE0YhZkdWOxNJtY/hMgRcAcoZ8gZBMrn7nhN6t/Q2+dV7vzBBV3p2TP6
Ec/jdYz96Qc2G/qZ7FyF/EOE8VWa34re+hl+2iXI+cBoM64Y9d1awsexUQ/+k2Z2
/Dq0rWThOeqrIV7L01e3xGJzXCCvGmFRz5OdwP8VydZ33TZnMBnweBWNTjwHvHCy
pZMME+7T7lD+D18/f1QvyD/HcRCFS2vJk0569D9x55U2oywYZ9NS46Sje7J8CY+h
rUkfFWs93tQyktef2bxAgI51mDoQVziImDjRysrzfcRJhSbSEQOVASs+rYCqknxI
iCSWRtuqW6jyu1IBKqFQJDbGra+3SDdltQGeu4R6YIMT6Ye3pYDqkkqnkQQC2I87
I9sHkeCVjGRY9VoWPw1e9RiO+D+o0hoc1KtQ+au0ryhJdpyV2dFLd8FytZLkZCMN
9uE7JEfWUSIzr30fjVT9YmybpxeXwJSyRpJux2a+90t4NXXTIvYQhTzKM60e7xa3
4Hs7eA84IyYmwpawzQtCMJRXe8nhFx/2NAo7maBpMf2M56klavVsxubpfBhZc34a
qKxsFyWaSzgQsDsi1dugylg29R9gXDVGEHS7yJMLaqdXATJNPXW0hZS6CVMCyxoZ
UXHWiGxvAokXvSfxiKkVKCHfJcSyZfeprbM9WxBWMMsV/zKeues8njBYG84H4wdx
fGwVCepAu8IvYLc4kVRuos6g0j+vDUaJ08ViXUOVS8StL3IA08KkpdijI9jOnAdz
1MycQ7KJ5ilrMQiMslDsdX6MUtkmz1E09EVrIKSlKuxjwhKrFxAS+5BQyngpayy2
p8UGDzfe/vx96dQ3KrFrhewP2mBkryohV0kdBBOyz2xmZ2jMLNjs1pLr6CJKcEkj
4XtdyOyO/kAax5BQG/32+HXjdT5Y9nU6efnzi+AQ9AHWDbATDVONnDpfv111qPaS
fX/pvmmc+Rqg3/df5ElfBBENh323ExXb/mlU4ZN394+rdYv1FWT/3ubDby8kbR10
XbyuVZEE/uXgqxfAaJ5pvop1y1WUWbKlpaX4hcX0hfRox92yAdfAJqPfHpTS86fA
MmK/sSjQUsgYACazzgHPNYP/IC5cjEYiFNAZBemUF9A/s3f0HQi1aIKuy/u1fSCX
bH2IS+q727FB514DfEt7C669Tow+HFVusz7yi+xUVoCcJ5WGUoBxCOAasnrLQ405
u2S8raZyrqHoenKU67h1IN539R/L8XwjPVZfT1Kdq9XU1XyxIAHgW1/ZpwlMwn9k
8G9QuCDTMh20YXEBiwPWUY3Vb8uf8X1EESHpqQzF+2Jpv86IvGMxl/QOCuHsSRxF
vJvS+MfRYMk7tDHYEMFEsnE9i9imA5YUbeTnh1EUmU6PngMqXSQC/mtteK9IWjye
eUN3BZIpDKnKLmFFiihzPjIiyka6Fa+Kuk9Dk5m4VhV0VxR0e1f1dR7nFZzyLvLV
ij3dEBYtmp95nJf9H6sGqSpXmx3DnbMJXuVQBGEk2K3ObddDSW8WAjAELnYQ/Yy8
3kb6KMjm2NKzYTAFyk923wRyiMYFxjLtZH9gq4Oct8YkIDizZPeGDR+VeEzX2IZA
sIK4MgyNZmZh4jAeymmnQQUYmfEdZRv9SJ+/XbcC0H9wnEAUkGJMTwp2/CGXHmlX
lh28Q6ZPzro4G5v9g8SjzSilwZqL9sSmmZ8nwd1x/edQjMRxGD0lNgQQophH6JQD
m0rHejqfIXsgT4WLwZfGO7KBczoT/8P9OdC31wGtvc3x1Z/OeqqgObUEd7e3S+V1
qDOmaoLGjosQCruP15DkdATA/2TZnDbr5lexmklV/9AXbPwWstQIfU07BpS85jCI
RmrhHShEPGSvJpOpLEAllv5r1r67tAv+bcVtJDI1D66hyYOAS3J7hLKqH7rcqUwm
pBXlFDMD/HOi2AEUVFpp4l9YdqTOn3AMMJvldbgqfwYtxgjEXS+PzZU2uMfKViUE
FjoQeUI1mE1K3F6gw6heCV7wg1M6dOaTxgifJt1U0SD1CHtzqiBhL1GT9PTlemez
F8Q+l5eeMEAzvcKieiZcBxnw9NIXXjl/pYNsxPnlejGPSVUru4wktPul5bQrBB4O
MqhqppqnSYitUt7OZc1s9N93L+Y02h1+zdVAEhJhCmgeI0mE+CzwGF4JsIzqhOja
WfqvGClPEtCO0rqnejMeNUSrgiWIK9ySsymLA/f5ec565/IF3qX85Rte2hB3lR5t
2bJ0/hJQklSY9EZnmpWfG3jDWsmyO21sMIXfVA/QNN6IWP+yRf82ZNr8Ucot7ApU
k4AzUWJaLXxzhOC21w85lweBoE+3fH5f77bNl5xN4jigigXuyY+KepajwXPpf0cM
jHN5YSSOEq7C3kD5WZ5n0DWOa2dOxbwzP7Bv1BJzkxpVm3VU3e0eUlTzvJ5Au79z
4OA0TmEkrOVX1wSyTL0WhoC90YHTNDYWWm2NOxqSlzN3n/lyxmDoRzuMHPFiXkT2
Q/rg38nAVPBUQ37A6H0/2OD34P7VwYmI4Af7SHzhhHr/pGfqC8qWvhScakHrvRgJ
NXWvA5zYv2FZ5scaPioWsQwgJmSdOM1DYleps/vi7EPc35YZwxYQOvcqCtgyBmra
Lc5E/EbyX1x1DSla8Fbum0AmoOcXHDPdgRFG9iQVK475NUSeSVMBXebbVwIEcXuj
0RGNAzLGqqbfurwewStBVn/ER71M5pud1JZtN6AH2oy82SAj95gLGEYfEQHLWkQp
+OSMwvIRoKnZHVTt2YFaa7nLWcdqXMBzvu7NERHXmsMQQkoZRK9s+/g1DdwfAsdV
fDWlf+fTuEmNc6J1Fo20D2wENaVDzFZ2gj3wAzSd+oWrdsCDGNFANluLyGMjlBVf
aGK6LMj0EAy240A5U+gYmamgccKkvPotf3tDAoAEOBJx2wcu+54GU/0N+4PMpewK
Ozr/XlgKjhVqp8wJFChYFEfBMzzcN6B7meo3kYBirx2P3Rc2lxB+ELaAY0XM8L41
u89F7iQ/AdB0EYKeQzWUwwx0fj+fP6Nz0czxTi64BqOlQayQlaMNYtHvzJHoPF69
p8AqFauJftnVul7qRGsuet3DY1A6kuji+K5E6is3LS9ks+xw14YPq4DXE8asxew7
krMzIL4wGB7g0j5r3CxKlF3i5FEQtWuda0kGxCvizZW+HfPhACBGW1eEV8WuwzB/
xuv19lohxrxu/ZyeibEenHjkUnxzZAwWvQEZ32x42Uz/3ZXJlAdEXW/V4+3UOUZ8
1pdFTwOioLq4/LzQvDZsGcSvFTZ2lBYs4P3adC9SHi8cU2MgNtsa7xH23IYQKgpM
QYsJ2l+7c69q3KFaR7vqGH6lxULUQZwNH4OeREVIIx9PBxTcnGNDpKFJSA9/NJhx
uI6/ryDH5fo0sJHeUvwkan49YkqzRgxqzdJEQhluFtWn3FyayC49oM9qbXLlF8zW
2XPbU92A3fu54b5F5j8oYwQcIQf4wIJeiBZneJhSsWF0SUhrmPWI9SI0668VMon2
Gug6NUbsUX+Xps15aYl2bthgvDLH8hnylam5BipvafF7g9IPeFS1oyEOuPg7O8XS
p58XQpKqtm3iRgSwBI3GhMB7pdbnmWL4vlFphbvjwZDNIzTSB0e1IBylJw7odgYs
bSIgYJxxQZ4pcoJkZG/3P/05+14TxoJObHc8RSkZH7oOWwzWWSlRNPLPUnvrEicL
5UPYUfBmAtFos+MJMlMHD83EqD8Hd7rJBhqI8oRFHU0pgvTQ1JP2YzMVW4TRR79h
tyasF1/ygj6+nK3kLJzHRrISqhp+cXnKP9y+3nyDq5hS93KlyV2yzBIJgr/Tr9Q8
E4t9JkPJ7O8YavKNgP3rsPr8XrKx4sMi1DoxZMYgfSoahcPQoHqrXbMBUNkAGk9P
/89RlLtzxkVsHgJOS64rn6xU0jvOi7E6qql+z/itWu3XkBPcgvshuah/0KPXwaWq
q3+wOMCQfeGso8tuPx6QwtKwzsIRFPaLhxw5x3zNZ2uQEBev2nThehKP9IEkLdJT
psWXerpiSNI/QKzIPRf6+j39KyKN4nhdjU9oIwsVzG8RG6EdMInicTLHJoOWIMjR
VORDk05TSGZRgj4xwc5qxtaW7nj3BoKWSRZTvc6fWWDUdpU6fGa6BIcCHqBxPKAf
VU5idmnoIzVtD9Y3snkirsHum79nh+PqTI6lmcgcErjtMBrYmJq0PS1UvdnUCuPQ
M64WrT/+No36E26XmmbNMDJK8K3Lr3YggoyW4VXgI5y7ZfpS8hSt2mghx1sabLX+
e4VL4TDBL3VWxEzHxWSs7J9/jLNJ5kvoJRNwyflNRiZRGZ04VMwlSVyP+QwrgnML
GY6QXXDq6FdPLHTL8/AL36WY0asZcawqbnTAyk/QfSil8fLE2xz9NLWsYzULMD9v
cY7OGVjJJEHL14M781r9XERodze9IXBVdsd7ijOAqAD5XJUG5HYNR2bNiEi5CI5y
VOIRW6LZUC06YlD3so2wn/ClT81BbeEMKKvHQ/pV/nn3xaYkJxKR1RPiy8to9qT2
QK0yevjicgyGnMUW5zN1Fk9T2i3CMUBLt+1KcmKov76zPPBPxmpILmKB0gM7KLU5
xur7JtpgfbQ2DhmfgEE57X09OD9+AiDyS98q9XciGKIVDgrpBOgEhaQJZQV+GLMc
VwgYLYeaXaJV1NulBQ0WWBjC4rgHgjMF5FGZjA1cTabdkMCIW/dTUYt32IJlyrh2
a5rqJvmrl+GsU2j2HXcszyXuw5AFurgPiRiclNB4a30r8PUrWWIaxSJWiJ4608r8
6QdXhGcvG0SSrDjHBTirRsEJ1slpWpH9xejaGbRUz9t7CuCkdYdnSDRvfQjxUPvL
mYyMdlIFDFiJd9AqQOymkyaSMc4ffoFUUjYNVhfszlg0aLAPxB1v2jnYLUu3ya5h
Bd9+3KhcdBFiEwpciMBXpfi3Oe8kGtBCdJ8HhOfbq8kkeF28UYeVx1KlDEUdJiXn
OJ6TbIBrUIZMeS3Ky/9LGE+q1g9OQB+T/r1H6ZZUyJWuhk7rdqfcvn0YH+aC6m0+
GGdWP0d0RPNUeL21gD6DmLvW6lOOMIJE5KV0bay2yYvWL1upqu0lKAmz9ddKiwCx
15TWKVjPr71ch/9EuZvX98QpfDuO82oSlCJPyC0jBJyIFdEXaY7BRoDNaIFUlhyM
wCWKGMT3kvrOTv6nGyRIKfUzyqUImHgqsm01fFZgKZp5ZqgiYP7Iz98AGSkvcBUU
FLhChO23LHTI1xpgNPhgF6deASPspmjCOGZdPVwgu1TRtVaSnMMqt/TTJMKTSQF8
OR7iUVira8I0GLhMbIFkwCyCTNkXZjOsSkdB1VSy/7cPS7c7Hr3mYmRk1m7HXoNc
RhTAj9fbMApu75AeUJS+JxPkIuvte3HK2ICzJsXoGGQWIWsLmGgF82EELt/TYnXG
NPKvovAPchjkfdRZ2PGNs2bMpdkTkhOG5X7UsV87caJMn70eM1kUh5ad8eJnHu5d
aNafJ378Cdy6AjOab7MZQoCb0ZDzHFiCNET1T+FxABX0RLHwtntq9s8nlTwBkGSu
FZnb7aW4qOR/z5zuaewi2i7mtQDC3X+Gqk0/1XFqHmPsPWXlueAlTv8uer+jSbeU
Wst/Osno14g20IyE7FcWN0MAFB6iKOmerb6a0VIM+2tegNT5guA8CskyrfQojdxI
pVH2eZzTt7nsypqsCXdRb57xdWHMzVl0YP8+dmYpUoUgHmd4zyl35Cm3Qs9iuQqj
COi/Q0LFSsWUl3r8+FEgainwG6AQoppXcHtdhd32sKFnSe+TelubwYRUZvUd1Mcg
oEyxCGwcDD32CWw09xxuRcnY0tx1D+oxD8Q86ebabk7Ko1m7mCl6H3sH9v2R/n0d
E7JSEHJNEmgrM0MObXGvKIw+8O3JLvGUNF1nRZlx0hWf8yo08Rw9Kclnjl61gVCw
y22vqpCVUcPDYmNElRDOlNjn44Wy/voqqeOyRLpolEuunfOBaehdY11RScFCTrKO
WBFU2fPwnTZVfkA4PRwwAXGSDA4VPBKa3Kgb9nhCEi50QFTk7WWZX6Mc3DNAPM3/
9NDDWvE5U8VrBrC71voL2znXGWRVYZsar5YzdBVuN0YlOtgNffvxpQBMCKrmKEJU
Rh0pqp6+MXTtkoFWIUhPdgSJ3/0Inyit6GCqGVU8Hwr0bfqUUq3+Jo3zmhgLcAgs
CqjhB9UllPTpAfd1IERc6xKaTmQq7HMyHwf4VTQHzhs6k7ZjViBdrYZWbZynuRB7
twrL5Mxzxek9+Lo1/sF/VYdHuldcimuYzkDdo6fAEPC90SKBCd4FQxSYnmvW34gd
ZV03/EwFA6KzwBNQQsLjTi/hRg0hFtmAZkAUxnXsgagixj+FlFHxjsFEIc67X2KM
gS0GlCUMDB9dyquJmF15uoNcRqqjlExRzHRr9INVfpB3Lm2WBtVw/O0zsErbBgCJ
4hsAZw0zTOu/6JvxiRjQ6n9tVJ7GEfnWP1C0KvpT+NiwtWdIaVIQddrvF4M9Y9nJ
bDWvXG20hq+8o9KuawAL/YtiojdsVMtoES3d3nMYSY9x8eQNg5xZBrAZwNRGrO4X
MIAOxhnVwFydoNncgOBoydM1mh0bRDIXwiPbT6QX8qimph7XLbQ3nxlmjzbY86Lr
GTPAtr4zyWE96cwOB4xNuJ6YBaEvY9q+vo8RKg/QlL5CVPXn3+8yIBSG+kpWgpWQ
g1caG5mjQL+kKX3b5Utu6hARKpR+9gaAlKlU2zGsqG/Hy8F3gMonbJGLVZek7x6e
R0k0GPbJBdrTfEy5Fap6zZ8oUVgx/fHIFH6TinW95R+PH2vFY/ZBrUsdrP9evQG0
WtwnLo0cm+1mGpym2B3R5XHVq/y9NOM4k0I4UgAhRpMeMUG7UK3Lg4fgX7O/0NmN
PP17932ET3QNCNGj8nC3SBGjxEIEQlOJeFpIxR9U23EGHJGXl9A9aSpHT38mFfHp
T7W4YZOxIehsTaoddlSVYUVOGlY4OOSzPeCARf7gWSShsJ/O23sBq4F1C5ckphNK
B6SUkiqUhl447HGsGnndaM0331ZdRXzyjSi1DtavnblGtLMBEpDUpiIMDZA+gc/Z
AkOkKSVa+oI3inCizBUiTzIBkRDCOMV4Wy2/qF1wxMAQNoltlS+M5/Bu/Uw/GN3d
7tStLFoKxJ3fTBXaTyQ3ocpmXVZ2pOueIq5zSHyJA789sN7OF+6lvMelTdGgqVnf
D8LQVv/pRVKy0URNPSKIzZTV7yR79wj4vUudmlx3x4Hd+uDb8414JG3BwY1P2n5c
F2L1sVpkuLx525uNGOjPTf9UJUgBn+sp5kpifXn7VIsu+UKySFv4qnuVKQ3SaQJp
wiRPQfs4Nayn4yjiBz745ZwPoZOt4CeG1u5Zg4Lo8ssmNlIuM5Gup/9ppOMMAqga
J6jq89ZykpBxMR6PbwzFhzAsaVyP24rFtHITIukauCDh9xfix3XeRKhfsoWtVygG
FenFNW9vUDM2aKKFK3osZtKhanQi/ocdV2POCB4VQwEOW2YzdnT16+gCkCyNo1OX
hpch8uGFFT8lEWFAQXPyoww9xVXS9C6n/QZ+kMFwFvV8WClAN8xgOPHxPbOPQZj6
PTgDBTUtiD+LuIlqHNekQyTTBsZqtJOr5YgxyWxpmAb4jCja3PpE88iRP9PwDw6z
EG1xleudb3sMrtk+Jw/ZutpJ9ldBOaJbe9qnmrKfoQ+0joDmOG8U4otHJtQN3pLv
W6IMZkY/gsDBBifeQ4SHP8ICkdxDyGQuwMb7XoU8v4fPvErkOtVtnvEpkC5UDaOg
bX7cR6HMJxdTpsQoIkl4K9HNvW9TbjHuNGdIjQtlnn5gtRK3t/i9QjT4oVx8ljai
1ChP/o1HdeVUG7nvymHzWdVJH27dvKEZlZN5o+waxzmwzyJEUWw8NGGbOnIN+PbJ
cCaWOgbLyaIvJrJKHhHtWgP9n0xUU3nr7CourZBuMeH8NSdh2EFz4t8XW1HclzWW
yPMw9ehH+BDg9/gMFLLyfH+o6aBppq2uQwO3t6HXeSsDDCgfX+Tz7RDZrFmhw97f
0/+z5+Mq6be8jkjkTbbnnqQRt15NyBn+t5AaZBbENMaociht1IJyPDrTGRTSAJ/3
q5NHPcyMvz3z7zLL8/Vh90DOBzn/+2xN4+kfiulqcXtMFicmR/f7UbinPBgnslR7
PZdJ0c1GU3yDftqoc5Yz5EDu0QooByH8hOHDW9NWetKODKhm3sxryjktYcwkrHg4
v46n8mz4oz2J0G6oMVdrppND01frE5UITT3ECrHxCEP8KGdQ7uLitq858LFTQNaJ
Sgaup+nsok+9Yvc7KBj1TtrYsk7p3Ll5ZHWEBu61AmqcXQGcm3O/pne0frb7Wh9n
z2lpHXOcUqqcbvLpSuHt23f8E+3PaH8RbqoYPS+WIhpoNQ8b+ID+EVW+EHPaeG9m
qThvhTsUuc+GXEFWfJaOK4IVoUAgiwPENk7sK/TONL1j+nhOwZikYeoPjB7DF2Dl
yb7/PB9YkHa7/oYVReqxzQWHIY+EdS4xT/pBHeg8K6CnbVHbNqCf0lYZx4C8K7y0
sFW/9+FWh4W03UNEcPVCWapMdy6Ji82SQoJPuedHZOgLJQBMoPNCXqCHMXGGNfOM
Jm02LTe6+woeROjV5ukeVLuQJ6hjrTz2TagT0xoJ1sJyunHz/0rr4JWJYJAyqxoE
5A98D1EyneurPmAINAD9ZPRvznWOgR898BIilKxcPSUzQ3Yj35sznzBeGqMwJ8D9
FjpJ6I3keDeaypkn1nz4vJSxAWcQzimxflyJcJWHHy2zPkfUsc5ZHlKkOdZOXNql
jx8Unwgr9NjB2EAOWeibYkEKsd8C0pWjDRINlOFda6JJtaI8QpcWZF1UzsPHrGPU
OB7uHsxdrzJ7TJaesmfOOxYh8bL9G5gfU6QPqe6EFvpE1fG2rhldnkX1qYqXSUwg
XTfdOL8c26/FPVaM8cnlHvA5iDuCTqGwFuozN3fNtOAR0s88uFCxKwculie1evtI
rNHdblWMWkzlk1El+xY/i2BXB4Oo2u8KOv+WWJ9u3ynMwL4YWYsq4PcKTRrqDZbU
+TLjCTL622fWAB7V5Vqk9Dp5PPd7rr81FgQI/y2jzquhAVCx1gI1s7hOzC1hLDIX
MbNYowDnUyJLnqWzQXDWz687FJZy9WDdFQu7wBMPt7Z8g10HenmszWxfKLEAxK1u
KKkSX06Lv4QwvXKccZpf46gHutJ53t22Jo6Nen96wrOvUbl9F9mVjdA1U8yAIh1y
EWrPSd7iUQDZ23ztvJ6agOTknPBOFoyNXwTcJ/If7ScaizY1C0luAo6uhicKZ+2F
D2dvnTzcNCVr392IAGCSpSVYJwYQT/EI8gnDyVJZzTi3+oIqeJrfB0A3pX3HMEZT
OPH3RpK1xFmQIRjJJbgg2GiCsyXHiDDc4DIw/gFJho1w5HGgnTxP3Il4//EN5ENY
Z5vX5vnezVYOTUO+2S8h2Bv+nBQ04NmCZMtpR+fdXemvhXqTnix44obzklTiD4+j
USYZcMNDWrBC4cA8EXVRyr/w8as1p/yDci15mZz40L15E94sVuIGQVWOo2uNljCy
clYCkWTjFEPbCtbhuDYp7xBSC3RPLG7RoH0UkqSxqsdZIIr8k0zeBGK1qo5cRrTS
xip37ngD40ELdlpJdbECDBkwMIVF5k3YlX9aq2l5QqC8HwuBFiiKLhU6cdPddnwo
QYK4TZElN5WRbTxGHtvvKEYpr9uNrTCET5afwGMmQlg5s17ckMyTbagVyx6mLr+w
21erKFO4aqeWayXmBOeoV0ZXyq/+ZHhaQJSPUc+0M+7fyM152Gj+AjJxSRrJnCOz
fUJQ+gsC3OfmDXICXxgmpViIZIVVVPyqG8ZP1AhcQ6JaWRpbAV6xztT5+CX85t+B
Yu2mPfNKPWkSZboxAweHrAcxs0mv9sO9ZwIXCRt27Fsfszs6UtIaE376V/BTWoDz
sQadID2RG+f4yqyXTa52tiBd/mt6f7oUCXr1M/3v95rlYmRSNV2Dy7+BwIUkhr5R
IMK6cQLdYRnAr/BOmkWEJqfwfxSfctNKKQiDLWQxjWwgCSYGZWpf7Q3PSWyx/k3Z
+ycz1B6p7hJ7o8f2XCGQ9DQ0QjUK1qR8az90z9dZaXd8Gmw+B4UrmshrlFE5ytK8
d9Xim1M8GRkVnV42p1Pu8HUS9TLxVDY7yZYYV84s0k5463wu5cb3OZYwzly4oRFR
D1gXQuEibXhC/YJ0ulM6lqIxdmmhODNob0ZaR2+k5ZSbWsxgzVvNp5bCR577ET1u
ydG8ZyROWJlkt0CGrW3JfMyjYHbd9zfKhUWQ3wPz7UUHz+U1uP4Vm+sHLvlD7xPY
BQEKYv2ziHY7rDYIYzuHr9LDTlU1UoXPwjHa0Uw/ZrjxFK5nTfK/wQ2jQlK7e+q4
DM/hWJl7gRoVThZiGfnXZEMI7kkWtvLn18RUMaPRczf5UdPwdaaZxbENs45v0ktv
MPnNYToVILDMfmKQ2VP0D5p89mdyMBPJ1zp9Z/RbqJcgPqysp+avuetERV3ImPXm
E1bRoP5yEmiBVjZ9nOc1e/NRj3Znc5Fo0SFh3nvewfitF3e/V0T00dLbKm5dB7qm
NudnTaPwiN7VcOo+r1XwONQ7cyLF3D05Ndp4mVhZTDC2KycCq4g3Szr8Em7Ax0pl
q/wkh+DCjog4f67oPxtm0uFspIe3dpDEybgOl1wB+m0v4eMnC1+qiMPYgHSWl3pi
LS0xPW07dWE2mDkCT6kuBkVz7G9IQrkjrhr8qoRUPxWDtZeveeLl6MNEXbO5FV5C
H5EkBbo1Cu2EZsX9z1y+VUnTa1lJLW+3IXBOv3NQuprshNpWhQEKAehvOWXB6Vb/
OeTDnvvtFXOnqwV3/pYJNCFGWFcvCYRuTo7SPPu1V1uxMHbG+3jXeAr5cIkFVk9B
TwutTsXyB/aHwWib5iTnak116EUP6b6oL9dbvTE4mmVVTAaPYS6vnkjv5vMQMSKU
26ejvACFFx7+Jo/KyFjqLP7Qx/Az3i+SvCmmfV6MmqKM56FpJ8RbMyyrKLBszf4t
CLbzc4eRhnzH+xyPXXc4of9BEMOk6Y/v9zF+fiiHwcNYsxNPWosZzn70aHn6WaQe
KnUKEdzwT4Zvcrx3TvBISUp8TRFH4Lo7zcZ+IIkWBaVn6Jh9y56n5ppYa+2f5SJu
JEC3ElBFQeyJ3fBKzCjFD1lv9uJ+yN4SAGPEEc1S0IJ2GyL7qoUvn4i75D9AexMT
ZEup/Pc3YkK6L9RA/x0+f7UqRydH32T9NRvz6k4Gi2VjVGpNAnnV3hEUMDSUVUYF
vo16zQqt44OjFPJwyVWZlTL+mb+xJ0zpRw8fDRig04dqI3cEfbyfvdA00+RD00vY
EZ6B3xDSD6OaJbmcV3mGWRY4AU7IJxwQUF3T9hqTXIjD0b+DKzw8QYPQnjjh3Xv9
S8JPriQtOQJvmPQNpD7c8PO5U4MYvjVNjpzWEIYRqgO+1HE11MwE06yBaTIig4qL
n9aIPa4gApKmBOQ4KI03nEXwVD3HOh2ZdP+xBZPJG7kWI1PlMD3AoynthZHZzZGw
V6dtPGCML3J0GANCRd/UV+dCJ+AgREgcT6UjgX1rKScGvjUDDeePEwFkKnRCv0mM
+lnETTqe1jb5s6vyRmNaqIhIQ6ghHHRqZ2a/7HsnmjsKYdCShIUeZ2QpTbXS9y1w
NQ5Sna5xLOqRrJAbXKKn/OgLeWth7CptsoCHOd0J5x+Rz3VxWy+G66tb2ZX29AB3
JsSs+RUXYPk6uoq4DxOFv/3UCjYci2fFURjs/ukCFQDm/OnvpJST0OorZjbc1nrq
JOmWCn1Kiysls4l56Jdk3YOv04WjpZ4lmOHknM8KA8jzpeZzr8zu/j3kFvGvcaSt
ZeYEequFdaFel/B83tyQD1VBwseCfvEZW3OFDGcDKBjkGvLANsyslJBMTFWk44mf
xmat83UW4djWeOSytrXUHtJfcNHXwegDl+tEM2mdLrQErRI5X2fV/ndXNtH0rBO/
pHJ/zTnpUupSnK4Nh1vsoEZvTo9zXWF0TO+g6311byFx03N4g0Lp+QZ40YRRR5CJ
prUi26J5F9A4gWUucKIeOnwECl9ao7SkSrfHQxpyxDKZ2+/IB8Z03lSY901Fn5PL
0fb69n0DTLB3ASYV6YvOyCt3xNriBfrZKNNc/ysiouKZC2R7DmG3ceckIjbfrZYV
qobIp9tFYlVxW3s9q/Vx0SP/9VjBzzX3KlskpwzXkEc8q+3B1dCSF+kJiIdyL5us
xCOOq9UYn5YcDD2be3qg0R6ZcWXLNUWROxBve8v9VfyRVm6SQNTLgh2/HgYyXMAo
pRGFTrfXbF/pxQGZ1kReQPLcuHVYHXbQ6KLJDz0i2NCKlcjXvi79EOAs7ddCvcdY
Bey+Lo9xSFPAQ9Z6jw3O8WU/0V58P31pbVQLvhDVPu7yYPSpxaq3aWXf/qKF7T9M
eXG6Pe+vBB6sPwuhKcsJCkoAqcfbYaeFglbiGK3SgBueHOhL6hCmdTh6t4Pr0WWc
um1pcIfKmTBAXvBVFB+2Z1SnhjHLO8/7bW5isidhKONni4HuRPqDSMfpjzyJhu9M
KNH6VMSp9m7ROSZ+T8zStCFUZ3vqz4U5NB1YWh15EhIegarakxHbY1nn7WUgbhK6
K28bH1pvLd6pcUdV+PuyIEElsIKY5qcy36KhEtw2cOQrDL9bseW4eHj4rq3ZrCdS
pJFfzhnRPg4Llh0oZjyFqQ2AP+rko6T3xUiB/jTXfZNUwYTOAHEZcnjWB/g5qFT1
Xh1mcsA7/wbuqYtuPppBeaaYNHuGUOv+8t4e2rzQdZ6e+sHnr3WWFBxehGdXApdv
ORTemGyp/XQL3RWw7wrNkVopl6933kcGG7tTRoU8a17/XEQefzwK57YeGPlUDtGa
KkOTpVS8j1adApSS7ssfKZkXcXrXKgrVcfjRzdCcVggr0GRaRPeubnt3vek2X9i7
VpTwxoDqaU4MDwiiBYTLJAwd6ipDBH+17EafnpPNLBQ01Ix+H6uva53cMRPKC9nZ
8fcdLa05RtEY03xfOBE8YwuYZiujE2GKcKs5m+jlmi2dZR3wJfDiLQ6gMGTU2AZT
gbkuZxBUxyB9G/lHoiNHXbqYlckxcztCrvLQ+8ZaZiiqV3K1Vf1enLftLM3jMZwo
b6uv/CjmpZiNvtjZLc7d6TZbYVuYno4rcax3Dtd+bQp8KsJe6mvwwqoBtzhjlt5X
3R5Cr65h1Fwnk0nA9lKj6D/YDnZoxvZjgkTWf4NNyLOoHkUw3Sul6EoQrg1b7iIa
kein7LIQNqFnGG+ONFAPiySbS/WIvaT2ScnWNnv4cM4XSal8KY0wrnbpPxxA7FCJ
u2Iy08rTnLGhG6Q9sahM+JWvtpxiYymradw2scHkygRrZwM8G/48Ng1FxfAs0ej7
DfqizZ+WxqkzkvJKklSCn9x7CIi9GdsM2nPu6AiqNu5Cf376BGcORdHMSiRZewfl
WPvUQF8z74+KhuGcgpw9oESvxTSJxjNJDd1+f9PHV3qrPoUp2cSI9MnyIdMAmsSq
YGhpoAtAAGlMsrwZRnYwc+dcucmfoyGNlfAhqqHGvmln6PPL62CC80tM+sjSz3+8
0BsOQQbQ9grPVB211hUF8S/GoD6QTeX9VbZAfd4+mlj29U0LzALXX2wFrIy5CeN3
6r9SmkY4wip0zIxhvcZ+3RqVgIxKOuLvRSh3DFyjjLTZtC70luQszD68Nha3zn+7
u6Fvn+WQyfITPVJy5ZXPGEjlLUscq5isLMbYqEZAvg6gxYyFRA3Q1eu1bSOIQRZn
TLPMUxWM18vqv40PYdqUwvduoax659AygiAZwlpMmFji2Or23KVR0qHDvVXOduZ4
FLZ56LHq8Gzgcbe9FEKp6Orp37VkyZSS5w+sQklcTAfaLurNde84H3HdQpivUnP+
GVZ79ZNejiA11UxGJjf/RewvlY81x9XDr/AhM/xfXCIwcZPeNII0lGKWV5BZYZw9
CGgCIfm7FzzjadQ3zUj7rP6BCsLlMeneOfomU0nm44nq+NqwTSrO2t3iuRoJvLeY
ucfA72OSaQY8XI5dhiXBDtqLaT6MFmq5oD0BZ2qiu36XNLxPZjjiqxgL9u0WsohX
PAmR4sYD5hOlALBUmTvLLtUonG0UesR0wUfqllMBGuPNR7oslmH6VP1T4r0p4UW1
2MkRk8DkAZjh0cCjk/5djEmvyX0TtHRVEFt/7Y8jzc/0ZytXCjN7RgGnZ1Hm8U44
LmRAPdBPFD9qE7jf8vl16IacbLwle51QAm88Zqc9zEJKAeVLb9q9tmIZb8OTArf6
ChqTCRiiy+72YxIS5c2qqXhbQiJD1v/XqNyTL+xT4kuawVWpveBeV395dywJxe4U
oroBpnat5zcMWO1E1F3LaMUnbHgbI64HG1FXJTaLKbsOmXDhF8p5I4m26YHazPD/
hltP002+R5F6vX1wrWGrfr5pEtuaoVi6U+BmYhxDGmrmKi2JRTLCCs76Cv3+fPYP
ZEaxkas3bOtnGd0t3HV5PQRrzSnvqKDXl1xX5i1rpHAbJMPc2nL/PWndvZHQWtfu
my5vQdgkhX8uGzHAlO+R0JRDRonxqGP4/IGDy+/sj8XCa5f+tnZHSF18VLyhwua9
ldpR0h91Muev8TPJU4Ak38Dv2lnoG++0C1vtGw84nG4X5WZ7HWLoRYtFAtnhoL9l
Iin346Q9m3pdAuxR/eHMwkEzUZS1n0Y1XxEP0gMNLjM7IkSlO54tcEN/E+bAsu7u
EXXWcNbwa4jYBEvlXSbsPEwHPOs+5QBpIoL4Sb4xgL3HZ/t0bcat2Lqan/LgUOee
DA7NrnJ+Uzq02QjZk7c/0FafG7+ptolYFI3rBMZvySUhTQq6bWOzDJrMFf1hxZAK
vXzxFjpgX/VVFoOIpjpw3Kxl5sr2HVUaio47JrWpRkMhpOl7RjoT0Nyi9ARjZHX2
u+0O3z08XijVk5KHvf36fuynxCKPg3KueFGpMe8CbjbfEvcn1+RhXHnLitUfS5xq
on55x5DzPpT2WWVTebZTVNZ5NjWum1XCV2rkg+V+44zelq1MIgQxaD1kdGDfs04/
9FjgSX/+2Gd2j12tsD5C32qy2RZJb2IFyKxlDMccHj1EQ9mW/8emigFihZGwD2Nt
QS1pbnMii8YBnPkIyOXYAAnODsHIRpCeH8By7sJ4k9TA5UnuricEU/tJfb4M9A3K
gI5DoDXnXl5QMAZp4s+b0UDHkrJfbNQI9oipwFUlM4iOjqTkm+WhUo6tAT+GqeT4
yID45+pEdCtnEx5bIlM3cm+57b0EZBdm65Kj0tv/nzIgXVdXdy/qdMvbV44oBU70
BobStiSeFYyPT70yf1eGFVQD21J7kbddnKYpCQXl9pXT8Sz78V7Yawq9OL9LJTHF
fBDAP7dQGYUU33FxevrhOnWYWFg8jy8roxSD65IHB72m8oZjlR/YznHD0TvArrt3
LFHAsCFu9wWVUZTiefjQRKbwNobfH9n/kA4pO40lfPF06dp8ukwQjdB12vGEHAzZ
OlUzZ9OsRW3xbI4jHPAvCtNbzhqn1a8eexBnp0BJBFs7tWMIC/NVHit4nzItEIAH
hEMkQr4E6YFFeeQWYIAbB/3n5vist+lrNFE5ddgL28VZwV3i1Lgde54ypAiMHER+
MPTSuZ20zh2mrgJbZvhR8EPsHdo73M1p1GoF7zw39tWcolQKNZboLF5yM7Lvz5Oe
b14jxIWNYGsz6s8HZqpe75nmYnMQx0/10KPxIz2PdAo2bBomeH/xxFMQzKz6zxVI
xtfa5y7UmDNmVOu2po8i5MeskU5k0hOI7wQYGoprf6U5F2HXBN2MwqldVRKkuQ2h
wYL8UUG3FzEnvgrK9MHaNufN5ovkIYAo32/Zh1tXsED8v585DLLhx6SNo+G5L4hR
KLISCaA0X8hGf+BiEHtzm9BLNUyHTeKyh59uNHFlnUQPYsdBJhZ1XmfDzsvHCUx6
DL6hl24zHJ+i6H8Mj9sjWalphsinKSPxYu7caOBrDQsa6gsEb52j7YOk5FoIDUh7
UsfK3eW000IionNSmiux+xBVdnWcao++poOSQwMmBA5XxMAKaG0pdyphpB6a0l+m
P50roszqa6pXGFoHJqaYUnmfIeMdVXhhY7nm4taOKixqk/zq4ol538b77rt+VVT8
Tjc6RmhrVBS5oJ/XerMHxZcHsg651AEwMq7KhgyqXDZsQ+4wLgtvs/O++JTw+wP7
FHE8mCFzMuR4caiz1O8+I5mNsXG9LMASt/xSFTkAAixSzc9cKMtBy/jgwM3OLrkW
nGGdExL3eOYynzDTPGJfI42stibjxuLRmyemPoJbDxjv+aJiqNIpCYuac5rLuj6n
CVdppMAjd526ajkNdQQGG559u0iquZz9916YgqJxj5y1/VnZ6BEo5TYDb0mxg4ce
cqY/bqD7SeuxK5VpnqjXd1Op7qgkQYujlVZpmj+ku0jSCATJ5sDk9u4iKHvNjMWm
X2JuGBMt9nkxLuod87zV1B8h+Tys/nro2AGtVnUA3p+Wz+QwLRotkaT/eBZ3wzTx
Szv/YLG9wM5XpMBdb51jw2nZdqOybCyafhV5KJi7tz0fMZ8+HpWtnAsjU1+Rkg1i
2kFLvWIhU5CX5y8qWSanGzWDvNxcAvf5cWP680KrRakaWh7dKMajAEZQd4lkKvcX
qoOZ20YedyyDG8Jqbha83caeYW2rkYhx90dXyCC/pwQUsNhxMLQYskWd8AUSFzE1
YBMwgh6q3jrHrZEwVQC6o+u0YC8poveJvj3maNGrGOLEElgm82HsDff9KVyps8fq
oHA3enEKwn3H+XyoROymxN9Qnt+uDfgiIzNBQ8Ff2XMMns+Jr6lBGO27DTojDF+Q
yYIkS5I0gmm1x6p7yFBSGhW0V4AMsj+mZK1NF6PJjSuIyR99AZARng3+u1ypna5+
LXk3nzg26eqRVrf9blg9BSEf7nuKlcQYPRPgP5zQFu0F9MYNg58NnhIJlKF7ewLa
f8kU2rBVor0vYBkr/j65LdZWYNOezfst08U1ow1P/d/3W0jT8z4YaDxSB0Mqyq4T
nrcsMwIWuHWAwOPQ8HyGdX8jglYFXj3q09jV69zJ+jFf6gxbzFUW8PhgqWh19I4m
8h4/TttfHuuuvfoqy8aa2WNPq6knQybg/VCsPa27jHzyYS3a2yCZSCXHBMlQ3kFn
b+JaOxZiT0LH+e6UdhMOe/QBmVc5D/MNjOXRX6gNd8malTM6WjhQErBAEtMCWiMq
CkU5oNus4N0xTVFsj+RZNx4M/nzFytSnI0gqwHLmjm1NSMSztuzsz3oBOrrUl53S
Ee26Cr/IW6tvGLDqHDCcl+zjU/BeebITwm7PRhhOSVnc/Rpgs4bE6cflD+7gqhQT
ihyioLBRkWTdxQPv8IlG5gnZ5zLFNM/CeIpDR0uu04cGJ7ldps3avTsuPF/uC4ui
TBLl3n7NRC8DKhsO+S8xFsrAyzPUQilTE8k+xPwCL2MSEfIaaVUAMfJ4TZHK+7NW
kZyDaubS7ZGA570ovWbZTkG/M946qUVMZHVsNtZUT4LAKVKIsDC1JMGulGlhFhhy
sFKoe6pGJecZIQX0x6Zudwkp9sbIK6M9MNclBdYlNonheBuJSsE9/nwqHmhPVqFh
tJbMLdzFVosujtKSFhKq3qgh5leYoyxytqvcSCiWZOAnr9rbangv69s5YRcUbpqg
JmxELmDkOjZOVyQRUyusfINu15ZPAwh0F7eL7B6eOEUST9VrgyxNz8ogT8BkuvD2
X35lcng+nURngY1Dr51ycAMonVp7+cfo5wRjEPDRqXnldPsbkVrkkd0Vj6Y7mGeH
K+ARoJdU/GMWyLbZKtUznsojaoeVgW62H6zOwdVF5pRXf1xFngOLnqtZ6C1m+5RC
7fmkgjA3RvzMXMLflv9bUSbe4jZPjKlS1Y8FLbrzjcU2VoF4tXt3l1/T/9KHP28Z
eiB0N2ZjrY8O5V95TvCS8KPBIWhM3C9107trG66b8/mhbVh0KIbqqkcHpfGsqeJy
+oAgcyr/aLSvLzdcyAlTXTTeD8k0/64hhUPboTUODDrzNi2psQEBanlJ5/ZNcnGp
AKvxo6bQXp16v59LQ0GiIaIfQvPXXUQiQQ6w9alk7783Hnx/oiESDHucv1ALcN/0
LvaUP5QhqoqmXhI6+J0v1nDGxGM5CaNzthgcj5TXrPST6z5Fs1x27DLp0k/ZBUfe
cK59ufLn47VL16BABuC5nW/vnqybNeeFeahhrU4oZQavB5JQB9/xUA7T7ggY5inT
8+cB06zV5Oske6kFOPh+1dEL/6IfAz8Tfym9lHUe6nVATck5ieuvHBVxqrPAuGOM
gIb2xTt5tUaeXaBFQq9l+nSXnopu7cfulyclyvigsAdaUvPB97DhqezSZD6zfvCp
Gc0LABttBlGZYY1PpUBv1a+af88gRZLmzsCO/yizIZEfPuohAr04NV6UXoY4d14z
UBDIOn5fM9oNvhUGzAN0VrTKyd9RcnDfXq2D7/QvH5Wmdy8Xg1Is/vYj8vT1j1MI
fxr8LTs6ir+CIKimiLVHwAHG4lKneoWgXPsrA2x2aqJN9PBu4Dv88d/M4+/USa9n
7osq4W0Rxee3PaPguZ6AkZh7CrozYiVwBVzFy/bx1vky9kYKMrfEELispmXsmoPf
dxT5yJ9q3OzHUo7xKvaLV48/WM100vK0imWiCGf4xExRjxqsnBVkZryR10a68nMM
YcP5zKsrOece3kc5RPQwvvGyV4yYmFk6rtKIG6Sz4nIv6C6KG9+xseoFLi+t4J/4
uMEvv81uhlnT3EyRC1vsHqxtCMa4wY5L9UokHr4VKMAzmCtanAXmiipCHub8X6m/
UCMXqfIvYqD/y5xIQYiFQwGFR2JG4HNZqd+/MBKelSpkn67+cksPNipXB4xPlXXm
0Mnop6GM7DedaKrp5FlJz0b/v78a0Z9ROubpwAp57v58qdwniwAcifCyYQJlao3T
iIWGokhhxvP6sfr+/HJRzw01dV1hyGcrZSg7T2DTxFdQ12i2sO12udAfsEq1pDNC
N9jLJiS8r7ikUAZtkG/KY6Z5h2cOuSl8tX/huu9QGqGwfMMKFeq3w1KQEX1LvYYg
Hkfp4is0Y7icH6a81QPLaPDqaT+MsBnZs0TU9cCNSirPdpNchuAcFPU4OI0ZBlM2
N9npLJ8BW1i31P7XoksMBZL/KyefBhDtY7d2RsMaOvJXCb4D5AJKfL59vIPgEfbV
woiORq9AV+BsYKhvYPU8svE7dlmUw2GVSexNOHvVargbJTHZg+HCob4dn4SSzYJw
iAyh/YjCpxjeGntFxP2Mj19fVtO+sPdllGLJUWn2E8Id5j/X5pgikhGzCozACV0c
ksWK/Lzbc0zPUT9el3q/w9dJh3u2B5JJ6zvtfb30aZZEB2U8hV+3kI/LPItuhAMY
2TLxeiJMX+cAqxNWEMl8xfZwcBMAV1HQVx5uz1P8zQiWbPv+xROkeE6bYZnPz8TU
j1SW8sru4G/R7xyQh/B+CTFHndIReZFD7MiHj0rurZrUSbboAlHhx9+Z438BU31a
v2Jgzrl18DDGXFe2kJmuyrP5XBqdGn7V0mivlsBnUFIo57gd3TCcKzW2J+xVqp+S
zqFLhybuclI/g4IdgI0LO9VhhOEODVzqNLxTT36FU2hPHWvkgnq6TCl9FtQp6QZK
GID/fCAbuPhhLNIcCN2dacxEYxeF3MHHE9cXQVc5vjOS4tNLR9relHcSJlNCx9tO
2ZyaU7zRL+YbclWB6mS7hzSi6dFcY6qJG8H0KnP1gFBnIUmj695ws2rcr+SyGdS/
+8yNHazFF9SMv8V0XpuAekV1WF2iMZ65SPeb8Qvo7V6cm9HNjOBBKUSzuRSWpVrC
SC6UXHgUN1TRmw15V1DarbUr9DDzcZKyFmIBmGV0xR0UveHjiSF2FFG+s+8H1rFl
gKuXSchsCe38LasvhivqjA2BkQ0VWWqN29R1wwpIsuv9hya30eIjz4m3O1iOcy5v
JhOdFmKkilJCZHBGP9ZeqC94V7W6kDDh4ETK+3bYvQIwjBQwJCaS3sU46PQ5vSIx
rjjrYb8QGv/OPU7Z/pa5WzSJmm8vzx3KtwjtboxX+3aG/4PTu2Z07VlARaKEYL65
yx67gDCEwUT5pla2UtxiD8RA1qMQ6287uogY6jmrM/2KLXTMM3oqSFo+E+WzgIeZ
a0MpAT3EdHkjX3Ot6yh4EUqaAMAzkkr000+rnrcfqLQSOSd8qUwWuF7RO3XZI8yO
4u6jqQlveQlfFH5Jwm0sk8to9tAYOmVQTck3OKq2EqbeBCFGFv+XKtDYyltTR339
tMJcCRcDJTKbLEuDRFui1oYCgJb8dVCAjk1vs1vpv/wxEO9gcu1+29YEqtrmbR02
xW3+/HsgRo2Fo5JcjJxQ7zilfZZvCko4cWhE5u4bcYL3q+ytnj8DzeQnHc+qZrTB
2AjvZh2Y3Tvu6ikBZ1qRAtguakb/grGaqWdpn2ON/7IpBbaoPDbtlZLKRYTDNPsh
L3v5oTlhbCUCazDsDLJGAPi0p1lQximyQZFv7YNd06bQniqvmAnW4g+EIN91HPcH
4LNKPKD5FooEQtH2FCeVyHOhgJ8g/wOCjSJYydeeGb4AQNJx3H7haqe2PAPwJtR8
minLdBZvcQz7SZa6IIF92lM87uMFRXtd8/++Gqd/5S/irnktcOMKaPStoNCQqXty
FNH5jgTcv5TuYdqVhdV/IxoS8iiNvoUjJX7aywbiCGAXUJz0blCQNXc0E7lEoyOT
EEvqjTUA3kpYMoRO45gCMp/tLwrbPIZ3HrUF28gM//6iap+gyoIDNwB9/VdpHd4Q
xymhMWeKc1PeensqOWlEwpS1nYPgczMe+dPIn23JStEMfnnzad9Bn0nYGnyOEig1
fPKXtUZCRjCMMYs1PioH6ryU2bW/BQ0wNAn2Ie/KCfd0f/ZmsDpS0jg0Imbc0Ymz
ynDKQTAmyWe4WYWluLpzKG7mYWZnP7Kz1+8HcLo+YyvWSgEths0B6K/paqUGj3fF
RJX89z/RsAev8hqGNJpP15iKJJ1lyOR/DA72AaFo/Feco8qt/dvvCfah+1m8KJNd
QpazxC7By/3j9SCyuCXZUYCL3eM/8dVQIumhC3GIJiMpcpTAyDzfJEEjC7fSIOE4
bbM4aEzDuOv3tIhbs6/8y1yvm8+/iTqt7eTXtMguAwX0IbaWu3iExSm/TyClgp+W
hTz45yx4VIIiUmTydA0UNhmoRDv6aomuiWkw32Un1RiUrCwzJffysdpG0KVfNN/G
s8h2B/EWhrPQAcA969jogEoPT5Wl7blo9TuprnT5kpmCJsyrCfehXsWAI7avFqF9
0yZh9OSuKFMs6OTRJK/feEonSVGLdk57xf9czOje/ac49AryR4A1qLxYXuH6XmOz
Rl+CXvqPTpIJj7hMubeVj8CHpvHwpjd2eK4s3xideO9zXt66ckMvaArydWZ2iw+F
PvYh5WzT1OpBHu1QESKIRkcxyAKgj7mpI5B7FbWLm1QbryIeouC+xPSCmkq8mvJM
gWaFEQwl0da+DkLzu1piCzp2j1MOTgN2EcUWa9iGVzUgBk1N6VkOYp1v8OTHHrKK
6AqkGs9Sga4nkyK5tQTzQxRkNVV9P+NtJtj2OyQJjSzfBXNHTXYYFsmj+Jlx+7HL
D8vlNEbNSbG+gnO/caX4wPjf2GgPvKPO7bQnxpH/g6k/8Hf3YL3aO0aNoUGmU076
neF1Mp93nqw9KESNqEGORiz7QFDy7XaWm/Uw7KZjLrRe4RBXi5Ca/lr7XqayIqHh
beRX9jUKQdyp8ojbSpvo0Fv3OsEJ3giqEsdk8gVjzhHj0Q6cD25YUgUc6NxnMSPW
gQgZC989hwwaxsnwF4AKG8cBYNXlFGbvaV/OWwWFE9H3tmRBYs5ORuyId67X0YG1
Y/5qzl/GM5lYdYB+hwHg7WnX4EuZ8F1IBTr1vCuh9/Qmkl0OECZxxZxfSkfSEif/
S6C6MyBwGBGLP9ZVmfayx04G/5PN/MvTx0JrOnsAjl4DqI4DJZ+V4Uop/nVe0SKd
MRYAS8qtIA0tgeFn2U1f/wSSSmSn+XVTNZAQepKxDngEmfDdx5teM2pKVjJ12Z5a
KKrDVwgx5v2BMqwsL3wUkql1j7Or6J9bCxoAqMnM50hmOyFbbACuy+K9bJRxMZhL
p/DS8gUGiQzC4RtNw2FT9sEl2jliUwQWl9VivXJ1crILqZPOUQbLOmp2T8EkoRbE
OygAFhq28TlDSaViH7bkpHvcirbtDMUiIF+DUTs8X/uiqalMdqeqgSIOVsU4q13Y
KaZ2LAdRn8Rj+h2VqPPsq7YIydSLGbxZbNuQ/AgB7E+OOzicp6gtX7cfrxj8FFIX
2ed1o4Dvft0Iga3Q6zJI2Dwp6LKpk4JamRUeoXc4NmWkTJGorDQ8Gw8aSk9uWgg3
2zJvmHx6G4osZBTlRes26gftS0e3PRw2GnM8glVKrDjK4ODAX7I1lx/GclFN3RQ+
1vQlf9lJB+DqnU+rEpJ8y/KCF5XnU+sL4IALBpZzzpLGoTm+2Tpt7bTC0/AbUdPX
ub0lXz8rqbizvWyjrT0nUvHCrQ6fvCGYhWyxbO8zfbJZZyPZcYyPqsCZHnZTs3kJ
YkR8ZROMfc3xgmTfRh5Xb7k6ot2VrsQWvPJZFDUWBSR9s4FjuTeOCSrKiYFEIQst
Stt4NIA28NZgRdFY9wJrNGevy+QD4FD55Kp4KFVpbR2MHq72t2BFsx85GkEGJ6xk
/XUUKx3PD8uOy5b3+iw6AwG2zJHZuXZeVPsRCSm0noXone0/vbz1Rk1W+un70P5h
3eNrkpb/e/FHZlmepRfd4ZCOI48w9GEczKTgV3E7GaLoFOqOU4Wj5ntq7DHizF4l
dBVF0Yqz8cluMxJ9/C+WAN/x9iSEv0cCPfya2SoYjP3uDXmEHZFe0Avp+MDSH9Ra
9fy/Al1+NyoE8ZUaMnID0YWsutLhocBJyLnlk5lE95zbhIf6pcu6ub7guei8Y/7g
/lWj3DBFm/7n7XRtS4/+Qtaicu301COj/u8YS0KMVK3//pxY8FET4pcl983Q14/E
TS/wd/f1SARxJeu9H1eu4Hoa3TXbhVg5yAXfmNeydaJp9Dli3y7+KLj0agkKREZy
bLHsUJY/nELgh+/nH3onboH+FDAtFtJsoCxuhRrfQ8d8MCrQuutMFJJN48lIzKRf
spuM/B2nI/2Te7eIvWGk1Y251o69+vKdzjndkxghAlaKl37l9RQIeW8REyw8Rgfg
VOJgNmKa2V0Jrl87onN6fwUo/vkLW7DhQUN73G+EevosnpVR5ArkrkBV1Ml7wJrA
rfL57eqAJWhGAvBSLwlGvtrU9k7Zb+kCA5js5VlsCkuJha3q7T8F+OCYBtuI76Ca
CiWE3hHkujjV9ZO9s/og8IIChMOrIj1eJr0KUmye3jzxhOu5yko3B2Td2pwUTlBm
CJWiVKcVX64mnRLVFYq6ChYgLNVOgDEUQpLAxLTYMhK5QvOWaEoNU4rthPsVVM67
6iVfkM5fMJhXOKhS/JPFn6dtC0AIVV/Hv7nVxw2GKew5CsAQ1k9Dj4G2DHvzGrH9
KuBU5EtB5H1VxuRFNXEeMSFEsM+Gy0ShX0e15mX1QYJE3YNLW1vplNI0DoJ4I7HL
DRZ9kZnEqtz2qLYlVwQubeJIgUyC/AxEscVlhGuF6dvIulgRqR6bMBXpPNVfztCN
5uYTK2Ep7wAF0LQo+hOTw6hHZA6Mp3krn4icK6g6yqhu8IQ9gCo5pt0oqF2m87fk
qjlhHHMAh+ighXPsP6PnW73t6po16jaxJdcWFZxNQW9wJLKK13rM7tlN7+dPdOUQ
75m/QoVM+b7q7HRQ+W7YJk9lNSOgYlJP7XPKMFw3dFcXNBT/OR89hQJrLJZ/+ih2
q/40QYoaucY1R8KkrlEdul5erViCshia/3CUU437NFBUW22AeaGgtAM8fXUoxPMO
pARUp7kuG+guoza5D+yElt7l+xFk218DnZzFcBqvH0HHagh6b5/2sFXQgmRfNyzb
msmka5XBz1/da5A37udGwZXL3b6MzwaMse8oL9xPJ0SnumzuECZLE7Lmzif7/hzw
FPSWv8V4ceuez79H+uhUWjKTTqp9A7Tu/RVDa457u++0l1kKJI0fvznNfeQvl2+q
zK5bXNOU3deLhgTdS0kCqFpTahjF6BSl3Eh4c8rMFWbq1TF6BmFyvBKER/qneP14
GBTYk/8BJbWEYkc/HSlohDPLPZiwODP2AMpmXyY5IOVzm6uRt8IZSeW4OEqNqqiY
IomcGGUyDhU+ekqwbImHe38oS2/tiSmuV2ajN2VPqiNk0Zfbr1EHGXw/chmboyHD
Mco9vTa8dbl15XVW5xKoNLv6v4gHYgGlYD+aSGCiii7u8Tx7pltZ+cVp62TSuKch
3s+Rb3DL7qiQS42uXbO4U6D5ZdzvXH17zpFSsGGTtwZ3v740cHktmT9r4tSpw9ks
kLX8uvSklUhJd5WZSuxE696XzLz+EwFBGXyz1qH0JUpy8Lo98Y0p5woXNH400k+S
dnJsTM7m5u6wjWhYk+id5zBm05o9Mux/bbuxMjOPUlHVyhAqRjvEPsga17rndAln
WvrWHC4RKcb7OThD88Sc1T4tqjdtGBIx+P27ARUOK/QJQN7HnOOD4+Gm5PhcpfpS
79KTpZwgTO2MFkUOWYPdFkMkn9HyJBoz9UEmE/wnszX9CWQMs7NZltTijgsd+xmN
PZpp3sY9rL5UEtOeW2YUCDk90IHthdUf8mDm/Fr1XcSzlncuLmODwwvlpmNs9kqQ
7JpigSDZpBhL4C85ryumHwT9n6eo276VHV4vmmq3Zn6/Es44BQVN9Pznb0DFRH0S
j55J7lkxfgrruufIhWwHIeD/k8dIHlEBI48XrfN1HWDqecK0B1QAMwCgctaRgPLd
fh0/RkD0Yl/Vgif2gEaHNRv54YbCp5IBK+W2bE3mu6LyZDvzA8nSxDZN4nZO2Ybt
QqGmfDoloQlgbxw5M/yEmJAXHlIwv6Prvdy8c8njkQCSHjbqw4j478bNv6TXk/JX
p7YkiKSVXmMwCZO4o9OQluRUmFbZi5bTgi4c+qGzzByxcZOY+xkeYPG/RD/FrRu5
lkkoAgeHv3nsv1hDdXJKfyxUJxu9WCXinOwaPoA0cLh+cl2SrEJ5q533LMjFFg9K
nFLvAMA0uK+JRl2vXeXo3op7dW7muQcP9GD3knaErpmurneUnGwPo+fiLuVhq7e2
B53U3mioBA1vksVGHoDKcmPkawSs34XUccc3cJFdNFnilo7jFilDm49h28UYbih8
F4bD9GiCJ4lXlsfgo+Pq73cVlsAMA2LuZ/ip+t9TYw9V6+39BkbR7pGBuCUVpXH+
hVOEKma8d8HW7Ilevo/8kw6MMUDlTvwz9LVofzX18lFEgn8cJfnCD9t7CUkZODRv
8Fms9DmXBrdsJsDl4iRbcCsoXcSNAmA5Y7I7q6E8j0Mgy1d4LAu4KPT79O/RLWoV
J+V+90k8WRWaJa6AhLqXUu+PJdb/K2KyIglzDaZnjqkAcdmgwZ6yf3h00m5ktPhY
xbc5/FfK+FB5JIROo6/nrkFa6QQGfOZqN/MUC0LsR9Fr24gZdQeSEpHrHYIxkD1F
EL0+VsE8jWEvY3As8HNg9/vj4XsckUJi16fLWBNzg1NeopoBs9uqgWXBQwXtv5ws
IPD1vGwZGKNI6XZQsLCM4Hj5ctDiKHhB+1x39VlqG6p6LPNbkW5mSMxW3FrDAVh+
s81HEbSoaJ/nSf6Ao88jrSLjy07erzTpImqsQkgh/6KZikEiSahIIM22da8y1tri
vDxEk1pcUH8bQM3bDYK07JmruPjWjC3undMIe2uNSvJUQj1AMr+E1J/c7U1/Sz4a
0GEflFFxs3bnxp/apDf82Rr08uWpZ/D9Kdo+NPZr5VoQWBPeE7aMKJw+M5Ve8led
onZ7gx/t/wMa5AzUJZ3PohmGGpACFwI6MlM6z9+yt26EeCqwP9cJkVDGFHGhBuTj
iXbL7BQ4OroFo8aOqeP0/sAWQD9gUtI4K8BmxGt/X+iOHFN0Ff+ypSKeJ0pJYxRI
P0GQTJXecjRjIp6wzd3sQPFC4kHqCdVhUmDmbvmyz+PpN56afn1DkK5bFxvx5H+7
nsjD7dQMsKBbebjlBoZ5+q1xi+0BfZicxLwBPXnCDI1DcGjF7HDx7QzTDpSijjdD
6cGNDaQcvD9cXmMVGiLd2xwo5fTrSAlrxg9ZkhCoKtnNNXYcm93tOFjnEJ05gFB+
v+QnvSzroqEuMzVVSJywPjO1lYUklxGo0Lps9YNwjg+CCMFhubFN1yXpWTTTajnW
A/C5U2unx/3827tkLw02403ZXWUCbZsBqmEMzWKPysrmq679DMAVoeiOdWk0Xn5h
yFAaskklR6LLoLnXNd57CPpR43Y2wmlmh5gNbRB2axNsxV+M9xKeAQyOheVl9ox/
gWVMtJTtMn6xuNnqbrQmRVV43+n6ZB/l5r4uY8udm6dVy15CrBH7eUqJnwv9V6wg
rg4QQln8UuNtPRQEGg9bMKuX9JsycgTTEAjJLPl72rpNIDVsn2BPeEn6ZXhjyMCX
lNAkM8vPCoHZO8K21Ls9rIhlk+NYEqIBl+uNH8PwDFhj1sN09S4LwDjCZZYX70Ii
yDKcxbgvlhb73vNPXeE7ISze8IId1lJzqJBEnPZZG+xbmnViGO/ErT2RiOudJLGm
juyHkiCNnLyQrum8+io7Bhtug7SYdQm57qzX9o5ecTZq7fx/Sbv5C7UkNMRimrXn
alt5CXsczUoW2tQs7FrOYxydYMFKTjbYgjPrBDiShpcCEB7h/S4nPnYc29w1UGk7
1AWgZ+/ArFUOzOrNCBpnFGLjDjMbQtpmVvTBoITt5zk=
`protect end_protected