`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
ddtXksX2+yylW5zu6QL2Lhnb2d1sD00763mmSITNX595NcHTEkwn0zB1Dry37fOW
FufOhVzEJp80NC5qZ/+F0Vk7Ik02dIR0elf3clrjeJRK85K4e3Hoo4xn7YbFUIms
l/8VZSb14+JVGURjfswrIyCUotIzlzVYZ6gzoZwDXIi5gQIBf/gI+KxNXPaKV+PQ
Ufys/12rjO6aI/pPlqSm0hCvftmBcnezN2hk1UeXgOIuKZnogjOsf0iJVX2aOOWE
6pD/psybjbnsNB6kH5uFTA5frkzIzkzl5d9+YDm9OyC+k84E83I/7/j+rk4L2dah
QJOvksSIzN867/4Qt8qYTQ==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="MvBXkzurAa5VTw+1JJ70nePUfoQXBvZOku/SMmg4TwQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
oRtzZL4VJ4iwysPsC8SXYCzXS8Fw2gtZTOskLcDV+1B9Nzn1zTyNtlo6lNICRmmK
ZRVu2BmCc2G+fmzynYlNTnSa7C0Cuel6FYpxCBlOuk3OF2tzAmLAuDyOH3Z1Yjzk
a0aHuoCdIRKv7BrZCdALt03JeUmXKPdOmIlkVGFl8yw=
`protect rights_digest_method = "sha256"
`protect end_toolblock="Jn9CQpRhJt4rnzZPRk+dOpzAubz7omckX1MrFd4p81o="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 9616 )
`protect data_block
gD6l00tciPUa6pDNTk/+t0OO0nC/UTtBwLB41d4inuAUA3i/ALrNyoJVcBnAmEQW
ptbcNp5fxEUJjnOxnedyZEuEBxWRieZFQnkRdF269oODwPbjA0cHbnv8EZVl1yQV
FLEd289fxh5w98f+m6MbOsCIjK9VWPD9+tL7giJLpkCMiJLTLyrYq6ckv5rtGeof
r6TUHgmgzJzQcyffmazIOqUG/sF9QAqKgxs+WMXn7YClxnIcvpTiZ5l2tfFQ4zAR
5D6xarZYlKcu0lbvYiRYnuFBnsmetPlHXPXknypETi5J0v6gJCcB7b/z35zwvpgJ
RfgbEsAPMbBHwGh6khojOPSagGSLJY2BnnqhNqn8KeuQ7xEqwq0KtzVXj07PTeAj
sxpnuMkIQo/gFYeR/SDNEjy4sq6WR0c0VXjTSD0djPBNMBN8v0fpeisHp6Nw5Qun
p+a/YOLnWnNUNW07O27mmBJ0nl/6nB/8g7tzka4J2tByQ/H2qFYgWLjmMKqXLyzx
A4cgDB6SzygJPvWAQhBYImYeBiZD8dhcjU5DvpRPF4B1VtN/9u+Nn0UOCnAaeK1n
jnqCWgU0CrS5wQZlJae27T/mPsxyfIxvF5i4uPFq4XmnbndCEEDoxZEQA7VN7grC
6ua33FcVKpPo/WP44WzAvAWxyVfX68U5a1BsP2XQ45dn5mhHdz6PD38MnZzJMHD8
ZIAP8oC46LFq34IRn8T29T0jiS9+XdQerB6Yi6pKN96Ys5YjZCUIPamlapUyGSLQ
rN1NyBOL0E5ypKRWeRf7lKVM2yNOgR1ewzNJhn1vzdbTwQ8NJe8QgDsHSS2o8FzX
5flupASx989oPb+r8wCoaRL3qL86Pqe1X59IpmcFYsUom3l/qWg8VfHDuJEK+yBW
GmgieK+rNgFgEitdfX5AUbkruCfAiUBUYqLR/G5qquEjN6JFXm+uTIpvcHaJg6L8
8x3gCt/Iuw+6REBDpp0loECphhEOg2RVxfd/gKOGyjipLSzatIgJbZhKexFrWrpL
rcXHEEW7toRyyYPvuoe+hbaWQ/ytTJOhvIMwjEzXDOjGmjpDcAkFs8DdhxRCTT9p
ESGIIxXCJFIvEenAkgcmEgOn7h8GPbMu/g3t4gDI1H+H+J8z87tdOlDCEnul7bkw
zYisUiHePyuFl3+WmV8/aFmMC56qowfQsuhI9q27oC5T20JGGyPdfA2eKKkE+Q7U
TygzdPMHN3o39w9N5XyVRj4jJVnIo7W7hlkHEc5PuBuyXzQK96jTW/uNkU63VPqs
xp7UB79gD/6N/vXOSkft7OajUqDVdPJHUcuOvfwdYKmSY2v8zEslQ8X/7WlKxRi2
coV0O0ieqZ4XTxuW2KNHIHOviR5nbFb3/+FyVDmoG4RZIatm6tmiIA1NKJi7szTt
A04upOpUyMnNE2T4iQK4bZ8JevmcbAmpHfNPwd1S1vYD3ZQD6EmX81G6SQue6eKg
3//obHCBjDLcg1E9UTbSz4gA69JTr8AA+TtAFyN9HyzNm2EKNi0Huo0DGHAztTme
4+hTUFWoFazzbFuc2zfkJ6AX5hVCVSFzy4emcBrtZHMCPowUqAZcvu9ooIEUw1LQ
tc4hICNg/uIt5kz3ojZqIY0kpi+yXmnbV50J6BH42TkNIs/kwGHfxBZ2DgTsR2si
/E3GEc+aTxk9ozSV+i2dgzjQpmDFo+YZAXF+emuNgXm4E7tssz4fOZ5JxzGLV/ds
pgs1ZspmDFVKkE0R2SUwZhWNotIGK2JZP5hnj84HYjkl2ng5/FNu+mdQnPUoBojg
V26vQh+0GZ0LZugJhxnKtC53x1rvWLmjkyIM+YxWEcxYVj32WxIXtTrzusaausUn
zAId/xltRuyMw6zr07cJmgARh8wRn+8/sjX96ssCwSKkLj06dTXJRXBojMHG2CfI
g1Bj8yAKN1mfrBhVftEf/pyuU8C7y2hk3H6JHnP+gXfDVYdiT32Hjgof/BKNb4BT
tV6dlVwKtElZE/2C1xEBBYxfYyRWI/0HUlnQl2ThciPgCs+KrIOc3ZhcknKzPd03
e5U1nGAZgM9wFASc132Yf0QUEuoS9fMLUXlL0ZYEPKfvMuxdx/P0577UoQZcW3m7
5mNxn9OXjoaMMX31EnWR82rhXyEyHrSVz4dgUA+2CnMvpP0CVM0qpzX4Lrx6qjMj
/2k3rONuSSRE4jlWjJMKyIKSbknChKyxvmsmwLn9z0M6p/ysDzkwrsph/CAjH7G1
BjcnPkafohjM5lIn3ABxonaQPFiX+37AOm7QS/YO4hbHcBEbR34BEgd+JDJmdJ/q
NBVYkZNW07akVKRtdZ5tDIK60z8i7J94vNN6HhL55gPIwiM93CWlRy4Lak6xEyrm
VAHqG2F1B/h21Z4Ya1ZMlkV/ff/LRUHaDbPOXTY5DWNpXxJZGu8hHMMyfDAf2Z5w
EjiaACy3opgG7CfKlFPK99R6xG5HkBgnbMB9nVbEMJ4WwVpXx29sp+xgBElQeMsZ
SbLMmQszn4ZZsj87rEFOKOSsxyA5H8goTJ4YhNqEbPgz+g6gncDYz/xxcj8QgQhC
dMDlbyLuEeJD6G9v4dtv6tdohzVvUD+YdlyfyzinMTJZ9G9jw01hHsVEesQNsxYi
VEEXpqm5vKbvYLMqAe62LfdXgV/NLfXPOa4uzYk3EGBJjm5DrugRAyM+QrwoZ2Rd
oO7ME2fJLXGPskTxjXNTvGhRPTq3GkUb7Zke+XHM9sy2wWpOSZitkxDNdeYVbjUc
paJQKmIEeVaYagjTOjdlgNrsI+cdfyaWAOFPmSHlOGKdk0KKWHTroKgAS6jgVVuS
E69M8r27FUm2New0HC/f/OBTfKzxIfmV8BGxh62qjWDpFmZ2jpZXPnFjxK4DqCbb
N9rVaTTZVvtP8QN/Iy28Ct+w6Tfk7H35vmF7BbO1IrAh1+OWjXBcDILtL1RZCRUD
AgaOP4x+bKzQ8SSq9BqKAUSUHR9uxL6qHqOl0j9KTtVH+4r3oQ8hFNSscIckEg+5
P/NvclcCWiHn1PxqPjMsG/n5ic6bZXvVt6FoN8EQ3XH0OfzJpHh5PNS/k5r1inVH
oMNDOvoebrJmNzYRKdru+D/bZY0qJ8JyRQgoKQAbPGvsIspNubzuM00XQnfDSa7D
K2ZX3fPjTYPXWFBCdl9mveFLOx/EGOCb0rjy91luZNfDA+FcTxelregfnOVZk50e
FFL5XxhjIOHqi22MCeTikUPHPvaz6IbzwruPC9KY+w8SRJ2BzUTKVQi0CMcrdwee
YzPa8suA2zA1YhE74O0Howibt6iKvegnvxTaxuEXX7jsA1Cra8tcmSv+qmHqZzkq
kWLhWFhgv1WVjGZthSTuiUVRnUVwMnj42aLf9unnow+QcwKuBhuD5j5Vj7WDTk8r
pqpNqcDZRrgIwGvJFsvLWQ/i0/5tEEXUPj2pU0/BUVBKuNmkIY7TpUXrhocNA+W7
/DmIZKDGcQVpAuhrmxx/gc6B1nAWE+Q0ki2Y5jkY46LNd+VuZqarFBaIe0pm2mr5
/cPQbeTQ/Gy39XTi3d+cmKavVcYvdkjauhA9FVAYj0FFy+8X99G6cIklCslDdU6Z
HrmdW7/XwiKbu2Z/IoQBAWZzgsNfdoWHU5GCpSiy/4slWjB9h+yOz1XP0bKDz2KC
gNYtuGYisYppZr8yW1X5GYTaj5oUEyM9QWaUKcrVntwMDKcRgPd+lNfRzGZ/mkTO
s4sCebDbxrZnPS9nVC2khF2ox3+q2Y/oKPfHx9vtg1Ljv3v2cj/ZuixCaCs5k8DR
xfrEqHyGqmPKED02XaL4vwNUYTgra5dcb9xRvZeK4SwCjDDxCi5a1ZZFsS0n0MgX
ntv0Arncf/nfMtjIYBmFRrI/JG0tKNxUUbI6TXFSzHyRJmNlICktDykk/jHRH0vs
D6YOEfcV6IxVxrQC75Mjd5jwXKBCPv23sKOjPFhR3mHc+bMDemrgBA6T5Kwpl3rE
4YdEX51gsA5VfPWe7b+gThPYjOL23pm3Q7/qI3CCnhmO2XMQMcER4+61qUvxJzWE
LcFAE/mevbzcBIOMaPPAFe2pqJU4i9U91PIjnJ5T/CYkbz2EPjp0rSEsJ+JMgo+Y
FYKgswjdh9XpvVVLLG39mZfr8T46RpkgoW+kdx/aHRBIgWB3hi+dScTZEGmxN/lw
hPfwh/T5hxIgkzqV2Qn2C6c6w8JKz04IdENhV7Hjuo21rCUOX3uHTsPVVuHiGP3p
uRFVQ8Wv6KnIMAlT0pLbGfmvP8rzXAODgG/Lq+RPA8RfTTaWL3fLQ/7BA/97J7su
tey7/mf5L5rVpKwP1Rvh0ULoqETZAz5PV58CG6pYgDSUu3firXeLJFT9ctfbIqLx
Yve2x3okmELVH6ZYTcaa8nuqJpP0ov3D4KU/NniZEmudA0/icIxgUbudu9mL3I2L
qzHO2ZSaxdTe70Xn5xb8arBeJHdkSmrHLw1flq+TY/dp02u+XNX/xLyDlQQ1jcdv
iyGxa4qckctPhnQS9go84RJEuB1s9FxUj/cmU7WnJTsIjH0KYgAoZo8449kH91sS
5N4XFJtk3xF7QYfYpZMISp+qdE2a52IqWj/ceBNTr97Mrhf/C0Xitr+iVPVgy+wE
br0BjYGCbyLoPRdaJR/ecAvxUOLhDLOxgGTYwAGnqWFVOBuGXYSHRoAqOuPItR1k
0EJzkFl3CvuBYbm2yR6oknytBlBjKn7jJRIPfVOu8glA+Rwho6dtah87Jb5v1TgN
5mur2N606B8OuL3ZGTpZuqOGeGkmNGGcMbSsg/STXKLcHr0Kby5gs637cU1j1Lkb
Ct5jxdNJ0UAl7sf1wOn9cs2KdtMiK13Idmb7vyE0Se07FCKOLbBV71YD/FuknIY3
1LXyVHA44Ia/0J9jtHoWAVCcRTcKrHM2/82ICOlpanIHxJujzCcI5FNRmAYZ98Ug
L3vfJ68EytbNDSUHDA8cUwsnTpeDZWJBoA8AB7EQYB+QQwnan8/HP5Ew84xezg+/
lfzhx4liOKkxeuvAjMTrdsdxhbVHOsHWblXBRywX3B5waHSQ8caZZ+YG3FudlegD
So/QAjjDebIUzowuIk2kmXyZIm4JgJculSbIaAplnkJOJ2F8yt2dvzwfpvdavOd+
95yMtQopo1tikQhCL7EnW6tQiK4G5jBg+blOrmuEhLQHaQPUMAOpXtJD6wAzw1Rd
JSmIw2dJ5VGl5MiBlWqI7FywWjSQ6ceWJ27NH5d+FgK0C0C7fR7lQaVznPi3D4Iq
SPmVQB4aneZxJg7ymFenw4NGC8YXFrGtN/5q77/mkxM1WQJwU1BjKQ8DOGTR87kh
yyN2S3AvO5zj8wm5YsN5/riR1tuOWfKUXXmooq6yfF/4qHfRmxaS1utYv+a93pQK
KDtiACB208PpYcUEdf2Lu72opAUkrwnrvMBKOOQdwFKA8Nohz9PcIZQTetyK+nrU
m9vvQ44/iNT87JHfKxgqV/m1zWueaT4Zvy18irZ+CcExaDqzle7EJjo0j9Gu87nW
oZK82bQDwbPblgvrIrvdaTTOw1UDmaQHvmd2JCKfj/RcNh4EqccrCLiL83y8YRF4
7rspABzY5JycQ12CUqhbzln9M4N0sr+tfK66Aw+TPZ2Vf8AMtJJF4tY1Jiiu9Ahe
JJruek23dsgJRtrYfxfxysiToaNmV6Eyg+afdh+aF3fYEPcy7KfJiNw6QuhIh7zT
K3m+mMzYTmOnsM/LcIa2INDeklEtw7Pb47qE/afDp9LJoS+YZSh1LckcmOHtNEbI
Ts2Z7yQfBby7gwz6KpfwQDgq0Og8mw/JMDMlBjxuYVZ05+ycufIvItgrzO7wQabe
xIvq8JCZ2rNis7/h9g41UiXtDWG3cbEc4n85beV81H/Gypsjc5I7+I3gJSXWwLN8
Aa6JumX9TQz7+Jz1Fg/ZbhwAoadrUbnc6tC5mKi/ZlIw+lB7A5qEL/uusrUY1d3e
7aEUdl54+BO12G5/nOP0t7/W2ElTrGw3/RSSCCb0ppIIleuMgBgfr0jlIhsFtTMB
2CUYBY3YPODXpRii4ehtN0t/rG7Cgt2z6Lr5o0p3y4x/Qgo+GQEf8u/6DBn/kLkq
QGkqANW3VQK9t0h0y5blwiIS0ueRgPqtJiuIC+wEN5JCEfQADwSRJQ6mL/39GVJo
KoTSh1+7462YHUOk+7YE2R8gMZMqPcDaylg72GtbzJpjtE7Yd/lKw+7418WGKaiu
6BSssa4jPdpb/jPxlVZikj558DQis4oNzWB2TEbPuV3nmf9d9Hyt7SxdemUeL6mS
jOeFIEBvA8rLx+xcYRBbI3h5zNlNuEztWZbeiqCqbBO0UZ3HIiAs8ycDnYZxdTCe
ANIXNZOfYG440cbKq4SvpYvuiFGQJhcI0gT3z/yMN+tdnCu84VP8kfsZryn35MEf
ekyq4yRZxiYXMzj7GEOBTZ/x26rkXVBufAhtX+MRmQ7meJ5dmUu2NjhiyFvc/jBO
8vCGbd5wHZHQwMoyfoGfRRPdJi7mJhZtsJtz5WQzDaMo2F70JOBFIB7VMyVNX4Zh
xwC+1ACRgAKH8XPas83fIZJTIPxJNp/+LR54Q3EyEvMDXzu17Q3HMt1s8c3T0JAa
RuKruymxvfGd7aYH7NEtsy35r7jeqbMZaHeVVPrVYiyQm9CrsMs8t94H8KPPrNi6
sZIWbasBklWtRiqO8U10HDB/jJEd1XK/fB3xrEUrjHKzPmwcYp9KJ68YQNwPTxyw
/Sv78psCU7z9C5Bibx6V3SODEM0Gk0DS6+liG9ZPB5I8VFDUu3Z07/wUmmcqwKF1
r4lk+ig3ZVSsP20cfC7WBxnpkr/FKG4T0YYK8TOXtOIsVEhxQ/zNm4D9EPRMSJ0p
NAylr4XOEonEU2nY9waJPvGNqi/nE6nULuWm3drcv8MAth9kz8D3b20/J52JdjDm
JBvvmZYicsl92WnlrEfDyWa/adm3IcbuHhxgl9JXl2JFlTGvmpNMahO4OTzALeHy
YJnLoKhP7ZC/5KsqCAgvGX1EWOHUSID+UI5XQj5zqFf9T+iCeDEjKmS33pj5kmIy
TQ/ZwM0GAGeXvlY121tvkcIEo2Uevno7EQeODaDn1Qs7/FfEXiEK0qBIkeq8w8vi
7F8+XoaOfMZ2Nyn22Ue9m3B71oAA0111dI9nDD3i1PU535frFHPbj43SUrSJTPNu
o3PMfVz4Q758fXc1yd8ooIRyOsAP3MpFBYn1XXuWKm4YwnYtQ4IyDYoSjMbuVExe
wRpeGfMbCGVafzzljErcor2BcZDn2mEHckcQ3t+pHHXLEHXCLEKxJ7NvYMipDah2
pkdMqOTbpvJrc2wtVoV/Jn2E6SOf3gUmWnYqbSEPAYiB3Gd9Etj6OGOT60zXaWnp
JvXE7nULkGd51p8ulSaLo6TDRbRHLVJPlDjSaMGp/BOMa9EB9U9vPYwjwSj1QIAT
A3qloP0520VN/v23z2Oq8Sk3bboVzKGGEm8F7vCooiK77cd8MkTupfPAOT7WmZ2P
tf6JMugAUE7/MsFwjHIA3QTJtCLMUeu/oYCIyNPwAmuoOqIFc67drR+rrT6Hv0J1
ZPurhovfLfKrF+htERT9KsjcBCtW70KCRgsfeV6/r/MohVy5DLFQc7h3U6I//NkX
fqHld6wNyuUlmrlvkvCDKTqCAA87c/5/rftZdO11A45Tol5Leu98RjACwHNY3/ru
JVtkWlz5+K+u9EwgpuWk5Cf7Mzh5VS4vu1N/OWw2clu5+EDtE6MR7cNcw0IE39vn
urd59C7qQAsSR2tFzYMScCDOTu0dTFKjgDsR2kCVrf7D60RcvTNLK+im1z6JjKHc
ZDPbIMOUZlcKKpF1OrPf6bCl/dVHoY/7eaeYUcfAPmuk0VBwmhrdIlXfMS4iD2bv
bFPXnW7Z4N/ZaZEfy6CvkJbFTnm3LxswjQRJyu7ny9eEt8ucBkuTzRZB0m1v3rso
z/MAVlW5/1AMtqv1+o2hVwNsbcyHHc+f0idbZu0p89zzZYIHgjeZ2kUkB3yzdxk4
XYTqP/0I14ReeJLcavbG/KUAHUmycwDwv1RncnS8+yM3GHEG0f/iGbyovqB7myfE
qEOlY6ASpSSDG00p7lj9HW4dnfq123KN3mfZ5wD5LQf3yWjKQ+rd/EXpP+FmpeCf
HGpybhxn36xQAMs2SPVPbnH9b/h56DX51Cx3QWxayLYW/Npo+XkpqE4w3DZwR8G9
rGhoIF4mE4ojGqCzubfUXPc2QuRAMUCM8SoXUtQtMfnRTQRRiNHt0Zgyo8W2OscE
fQRKkhE7PTBKD7cQf2JODrBqsS1hm7XHOhZFLVklnzgjIll9LqbutYA1iVns2RhF
NQgdeuWgL5VC6kwOc2Sr257UVPFzk72BggWa2Ot3x+WKc9nuF9Qsa02E0Qr66RuR
iHU+g+CtZoGDEv42T6796yNZDtXPqpxpauE2QP090FBeDFCA9LQZt0FUt1S6umzF
aAnC0uKqc3EbYA4HW8OmbfQVSu4l+Dj1n0D5WC7OzIGX8Za1Krn7wC90lLUvbVRo
bd3LQ/jTEpKsJPtRWtJvIdDV2Rse0znWcG6hOqWkB0dCyDJoLmTwiri4wvN6t6oY
hs5Su9rGBoDdDgdQKov+2rzpq8CWRFuBaTtH2h7k4+gopun+pRbBH3szH2dY6xFS
7P2rVqXb8rXC/HoOgRed9ESUMhkzyZco2u9+BM3Z4FXHJ4BI0L7516YbLQj1b0KS
1ETe3sLDip3OHiRmpXiblAbDCe3/CelvsZMVt7pfrB6qTFQEx7WCdd2DMpWByeIi
VyvmozCKxWli+Mmu7I73KoY6RMDSai4ZU8pDGsVOpEPOHIesjWBSgJzViSwJsexO
GowxItKORTvAtOFQNgWyktrB3ONdEhyk7FF75sFK4CTeI2U519Si5I08GCAgrx96
a3+tLN3Yaq/CwO/p0OhUgi4CkGTVmId4F4GWTaeABJ5nYkjQJUT375pm0maTdj1b
kPolE6IO3RBUd4/85Z4hZ8apqcIlrEndE6+VgUevKNzz4LuDnv9WVwzt2JWN9cuA
skk0Sq3uccxsmzKDFBPsGyqmkj62oZb7qNAGiD32cnwsXMJT7lpKMTEkdPDr5utM
fjXeOH847W9lRdL05kPgh4E86JvJnqG3HHwxhaInPxOKu+Oa9vwIEILzh1F3NMC9
R9r73VhYXlZp4jeu9qezOaDmpKHPELx7IOnYIAus2qJb8NAfkdh2rw7Udqdgj5lK
WVWRJzU/E/1MsR5joiosefFLeZ0disFv4l/yjh2xJfxNQlC7uqyiUJTQsqjgDOog
gP/B0xs2zrQAeWS6scEv6bGfYqUwoJoofMJfRHshv00dblPsdi7goC+HUk3zUn+G
Hd/JjkurQkU8MKWZ9riXTRNQb5bLsE3PGVY62NqNFnM5WiWjUr12xQ2nJQcettc3
NP7kFrteQYp5F5sIi2rgBI9c0+T1NA+aHkfsm4Zai4DMzDB80cF5SAbxnDURRlgC
iFWzmMaML7lK+3VJgi0z5lhT64+z2uPVU4pUU3jw19Ji/Mcax+/7Ip+846nblyck
Wqgnf/3Fg7eKevLwtuE3e9IacPISxpJr4TCm4GrrEy7hqf+X+YauDbwNplG5lRM3
VWCjcXO3YjB7RKrmtPBDb/n9BAvVjJIT75nvMUM/dgESunJ5FEs7bpEOjJud1oVi
ArO8QjrZWwZFo2gB9N4U8Nu2ZAu+xqqPy3CSBFp1loXuK562A6LDRBw7XSrMhmAV
5RSLjprQ8Vji0tO1arK31QTrGaxG/Dqd+cncROcdV40cqOkf8k0m06G9t5nxwGUx
PFyC6DV+L/7ORtoBvZEIs79lxZ7L0wPljoK1lkJF4xZQcWCHEMCqWvh65iU7bWNO
FesowKRPl0Bw3rh2Ei5O7NlbZyN8k+I9WYxGpA06yD1E10oheUMTPi+02zJYl35E
Rs5YiLV638nZzyPRGOTahQ7nZTazV5hET6xeV6wcS1UwTI+lrLz9W3xPcLtpRqOj
Qemzgi23Lxyq/haYtwWcGQRq7/PxY+rOaRvqYeuuqBQFM108Bi0Fuyf3Gy/BZ0gI
0lOJfVtXK7SWmr9Bo9DY7HZiek2LkCWRBWeqYBtis6z50x0rIfVH3TpLm1BHeDCO
q+BEOZ9YQV31TDM0+o5o5Fuo+4onGm/7DQUCbwWqc5XplBjfzlTUc3dV6bchlb0v
7nznf7NgATA1Trt76eajGXYNpsQ40C7OxwI6Tkj+2W0Xe3K0mY5YpdcfyCwRS4KF
hRq6zN1D69LIlWWbpY53T+1QeBMJmhjp3VjFZcj19o1qd5WznSqpWSzk75d64Z/K
mRK+0UKEdKQUA3pm6knUxAA5DyURjynm6ni/JwBDrY+v984+V4V4L6j8fskjehxu
s8ne1cV/BVRFrqk1IO4R+ssRW7+aBKtmsNdl7co2i4/BmFi93Ar82YcY95JCkKk7
pKArB8AOaygyScXbnzqIbOnlPxs6sS0XZuI4MaDI9VzZBhWmLMBD3T5SL9tMHIib
o7v9EsQGUjd6DWSqUgz5l7EA/OUP38gUOj7dwnk+kJWP+jif02r4zZyJRdbAF9FM
1yabCNPKgdBr27dp54ThV13/v97heZ/rREOu+8xRW9O7Ee3mYB36QsOPk7iKMPdD
VjrMRFX05uq+OrOFj25prHqULbscSEH1+twp4a3x5lljSL+SYJvVkMQiFLrWrZAR
sEC/axyFDhEaSQKB2swBTvE/tYS06iLjc4KjVGQmLTAw0ftViOVV+TY7WYmyIXoD
CDfDwEcUHUXbQmSUlTSO7AJQ/Ndcf2F6EAsaqKzDFtVprYX34Vj275uQa2Oxu/tA
du8ok94CAb6G4Om6XzE//m1oxXoQrWadKPkBKrqmGuIkeS7qrt/ZeAOjsNBZVFPu
A9lLzD4/VRUQFbf1uMobd6wmhDYWDG4tBf7hdpVH6U0VOVt5oM8AaDRRaOt8FRBL
DbMCwbCdxyxmnU5v5yALL97cG7z0wv6BZEy2oCEY6FObI9OxtnWX3NaQhPT6MWFM
wOoy2eK2/AKkBysDEUI6+EYLA3l+E+f1DKj3z1FcyTsU/9ZR92b6acrcwQJdu8tT
/161tcuQyZIIRxd0u4WLRR6eEqM6QaBBKcz3x+tkCf6DiSqUIuXIpq/aPyVpOJrm
PiY0xBwsm01osXh9hhYLyztGbmIXqo+NUPYypub9YgV/1W3pkqX4uoTCqiT6K1in
q+woKJUyQXKOltQvdWzewm90T3i7i8iYrNNhzJOnLO8IP7zklUs0FemNqz2xUO1x
l99P0IfWVTfoqunkyE5ogZUkIlCeVKniNuOD2jTnRH/QpPG7vdl86EJ6YuUUWeoi
0d6F1Py3mJ5A7LdUL1Fe9PIg4s7Y+xy51/8q57szj8sU0Vepd2EUTpEITlRePOr4
K+Bim6bcoJ/Nm00mhDnze6koJS+hyZFp7CM1CfT2QJvp8ARUydyGP4gue6o1NCYI
1DeU664Ju1RQ/oGxT7WU82yJcf6zsjs8Z6mzYjnx229Y2njvyVbQuNpOMQFnQ79C
94Wbs2/rwfcxgOxiaZ3sSXfMA3dhI+ZPkrL1z7Ri1UdPC/qp4B4CnL/QHolpJ1vq
lVbjJuCX0IJeqt9EmevSCRi8RT5C9aw5EIN+jnOD4CsyvD4Zm9ylMaI3sKWfNpLk
dwZgcj7PINQ4rhZ4QDyDWF3dZuvlJxXqGDW7yFdfcX5bR7JiJT0+xyi6ydcSRH9R
+9gQA6A3DUx9I/wGV5A3hMevjft0lF7zz65CxizP38bnfiv9QqbmnN5yggTpWrcg
L+MbBDe9ZoOwuMNyJuHcMjxgQVuxZC69edAz9jIb8mnfZ+ewec1cSBdoAgkKHQ5i
SohqA637hZIuWYpj05RYCYE+DA1h9DHgUVUdDAx+CmUsvGzmruVcJOvLeEV/8Gcn
fa8SrnKOn89V3dMRk9ofaa+m68wpPukMIPca0svQO4hg5NVzDPs8ZYZ8ABBBDGK7
akTM8p6DlNDeJHXBFe5qXQBmq5HhQNSeBClomm5SlYPu1Lxcv53aRm19QwxGZ5Qb
oKORmB8m5YQcuSlAe/Yv2j8AttRZRAuVyzPFP19SDwIc4eZIXunrdTO1mOarzlPy
xwEVLFY0XINK5sO/TexrD9W8Rox5T3UetT4Z35I36PdbSotFlUFNoqEbUSSwAH/1
XRnGoPNyWYKnl7ni3sQ47Ym06yN0q9BR7y6BaJ7rxkHUetPwkeUZw2jBtGORPdUJ
h9xQ5tzYhqx36wFzbhDGEWU1zrLVsHkN8sxY56KLN9gXvWNWcARt+MJJGp1EGF6N
cZRaE2TB1dP+7I6J6XH/7iqxfq6pY2xwMyyXn6FIXT8ehGC5sIR1oqk5JyDgf+PN
jTyZpeuFLc5J+mG/7ahTxKNN+oq7Vt5ocXxw/KbDtslnLl0slvpmC4MhSQXmeElU
mONXa2gG5887nVYDMHDID3cZotX+/OfChvWSburO5zYUwF8Fk1BtbnMGGLou03ly
yRbNUXeDAo8unY1ua5jbqGzAHqxk/b3ic/p9mv3BDAnEftVewXx0sfKUexf/xSSU
yMUhHL7DojoLU29SP9yupucrnwwac7EyERupLPzAiMsoagubJ01xYnix1d3aJE1P
1VhKbCjfWRzmw3wTwFR3Ou2iGdtalVBwxD7z3I7n2vx7RuYXg0c2V5vspt4BA+EO
n/FcxAa+F+sUz2sIzunP2MWI1awQ1Qc405wmh8bda0WbFlypEdcf/ITXcESpELks
Y40d0amrLvGQrDMLBMV3p4Cs/TpLWwsv3lXsQ1cQXX2nwE8Ms830eMRuZOQiLqru
xzg1ngdWNRFzPacV/1yl3A==
`protect end_protected