`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
ddtXksX2+yylW5zu6QL2Lhnb2d1sD00763mmSITNX595NcHTEkwn0zB1Dry37fOW
FufOhVzEJp80NC5qZ/+F0Vk7Ik02dIR0elf3clrjeJRK85K4e3Hoo4xn7YbFUIms
l/8VZSb14+JVGURjfswrIyCUotIzlzVYZ6gzoZwDXIi5gQIBf/gI+KxNXPaKV+PQ
Ufys/12rjO6aI/pPlqSm0hCvftmBcnezN2hk1UeXgOIuKZnogjOsf0iJVX2aOOWE
6pD/psybjbnsNB6kH5uFTA5frkzIzkzl5d9+YDm9OyC+k84E83I/7/j+rk4L2dah
QJOvksSIzN867/4Qt8qYTQ==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="MvBXkzurAa5VTw+1JJ70nePUfoQXBvZOku/SMmg4TwQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
oRtzZL4VJ4iwysPsC8SXYCzXS8Fw2gtZTOskLcDV+1B9Nzn1zTyNtlo6lNICRmmK
ZRVu2BmCc2G+fmzynYlNTnSa7C0Cuel6FYpxCBlOuk3OF2tzAmLAuDyOH3Z1Yjzk
a0aHuoCdIRKv7BrZCdALt03JeUmXKPdOmIlkVGFl8yw=
`protect rights_digest_method = "sha256"
`protect end_toolblock="Jn9CQpRhJt4rnzZPRk+dOpzAubz7omckX1MrFd4p81o="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 6240 )
`protect data_block
gD6l00tciPUa6pDNTk/+t0OO0nC/UTtBwLB41d4inuAUA3i/ALrNyoJVcBnAmEQW
ptbcNp5fxEUJjnOxnedyZEuEBxWRieZFQnkRdF269oOfP2aM/XMhFuHWiUUt9mnd
s3UC++1L6YLEBlEGvMKCKb0SPxhqOxdg2G51bE/1kjzRvgWvETQTOkWYpw3hsg3t
7VXOCLo+4X+AI2FeIf8hDMfmo0rtp6T7lIXLzoHq1FjfGun4Ptdke4+Z+pMsfOuJ
1jMzU6FOdUX7St/rNVB9sR9bmJ/dPABjH5zk6wOhc9g7G62DZcSeGTOnYpC2WfhM
YoIYX7jQ3dckB/E/wo6/+tWKnQVL7ZnD2HKuwB0/3JSx3ugThS15rbDKgV1xtibY
QVe+cuUAR1BBJgeJlYOyybpOZW5vxtcvF3qZrREX5w9tVEYWqZIAClTnHgRXykxt
lDkfRmKdIO9vIJpWN/78hh+UdMou2c4Y+PfsPDSrPJG0wwPBXM1k0zAZYlhQaOKA
j/HcNM2f3NtBvQXx+aC7FqNQDGQCd5zhu64Y0mx3iGK9HnxKfHrhnXaJnjVPuZVR
KC/DK/U/JZnwvNPntng5WRAX3vDY2EuV278fgbpzRb3hfJ6vtRMOhCPzrdoH+grj
FBZ8QjksL41x6byrgyVobOItbAWO6HLdJi1kwo7jP57wp7hTzPbwm0Gvpv4mUh4e
aUsjwqGy1oleifNJPGN1kpZts44+WRkaf0f1SsgT3jj177KrT6UVlrRjt/RaD0di
gGeEClm5xbeWMhyN0Q3w4jamquhAf6PwZvIvr2/oN9WO8CQy5HaCFQaN4u8F3dZp
er5Ec+9oif5CV9iT2CV8xdOmlk/AXSMpeo0g8G5NW6aiucZ1j3IFg8ojtXEcb0BS
+Ba23isMvZFZa/CREORd5iOz3B0Sh2o082DmcyPZDBjAzjQxdYIJXq3QFbvCaoKl
URK22R0pixe3cdPTLxuqMC7y4+mMwmiVqzco48Oe+wtof0IXHLvETJbys6AOrqz/
emYZ/JOd5t6oXB6mqDMVRsxkWpjORpT1L77ACZ45l2Ck1mXeTwQ59S+9qiuegECC
p5lJz0iUJRJ46Czmqfxs6fbrW4y7pbaGDTV4+gWDsT3CJPznAotvnxbcABs41jO8
o0tqB8d/ocIN/KzocUIEGxbA6pq6EP/tfzxGSWe377HIQ2xVpeDBQiYoP/7oveIO
x3731RgIghlP2lD0gnYrwJTrf1fAvdAoGcTpaE9dNDzDMzpW4yADIV4qj8eCWXya
RzM2ndn31pU4TpWndgPKivsxFeT/9k8jeLIVf3GVibsAk2LK+Pi4/S6JO/RhaO20
x+7XqDvGr8bzOVoOSCBBkoZS1ChDkjBsoaOu7TMluaNJmuhoZN5b7s7lKxPvzCUh
Rnrw3ij7tBZjM39HIqk3YACiw+KtTmBcPPNu6ojFfZJ6EHSZqRt+eLBprmi9cef0
L9wezYejLajQ9JjbKnzKV+4Eb/OhGOOsemz7mkcAojrlYtF/n3OcPiqiLQRQ4C4S
RZ5lVfxzqTF2125MMoHG+f7Ai0xTVAMb8+TiKhegwccKmc7MdkNENf8vV9fcXYkC
t1vFgxgziR16v1ndH92S6Y/N7YGsdSzgv+TWCTYnrFzYOB53gVjrsKeG/HqZBrCI
DTNwPtP1zF7rjqAH2x6Ad7W5rtJMT2RLrQa/XmCbb8j8zHVbmdtbH87z9/IwFhZ+
2GrBh3PvRZSlR2F7TtOBozizh2YXz6N6XaiTU9W8OeqOhsZg6cWGJOfRrqTbaWRp
7W63qlD6XJkgGT9pYp2+JD5VyP/buLCR9BKpS75K3V/aSYg/77OejnTshXUUnEgy
+OvWTGY/o81Ea+odOguvaAdtFMB9o9+aYtpqnMI49mOXZeDT1fDH/8VSVDmU6Meg
3kqSWS+DonHvknPTp3VR5/K/BKRLjFBRl89IMfiyDtKc1e0Rc7/MWCO5ytfMmhwH
jUWt4iCrtkavpxTprI2z7AxlAye/GPNcDTI99WWFHwWTAG9TqywY+Q9cmfkPJ6cZ
VWYJg3VqcMATwgYOqgR7nofwmwIh740bjoM+3HmpiY0OoREHIMMouU2fLVPKuuTA
6ruMLnCB5E3j1/PumPsN8LTgiflbMYQjGpHvUzOm9Ex0tuzLifA/qNwQPcbhRR1+
F3qI3uh5mXclnIZK4+rcSRQunonnU6FXvTFwTAm0UEMj40t0u7xm8oe3bptHk9s2
PJSTDy/AullHJJ7EZ3cHuM6hXIDNMg79OD8u6CEYSiH6Mw7NkJTP0c1E0Apzyc1s
Z1TxAA3Tr8kv7Pv8kx/1oYmzZmITLbOCJsvbcfUO7Vv1VY1BsIkmNlDCn59NJqlu
amGwwfhYdTnFzINAcHHn55acobM2PW9irdqoXjDsW33jk/Xdgu2Brw2miQHyUdqo
ZyD3i91LVp231c41XEzxhHRfgdPX8wj8TIakyy7zhD9Yx8oPmk1NenJzc/wzJMpZ
ZEBPUx1m56KeIbjA1MdktXl6p+qOFCZyNkFYbGGBK6PqgFgYaCJgeVITUkJcVpTx
sqWmj6iBi4VGaJ+uvkBXxcLrc795un8hXbEjGJDZLQv9k9l1Qv2wWH+pnryNJmV7
rA069por0h9FjTgBLYtG4uVo5jQ3o9fkQGeYlLh3s587KfvNXl8+WJfATxuWcZK0
bVE2CSlgCVvL5gNBeHTxBb+hrV7ba+DlMbnb4ADEJJ7SntEHQ4Q51PZyMd4u+AsK
YhLHEeVDmOJ+73H2JDTkZSaO1k7czPQITWK6QdeSqo+3p/DfnfEhVaE5vh/Sji1w
Oaw7bY/rpvtKIt7HYyNwn3tpp97+mDk2n/crxXzkhpvnGRFovHeGYPBX3G1IP5gN
ymfsAKrvTL3H2P/1KOtS3T7YrZgEB8DQPKW/+ZxefV3zq7+t8wee9+9an+kbOYXS
DJEQqBBxG/pKhsg3m6uWaTVbRMjloEfP6Yy7HwIiDJiUtI/wlTNyrbX5etUejY+W
6aB/IBvD/PAnbeAEcsHG2xDnfe+yBAOamPO8Ql0fpaULrwSLbOitlaIFvBe11JHd
jzFoM6ZtfvZucjRDFlxo+1fAuPwgh7He6EItLp9Q80dYQ9FXHAKoi0GUo5HdzMCt
JxlRbpLTU+okLBvrlcf4U41+JG1Q4buGsQLsMQu6AlXm2aJSkUPckm2X9m4nepVq
UTFD+dNnr/kdtHkQe1hSMSDlUfP5U06NuVK4oCz+ocFxm40FvNsoEkmElKGXAXed
mPTK/FChwAouWXz8moOewzqzCqVoV+rhHgK2/25DPDuakp+5pPrLnYHjn/bQyxxB
3QSbxbHM03xf6JR39UkDYdbtbJeJswhgtmzgOHYDV3v8TEwvC6SALX6BaUTRj9QL
M4GEmIV0etf6t4Sgpaa9KoluZI0PKdcngdcXqrVotziS6xWeXYDq3tm/SgRWD9cu
3BG5n8QMO0A2lcxe8Ys94JpcyIkOooSo/ZxtCazWQ7oEnJjZz6C9ro8VyIGvRrGN
UCJnGjET/RWH8syVR+4YvRZZNa9jOuMR+htObpywZ79n1p8/I+TDIW0/IUS0jlGp
B6sU7nJlvLtoF+24zTukK5ZrVBgiQitNc00MPYoVnyhXXDfZxvt+kQ1E/cLmHvi6
DjI2ZFBoDZ7C86bCE+CE5Defqncrob23i+0uA/yaFx6mA0tw1QKudhyqv9ogPzsG
k7OVSIxrSylxH1iYUjBDJkj81B4DSp5TqCJMB79Zl0abgS160KVozgllKz2rJMMI
4jq1Wrz1x/L0K4C0JuBogmmZcZ+GFvYTuLe1xbdJf7Fsxf6ZX/A5kLblImbddw42
FpEoAJSTgvEvxOEn8oxnaGzFc4if92FUW4CG0TqhVaNU1vSBwedYfqkbltwKxlgE
fiM7JBA3MsXoPXde/J+vUZR9ZkBrPUHGMYjVXT2TC4Owpgbna6Ac0y6163QNsmiQ
PZlbusiPc9SzpLDlFoNqclt8ozUbkKMLppOdE32/G25nfns5AGu3rW9roPhP9qq0
m+gSsjcpatDkBwaDxCj7TspbnlX7tRtaEAIae9rAPToaA0vhWprA9U9A9SpgN/ZB
X3BWuxALktPzpsCOv6mvdjJLmCQQMuWZHmRnKnlbrXXNf6+oExJ16OvtaT3jbMIu
xrtm6Ji8Z6JM7bpscz/uPxvzhqn5LsYl1KBmzj+hZNxSOiEew8onyA2V7PFAh3OI
Jv7S6UvMm0Y+AjgKFBBmFSQwbul5LOXxBAm/Gk4g6TvLC9mjIqNa1WlXtgK8uy5b
/2009f00f00Jrp4Jlfh8kxzJpuikAV88/kgeC6eoR24YRN6taWzYwXWVbai/C9nF
zdALCDrbr6129JOwmNNY+8Nt0sM1G2jPBqM9yhJMuw2p6DKNizyEaPt9K4SyhOn5
pyMoXyk6R+ZWcQC60pBRjuXb4N33dX4bVPlVcc+0xDqkhhqDs9p0G+AhNZcKKzIM
MqNNYEhmqn5y48+xsUyhDGuVVSGMwSuM84eT5KUb5Qbw8uxZE/pZcqxnN6HU4fj4
YwJ/dSZMfyUyqscaH5xKTv06WkOOYIY5bZTV38jdmy4v70DG6tvRi3j5CkYCvyn9
vWKmDeb6rk3DSJ5VbzaFXCE8rsMMfZ/OPn+vKgYmwat6/2o4acvt2QG6/Z24LEmg
+cXAikqNL7Sq/WT0SnmBOZeVtD4U0myeczgDELggGv9TZ2fV4unT6fzWobxd0rae
oSuDRM09HqIRK5h4S9BThteYFl89YtgKmYCmvJsOp7mb7p4Da9WQNSA8YS+3XboS
9kt9CFEEUSzERzOPDe5XU7xDZnGAbwMaD+dcdZ7jOhdxvE+XCN4WRAzWpiOVpBET
+A71jzXgM7T0Da8P+72YS2RoQagTZqT4yYeLAt/btKc+ahaxbmcBlOPh+nJFusun
Vb9dRPqUMbENz1iNID4benolmTdyS/pgS2GrXt0AdlH3T38leJMXkKjSgV3jFQJa
RTe2Pm16WOte8e9d4xMO8YFpmMKp2QuIrlu0VZbp+jgHtpF8/0WfNgVlOttmWw1v
yEGVrW2uswoD+6lMaETJdV1n7+xGTBuf1X26a64dxBma5fy0Zfn7TBuuJM/HKGjH
Oxk5/TM+pvnu/OLxkxw2I4z8U7KGFTbVmYu06i+BBCGNwd5QPxgJMYJ3B4i1L9wo
k2zzeVip7W5F+CCfvMJRYBhjYpbcZvT9V0tshZq18qgCJOwtpO2osAirVUG8YACF
b3ZCk06zZ0AxXTliEUQRrF4TalYqRJHl/AedWWZcOQUyUeYuFnsrbPOOm3FRIIrh
GarRsDT8bz0wuuhV1q4XHf+lLWb+VEZLcCGv25V06ihK2DbcVlmyobXG34RRwk90
ah23qrVvnTRUUROO4O3BisD7klvbbDMtc35WQENgYewPigW24Yp0fvxGptxh00cg
CCYYjTEADDcJMgezmoXeGD4BIdr6wl/gzZ4f8XmSwxGgivZkw7ckgAVkgIh4/4uw
0kBKd/iHc29zL25AJBI76agcIzPgQlfqyHtsAO1qiJj+2iT8sMW3fWd1t7jlruRS
8Uisd2p42ZXGplgGk8ZquzUJi875DqzmHfcBC/I7T2okpoTQyGVj/SukvMOpsq1y
Jwvn5Fr4Ou5MurvtjILdxaL9zHTar0L7vaBbWG5LoJ9MvHYUZsDsPDgZTUirScBS
He4xa1LV+h6oXsIctkjYf7G6H4Ljs4tpFBtZ6mA9U1y9/3Qi1+lAiOAONBfZztNz
nokiMwPH6rcvpUowpQd1u6aDChCtLfEHL2pFtFEI3M6TClL21/Fa9dgqYDvrR4Cd
dkPOYKHccEiddMdnTyMGGX1gnlGCZCDQZNI6tuw2ZjkHKH10c658Cd8uBasR0f4h
pf0PHapyu5Kb6OxD1+8zJP/4oQbGtI7pG+zMKCaejr3O7SMOBYy1zTqRe7aSKMSD
d30TLMguwRI9AuONl40KrmCahZOq1HMDTjYBfzK+kXe5g3KUoajLAIEN70hcF1Fg
/x3NL4t6ZDU5pSlDtJ6fdetKVLMxZgYHSFGr/4fulWhX+DzV3SaEqL7PMima4/kP
ZxxzAGNOGMRQumM0r0An3eVQ/YM5uIurwguVQRl14o6IXG95p7dbxoc8EP9A1twa
eF6yq77CUyqBbSbIy0+4NhMKWFeknaKwNJVXIyQBixIOzj2wpOXueE/RQtha8emE
JwRWkdY4l8oGoJWKqz1M7awTmph02Cky2VsHqHQcnCuzviusk5hnAEFLSJE1O1Nf
aiVBl/cGxhtow4nsckfQCfcIpTTZNjBIfoZHipXWOehL7gNfUj4BS9txDPxutTu7
kstKiRB0Tx3ZkD/vKnZJc3MNU65C34IXISq96gYyl52CsEPcL8wXhME0qx2IVaGC
DA3x3q5INP/8rQKdxELfL6WDGt1RyRO2mHuoABrxSKPdodymgt+tZOTvj+sOOTU0
7V1N3WrVlDhN2caGeLglpaEAE5S9URjscOprSKLa/9IYE76xRnCKPi25poonCGlD
S7VX9aK4D8iTL1ethkttaSu9NQJasROZ1o5kHwkwFeU4/JMnHacPkL5/BYEQdcVz
ZSC8SDVvH8zxP548szH7RUGujZsOaPbb7tGmDGKsOOhnwtIr5igbjn+PZFkMQj0C
tyFpmbINAguSR9s4yC+XTic9bo7Dwre8ctV8rOP+hOdP0DmgM/RLFAD1/uhFc7iL
2c847Bi4PdMBjq50cmwiDOQlasMMgYtd8ZstEmci03XdA8TFQ4DtDw2ESGosYW/x
FZKRQkkaW66DdJjsFaJhJRC+kbrH2lJyzWuBbobcueKSckO+VmT4yqHc0iv3UJ0U
h5HbB1HGBsXPMdQR/1lm5Ndrfusxl1VK1lw0DzuCSsgVgoAEHQxKYaIEXztIFTCg
zbjRwlh2wNKWoEcu1RcatkZaKlzOWm/YtxBpMS0vwx3wGrJyMpeGX8+Ck9LlZDrr
XHg8PEXT9NzYhBkZt4Pmps4KOI6sLKDqKoh2BNh+VM18QMVKAy1wLh6Vint+Q8ns
B1Hy1pE3sY7+hQVJ6D5f7/cn1IM7uoPgMPo4GdUtvRg+QpOS+wyhHvmMj6B39t0T
WOkAtkBThjATAId64CTnB7Vb4GfNCpMjZKCUen9vSfZbJ8Tx2+P1RASf3120xAiU
d1pn4ytU30Dv0XgDZm/wQpvlIsgNe2nOHjcYCpjRe7JTgd5FpEg3ktLFQhKrR3CN
XuIC6x6QZ4QjYOk+0MoXJ93Wm0r8ZWcuIfpXr48c8malhrKX/32sh9Flytt15MgW
ysFMT/Hyqn5rjzNq26Fv+rC2MA0jIBQyJv1X44qhND7Qr+zM0q4p4zywLABrV03L
0LyEMWRcgjd2kT81QMDXMIh0BCQVFJQlKh0Sm57N0qpqxTy1GVqlSdMkmlEjbV/C
dtCxVLHqQAk+CgD8R5KYcaWHASm7sPPPwkVZWj7UR2miQL+CHPopV9LKc/GMIefX
J80FWoL/50pIcu6Iz5cwJsgdqGmOTiRkujOpUUmnDxFLeUbUSHPouk0cKNgweNYg
beQxnaW5YTX/GsLAM9xf0OKbR9WgdSTL5vWKaXMmAXQ+BS8iW5IT1wcJpQUf/Wzz
r20I6lUs2R88MTTz7OeZGjQrOhu64DQD/XXVeeGs4t+5jMj2SFudsskB6abZ/Hj5
95QV905mLBy3Pug/rI7Ker1W4oSP73RBNAiFkmAX8mws0cvhSC/t7DsQ+08aAv1A
DrYIjlDikEW/si6QH11ccaiStUenrRR8edSlJtdJwMWjXQWyf4QBFvac/tKr7n9R
R7C55+Umj1SqYrqdfeCM0NjrSZYuF/3wkLjPUPz35HMZvLMoqtg84r2cWSo4GrGI
ukiSqRoslETEjx/Qw4WVmK3AYgicmyfs6ijPvQVcjtU+VQDdLCM3V7oLs6c+uYi3
0EITFpA3OrKWY8NADBnEL2Wmz8AbJMDXyiFjy2+UpKtEI0PM0bQiT1n7UbdbPqnh
yPvChbW18FC85Y+zhwXmUFLpPvbCFPPgWdV8zrd9TP6xYqFJv2TXy3hjx6J50MA7
Da45+MWjpZMsCqGzzdpDy3Nz4bOPpHs/UlZyiw8P05DSUXuCJWf09lpiGhsDFRCT
c6WKs1q7iVEg12EqI6A90LVxp18s+Z6Q9VNFlqLWxWo3+QwA9/eyvPdfkSRZ7cXk
SD4teLIXw+Y298zVIMzEbAJ5J1b0ccUB6fg5Z/684D/+ZgGT0e67/hE3Fg3sEB48
S7ViFg83oO4TzrzLJISOhiaDEzkXnWWovj99MUyp+okiPoES6i4pPgSDuWzZTUyD
`protect end_protected