`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
ddtXksX2+yylW5zu6QL2Lhnb2d1sD00763mmSITNX595NcHTEkwn0zB1Dry37fOW
FufOhVzEJp80NC5qZ/+F0Vk7Ik02dIR0elf3clrjeJRK85K4e3Hoo4xn7YbFUIms
l/8VZSb14+JVGURjfswrIyCUotIzlzVYZ6gzoZwDXIi5gQIBf/gI+KxNXPaKV+PQ
Ufys/12rjO6aI/pPlqSm0hCvftmBcnezN2hk1UeXgOIuKZnogjOsf0iJVX2aOOWE
6pD/psybjbnsNB6kH5uFTA5frkzIzkzl5d9+YDm9OyC+k84E83I/7/j+rk4L2dah
QJOvksSIzN867/4Qt8qYTQ==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="MvBXkzurAa5VTw+1JJ70nePUfoQXBvZOku/SMmg4TwQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
oRtzZL4VJ4iwysPsC8SXYCzXS8Fw2gtZTOskLcDV+1B9Nzn1zTyNtlo6lNICRmmK
ZRVu2BmCc2G+fmzynYlNTnSa7C0Cuel6FYpxCBlOuk3OF2tzAmLAuDyOH3Z1Yjzk
a0aHuoCdIRKv7BrZCdALt03JeUmXKPdOmIlkVGFl8yw=
`protect rights_digest_method = "sha256"
`protect end_toolblock="Jn9CQpRhJt4rnzZPRk+dOpzAubz7omckX1MrFd4p81o="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 16608 )
`protect data_block
gD6l00tciPUa6pDNTk/+t0OO0nC/UTtBwLB41d4inuAUA3i/ALrNyoJVcBnAmEQW
ptbcNp5fxEUJjnOxnedyZEuEBxWRieZFQnkRdF269oMbRti8qxpwa7NNmhA8d4gk
LwK4JHGD7Jvw8Slp956GhBlsJqpdcSkzsgaWHntgZh8shlrWz/xn9YTP7vmzbPRT
M0CKFPbc+WfXhDdzBB/9dsEgZ4lUXvjqff0N4mTX7scKib160oFU0auxy/dCsv75
lFkacIXRG3+qfyWQ4v89ntiiKrpkXHCtSRGavDGM3adWNXpkancOx1yI/nQyG5Qh
sAYKvCC3wx4y0+0sAlHxityp5kKLsmY44Q7rO6+Z5oWG+QrsucJ4K2lDbyujWV90
4yecAjKUijFuYTXzAIA2JtG6bCJaiYOZdvhWJVUkREZKgXtamaluxsxdgs0OZD5Q
AS/A+wLwi32MmHaZ37mP36CAtyTD8jTZ5nEIkSEtopTVRl5P8Bxipq1Mo1jDr3gn
Rq82pNWCMZoQWmPVROosVmIlWh2sByr/XimJWoGvkv9hsy8Kjg7QhwvaVJfm1BAz
xG1y3ovzJa7VNtPpVpJNF4LGWQMCJNmyft0GnEMGJizcxnmxjqVjR1vsnzek2bRo
Eb7LDVgVc+6/pylodos58RUzSufSU7gWZB3Q9HoiULUVwsMydZuchkeK/oH3MJ1M
osWnRBpXbJHcV6Ta9SzEno+ePGcA1RimsvJ+xdo76O6u9/LKD5DjAZxkeqlv7qKk
QFFMOhOnsOVs2Z3nrXFJHoTVr+OIneYbARuUkYWQJvt3JAPX2KZMOAL2jy5VjW89
BciJmSl7Cl+4zVAk/Jcvx0ZzpgXdMKItCggjwbxS+NcVs8psF3PBF+03ucpaSLxo
nwlJlI/65NY9YnP4zlNDGYU+H+VSyXRbba2JLGKL3f7arj4pDbmoZx+tMbLTp5EA
nxkG10f2kfG2+G+RlPdwa4xpoGV/yuleqC31lSAARkIh8HwT+PLSoMGljIbYi8cH
hEI0ZLC1VD5I/g6DfSCHqEJog/9cWlNxiYfKn847dEm4qsenLZeEMzNMw8zdgmdP
EWlWoxxfVNssMcMGmHZEY04iqMuItLgBWiF1tkbtdiPlahTWq67PsDOW0J3vSx7L
VYHz+ZJLpCPDrJnCPEQs/SXJXhxHwWz17gTSYYrf+XsBiJLvF5QDrWU0AvYLclWD
YTEr10HTvZlEYJ+LO2KyVuq1mPk3sCOxXF6nId9cVsIwCpFNZcOEZW4FWOhdyAp/
wt7UwwmpHLrb7pXbGMjBytNqFuFnfEoa/J/Wz7FiXG48g9MXScUSWuOuuVWXkwBF
F/VD+73Lky+G8mwbRNagewf7UUBj1mnvp3HIOmvZWi7RBYfKoS4Oj/FAiK13yRZ+
9hTPuijDnPU7otWtFbfbxYO7wCWVKi/7vRStK7w6bkM+Htu8cJAjmdh9K+D7M36I
RqtW+le3vcoP3+1Yfi4QF7tROnTwbeDEmTJwivvY2ZQD3vT3q7gvBldK24XNHaX9
Lq6dE0GC09fCiFLkA5BPf8dy0OgCG1NCIQz/UWhO4xmDl1KnkOL9/FIRXB92GHgK
VfqBtaZ5I+3pw5+SNgIyd6ff6kb1j3Gpvck4n5qjFPVOQIF5pzrQrgwDj21eMXqP
PF1782SKH9CJQwpFjkJUwB8y2z51FpmtIKOynw9zwK/dAZlDvmiIkQtS9FxA6E0V
DxmvckxIJ6TwJYKYU+xfRzMu2QVIxF6Ewyu1/U5BUiA07jL/pnLCh1q4q07f3IT6
y4V0nsVCyZQ9MTHCNN8b6KzfRBG2Z0XB6uxwBjQDuL2qMRlcl5H1cymc070/PDy3
Ctan+7TUUcaolA4V/grka6cjcaxPbTAA/udQjcngmbMUIckYaMPjW2+rudqi1HHv
4AUmtP+zcuBH5jDScmI3BCrOKF0/4wh3pWij1ZXkuVPsXKCIHxpLuURZ4n46MJzi
/l/9LKDXfFzrGl5OmAbXB8z/7ifxzxQmK+0q2gI2LBDr9jp1HmteFsiqr7vj3b+1
NM5aEMAj4jUIOmVYAlqScqBe3yDmnch6j1mlWnQommLz4VTrGP4UZVAeUF1LPnuY
A8VB80x3nWF/+nduLcX1y4fi4ite/KQJUzxvhrJTeF1KyjauU2Eg/HRoeDvttnIQ
Nuu76nu3VHmAzVX1CotIqiX75uKE968LCdTqlEa29+tC0KJ8EprQYd6YlshhVzzg
Yuz4+J4O/iAfOsmByP1mjdc6oee3Rgx/sUPUanCwuh55zGzuABEWspgvRZzLdJeO
AxXTFtwhgqAIMdvllr4TWkkhA2Dad6Qzms2oIAu+AFiwLDwRgZXPppKBJy36KkOs
R5rQNW3aHedz0rXG+0Lqxmx7V7w6iUgoySSGUDgozUHeG7cELf8CSKJLfO2XT8Vi
iHsCr5eye9tp3FT7enbDynyZNumROqO1U5fKc4LJthcxFpN//+F9EXxaplbHLpjb
ncIvy0J1yqKWN6etf8w7ApZXVOmgpKN4TYOrZ5YzV7gA1zZpg36yM/UwGiGk9fGd
4kWpYUvcGVQtJq8YMsOnvIhztYIUlEUlD6+EvgVzOPA5Sgw7Ji2S88Q5sqE2NzSz
jK+YSlztcdNEzrQaPoO3qs/GAjeXcY+8/nYpiq5MEGgH4Bq3LNP9DP9C8fqaOxRQ
L1lVQFHZBtlNeUyeCWIoeEohtmYcOfBFpnF0zkU2cawlccF81PxR7y8jb46vp1uk
vp6IyFPKXtgo3wNAscASdNgnX2xGL5ERyh4q4sK/xu3bkVUBJHnag2gA0A1lwIz2
H460P1/t8YVzFBYYa37rGhcxZNcnuCcmGScMHnWhXlQmJ63duDSrEy1YHK7KiXqT
4iUkXAUdM9cJiovPUH5TBNEfnj3M6N62XhkDikZcGsgKpcxj1HCOX2Y9QNQA/Y71
ccdqLmb7DlzZbrrK5b6nDM/zzEWW7E3iVHgGYTN49suKoQAXX0CdNfRNV4TjV6sz
bQTWszMZE+YTs3sSmnx/whvCW+TxG8B93n5B4jfH22i7l96drOgYtwDshxV8jVhc
4vJ2jIVZFKlghcgp7GFOdYZwLCa9sc3JiCbUy6Lp+ri8fTE3tVWbS0AMmZ03oVm7
BcRtRP/V4oSMAWWkNObBuuwUBKBROJnhEq3OEN7hR68nofCUriBdh0FXKsZB8vUt
CXUCRddb3XTVIfLNqCktHvDf/EJ5L1FcvbM5tXBtjTXrdtjF48r4P8GEupF91AE9
/jIYHqyyN9P7ookv+STkPXueXMDFg5q0xmRCRySQNdNzRUyS4aFvGP2LNNJwcl62
kBcabEFqrsJLyDC5e39UbIAbELkdY9T7g5MkqBpFfLdyQRPEibVOmhMuEvsNHW+U
Gy7XWpcd8BoGYoo/SL3eBGK/OEKg0OKOlFyUOHxwGmiMMXuGinzRrvNfu/I/SAmY
vbKN8AAKfbJqI3VDZ/YnSILJlJGx3L4DibuhyGznaxeq8PL1GRtk6rblExDpGUOF
8Y1eqvYk3ezkfouKDNWmdQXmjO2HNEkUIuUvVSuMJeYxfxcv4rvZubq3K05XUnkW
w9MpbjuHvTF3luz7i/IEDrG/apDSg6W0eH6hPThvp+s2k5fiEocpBtWpyyRHbSkf
NcxCkEmxUDB+e/iVyaewwKgKd6tCLWM9CS7qyp/vmj4jFDey4eQadJFRFokwFsUI
MNJOV84kPIxjoJOstvwCekEwALiwzy88JrhNGe/vPUK3OSxT+e0cxHaAkhV5DtRw
3NBPXjkYB8UT8pF6hD8qkHaQRMe/pfk2njNe3vbjeXT41vJ0LxmBEnWTsGTaUcCV
jlNi693GGW6CQu2odZFTXDxMMjQY/w8YkY1wo9ys41Hlpm3s1CZuqOmtJ8WOF5hK
R8oEXno86cliMX15ZizwZl5GzLs99oWum7bLuXKNuMubDHojQnpFJkwyzFE8UyrX
l2f9jtxb/qe9YZpML5QCgvf4pk1uyjuua6tVXaDku2XCY0QRYo4BQ7BpPXq8HmWI
5anOdnrqjEzdMp9g7/yM6ykVqNI4GT2VMCkU8A9lswMlC6nS9zvIAPqrqY4jKtU/
DsDTmdAeKrjybi+N5//DX3ZKDTlDy8V/J0tT5d6Ih/aLJJ5j66aHHA3AYPec4kJB
aZNQ5g0YCJLdGjc+3KOhqxD3idKEy6NiXNVQcvhgMoQqU/2O51TKsPftrC1r1KUY
5C5u7haUro0IkOPm7soWngh0LOPg1UtV9bbjsBNiVYDivF44NLB2bQA5lDbrl+W5
XoO8d+y2Eh9j1eKSupmt6FazW38SJyVGovn/7CZbGymvw6OzKP6DWkD0x7dohKiy
YzkdnruV8THGosSytEHM9zAWCtrJuxVMyJO9kWIf1WlzTnRALZrE/YIk9fgqWLTW
6oqeTn+a4lb5uZx9/nkXrw01bVSX/ltD2YY4131gcNbjtaQpFHLEbcMvK0ocn4Ag
O0c/xb4VaHpUclRAHRDrj+9YdTX9r8VuVX1Ar84tP4PmBBXjf6lVL3/N8KanxBYF
ceItg3sQFHD/70iiTJxUTD5pbpqbW6aTwTaowKQ/kqDf1ZA/7kwKVScLy1uNqYxw
ly2SIN69hq1dDyMKHcmsE3YGE6ES1j12qD40XjG1zZzkUzhZvmh+A0mAiApBEYK7
/00vta0mU4PyDb+YYKPhlxhMwsPUMbWSE2XDYJ0YdzEwGkNlMdbInwGSRCoSF+PP
a8PCcPn1KmGFMmW96FtK5BB5Jvzmx4uGLCXGFyTBn0ac4D+LcTnPcfuWeZA58/1b
9OG8s2nNjga4vPXP21h1lYDKMHVE5DBc6G1d3eWL0iM5g9b+VWpyqKLG1mohIS+i
JL5eLNVb9dShIHg2cWpZ9oL/ZQgHmk2ljWDJaxvj8GppArNCnOhO2vW2V3gFwimc
lnpBqohKVD1a8ZycLZDQUh7TlQe7AQlyMvfv1PQrK55dZboMfLbUvQRkeC7m65dj
Yg9z6aIcEDYtvz24m1aJ4zT5p15X6lD1mjuIq7h4O5TabimJ8lTogH9+5JUYqCOH
+62R//k800VsWv8gbTpd0IcAiP9yrnS0Ns/KGG6XPr1umaT9PMhQfQ3bPciDjlTn
H51gQ4dnQkHxmgBdIlqpPNJVcXIK7QKApMGadITrPyEF1UIx0OHxq7lSeSloULDK
11lseqqJamWyAL1+O1V+rZxWv9Ao8ph+fZ54pDRu3yxsTPL2uUgM2DBOT/0s7kZG
MejA8gXhMsSds6RKGF/9L+Ci0bwJOSnTzufYnU2aJtu7aV7ZGZL2Bj+EwLUCio8j
co8jbUC9kvS4rHB5OFf05KimUrctRdaQKwfhFXv+P8sAKITmYpRygciMKnoYqgbd
HuABeKMb8Kc+ALEV0sfgqB3Sl05ssHRm6MG+jllctYJbOvT7L6qlsHYlCMhW6S06
51OJXQCyCKmSQpbgycnagmJatXHnSNZrq+YUEJyoskbjbd1XZh0l0x5RNuBzGouH
G0gm+HAb6yili3+EMq2o8hJczKFQxVMmROl5RWetpkl+iGnc3hS5atlz4uznRjeW
v9dBcwIzfOJcKCHyCb6kDzbvL4lxRMY3XVGbhW54ppl76aOV5T2UUG3a6W1VEaUD
O11eVqq7r0hnWXxycUXyWTC5r3+dFB2oh41SYZNjarZM25/+YdqO0CyfuZJZW6Vb
13gW/KqOcqBKs75SF12rQNIYqOy/DB8v2FMhgr774dd8ywB2xUdgrwZHAibLIx9O
q5/Ts7B0MmciPthz14GOVoLSSMrjyFCjDHPVxhMHJqFdJ0a0d6JeBl9pfg/sqq0n
3svcu1VpWd/VmVDuteEQvEz3v26uReiSQsZtIDf6tCIG6dqpd/+5heozLfQ4vpWI
lP65s4+7RRwgR8LSFA7QVv9+TcXZJ6ZZFptzODuhTjCEQLQVRmT9UqmnR3v1zycs
sh76TVbV0tbStOEDouZX3i8LnNX0t3p2AwnVle87WUl7flTVUO9eDVrlOeAy3VGK
5kELyy6sDLdKT0hX05kg1RFVuaFYtvxFKOBu8lwv+suHFr4zdXuX76KxT6COOETn
eW/BhJRVB+Z7rpHQ0fgKATroZHjmUSni4pPdKKoV8fExLCgALimKAkp+Nhy+e5jy
9Z5OdaFxLehVVW+vwWeQrqLb4HR+7GabU3yE3auQnyGpNxoVVKGCfBl6du1ple6Y
XxHJ7zL4RxIrzwquhoCE+983a56j5I+dFR9Eg+O/kN2xsHdR2IjjMcF9YZkAoC74
/U3+0FL7sp/cLhHevF93pUBIWFcwrO3RBY5DPJrSNcYuZrrnMuOwk/X4Tdk/K/EO
jKN4AhO5/27kNZP/BxUmSMNrN5SPPMDkT6M00r0d33wH5DFTOtXAJXNWc/ymK++c
SMZLmA8Ql+LVbZGJZV116FG6yRggOEKiQOYpvG3VftHq2MwsqwwiLbRqNdN178B7
62UY4JourCuyWgFkGiBuLnpVt8lRBBUJ5jff56Qez50MOBfTordfNH4e4XaoxAhA
uwUKsyRI6HtCNQS7zyuWe14HZK4OXOwoIipfbfodaRPeuPd+aDkp88dVoinmC1UK
SSg9xHZA1DenJ6cIXnjz4sk4YOGNz+YO/T1qkfqHs3CjIKUHDtbSN/MxzYlqUTbA
ac/ixdH/cxuVvaUZVUlz/mRqiORCxg4IFVUTX2BJZTOdvN7JtqiA7tzdvNnb1g1N
7pB/t/lVHojAEFIX+dn1mF/arH5e/UidhirL2RII2yA4s2m/SoF/xyvQKIVkIVwd
hncpv/AT/6nqHbVex/VVdvhLWPA9PwGHWY2rY7YC5iKo9zBPIuqH36yXe8WnBh/d
bsEK9M4wB8yApGLhsruXCGawAuyOYUTk4KTY21bAljUyy/nIzMbUoKNlEdd9ql9y
JeOEqBJQuK1J5fvKNr/OuNsL9YJGE2kPauKFIALbd4hQg4dGjrBwhbnSJtm9TJax
WbNgT5kUhVzddBum+33fi9PujtbjwPbUIJCgFz9CxJAH2zHqSxfjQwXZxSNNQamq
LgUIUXdtY6/iyqFZfaoIy8LCMr7StH39KVeAe7OTbgjeYTbUjCaM8X0jkhv62y73
TzujA9PklkfPstEu0/OyQnD6yNaNWjU5s8BL4QR1bVu0gT9f6q06Dpbvg6ElBMW0
XEYNKCYSkpg8gE6EpfNQ5c1oxNjh1JDdRezhT2mpfnRNWqAd978X0csQbE3aeAkU
7PY8l01BDArJGvMXHNScF57V6+Y9+gIUzUgol96ItNBHMXqBQ/SK+u0+NfJQalKJ
agO3JmTH7YzMmqpA/zQrREEz8//ueU0RxtK3JEEO6TBDRsK9l+M0dNZFS8Jqapd3
Z5X7JrBDGt0qq/MBWJegnSHwHPI259QDeh+54L3L/bcF5d5zNWiB3nvk+0VfA6VE
ZqgmLR19Yno1GqAJ2x48MJ9wEXXCpe/0NOQCEXQBd0ehbBPhx+KEB9URKjkNQpCx
tBkYj2tzossXxo40VH0v3lO8wdNixLD7/YJJEHkzFgeWVGqVp5bxaFB1H3P/B3Gu
uYMyRNhL52bFmt+u1vMLGME6cnGzb9nwG77iSnFLvjeZH6BUqiumF2cWaboffSsq
9JZmckjA/70SLWuCK6RtyWCor7HE6GK+oL49zuirm6gTQECpDxEhj+MZ4+DwhSm5
7nbl7gtUaVL6V+GrIsbwwKUPS6CR3tkPgUXOkp8RMojzJsKhDtZTPhOfvimNKFRH
Z1xhaxn8WL9k67d5R3oDfq0zCfOk3lYPp3UFzCHF5Yf9lD5O7nyjtw4FALKEvd6Y
JxI/u3aZzX4vH+w8NpSorHDj15gKDUZ0qSF6sZeG69BSSufcLt2K09jBlj9XZZ3d
bDNCiz8haOTnrycWrKcmaFgRHFsF/xk7TJl26FWHF1kptPkLTTmmUTrBNNbxN0uj
OzeX6cbfFVu0/mfZJYNXplv9GhAvYmEIjZTpYQKUwvxSfFMxWIFTgA7mPaJbs1x9
zNh8oz5AM3ZI235GL+BFBeT6xFzg2c6Onz0F+FsOEZ21uQaaDS4uT/RT7+V6A4XJ
ue96sVUFoCQ/nvUTx4P/I+OXY2Y76l38/MPLcyAr13M/yqIDhN2O9o6W2XVlnQwO
Mg6eajYAnmZIUhQeGB805/0UWXGILIamVkW13ry4g33QGGz/RRzSp1HrXHOG9WX5
R/CwN/GiI8ZwRtzaeSSC4RS4r1IyXi3grwwd/vGkUEOXuKvgIMIFzmuJZq1YTG59
TDAC1WU4bRBgyDyMHJM2JtuEdgiw0Hoqymwasz702sVoYxROZgvc8l8jzslrWlqo
pF59E3HTj9wfpZ+yK5teVtH8VyibkFE/yQT03kPcP7wYnjXaTs45BhYQPuFwzojk
PpThWaNLuLMALi35fqhNossi6dMAqfUY27yrPJbF0JqRQ2m90guVARApvAbYIqpL
7LXL5XcSG3N+fnVqGHzoTfQMN8bVp37scknd65lvTKLzVR0U8qm4jNpiserFpMpK
QIKJrxXqGlaIXDC5hB+PGXLkWWqKfUYQFd5vly9l4e8h30UYwSVlfQaJ0DO32Deb
UET8sZMsxCkehUciHaWLx3Wy4tU6ij8bo840zfRRBH/Xdkb7YDQfJ4OnYuw0Tvjt
v2uVGBx/kQWtRBlacSnHmhyRzL20g9pIKQmKCtEUiZIGrJN5UZP1XOmAjzLCU2Ks
vDwSYy6mBwbsV4My6/9bsrE6hZ+r4+87dzKEC5+nbUPWKEoK2yzJKqIL6i8VonRd
wCTtaTzk5FBgjMUgtjtMsGMtLNofWWyhrjYAfcqfJlml2liyBXl9zTey+Pzuyrdb
oHge3esUjCj+u42HQ8mFUndQc83i8P0shOkD83F618M19Emt1i3oy99gAr4rm/CS
yFDvvbe+SKyCpKerxdvRlTzBNLyvLx2fjyl5IKoNdoZQZMQMy11WFzt8soh5M/vL
buTaLaHE+ZOnpGll+7aUc0XILQCoVtG3oK7DVVw5eDkN519x9peY/wnVS+iyj1I4
/B7GiE1m8XhqXMzl2+JhxgveUmMBHW7A8eCxNuMJBaiUYHYN5inekODjAcjlCirC
a3//q78V6HbxCajh8EbBLeVknFQ4rg7G6kGP/+BTFrb9cov04I9dTGFAYDxSo3mV
IRYtSMDOxnWKvT//B2z/fcy14fbpoTuWk3bPh8sgejcs3m98WNKAhCflZjv/dIMt
UvKbLp7DoXA9HavfocVsHiU/JaNbYEIBUTWSZbxfOPWEc4Q9/IBm4Zl5svUgXPq4
i6efUQo8GFnlJhoADDlgFaiEFrGRnTteMibr8Cze3e/zHQ1qJPby5lBMrdi+ne6A
Jpq4DABF7nifVthhzpUjRftbT8M2o2Habi1wNThLJZc2QH0EFzEES83iyLZixj5+
c0ngdOYrp/7AyM/60fXdiP38M98F9mY9de3ywB6Q8Ibu9ozABGVmtGBUwlTwGjZy
YJmG40TuV80LdUhHcODLEccUlulfXpAwQmnG4t/SDpnX+ugNigPsL1DPHAfwaGYE
aWAqfnheMQsM/9iU5gO2N5bNWyhFqfW52PfF47DuAQwxW896p57FjO+OO6ZLmsEW
UmC+uEN5FITq9kLqFILZLB8A4sbQr1GtVDb86FsT1/BMK0N5T7Ayre61G8mj+kF2
Tpd+V/iO6xMHAumWF7vbr2s8neQ4kgCItryA3O3e5v8rvAM9YLM/LxJRIhuA0++G
Zf3rvWSHQX/2iO/S9kuPtdHniNrRRFb0MqLWH90RG9PIjA2wjCHhbbwcHJW5ue8F
ceTSax+KoK9Fnp5+ZB34OXuBc0nAeACu11oMwD8baPjTQpeRtu6EvYvatjK0UBjB
j9Xj1kAxXuzA7EuXdXoLh91h5fehm1Jv+D8koP3VbzWxZ4uwDTj3cLTQ8cZBdPd0
fUHlRbDOlzGY1j4wi6BBwvaE9QcZEalaFLWiu51rqs0zC9TPd7+Kw5SLNKf02fP5
E+kJd0GuqdE4MwrOcHXANoJUTtFrH8bqW8mhnEh/wiihCGr6cm6niYzzTPDvGwjD
qK7YBHhLvPbuWyPOTVifUWxB1jZ4JB/yQCkB+s2BdnqFuVB95T7gA1kh5gxJHMx4
r9Lg303y5NiXk4/pKVs5sijArUU0BIERGr/1z84aynDZpL9Zw6QDtkZl8ZH3MHCw
9p6kqBLmSp6V2cbHF2I+cWwH7Y1swh/zsQJGt7c6bqobugCsKYs76CQBzD8dRL7A
Msd6pcvAGotEc5aqSC5CHM3GxeR4NDoQq+vUOIDKD0eKnpc8AbgVUsdaRIfi3Cr0
IliybWpyrCdYwbYDwmqu75GW8K3qw9KVFGpTosNVnCLZO+YgO6LWhzmG24dYSqOP
fdwRcnsZewCArSowBRno0zzChNrucjNaOZEevzGZm27mV8m4Hid/Zca1oWmijBkb
Cn4BSUodSLbxjT5rgf+F099JcCzWFOnItSvEjsWFtoab4AgwA/VVrrEuW7UePwGz
5X27q/26Aes/6vN+PpXT6udZvZ+4PUl/1YaPdEglWNrRHESsy2raeORw9ZrX5fWW
sU8MP0WmDCWMh+kzG0vMDS2vRDNTe/e+TULyVW1cX4GSjPQi1cve3aIbJG/yU5Qn
Y0OfpbHuEQuZdHRAzyXzKnOVdv2Aa6vthIZDAqoyqw49Ij2Ege5oQiQ5/4BhwkR6
pm0ySWULESGiNgO5V9ccJdzU5fISfZo3w/1qKs3I6ITVehsotOkH2+vDlOA/oxhJ
Yu3Z3vPGIfWQMH7xOjWe/fMhEURjRZbNar4tQGHX1fceDRKTpsZ10/+lqZXmWlMM
X1ZyjfdnjoHJWoyXclaFBYhShiKM4NmyHYMByG27r19d7rWRQjJFkFRzzSEq17sE
ClUKsGAO7hKVjB6DmUlHKr/J0i4SmiOz6Qw4bYnvtiNPD+pgbQ6NLHwRFYQEVDFW
dGkAVykVv+OnlgWwm/dHAn5j5y8E8UCpFvxkiPTR+gdeT4CAhDvrPj5Y73J/NKyD
9lg9cwT1SncG1Q/55V9+lJFm+RW7C3YaWRkrP/hjXJDTH1qAshk5aCeHKkfl7tXn
XQqEFDbiLbf2pono4NlUvtHKrJ+u+q/85CZCl7USGrcVjOKJHcXR0HDXY36nsBoz
atBSBBYYfic7V7XRsorSSKsQu0qT4W/kgUu5Tq2JHKSlK4yv9/wpO8ed6w5U2JEN
R+u+EeXNWOCMpNDgC84T1P+XU3oVpW7Hfspn3Hqzs6G+ZjusPqjiDoYfwcmi1Jmh
HLJ2Trw0akeLYyCF7iYDPLMRu4k1PWe6rPPZcnt/JDFsk/+SVrkqksZWqrUvrdaG
kDXXA4a4xw5n6XVKWZd/jg/SCh1GpGQOzWSGyD56yWnIcjP4dWZz8dmNw6vst1EF
iICeMToI5HQdCsLtLYfDjBKHAWYOZswBCZIFb+XxjjFjUXsIMQ1jj3V8aQ7N62iR
2t600gbnSL6LWja/qW90p60zZ3VhxwFIKkE4XZQp3gauCnC0e4kEhAdQs3lnzUjb
9CPqxDo4PEUDa11qJUwWFyuhLiVwZARUJq9GelQkLVY7f/CxSr3mpxbHxzBEXlsP
13b6KN1Z5LqIjllVkwfS/dUzFIR10tZ+oTJ/egCxOjv2HAz4EgLDrF0VorL4FRWv
c1QjXQAaUZJcfAyh2n3zIY9POaJW4uc15mQ70szRAwij1tDCKFxxIBU0cIwiJVFL
//AozNvdPX213clJdzJ2cD3CG34D978hUDEIsv1q7pjhsBzVCIeihXjvFJXzfu8Z
5AoF9cLgXs+GpwTihUXrZkcEZkzEKqGGd82NTEd/VKzuFToZ52ZUZVJAebAvntWk
te1BTNgMwI2bLx9Rt3JKY37GT6ZuhMWV0Vt9AHY9sal7Ue+uLvxnZjBACFlrw8R5
SbSDpeAHvqeoNAbsSAfS4mfKR9ZNpupZ7E0SbyEQnUncK6tuLoX93w3Kszm8W0Yl
sdwd6dvQCE8OnKsOziY718BJnCRQIoAozoJW1EAbET8D3RLio4pbMpxAByXyQZY0
EnwqyZDLkmzbYZSRndbcJmaoGtzh3JSIQt3YIKa3Y5vM64+e/hORWC+8FlfO+On9
R9Ma4lm7Xg40aByAVxCQ//udDlAzAuIjaPg/Vnt4VMYPtWaqnCdhbREVpM7TtJvw
bIsZV0Tx70r39+EFPn9xJYtBY2OrRpkK5xLiSdbqKmQm641jmkexIwJg7cEfbiFX
C9YHDi7BSWvisdFH3qLz/7AwyTQpHAD6myVmf1HSnsUIJsCioDpWrUR0UY2FfH8F
8CO79g+0lqiteJPs2028Q73nlUMA4q0poO4tgn5eVpheqjpGOlv8+n3ZMhDEmYvf
+J5690MbMpF268B/1yUzdASkDxeJ3iXihnjsGFKNBTAQlIYgVPSXz41AHq0sCbg+
MRm8eh8yJ3GJVvI4Jifq7p33LJM9SeItuSVsdoZGWNXPWSPKfpi9HqXP8b3hPUJP
J1SG3RBhgZoh+Pa0DcfqXfAEiSSzMKQZtLJI5talia42nCjxkiIZEpD8nAcFmFJ6
xNuGEygQholLJ6EpGLTSg6j37iNfICbjwGPEqfi8xvuWz7enHB6CfKp0eCj+4J6k
d2t4DNAB/o/ymjLeW4pquwJN4YroB7re/alKO+R4oUON5+hFR8sEeZKug3jqx29E
OtlZlT4a4YdJZqhWsy0Z14N74gi3iGrp69m92wISMgkVzkDDOpEbQa/hrqhKAugJ
bx1+yg+qlU20cbhvZrQKDkfavphzOiM+wrjZ/996tg4Y0hTUmhDfX0dKXU6ECYoF
yDWPu0VxGl3ayGebaRXNlUKARI87SWCrNATOeT9b5C1djs0Zhlom7piCD9b3k2xK
6nisJ1MMhbD2E4bDicObalbNKAniWFwcu8MDoxwUzu067zdqkeIa96q7BEY+2cL+
t9KxJmbVC5WvWDeSnS/dCUlIEil5aWRIkrpYBLjOIhLJtEI0WYwmwH1Ox0SO3LXN
wrmMo+e/6Q9EYEuQb+KTX1/faomBeXMH8HCgHKASzyAmmEATgoW43ijv2HvYuNNZ
wEgCObrcEeJc3hFBUiHvt2uWjr6+PxlBnPEP63rh90nYpCn9O93jZjoZjcmG/t/b
6O3hxQzB7HnOPfJFYOcdiQRvWEhFbDcIl4UtZ7NafIIlXP985Djf6uTpTvfQECUO
NmwMVktrXgDEY1AV04DvX6WAr8D6GI4Xa32L+q+5mRUywfvAp1bC81DOqGObvDhr
/bT3G8fgt1d+AM1rSxa5CoSQ+KnHizb9mwCa/aFm4dzVN6Bb0TrTJEsRyC4eCa75
EhhJwXbPXslHL1lVt+A2lz3Nw/EOZcmO1yYpH/aVWWBEfVBJCI1ym2JWOs2aSdgv
U1hxZ2M9uAfcyiPK+YhHTgiohsbgU20tw4n2HlM1nJSVlzoZtoWQ53SEkJdkWK+7
1yeiSNxbeRMymZoGIW/OZei7mOMWuWQ9tBflMKPHQkOB+QXpVqHTWX27JhRfGfYD
FPZIw7qtf014Mr6WvW03W27sOW8g7GD5BzYmy0ntjjBUx16n11nCKwboZwcisdxY
4WRqa9UplUlOBYXXTHIBK3/yyVU60ndsQkKRmiWyiXf99p7bmnNGBJH3lZLWO2x1
dpFdE/JUFHIavDfHxgyXdRbvuaeFLkS6HioCgGpyHT7QsMO5A/Lntm/q8pcUOUvF
P8e6PtloHrEk+HIX7p5CB0WhKLUzgUfWwYAXDW/533dOFc15U66uKEwQ6n4aWJ9y
OBYs2Ri0KooGqhWyZ6LFan7IGXUjEEbCGen8Kt0Wb//XfPc9v422YN80ILmcujRs
mtnYnpYcdhb4bkqDTxecDxxBKzEQZDiC6d7twwjyP9clxwLKb9sFBEcAt1iOGNDH
cqBPDRDqhZ8mPI09xbXx/6xsnsjMfCN5Y5w0y/UvUw92nwKtMKi8QG60nTKqaFkr
4LGtBB8m4rpvTRkY41TSl9pkEiXU5K5Ew2LLpH5UnzLA3HFdo7RiqdmKZlSLWt1N
m3zULZXlLqv5QdThrn6vg9xJ+W4LqFtYyoSPEjAJUuushVEPn+Rs8SDarZz80sXl
bE+WYL2WgADwnwVI7QGHzzxltPrQFxKm2IupRRhombsZmpXmlphrMi1s/ne6j7+d
NOTgxbvRNkAYtXh8/lF0+gvA7BqD+lFE69kJnlXUnWFeVDUAl8zCmkPlG2TlZQFa
bS/X2JLgtXjai9E1vBkeNVX2HzE1sSmXsvF/fphFeO5iGb73TGrsLWGi5cZ4ByJl
HvnnNXQNEHdnKN3QuvTq5ad8SihbeAA/OZdSOUbPMb6kBW13o4FVTBZq59rJu6et
zCJp07pdzqPZmb1athp9pdQq1Xg17Jp2kP8vuJCz/EEXg0OGLrCR/Ay8eWioRCR7
2znfZ335NF6+lwAaJwsBx1jT4yPOrTzC9m07ZfBQb2SXhZcm3UVLiu2aZVXK2A/u
chQoeKn8WvuY9FozXSC0HPwJSO6g0o6dWO1t+sqpIxCJKpomBbBBcCe6aYGcTqiK
xIeUNpEc2sYFH+wVO8UUC/VpW+a98fARkjxyhxoTVp7PmTivNjTPyKnEzsdegv60
VbJBRM68NLcroNRrgwDWCDbMcPaEOZ1HkRUbsSFtWPbznKYKGAlMQvlYbF87Z9Qz
y7eAVADn5zxULY1lnofuRX7vDmtny40IeN6y3r6LoCl1Bdf6zfhLfH2H3iC01f80
tls/p6ln0gwhBK8lIxj0moDzdDNY3n08OEciKrH6AmXd3QRPCCAtjnb38t1U8yiN
jcmpeMVYiSqODfo8/Uwx3SV0P3FlcJi7sfQlfZu2pkyKWmksLg3Ofnu6StWnPV0Y
+CVecyC1dGcUsjFDUHWTVCy1Rvgx6O388giWftRrimYOGghkD9UZMbS/BkIX1Uyy
57P3ax66SMA0SylHrNIamyhOclkgoDhAMZM1qaccWWIp1DvyPuQ2k+O0enHzul6x
FOZZdLz3YUTRBUzBNDsSimbcBeInKTyuCir6YG01BOcRYGweUHdsBqZLaGZqMK2u
rKC/w2t+dPi5q7+DYTFfXjfSInEHqEGLg53TbvembGKbPQMdVuzkjNIlaujxZFpM
La+Yph2MhTW4KFiPE8Zq5+Rk0iLFzaSmgZQuEylJ9D2RXK3etwLMnicDsJcXKxGd
7f2zD339siowMHC3lSHALSIxOZgJCnXDYBNa0gQIaLY4ezmJTDR8iq3iwf9Xh2MS
I1DvKthAf+a82z7SnkGW5Y1KI1rfmO99sN0vOq5jGWkmGj/WKAXpiMvroFRmBtTq
LxcUlynn4DbzRprU0zTZOxDZlAYElSL2m9zRiLxurCPhbMeiJRduKLh55SSP6LWY
j0ZoUBvnJ2CJ4+kFmrfynPRiTFlc9xr2tqMVP5Y+3mYZ9HdxEARX/yWgiDGiI/Dx
OwegMViZBhYsOoeGeXqBCcyN8luFYKZarSdmn4LJ0Xfzh9rtYEywGtQLaExY32dp
85q78LcPAmp6j3LwV1mpLQkvVGDWKKJ9mS73mmtn+FCZogtLXKztz+kPy2Sj8S5b
4CSsiL+JeQTrzJ8trRjN6CjKprjkwMAQvLQZMBtgab56hTaV81kxMjmwNioJ1Oau
fDkq2KrLzpa2Qce8/GT7l47LPitqKvzw/t4Tx2MttxN/AcEdrrvFOgRDWuXSqFb6
V5UEly/27vOja8C8yQFmX7SUJkIo6ECoOD8iq4peM3ohmPfRpO3gFHEuxz/HDwsI
PcZJwJAaTBrEbH8Ob/oQZm84qsfYcAGgjVXLr0+QRofE2FyQCXjXCCCFcqyhq+wg
+OwH2m9LkPTjNDoL729akKM7fCxFhiLLMDG/iZNjyZe94BpuDmVmOHlyds+hQ5lG
J3vTMqnIdhd8GkjpfqSd5OHMW+XE/OhnoNsDTRiXDQ4TsmxFFBq2sAg2xKYFWCek
yZvIZpXSE9H/OL0Ha5YGPzhl84sTiCLqAGp0+rX1nOetovz9mw9qrnGehfYRttiV
lCOBklyQl4OH2rg9AiL2fDCuWPa3gf7bNrDBXij34VswOBm/23edaff9p7LFL2Cf
8fjoAA14j4qvPCMdr+vJ5dKTj3OXMw3GuFFv/yppac2EzHPMGpX+3PUlr1/xSuW1
JgskV1uhrMPbhm9tEfygcGCSoNknalJ5adOW7alqv0Xs1W2eRChWqRa+r6PVVRVq
iTjaJwsxCSrVmpWalD9ETl17WtEsHqIsLZ9UIXWxtb9Nd0XqI2CgEQelb+etJabD
TcX5To7YGU+TyYa5QTcGNOtbDiJga6WM0cyDcdFg64QkuZRTJR1M181TPxzxBzeR
0NGYhhIMZ4JLdEKLQfrvhCranlemP7+1cLesvKZT0X+TqfxrDu13w2QyXM3k/8iu
0EksTWNlrG+j9KGs8XK8xO9D3LSs+SvOsMa+KGcHtufLtIRa/oMKbARuNgY1Uu0y
RxBUHpXzGRblyqQdQ25stExKMimC1ZIYKyhXo6EfeSEuvDaPxMmnO2Dy7zXoxEJC
BTzF2iD/hst/6Sbbsc9BbkACnm+moQ/b2pgxzJbofdjDio6djBm239lqVJGjJlep
UNaOhkriI6tqb2ORQzRv0TmyXAdeSdSHw+jk/0tdBSCUGHVKGWcE05ZlP2T6YpPD
ZeGb4lNUwop3KjYGHC/+1McLz2ZEkKgMfUULB//1YK0ojxqkBI7r1sNdMhi+BIH1
MA8Hy5DhekfITeC147G0ZRUOi+wEwotALkZi0dnF8pKnvtYFTlWj0Cq93apklcRw
mwF7AHv4Y351Jz/B8lePp1nuIRRJ//JdOOdlfOvG5DWo/2xiQFFkg/CeFkj4zhq7
GdX1NPjwN3zLL/LxK55ODXUJteNx8WFKhOv4Rz9GCLaiUgnb1wd2tt7Klt3xJiLO
2wTfG2+pVkeTevaShJPiEtuwLJ4AHB4RPokscfQrDF+l/6R0JVwls8a+/dmUuP1W
TUM+ASusRqvQCGbcObP459aBKea6JuphMTn9o5qvdGolV7JWbM+qJXXwQXHZxMVC
/32f5jZCNPYrUPnp8OhxPhl7zTAB1e6tG+JRfIvxx4Op42x782N1sg4EoB+h43Zp
WAGlIw+koN36KOypdiZhh/Np9c9NodLBJCp4/2eu8O9pUfWw1M6QNO9YvvUs9vQQ
KydrCsAv/yJtGEVPWC/nta9qCvMnjor9Xcmb53hAfFMNlLVG0REWF4Fm5l6U9Nv0
ii2XKr416wtAu9PkMzFJev3hsurWodPiu6qGr2Ao0SVk2IwdeotVgtI6mk3ZaGEP
cGOzktZW+UAYEun8YgGMt1LyR8BIgQLqdo/DWFhZzU6T8fOeorI0XknSduKtg48E
pvktw2HeA/hlOfO8TtcLvGDAuKxMdMvXI9KvgpZC7FxQiqR0h5xe4HMogAApipC+
SBlWkreQj1kCS8nmkvUUHIXb34vA9XNvGE/PH3okQuFy8bjEJcfkIKwCzYsBD0X9
N1fqKPpo1QCpdYtcedWfojpuMSJshH37iK3GxN0XYrX/iiud34wGnAFVbwt220Kp
Iz++qQk72XFDV4CGjAtHeAt/Bv3ro8T37mKAO84MPy+ZaGkUc+1rGNWMk9H2ZIA0
pKZss9pE9G7RtxMoCn1X799ykvycWD0NT/EGw3vglNFvQvYr/MbPl/7/y5HyUBFh
GXzAiOUlP1mZyfoUClcCn4i2MyrU+exUXJIxq1hontXA97+Ce6FOOl3TKL5ktH6H
4cusQLri0mGZ54FR24fujShNyxNgAOEWBjHRai0SmUqddl4mhBg7/Cukk7VXlPmr
3xUc2rK1YB+A1DI2sN0HNoeG/8xjvp0XUL3tK7ZQqt+LVrMRCHNzEW9cgwKSfmRP
v2fPHjmaUebWDyJIK2VmZEFfEH2cRGAsMj6aAFNTbmFfOkj5AMOiR+HFy259maAF
YzdPR8Amhx36Cosa6wsxR4+164mcJ7bqRRqkULOBM4In5lutJkHJ2nlQO3DXfGjV
gP7ZKeLAX1tLU9JbutGA3WYCYTQQl+KPw+Z/bV9zXVBchX/p4M45UXLzBZvRkWou
pIam8i5Xh8ah5NDflFiyyVl5lXCM3rMRkNF2Gzlc0VAH/yXTUqzJllL6xFWxrJr5
QyQlz1B2Mz+h96mi0QuvArMUzlceGl+uY6bVxXvQoPsUedESAuap7Ku+j+TE/yJF
ugEMxK5iXzqdBj4RefHo+TlaO33yU0WMhe5nse3fU8tPQHuFn8EJH4aktDvEiloJ
/2Lau8s6Nj3vah01IIsT+DmsUTUZZL9SLrSWZ1kapklBMSNVY+94wf2z2H5x/wHO
mEVSRCKsnATFWnxM4wBV0L0AiJiChABikgcmxYPva2KAM6IySiZFgnlz9ych0JpU
/NcRDzxCs18/KN8/Qs8+ljug7Zv9tGGlPd9WKN63fXsIIb7NPtXDRiBI08LFqgdZ
Pviz0QbCak360LZFh7vRfLs/5uva0ebVu+h9Hw/iblgHwzbBbgz6tDqSb82kZQ2g
vt6BEjxfjkGq7H5SOPKiwo52olZm7Lozpg2oHg1RW9i2Lxy0Qd7kQvanuD0s0NnJ
GVLLPZF4Bs6wbCEyuzYZUI1Tns7o9xJrNVKVE1AXVC9wzB/GklCsyk1tTlE0lYFe
3iE9HR8H+Fh+cfgBU/wSh26/7Xgmui277uTsq2NLQZ5QBTjHRouum6H3Kt/glqbo
hMSpMkbvA3XiR2j97VS7IeQJovHA5i+QHYMypQh6JY/fGBzVzuLcNVLfFDD5fEPM
XcOerY7/2OEwC5eYKhP0JnHrLt07w3WOoQ5NUiY8rmX3ccsU/EdvUfdmul55IMZF
AB3EHJUQIoAO8lZooDVRQQpSem7m31mO343/c6ny5+TPa9l0meva8PDXPtuVVmG2
Uzqr7UY5Y0/pkzuo217Q6f0QJ7pEGOHTHOo4qxsahUrIVQ2jKOHng0ceo/Rtu51g
/yQ69OxI5uqLTrJUiEUxQaeF5Ap3yxOFNz+wFs2WVC1kf9YezeyTK2EaOYn+SfWE
tmLkVrAClWDa9v/S2HsSaW0V1avvFFdc23jXN6So65LS/fHns/L5VQ2aTOQs+DDd
b8phxoX3V0lKrIWSIk65VEuszOlSRT53NITHHjbEBEwduLKvCxRMcvAjMuVu335k
wJW9ULtAH82SoqElTcB09xFe7tNrBqb5XIKb4BXpE6o8IsmihOn1pUIPvcNX7FFz
NrBFXKeetcEKUIeBjb41K4pnPUJpq0xLkAvShvB+SlpqQQ0XjHLRMNgpopA0GkR7
86gzSkrBYgFfufTv5PLkrdcMHtNKSHQ98SYUQHPTG2qlJh8zXy5grXrqNaoNN0lW
HKiybp6KBeFTPhvQMK6+HJmZ8jlT6SRRm1wiIuN4hn0Ehq7kCPvqZ/aTfuLI3dNc
R07LdgQ7n2Dfn0JkQJnV30UHp3yO30KQP4TpNq+ARQVEFDZhzfFmbYeX9t7KTcws
RahlOnXxeHwM+YQwVM6otqyDctuxbdcT/2UT7MimNuMmmP9ObEUxnh5juAyk8dja
kEjnhI46iO8oK3Vgz2swAIEa4LLyL2kWMSUdrI7t85HrDvzYzRf8P/vL2VhU8Kvt
g1aYDBBvNPsiZc8yUu0h/4J6YXuHQPOgScFxN1H87SdLdXul8K4/Kq5tBAzhm5hc
NNSYNiYm14f2YOWTUS3CU9moupyKz9PwczSuIY5Bnqw7QumH11bg6awlBase3eCU
Jf8vYBEpBOGgBwGPj1uKsFcNbhU0W71DRRqOosTlMPp5BCmFrP+HDp/iggi0prZw
TX9FrDURXAZ5PCmXTYKKdUI1lO7TsPkD65mrx/veI+Hc8r/D4ihtka51YYKpcV7O
3xKsaRpY/lQq/lxsWTBFnI0J6CK62SLCa3TRjCIx59jpXZrqxsvJWBCYJuumHPnk
BmXM3cqvE/BHF5ywwmmC/qw4nAXTxErICCMFq4tCw5jMUog476rtWRc0DjLxgIu7
IApqmKhxAo+wdULINcTVnkMX7imnfTs0T32dGKpe0PkoSJuwnhdi5QxDSKjIuUpu
T8lLjMkdQ3bvYC2wC2Ecov/a/TOhlSJRsxYkHubKKxMM93YbfnxpuSN0OV6l2XSp
D+XcD1pi8GEWOhdCe4c6Br2217b2Tp6msXBtDLyDe8dLRSwD0RsZMLc+64PZsR+X
PJkNlXBcb1DPBehTmuTkMTWtuvBAIMCSIKl5rS0IQ322CaJizNxRANIYvEzDxXRc
T0HDl/tCmhxYc3FpaE4CnvDOTfF+5SiXNadFIS1qGS4pBHOuaAGAZ2G7CT3GcCtj
A62UnWgXXfr3PxftYADypPsVQEn3pZ0TnJYNE9F9602pAiPlT6JqYNx6/iqbjIVN
VpMtoW4uOFeeavkWzPtrDRRYODjEOZrprmMLDTjsRedm22+c6rGZOLBbEISWG02v
R4RuLxu/tYHK3J+aKJv2WTQPGa638IvQwBYDuRqGH6n4uYXinjqeca7zUSFoj8/i
5c20eYYYLvYN+XAQjJGc63/Bun86jlOjTJ0EDbFmXy3iLrScGaNbpP36h0wQUxqh
PEP9rRg3eFftBcWW7+HHOZp4jUrHvXHfPpYua2lcFkfeURt9w/snKiBSBVAFgf+A
p6bUlonCTFXi/0yP/63VI82bOojyu8fBMUaLLOrLuIOslhyvTxDEomux1+cptIAi
gXPrQ6VREYTRKcOYSI8wKLP7z4K9sZBj3Tk66PUMwi/WEajoQ76+9X/w4/Dj84dS
CM3Gv5tBISuWm919tVMHCAVgpIS3eCjojKXMLH6YzWmab9zBYRg0fjToY7KBqwW3
hNXeDrkJE5aLiPnAr2bT5f/8HCTalHV0P+pmyJSdXNghdzVLvoUgM4HxZYgeCCT7
du+sihE0eTBBA10MWMxoWDJLRp5cYxt6tw+qXegmWPGxXtgzIxhQ8FMz5NXU6MI+
IBzemtIoTNGSzsKwNx6Ti+YE47aGHbHS9EWnSKV5VVtb2CZtk+1Svi/Te9lPUJWU
+vXp9Xo19GiEMQyCjNyPrTqL/uHrNwR9k7tmn3hQqJrqurQHBv+POcSJtIKsIEzR
oBHtKEhWGwpNvBlx6lmZQhtZTHlHfqo1bU9o/jAx1HnVTVtgFPP//vDjV0w5+kCF
gxep+SLtqqtqg6HOS0aFDDyfRnC7idRD4BX6UWyBh59pFsDfUxGpWML/bls0l6vV
M5XSux+xqJzuh7bMXsDP7MdrAlpz8jS913BkW1JDis6pOmqY0T2oNFwBrmxkoJto
kKuGj7X0BdRkbvTJGdti9hSrchUsLAhdwq1iFHYXWAbQ/CpNcXuDQ4/rVAKqLpw6
QdrVbBB+rfhYV6sZDbUW2bDu2tycj1BlAQ5+gNmornjO7pvP9mG5tGS3KD8Z8BbI
oc57qKj4u8rr0E+vXB1u/Ja1/HFwp28b+Li+GAu/1878f7iQhYaq7pJebqe0tUzb
qwJVVO6cJcEfu4z4YIiLo94MzXdztRwIlOK8f1ZVM23E6V83bwZ0hNvJ92tVTU8X
f7oF1aEUIyDb5yU4ttID8vdpUNvbSJqn18DL5w5g8VKoqE04syhyIfuESRefcxgY
TyqQybkNicbb/BMT4WmzNx3LfRhSkydBLw2Ds1p5FJcM+UyRZb/TMCkl4VzbNCwp
n91UDeDdEa51Xy2ZFZWdy9tSS2T7Q5ZYXErCCqqZ1Aeg223IsUExDBBudCInWpv7
eDDeDI5aNOuqKcHNds8DicLJ3onQa1xilV1o5KwR7tAg7ThU85Vd2N6jmNbeKwko
dfMRE0tTzQAGYm0RuXMAEFQZzHnmGajBe6qDIyF3nI9X0L5LE7/G0dGKlYXO28o8
T33lB7Pb0fWAjUTutN1J7wBCy1LwkGTFbUNFAdK4efsQ/F3jtbIwhtSbuXsmnDc+
/6IrvtqFuoC5eAlF/z3dppEiyOmkUIsBDSinCnfkiaRGIFbPIeoNWbCDCTfI/djL
IL90W35V6f3qpqxnY/LEa0bmMT4hangcliAqSq0jWsuWQW+YElhbdey4HvbP/lkE
ClIvAqpeL2Uul1KN5yaD+UOojjVuwbDpUdufK/+fsBqsc9bclWLOmGebejtOeROH
NQCteY/4xKR3Q8pOj9eYOeGn86YgEllHh9+Lf7Ax5RPxyKNpwL2tJ8lMTGk6UWwg
`protect end_protected