`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
ddtXksX2+yylW5zu6QL2Lhnb2d1sD00763mmSITNX595NcHTEkwn0zB1Dry37fOW
FufOhVzEJp80NC5qZ/+F0Vk7Ik02dIR0elf3clrjeJRK85K4e3Hoo4xn7YbFUIms
l/8VZSb14+JVGURjfswrIyCUotIzlzVYZ6gzoZwDXIi5gQIBf/gI+KxNXPaKV+PQ
Ufys/12rjO6aI/pPlqSm0hCvftmBcnezN2hk1UeXgOIuKZnogjOsf0iJVX2aOOWE
6pD/psybjbnsNB6kH5uFTA5frkzIzkzl5d9+YDm9OyC+k84E83I/7/j+rk4L2dah
QJOvksSIzN867/4Qt8qYTQ==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="MvBXkzurAa5VTw+1JJ70nePUfoQXBvZOku/SMmg4TwQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
oRtzZL4VJ4iwysPsC8SXYCzXS8Fw2gtZTOskLcDV+1B9Nzn1zTyNtlo6lNICRmmK
ZRVu2BmCc2G+fmzynYlNTnSa7C0Cuel6FYpxCBlOuk3OF2tzAmLAuDyOH3Z1Yjzk
a0aHuoCdIRKv7BrZCdALt03JeUmXKPdOmIlkVGFl8yw=
`protect rights_digest_method = "sha256"
`protect end_toolblock="Jn9CQpRhJt4rnzZPRk+dOpzAubz7omckX1MrFd4p81o="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 11616 )
`protect data_block
gD6l00tciPUa6pDNTk/+t0OO0nC/UTtBwLB41d4inuAUA3i/ALrNyoJVcBnAmEQW
ptbcNp5fxEUJjnOxnedyZEuEBxWRieZFQnkRdF269oNSqDyGz+Zxe1f63SpwsJ7J
F2Fsvbt64/pDAv+mTaB7jY3tDu88FuhwLBhVT8o1EqG7Bpu7WKhEdNQ+wcirYY5+
FGc3NPB5qfw6z8uzsW/CTzT3/4+ql9x5c/cq6vGjaHvqt1YzxfK5NRpvlbJ+eSFf
02jCmByc1/pplYjjUYBBQqAyGRZKFBsD03eMxDJ0COzcVmDvqUjchTrY2uvEG5DJ
V/CryrF7Xilz9q8wz46d6mXe7Hlb66WtHsNWRVhgwoI5kM8xzoGd5V34Yrs1VOtC
STtV+rfTRzEIyPrt/5PDkhJDsZ9ld7Z1IKK3vq0kvH3vdjkL6AddjbWKj/L2D2H4
6mDW9oR90dR9C2hYW1TxL/2Xb4akqE3IF3asdeyJlRvSpS0DxhFPg/VbbpUSlwS1
sfcHUBYw5vh2byVu6eOUu4MMdPhTGbZzz6hi+f4deGXy83YyA7vOGZfqZsLpyDPP
kFeu1/xKwA1ZfFf6iSKqfSr4S1iITBL3FA7h8ctkSYyHdDlPbfZBTCG2P3cprC6j
OXk3BKNY68G8FccwtVNf4GOBmlVy8YBpnSo54+ibgXfZEkepw6wX2HUdjBAyReHi
r7n89ODIugzF/xxMKCYGw6gq0x4vu+tT7NlN6QrVQ3hfwUC8wNDTzhugRpXqrUl3
LeFRtFWKXEGMnrE0qnpfJ4FsEDvX3OmOmKhdtLq0jw3hfCljtwX5OqWKTmNAlWnk
/DtlvPLIFVs/Al23YPrxYH50tMbJVi9+tPxsm7c2qpuI+WYhGk+bFzTXg0JR6lwa
YYuggPpKu39nQRkhh2Divqqzw+ls8WTZcczjCPVuB191xYAu2pBjJPSnWgYMNe33
lczV9qWWN37MbNQrbzjSZeu7M8dbjZe+lGLO1BpDezn5mp0DJft5LyRfZ91V2I9s
ejjEwubstbYwjmsD32jXB/4GOr+03vaiso/vUmw2UEDArw4p4963rKQEES9oUfIH
B256y2rrXN0A/esoqg7aG/no+EpuFHMIMLlrIun2lj5Zn7IXgM2nxAg+7vReTayA
Iq3zM96GuK+e9L5bcqYTJi/QKxSYE+oCa1a9ECJIkrKxS7EJu7xMfDIe2xD8I0wT
U8pl96xSj8tK2evpPMisx9NgGSdckJ4myYE5CbcveuwufMotPpVDonkNWiV+wDrA
lhfQm+f5MXsyaHdTkNAz26l3fD9hFQGCTVvC3HQXTFSf9wMm2sKSdf6j7JIGGL2f
MB+pquQFRfnDGASAo8S7YG8jm4XkxI7vtkd2HwpJsMbDIlVSMWL1zDfPc9nNIqQu
KnNmTUIn1a2P81GHH1OYSBEX6+lmMaOlUPW9WJkxDa3OHrR5vH5TCTz7DoteCmuw
xGo3i1hYE/69bHBpKezlUF6jUaXpRlzGQ6IQhgpqa1iPtU+JuV0C5b9N+6XHw+UQ
AlNjZLlMfOdTaIJUvHJb2F1FezcsTgmXLJaFgWCuYssOu7g10yRC9/iSE+VQkF7t
XMCv419mJSX4KJCOTXmj873TjY1So9HKw2JYifeRQwywhbZPk1XfgshNfbLcOa/+
Iox9VFeLkWXQk/dK8QeyoOakIMX4IKQTJ9HTxDB1v6m9y49tOhIAi/UHwOK+VlsD
OBrUlynx0y5f18ca1l/pEMKVLK8FhaFWnKQZFikekwl9qd5yLCTI/Er+vt2V+I2h
LlaAGCtedH3Q68QtY1n4Nzad5x+k0JDFw5i1RyHh25CQsutzSFiGTm52N87YQWJz
v3uQhN6mrCknGfVn1+OxKYpS6OA1adXYPUyTVtBqyTjmMD4uXiiGbRSP8U0H/vIT
FxeZu2esWjezFVF1fglayaIkAcwEnSRhvC9009V2RHciLrXqR8TvYOIrGvzHHuIR
TaQWm/SsTdqo1cFRqBJ5iNe79e1+hZZEyfGelEDuxJWvpbKtwzxx5qv01S/+CvV5
Xhm1GV8yZTB1+c5n2RaQzdpN6fLNaebrOREkokJZRSuBlt5lrjiCampabg7m8xCe
I4pasQcM3z8LrE2IocrZ08voQFLoW3TEjqdI9zjacWU3Gv9ckt1+krpWjh6A6kAq
UQqcNroMNZH2b5KazJHlQl5SXF1omPMd6JjJJAGoskK/fHnY0rH9ur6JF5NNvyK7
dLGSso17tGHO4FM/w0uHu39uBeylf33j0HEEhkI2tXR/tI7wCnr7xBJQjzqFvW9G
qfTogRFyu0fX14OwjhGN++VvLCuvzAwb5wUKdqD6M9xw2qGf46WWL5LFzYsXOJa7
uRJ9SJP+/Ye1nqXn90uhw3HwUmOti4AXnK92mQh7VXb6kCpC732Uxeo7hfbYcEJu
RHjFYJoXTRV6YtRCm+div3A0AsCSC/eWBMk5Snb9XRIV7nZ67ro0zf0mB3yWbaeo
MoXbW7cvuNR7XNmrm/+sgoJX6eDY3+THmxdO/RA2Joji6zAai71r2gGZgb7w7evH
4++k2378N27fkWp9MmGVQgBthw2sRFwJGp5Ykkc7r2Ls4B6V4+VyM31PQRZlAGTv
ylrgDi47GwLfpB4u9Zy2XhXlC+GDsYPsnJM/z3yWZYA8MreTlCtJjdJg97+M3sqU
QY5Okno0ln125XYJKSHaiFYfjdieZJp6JojKttse1fJSf7WOlyxBjpeo/q0JFvhn
ToBT14EbVfMYCY/F2OqHyvBD1IrF+P3WjgwJe1yitgfqaWF+XgztJ4aYqNVqCn00
w5magHPhnbFBErcKMNRW7NzIUhuuEX1DpSR4QJ03je8vCK3JqCAjKOD8Yj9Czu//
yn5k3jF2KODDQHZLeTkVY+dr3HYeTYJeI0Tw5BeVQ1af9uBBBQ6jWjwWno7Gcm6n
ppP52kuQtns/ktUpqdrUUCfAOAiMzJMfoVWEbmKNBHJYpHFN+r7jrU+Ew97PPtNn
q0OSw7+0ET+Gm6c5ekoEqxcz9hLiS1tc6ZiALPm1hbIUDaJwGtaKIgtGrF8XZfRt
lVDRrEft9kuq44/6nNCJanBMKn9uBmXTzQZbpNmzqoUK6+ph80NliQSQONRbWgO3
YzWXA/c0gNYp87R8cf47ZEr9Ynvf6pr29z4i0HiAc/6CDFrGaTyd+XrTMwyet2i8
lB9wdu/mtYgJsO3ivk0rL2Z29i/RKUI08byFyo/jKUYc1b6QXj5Vb5cjXsB7TQ2e
MSArxsD8zvwQwoGH3OShbrtYdoOZLwnCPm0YVy56YeS7Z5XOxePmH/FlsusyypS1
s+3+JI3l+PAVvaxSqFPhaxtIib14wIA1iWMZ6Z1ax3hpIIveJ0l8lxuhWyGZbSFy
1eiJOidy8nDlM7Bo+741jNN9ohPtHN1GRYIYYwFd524hlQPlvQDA9ClT12ahgJi5
ALqGkNlVqlRH/rr0GnIIHiOIbua0Og/L2Mu4YpBXDICI6RufZ2P/Vqp/V/AptMGf
slXatOursVdl59YC/DPtVMdH6OZZihIH0TbzmMbFBlfbGJ5p2J9I8I5L5B2CLT5Y
HGRu7djmQa46Gp1SqyfifD6+izE7NHGpNNJE9GT1rRSB8HNMn7pG4aKd18jrMnbG
6zY2E4oOWX01Z0NuCUS3ncpTG39qtKma1Hs1DdokwbJEIBP/u2d5UmoG2ruJG2RO
8kXbehS/U7BqDE54ugZCV6w01N3NePkS+EyEvmHDy1Ayb/fBYsehv+llR7McICNp
zjN7k3VLyWZgqjIUA6wsh2M7POyNy7WTfBX058JvEfeW54iBuv+h/oMU6S99TXTU
t3wp2binlq14UKkPl+6lkjj3TupniXXbtCAPi02znRtPcmp1bCNGPdnuOAkKGX1D
OLAWIGqNip2Amcw7a1cyjPFhNibW6cn9UiN4VannLujIkvWaRwfg5lDmjoL+O4EA
DxjIOkGBF3Nvev1i1Xw2i0J+T8YiJ+tBHR4Jj/XxE57ZDLUA2nAmjMf+pSR7hN+X
lYFDidGMvGi139AVoZmml1QVPGCjP8ggXTvmA6Qg37Z/IIHQpUQj+xviknpK0vD7
v4NFnr3tbcPRVs+38zY+BXJzZFZHqQWq6yV85RHDGo6whQ0X8lrLJynZ7d6Jn2AC
aE39buboXddOpswnkXcsZ4kWduCUThYbja+NxMYTBDIsUdV8Ostoh+xwgh34WW/Q
omZ3FS4Z1kBRCHEbBve8H+jOq9ZsRQr1I7DJWfgtJKsPChyW14TYYuszdsJG/MEV
AXrH19tIWA/K167tBFDst4Ve5UMKpIzu7ld22BKSPrdLqo8gmBB7fu6GRxsrnTee
asvmQ5nbLUzyy3GivLvN5ASp0iS7r7T1y7aYlQI0SXgoaiG4E2J+5CYV10CzPmML
Hor2wZm9MN20s+GemrNCDfi7wyw0AXLALS842yhzIlnV5THpyLKAeByt5fekraJL
Uf4W7OXTnPpJbHHaVfEzk0/AvPtYnzY0vxBegjP5tmMjaGFowTZl581ASDINyvY2
ZHSmU7Soha/kKP6H0qlSh8iFMwKWH8y4ADqBbrqfbgrsiRVtCY0dYKlUAB/6SLss
+6XGLT4hQT+3AL1A1/y4CmL5kpMQzD89SmJ+oiTBw+1uQEb1IMeQqiGuFpKQON7u
vbOk4ZCjjvwRQfqnhIKp09C6b5pXl30RstthIwIg52J+gtve//kclhtBDYNY2htM
+MPWcobEyU7JF/y9JqrWGhgbAQBKJiWaRoHuvNVG9/f9EuZJTf6osQGe5L6Z3cPS
EPPe/T4saG5U7DoX5zx9DEZeWUSyAxdPicm308f5h6Xx0SNS99rZrsCNfeQ57i+C
uiG4oLd2BIDB6/s+QeZjaqvlyoKuJdtr6gobGZKky0TmkWMq8GyDdbxOtprwARXG
cbObK8DmdD/OLfTKxIgqrZWt/kF/XdvmDgt4p+OhrggMisr2BvpbBy9meYFtgcxx
17HI23MDiBAsb1hyiVGhuIWqo6nHYvU+8EN/yHOaH1VobLdnVPx/q0usVRDd8KHT
J9Xtx9oSrCaN9HrzkA7hq6QLM358BIkTgfOHMj/rBczBFS+qPkEP9qH10dNxwhNS
V6DKY9dHe/251xv48lvGO3+ffDsbH2E8DRu11KIqMJvgtA2Efgd8IVJ1WM33RjYJ
tbtNnGfdLhGiXxyxzVMqhzx5fw/hpTJ6KhIUqyUPi1cy8RHQ31h1NvXmPa3J5ja/
1nNqizH4it4dmxDS/jZmtni+F7++CF1b6Bgm5UFe7jA+DIw28Mrt/GpmyGy0183r
KiwCsNwGx0LgeemnnaYAB/w98fQN8ryIo08ra2FJbLjk64VyOYJ1vhm5i2VogUmC
YHhz4ZDSb9bUO9mAhEY0LZL3s8gPy4UH3lbFC6auldNoo7ssDMyjYXGPfVXxqjqN
CflApZfKCkABz2siBBphPS81AM9WXzxVXlJWghwkGF2tFMprzr5guUWDgW4Uulva
irhkZ5vguQzUFKMba0DJgwK/0C2cTfabH0ICFdrkkCt1Tgq2Re5bApkrmd2zDCGt
pT3vre9fJH+Jk/dAYucqv8guNDxvPumd2Ss1WxvfnYgbvMs5Z7cIO2qYbRxcX1X1
kGhnOMWvoFsUhcvj29Bc7mboqSLCfg0jnUQdtzX5n4h7hi66xGx0jWdQVdrEr8OF
vJBywopPgquduGaeJsYiuqmgDagLiVAs3QjKF+kLOXVQKeLCbgI5lnUZDU/Q5rxa
oToVYla8NnE8ZjTMAilgVO5wJ3xVDMT+dNgabrOYOg1Zg0B+mOz/iFNgFkGA9M91
DMKvrVjDQkoonvAyncRD3aBozPVutPQ/hSbBNtfXhb3/hXk8ZcOkzFd7S/ZfRFIu
3FI9cEUkkKoGsI4nMgr11QLIDqQQS8rTwfawd5TcZePx2lYviJ18k3D7wyDojnp6
eCPQkwoOBNnfgfAT9bveCTSg/YDRDKlKQTe53TgKm44Gz04/Y1/yz2QqWt6cOuFq
BlwpOKp4BeX54UnupTgh989lT1Ub4kcmteG6oi4uB9aWcEWEBjH7qkW7m2Qy2ZQb
mi53wNMdfQBVSni4h4U+GGMZay/qP4DAZg+Ph2PaAyu/UhIibcSLbxnXoeLIe7As
6U1p3rTNUtrblleATW0pUhifXDO3nKMjZof7MRmUwEqdFR95zFZilM6m81lf/lQ0
SHe9G/kzzU/G1rtSyrLfdL5k8QPz3Qx2UIZA3mW0yW4ey0Ysh7crNdLOVoaBcmEc
Q+yQpVPtfjDV2ogIxJGeYCMNPRG3yddZVwEcbehFxR5jpV72eYAAXMZSaGj2RRwM
5kGEcWrSRsygT1G/e78PAcIkEe6q5Ao47YITpg3TCdllqoQNH58CNpeHYRH/7N2n
1za0UmbgxOAAV3AwaXkSNub5dqbpMTClg0Rdqckj9Zvmj4jQuLk/em2N+FmIo31v
1lVDWT/58eMalCDaAMFvRHxEVwMXJA9nTHxdOMgzigPrWBPTUB6Efi/ZkHkDwZan
suHJ30CabQoLBzA8Cswue8fwmNUeoIKadZk/n6YSLQS/3r2jTMQWc+oKGtRyko0R
haXjGBR2kpyjxNKIfGY3H7G/UwDu8wDLYyyktdE8gkeDbxS8XfaGyX0nlBwFhLWo
Gu2qBoVsRyXOaf8oiJ23HUBwq5tn1fR2pFGExYsZSdFdDaFNWHOfh1MP+YCGOIB5
F8tV9mjnPDfFTtR65mJ88H8+12QbATPnq7wWH7JK06BTBWoLs3BhkvS5q4ubHQJI
jLE+5S1HvTA9vXyvj0zwp0zoucr4tnsc8iXqzAAgpWcmKvW+4B7T9TS61pwJIzvj
U6ZgvfIWAVxdze+zZscEJB6Ea5RyOotXPrgKn8z/AhYHynlEIjxAYFz7UQ+ihlwg
zpzsKn3AH+VmZNTVZ4kKLHcflNuTWegG6HVojXU1FXWxfv3iOCIXzFIau0HUBtYq
C7YEEAxDDIeFyaYea3HcmOyRIMCCyqSDUnn1kHsM2gFi7oRk1X7I1T9MmhiYjcFe
VGDzsq2tklq6nEwo6iAyIXYTdUnmL8ps5uADn9/CKkDZo/9maM8iaKF9AKmM2dmb
pPvy4/77q5DgD6xpvcqrnaQznDT/UXyZAS8oglEXyHp0lBaJAkpT17aR/mh7D1I3
FwaqJzkK0Fw2mgvU5ch7NuuBGN3I57VZURKdxbxONmNfAZLZ9+P9btZaHinV3CBo
9O0qFN8rUp5GvMA+dqrNnPMQxEkuQS+jyMMU1kKdnjWfWr95nR0zrgt8Z6xP+LO2
ZGA/H5J91a5rUUirCtMm5Alycwat3QU228d64sGUgBMW2T2uVDHDgvdX38edTTpO
C9GYY5l8SU69F+1q79adOeilAPfQOcsuQWSU4ywFs4HQUAHPxhNBh8Y5/rAU5ddb
l6KPgZnIFstVb9OEj6rWdIqHqJk7xh5XVL5KafE2dyFIbCARAy4pxYxfAJAI3bpE
lszoA1HNccCvtgB7iouP7/Xs0V9icN+RPgkCQwnEgm0XdMI9OhZ/Y7my2bcifAvX
B14aGg36ZF3N90NoMJbNEJ7nQqwZV42KCYFsC6ry3F9666MQEi8ks5HrAX12o+2P
ZK67WhwZSwC6hvCDpg8b7NZnJ4do3v/2Dy7L+fPN3jsKHq9sV51d4DFfuuAD/no1
Idx/pdIjPvYbKkBWhB64b0ZTDQm4OUwPyOwMWEvuTVe4SjvWafGtJw98VlSHJk1w
GRdWDZo/9Q+TVOS9GgY7aC5zKFhTtlbuHSC+wrV8GBI+XALHP23zN6yx6D6nqFzs
2k3BNVwJTbFSEzNhIAJlxH7HM0vkSeqvy2CI3Uv+oJ6ZX433zd55jtjQKJJKzb5P
yQAZlACeD+WnRxXMT0E80/26gYaWBIUvJ4vk6sjz+2zw3dvIkLsDZgBYbmYM2oCM
eF2xhidn+bcLt4lKQ3Wcfn77BsqsoJaebi9fIhrxX3xE/8f7GxGIdPEDYiXMNpuX
SCtTV++6s8IRf+wgNNCDSj+eM5uHjToB+38fFtty4XVCeS5f/sKwNVQHTjzk8ady
GFgtvqw3qnEm1Ln1/QnwuS/da12/bDwBcwP4w4nuPtvYsjIiUYmgtR6bUeEe9+c9
2xEi0DiyuGzF1hxFu5d6B1CGSJIM1M2pmnAmgCzFX6IUR/vsiGENDD8y82X4uMQd
ZYw6h6mTMEZQPvPM3WjOrz93Bd/JMh6yDblilNwFFFxFlU7JU5OLBCH5lOAMe038
3Cqfle9PvmdyI05wKR62qOa6cZKWYCzkjOYoXohOh5CuvCvUQAtPWvFd1nESDLge
2drpD3v8y31HiZQch9gkWhJzENsZUpOJrlvzM22LgZkCLMeLzPMjO6iZkasvgXQw
g6zox0T0DgejlKFSKZU9aOPChZZ9mWbZj+8BecknrMeFOwHGMtk2XVtBCQUazE93
0tBK2Ww11uXICNznN4YvYMM3iCVororWAVeWDwM6QO2ZNerKexFghlNiS1sNC8Ra
4IG3kE75FawLXnpTZbgFwmGhY46J3y+4Tc6+9rHvbh+rQDrGnHL9dXCUDZnCb7il
xXubi4iCcZujpNwdu0Re5ney3DOBe4fzNdtNJ3dlKthTetLMwaGINkkIRq4oA9Tq
HLCm31JhYVnu/xfs2ObfjaKKH7A1faKD5tu3Y0QoCGtLxSgp19RGXwPu17vTLvMH
6hqHlsI/MI15o09XQRYKu+/R+8cuVOFlgFumud64on0gi0j5SfTatWmDMxGouT26
lEHK3YcCHEd8sRtEk7JKf471AltV60Vm8fd9kOBVCBTSCOiPp8iVsM1bJF5hhe/l
b0W1CTNWOSsMrUPi3kyA0W2D7V4SowGb+UO2a0BhDg4OzBMDA7DRnKAuWnLlHabj
D9Gg6weevbsM4cgR31lcNGqWXunQaVg3JXUjcCOIig6PTy6eYgFSk3jFQLXGpLDT
ELeBxZRZHcNunmiff5tuLj/kkIpGzDoskZyqZbwVFrZ2ZqyY8/wF3MspL9hLL56N
JWiiN6uyLymErlsnh94d5TfYIlgqhWxM2Vo/+QP07a0dAlNnN4MTCuAb2+amZ0u4
icWf/SjjT/tQ9MLXXHKMpCvKMXcYoZJGQn564AjBw0bRc1ZudtDjbK/BrjTuaNUU
Q2x71LYYkrHH1Z+80jH/naBSU5iBF22PkJpfSUPy1R2S4rCuwdzoDcHwRXupIqHg
z/HAjzEM2Y6fKn9lT7Lu7XN0kAQ5WQ7iX+sw918kECoDhQRp9nRoQJRve+6Mv7++
hvam4mFVBcMvSpUsGb6BOW6OOwVC6iXuCQJCI3okfsFF5AuFLrolI8W0IRGaZ2tW
0EwiAgs1SVuyYXJ+14ehpFPOgJRQ/f62PHOyS0KrcUFC4NXPXi9/60uEf25k1ikT
V6QpzYeLVT32TJZmIfNThwTbce8KcUV6d0z3NWuMhDWZwk1RRf5f9tAtC5yiGba1
Jq+za1otYtABzTprk1FlZ7c7MfIomKScByBxF73QOR8E5ioUlSW2/RmuMeZOIr62
BMvsoto3iPXOlc+uKd/54URnnshwnf74+RI6Cf9r+cGzX8HgT/qu6gAGhqXY5Y8m
2aiZp3iznh5tVu1wkruO1YfYXYIb6arVMKd08aUS5x+nJORy0QhJUYbzaIsLEqOD
a5osCRtrBLdNNh2yyXO5chT+gCaAu0y6c6gwL5yTPt/pL2VZd1zKZ/Z+Z+9XVJGU
0a0aS3vjgzq2yzb+S3Oicf7Dgba809+HsPMRrVbLuDmqc32LKKzi1kPw53aPK+oC
/lLRxiCN/jm8wSuxkq/7LPFcKNDfbuHpYkurPvcl8rLnd5OJMaM7qTUeFlZY5jGC
k6QTmWQWqzNHkGUOX5AlKBYSCHwHlGQWkryzv+KUlYqrAnyCl00+IEKIlGvqPAV3
JKJkInH8yAl8yJFOOsPHFqsqmuC6JUJWraB207FO2HV7olsOvXsbvIXseNQjkdwk
wemG+2+T3NlAqW/YW+kctyQGck/lYzGRsRKyXEdHBkOVIAMbFOuZf/CEI8rLnTuR
zAlP50nAss8/+HkiXfX8KQFIEe5MohENzgoMgtp+KdT5dEu8JanqS2Z63LAbZEjs
mckrKOS54Jcq87IG+vTM5SnH1gi3Lp85fXP3gN/kNhfZd29vfCgBlqbuBGHa8nf3
1Xd3ZT4GsA35Vjz4CkR9+IFtoHI42zRYhFVjn2bc5xXqzGiKfW6vyC2C8YJUxZZh
F4hAiEyF+aQMA5Xz4BeUEZRgKuPD6FSOOPggnSOLVrG+LtcL8I2sG0OHc95yK1Ny
RwTlJklNaWsAxUk2uzwkaADAKNCMWLXhwpvxpb2sDT0XDjfu5BqXYucAHIEVwYVz
7AAKLbasfJBri7Ljqk5MLd5Csm6PN19CY3W5aNUvXPr3rJULm8soWHlQvod7O9H1
dzgG2PK3zLTVJcff0IwefCkrf0m2oN17j+FNF8l6sWUu1Rmx+dMAjZMe4szVAP5T
9D4nzVcHbnjjuiPVLM+PG2XagwMVumhQ4CrQYbA9CJlVm2usllCKJqxY34kHK+rT
qJ3Q9qhzR7Eo26LGFUqSc5VxGUfkckUhDQEE56t9+vkr8GF/SCF1Fc3B0jvQ1zZS
kboZuaM/zqOHULjN3fU/ZJ1qBLrK4bop7PPMIh9SiA856FPHvzC62vzbpMLd7CVS
j0HImxcnmQuX6LBPzIkOzu9Y8NkPYI/aS8lZPvIOQrIodglO6RjDM07V22WBIlvI
dd3JtnKe7oG4NkszuHP53oVUwbHsqEqPKmQ7bwj/oHWmKDM7ARVCWEP+LHg1yvxt
/5bLZuzwzWYOeRVuSmaq+gYzbwoHEk00VFhRCzL+8SFRnpVAyjWQY9vf8Dp/lzkV
rSYvyTWjT/AVgyPiU7xaX9RlFOpyMSoz0vMF3vHjEW96LXjdwZ0OdEZFDXMan/iV
qCguSzD0ooTvd6MRAWllTnuWF5THZM0bu8bC4o86pUusS492w2E0gqG7yC/dU6eD
PgrznEIpHR3cyDPsvLwx7eeQS6SynYxJGIhcjGL19c+MYYoZMEoloQDLkkYuUwrC
WWpL5X6cE8wiJ0dLBcMnqiGPgb730OGVwklmVqVKCrBEYNz1b47PV/bAUemFixf2
j7XopBMJzyfDStGyKl7xp0GjiBSAWI1fAF3SE/L4w+izRclxR1x3NCojgUo8MxYE
Pqmxpj007TdKgloUA8JVI9TCHVoejnMMxvBePAAW7g9W/gCXYbgXoNtkTxuvIR6x
fw6wtrSJ4crQSrG8YZe17aaAdgACO1djpesazduBoIvaTc/aVpeLPe1DQm+FUhTF
ZCyXYz6HzKO+9IRc5LPqw1B4cAfy8TaBFDTsm5TVHr7dsYZ5VuylZDMHR6Y2GRnG
dRb3O/HqvWqzu9S2s1lPtGGxHOF+xM8X5lSyGXLnerITh498lcElE77GBXxCaxtN
0Ih1Luhwu2u01k4BaiHof8dKeqVXIMplq/1ltupuiL5qYrCQMieVBMUoEUNgkj2e
N9Vj95Uw7x4EFfliZFIyU6XDOTvH4KAl9XluBNU1iJvEPcWvCz/fdJ1+RLVxjFft
3hMkxtKTygVoP8VNLoVLxvzbI0LG4trOu3VMCYN8uJ2fKf+RIEY8uAN3/zO+PXZV
mn3EqQHD1eRX5IEzY6ex+Jrt4ZS2R0ETwzx4VchuvsLIvHhI2m0ZNuSUPV7RKPQU
X5ZPGCxmWhGGmLXvlAFxspkWfKDVBXAgtMmL8gd14H6eNSKzuZoNP7jnXi8LME3S
3llBSD4RMt7uogcCs5duVbhLNKmqaJbTJ70Ng/V+ZZS9xi6Yo3HTvwBXH2W23yX1
9Ie5IslTifo3nRRyBZ9NxMjsJjMDFK0wU7R+yTPGBeKf6l22eFLhTUXygZ3nZEnu
1BGBcpZb7OpE3WhbiO6ojCXWH0fNOr4GmGAxk3/YWnBZZ0KdL5BTDmyigEPeAcbm
8jnUNamAjlMWm8w4SxpYFLx2XPbsgrSAwuLxqI289xRbM/DJXz6+N9uBF1PhCtbs
4m2H7uGQoZHgPd/8SXOVxoJ+2wDDZC0H3qIkLb2j2wZuOh/Xa+t/cdBRC82gOwAC
IWK0MX+mGUacGYyCjhRImlk/xzhTphB/R+wTUa3tuyWnlP1IZAcoaFcbe7xiRDiQ
XCbEQy87VTsgKjXUgThyd/drz3KxfROj4vMGfG2AVFdGr2epm/Q2fThObwTMtI8J
x43Nh8p1XSWflaF/kV7MX/D1lfK82SmZBJKLvDYwIz7PRmhtRMGnDz4pwVDA/nCR
e56hx+Q/sYO11JQfBUN4taRf26uuv2V/DF+Ly2RbuHolh8knv43bho+oxTvJVfz4
vmXJtMI5OmYpPIVwCphsiSQMXv4N8HJskB6kINchDkDX2L56sQ2h1cIi+mPqh0ws
kTj4Qu6CHTGFHg7J7GRkkRfDvlqkgycdvtMY3vzN+vL+cDWrofUpFPvIkjA1mSMr
8KIGYlbc01zPaJ2YlbamlRCp1iSruXVydRmawvVuBSaTHjcI8RgHXslDLLWhmtvP
kHFBAGjb+r0lHGi44ttH46jyM5Gvzyf4pjYCao7/8sTf8NF86MdG55LWceeT1qw0
3y1UWx0FS9J2X/KoSSNl/PAbn2RwU4+BxXiuJndJgObMDqvXT9Juo1EeHYfhiH/5
X9nwbS0DHXOG9LB/kbDi/qIgX7QbgjiZouLBu/e8UymGrRI8GTfUvXwnyVsZibZV
GB4lrpzPUxRkiscHBS7ZpAExaAKaWRdiRyLtJWdg17mgacMPJ7EeiaW+1N9Qg3/H
hOsme7ZCUyv2HEVayu9GFu0AwImFmVU6Wh4TGDExIEm/Brr5D5KHxaqH3Du8j7M0
W6n7TzLY8Ew/xQgOUuk+AFEirqnA6W6fDxEdnxFSmY0iRaKUPUCmrupbnfvcivFM
rIUN0lRv0ppIhC5P5DTNMRQ7sw645QVjG8fX+xn3DFgd06WqAqZItcE14QQnLO+7
jQ2Vfj7AXmsAvu+2dr2TDyTRtA4ZxkCXXgshgPMX6ybTqCXJbLNIe+KzP1TPOFbE
61GYtC6+eA06QR8/nmdhd9juyyr6Lwy8GVlJwBDzkbmw+3/huskxrn5+oWQWRN7j
Wzs1itzAqKFwaMjOavEAdjlwGWF8D0cxkbJoetzYoAf57keC4Pi/s4HYyTgw2t4B
wRw3voJCQRJaADJ/mH5x/74SO+YvUxdefc3VpkTCl0ss7I9qICJoOnqffmqdjPxr
yWA0JY5cU0Qr8CUEl+sk3Pb8SOB/c3xlwwljXwe4Qm7e6ePlmnLHcc27tVV/Nxe2
3sWKGwcePAd3TbnJU+6nHpxkIW9V4LyPZJZ4I8qkz0H55J1zx/nWeU1xspmZiU1l
pGF4LJSRITq6COa4xGjoVhdi4qqxlUtVrh7/ye5L/zRbqPv2RTZW7xJV5DWezWWt
qO0R9otRxyVZOPj+b3PBiK987YZH35jFi4k1HdPu+/8GjbjdYQNJsE6iu+OVs92w
3PIfJRehlQGt8arjSNtUp5h7D+yenWpBroWvVmkcNRA+Kd4Qe3uyQ4NG1yFUO0+F
PtFrux1sOG1/W+5LMOfm/hi9wVUx4uZqqgoV/TBKLTf6cMdNg9sZ3TIJ0Ew8fe/x
fx8qahz+E3vcYpeDyLZrEoFnQc4oIhBjB6t6vNMIvX27xS/9QfBVe6q61Ne/U+yI
rQDakY6FBsJJ+LIlspRZuRzei/atoZxT7eDNAx/nCHo7qWrYGOZkGrQAtUKvAADN
wKExeBq2KiPrFonaEWFccjSyVVwEvHCmNkLSA/W3qCxJZSi4hDoP4d2ol8XIf7qf
BVsF6AYgl8ZBpdJCV29W3f7m4KqJkBrtm2Wvcy65D3N69XIPNxwSu75a25StkbEk
Ufoid1L0Av24z9BMZnGufDS4K76Sgs7pjNdwY1Qt4RvK66KBJP64hf/cX/RXXGLI
zpTOvhUeHjIa8ZKJw3KEVoTI7mH7IsXknTYzYxZ7HwsMllQIydeXDboZdYnujHXv
eVLuTgKRltzG4de47dNH/5rcB3owrjv94TslmHAR7U8bdSshJAp/j8nhVhYyNNba
RCpnBgK7BgkLlbH97k0oVUveMGMjG5xsYORnNeHPOKqQTRk6TSTn01LSTm7+852A
njX7R3wHikqnkC2YkE5eV5EsbZ5MEopoF7sjPSCxrdMNDBpv8NGFsgBl2WB7My97
kRkXqyHaWVXnWCQ07hwB7VCx5JP7bBUXX4q1d5ONfjfde5c9WZXcSMfRhtHHi/gt
TMSmKlTWq/UZzYZWBbbBFvFKuDSSg84qKHQx9KDJW/h7/1H1nhmhQYklMV3V3bAY
X5imaL/z4WxQLccGc9fP6iA7bF+/KOftLpBaqe5c87JUWgwv9o9IV7FWNs2Xuvnw
VjV8sVyhGejo12dgnjQbV8l+Sb2xUzpAsoy1qohNRfZ8cVmWnM4R4gZ3O1oRA4OS
/ad047GU5qLUARLj9TqQ8WmhdnSa62Ck5euCB3qFttsDVPzdpi1IR51XauleDSZO
TsKRDbT6ooE7yQTnKkT02MkPwCOnwRCkyno6PuzhetoAf19nYJymxyGjCDjZn6W5
hDS/Hs1oH42GLiYYDkeD5ogZjYDYYP14KlW6rwVQ3RmeY/SlO0TdIRam8Q0ZcRN3
ZKQcaaVZ8L99UZbH6zaibk5KElI9FnWaBCkrWj5VfhNKneIRjsoFelMvJ3Jr+apJ
Yl4PqQxmrXZ+Bp/Up26LOB9R0RU5EALE18OJv10BCGX4NtXgQp1c/lD7JZZZI7sj
nVrxm+13V+78N5afTibeK1VyALr1jH4cM8xLq+up3iSTkiY2q/3Jzex7A5Fb4cWl
LMg5O34ykvVl4c9C6pRgYyqneG/rTLBummvHh1hZMOSqCjRJMPALAde6VUGwkHhX
MdTQDs00kcHV7ZNb0q29y3muyXrg9AfiZ5kTmZUqLR/ZpcxwVJuf0ebdNdyTvQ5M
RrMhKvHvdePcbdRGkZU1Fs8mlniuLw9ldbDOrkE8ZKda4pPw2yM2JGcC9nDL4z1U
05+6Sw6Xkkrm7ClcNoPioueu/Rl2HfE9AfL6JVWnrkt/T3TI1IQVI8xt/pyiaGci
m/3nCwhojBfitAkuxMk7NUTg2QJ1DgdlkCJQcgZ1/atX+neEF55ESfocMnWQwbDY
n/PmoGtrZa2kPurhY+oICyQ7ZAoXohe8UU21N6EnZSZXqi/1Os0WYaxhX5jn61yb
ptKQOKmDBdWLwC8Dj8BwTxGr0dgzIpa+IbfycKy6ITLPNAYomF0wbVpVzsJLW9sr
LcRvuvqFvvS/eIb1LxpuVFWETOtZ017iIezg3c0nwPWOn2lW28MOQP0NhvWeR9go
6q+WLGso39KwjsElNF97dRQ3a3ap4vMfOi5/h9bCjXow5F5B2SXEMM/h0qoETdfN
DcY6nkiCH+kE4VTWA3VOJlpLFBZI7tlFq241R+DmT3NIpCWxe5cTQW2ES/+O+XUj
`protect end_protected