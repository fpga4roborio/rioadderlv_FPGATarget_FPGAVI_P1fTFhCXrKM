`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
ddtXksX2+yylW5zu6QL2Lhnb2d1sD00763mmSITNX595NcHTEkwn0zB1Dry37fOW
FufOhVzEJp80NC5qZ/+F0Vk7Ik02dIR0elf3clrjeJRK85K4e3Hoo4xn7YbFUIms
l/8VZSb14+JVGURjfswrIyCUotIzlzVYZ6gzoZwDXIi5gQIBf/gI+KxNXPaKV+PQ
Ufys/12rjO6aI/pPlqSm0hCvftmBcnezN2hk1UeXgOIuKZnogjOsf0iJVX2aOOWE
6pD/psybjbnsNB6kH5uFTA5frkzIzkzl5d9+YDm9OyC+k84E83I/7/j+rk4L2dah
QJOvksSIzN867/4Qt8qYTQ==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="MvBXkzurAa5VTw+1JJ70nePUfoQXBvZOku/SMmg4TwQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
oRtzZL4VJ4iwysPsC8SXYCzXS8Fw2gtZTOskLcDV+1B9Nzn1zTyNtlo6lNICRmmK
ZRVu2BmCc2G+fmzynYlNTnSa7C0Cuel6FYpxCBlOuk3OF2tzAmLAuDyOH3Z1Yjzk
a0aHuoCdIRKv7BrZCdALt03JeUmXKPdOmIlkVGFl8yw=
`protect rights_digest_method = "sha256"
`protect end_toolblock="Jn9CQpRhJt4rnzZPRk+dOpzAubz7omckX1MrFd4p81o="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 13824 )
`protect data_block
gD6l00tciPUa6pDNTk/+t0OO0nC/UTtBwLB41d4inuAUA3i/ALrNyoJVcBnAmEQW
ptbcNp5fxEUJjnOxnedyZEuEBxWRieZFQnkRdF269oPWCYOsMOa0ETUGZhDJBf04
ZN5ScIvIqUhthUOZlvtYnIcVYRIudmO5ZBM93Bi0i9YwWHENviEzOBP8/wQYKKMP
Ob2Kz31tJlXKWQukyl9AQHjnnnyPMmFOC7vFMIZMulnM7fJMA78aKrHSQgreYCz8
fx13/+OSmxyrUeBpRkgzGggnlAJbrpW2ty7P9AFJcqMP4tZT3AG0Jsd59z/2+vkH
ohzY31Phhgdl+JRVN73BDczLs+vm0J5vHb9nyKS7ArmWzPkBIOdR9GHkvrfUt9Kl
k06tpzbB67arQjElNyjIbC2zbnMqExBI7LMhdOYEc5ze55IZdV2RMHjiVowrqiEQ
WGFhlSbvl3Zm38mpNNLS65izqjUnjvsxF55VR+u0EDWirXnhdiBeHOrc/qqBi2Dw
Hy52tRzO3qtpYhyrNBw8SjKZKVRKHNMX+QzOBsLJDbaDo92LMCR/I0w+u+jSQIuj
iM0MhElaI0D8zKD2sJ2pslHID5/6mtS3JlkCUgkzCX8TqAjNCn/y4NGJxnkuLbyS
rJCwf1gGoC00O0DjZyqezftVV4wTYNo8dvBik7bUcWPRtLVmrtDUo/oQNTeaW5Ne
se2BYecgT+7aPdaoyKJ6C1pSXUlW1o/WB6PHpBkJX/QiWrMZKclchwfZZTOTmCqv
mRwo5sN2Xwug7ZWWkGdL+IWnh3GXjFicQucTPGRpQnTjbbr3ej/txGfjSStTLDo7
GJfALxbV3xd+gjLf1/3JdUmr8zLuA3ZZO15OGCQWChdwmKomUadRHU7tn3TE+ddd
rxBNjdBr4nvgC7TlSwijBMuUXXidQzCrMk7/CQ/KrrD/BkQEbRTQSv82E/kMucwW
JKhP3BefeAw8Qn5EFsIP45rpAUo9Ud6rcPlVSWLpKD8QB9Xp5qqLkzNrGspWGdhN
eNmBDjkVaB6w4lOtiCqH4C8fbXPJQs3WgEV0MipujTVrt/rQOrgszK2fYYp5H/93
4Jpy4s0I0y48t3ooq70Arlsx9UJ8MxDR+7kfGSneJqK8TRucBC76K1RHRREqtaUn
PIZ+g8oB09GzksVg6GvhFWVbYLYo3ET7+09grdGs9sjsTpQD2whQ03ED7eqeGRM2
vzFhZT8SWIzdNoLZrm4Xsh1NfwIXXpfCbNmMhisg6YIDP321rBipplt4z1bFavIf
/88x5fQh+R0scMntTjPFNLZZyvfLrZT93kQKwG5hQS1t2y5lBekzQ6zQpNjtOvYV
J5rvI5xaJ9qmIiA8K9e2+xVz1ppPnEgQmmg7riBxpKFRqywkcSpoBD0ephF7LjqZ
vSML5C6x+XEp/hwZL3yj47rlVOjoiq9nrgDYiitPS2Cb4lGjS0seRQ0Yr4dLs6Bx
ahPuML26orHkbxmgcbZ4WmzbrQW9QczSzqkWWSKqVPYNYxuQhxB1Q4Ltff/HJsi8
Hz359nZsiUi1Yq/fU5hSOSv2Lsu/b/uSH2U/Wk9Nmha8hSUt/45CoHfTVIa1cth5
WweO7bfeqVydM0SxgSXFUrKpG/jjYEfkp0IxXYpsVVdYcxVdLuLNStlfpf4b0RuM
GzNDZzuyURmtPf0AjhuztamBswJls/4Ojcfjv2otWZM2dDWfA9gsIgiYfBYMwiyC
iZbUY4FBziVKYWu/eESwhMQVczcUfzWc6Xfre4Tw3T8bG1NphmogJ5ZsEAg0J8R8
b+lnTDaqIiqTx6UfaJsureUo7Vzi/JXoc17Mr2i8KUSjjTUCn16PMSsvFx9m7PN9
l1chFl3U3zoOlokZWIp2+/t4rlUmb7785agz2oYtQzq8m7EJJ79Fxa5qsyp85lVd
pnsPE4P9PLCOMqAnreq6pD3TIGK9n0qB6R8UZpfb1KG369uywKc1utr9AZpASz2A
E8eStvOS1sgGRShsoNuvDKeN4qGAmj9agsIfKltxwOpejflaPn0ID+NKz5hL4DMe
gTWOaeLuJ+QT4KQ6cJnu1avZ3BhonJAYET8XSCv12ksQ1kpVxPJ3lCc8YlAxi0hd
afQFEiP1CJqAEuH4T1oshz/CJOfl14wSzBct9Ag2O+m5n3y6yDJoZecqoxVXthAT
K026O1Ig5Bt7tE/XRuZSUMQ/wl1xxMmrQj2O8J9jfwixFMvECh0RdQszgG7+g1as
sk902UFa6bzXzEujAS/p07NFbZpKwkOCgxDoK/j1mjXMbwJIk+dPNvqjHcTNpoTL
2nXPiYLB4qe6Pb0BzAaoYpxnPYwqBSetfmFMC53jC2OBOOWlgBGXqNry86M/xpwz
AfwBJSPaOR3bmhUTCllrCqU9Ps6N54gnjX/NL8uQYESWRMkCREvGdWe3y4xNXrv+
tMCg9QQIoFLG1RpVu47Xo9Cw2eIlVUA81eOuuqKa7e31czucXIy+sBG8wkc/mGFl
zsWd57Ha/QN90m0keE1RjZkqoLSUtXhN/+6aO34bVXB1M8K6BlPNYB8wBmyLu0Y+
69Ta5NpFzzqRepDpGG06guFtUhGVjtgQUbg/995gJy6j/YVOiFspiDQL4jXMMXl3
EGhY/MgIlFZOdq8WkeGMH0OYDjvtLxOGx8iyA9cK8Hw5ThJSK46bAfsdL7LxRtIP
HBCLh2wO3NwOF41VwwDcaAe+QXeUMSrVZ2D4CXKolkXv1JCZXi5MYaZkbobZpoPU
b/bcNl09onnZZ+OoK5DNrL7O1A5jet+CQ+x2n49A1WmZqsG1lvEzt4k5S4WHQyBo
Jjanr61KM5278XU3QxpQFTNBfCBOyckRL1Kuir2Uf08yiE8ezOYGw+2DC20vnsXB
2feLsFqRN9TE6jnAZ/vIIvdVeOspv62/G9MJxg0gM68PJ+QbIROIO3qpD57OtTdF
EuTr2Jch2ytA0W9vE3NTYeQHmxpl+qWqT8iR29vB5/pLWTAH+G1XP+GyQAJi2cas
5kBSL+dTHJwHfdHyM6qAYjgOvQJ6xwfwfrcJsH9TgwawYoxTMtc+ONgkLAwiVQEC
MlEPM0Mb/8TzJ2Tu69CukOeSBoIVGcYijDv9CoKsJsiHGh+RNHHCq8BNwcHUvGM5
qfuAkdtPebhRgOmI7qc1jzD/iBtBq1yBoCnkpF+WVEaA7HLWOm5VtrPUJFzrVNhg
qeZqNsdBc8aCkUMeuTOkea0wlh5qgQjy8wVOd5tultrdd2P+h4M/+Ek6t29oHXmv
lu80MPW1geYc+yZnguOI0rAe+8xMMuPs9SMmcCCHYYFHp8Z85d/ItlWAY8QYv7OQ
Wpk6c7iHB40nHYUEGb6ptZng/WcPC2k6Ds9SdhnUg29r5ooWHN/A+Gl9AxlbIm8b
YBuDaWKTNXpjrqiyTMK6wV8C5EFne3BZU2NcHo1eMpsESTFQHJjI7Aj86BNzhG3H
4Th8tm6rTdAtUv5yXVUlUaETTClPQH7w5UfTuYwIp3GUHyeubnIyo8byf3X7uaaD
PvBW5rl31vGSeZPCEcAufkAa84k+4N9P/a3Ur7N9V1WaZ0hKIpyWRvJTUb6M9N1x
CT+c/WugIJCropnFW0r6KVI9UJg5/oeAD63B7Iec6ylKrJ+nHzzCe05t+Suus/3h
2XHBorgcXsEOg0Rj5QnF9UoUAB5Xew51a+0WrjLAIMVK79046C56TXV/adq9zyBh
0iiXh7Y0roIPftc65RsYXv48xpq+5hH+A6naMYF2GcrAaolfCxN+H/iyxJLORoe0
dbjtLfffgEs+W5GgL5PT8F9+vxYeTKWrtF8oZKr5I7P6fMUguWiBmF0rkykY+Qjx
a5KNC8CqR0T//LDzViJeKYMOYpInEcvmWZ2b3onJdtrzWDHZH7D0mf/PqufdA16r
0KHA3AoPpSQaRWAQbSWFL+LyT9NIsmhZxHaAtaGRp3sS8ajn6bK6OLgVCiGYIWtV
ufIceS445o7DjXhjaA9ZBIdbA4iKEfJdvl3dqvy8kpQWKCeL7opODqRMqzKvKDbw
CpeBId6w8NmzepjguhjeInm+asriCkUsK6P9AZBrFD1q5xbijOSftZwlu3keNEL9
FapG3oD31lYWbqtnPyU7CQzQgnjKhAVqnv9f/VSsUpVZlzKel/bimCFLrH9SBNXD
yWenYqGrwFpvNygQgWwzRMa9sNIPYyPDeVp50+fl0O7iE8b2XMlxER/GY+cDNmuz
PvqPUKI8j1VmhLrCyiltK3Q0wctVAJpmQw+lS1CWKFl8s1HWrKWqsVC6YJjhSjbV
qbgFkRQL9dKnFrnlLKZS/metJFsfK1r56Bu2vXV5NCkQOgyiZeZcVzwW3EiBdZKb
cSscoYQIf6oTr+rnC2/dw+ZkETyVtFZLVkIXNLdqeImvcP3pL5g9Wm6e3JneU0ms
owb1ZE6dhqrKTThm74DXhtxy+NSrfqFLlROPDwrPnCjGsyUZuwbag4je6BC6CMDU
Xkp+fijLXvZ1tc1qNu8jtUPphVt8/T5eNuUzMVViuRN/pCspT8koPWyyaDNW3CtL
eTHOB3GWOHHbeLuVZbXnzMFHRBqz7CJd0Gs2KrWSZH5/GPqpbowU8M9REXtJu15x
UfzP3wdQesnFk+9jAcDTQcdGLKNxNunerktEQIdygrYGCwXCFiKlGc4uwCylv1N3
3gIsFVB5I14Azb+0rRd4PaTxdUAcLZvioAtcK63B0N2MNocICJ68pShH5AVENqis
b4hdet5zx2iQ6FMiY9T+YIgfOlVSlSONjg69FmmLdYpqGs2F+J9nrUPU9aI7i2n9
p4QJQxbH4CiecW1ZnfIONE5iDtatKnsarnUz4Bzv6KIU4m9uctWoyDB4PyuiqSxY
T5ooGeKjMESijQsaSWQ1xqV3fdunzVHq5injO5lZjuYY2acz/ocGnIYwGZhOKKHP
B3SNxHgQaShnAC90tXFuKqzYqQZwCH3WsEMxN7BnLdvzjxvUmeyUX+EQWdsx+RCq
wiVeg1plP8mlBTfAifEsCxXjKgBfb5faZBuWXGvBOTrtM8GteZQDughVst5oo0Br
vygHloo5NLHkWTrsemAzBe5S++vsEGGJYO4A2HvNoO/7zhiniQtwogPoih53HNJ6
PN7//LiP6Fm5WysFrkpbwcDt30AvYXNU8jNplrndz3rMCN8WIdG1qlaFiWncYiD/
pAjEfqTdzScI3FvDfM/N43M2D16VMX9aRV+DG35EU+0KwTV1h6lWYM+SiD4JvDgH
Dx7fODpp4ES3NfYciPGhV1GSt8xLvrsyWdkrUAALM7FrkWeNiHegvMhzchlQJeZb
3g2H1oqJXQe3r9GwN3H1zZTcGmQVd9hpUB5ZGxPM+/uFH/Qqk7LnNVw67ZVm+Bcl
GDzSfCl6jjmZhg4zyNCuYri7mKokXiZvX1P+415yMkpZbn73s987QX/cdkbLfWoT
47dAe0QE/xLxTqRttgaZ8NqZbkT5QnZ6lrpX1GcBsLbfAqZ1qFJ3TBIjcnEnOGSU
3iDQe8VBpH2Cgn8IcpUluaOZPWFL9I/3QF8/QI9vpg57qLXSDe4ZQUnrWi6eNb69
YBsQjTaXuHL9b8JtSNN3vaFa7R9WPoHZ6OTjU8y82fE1ZudwtVN7jye3wLHleCBJ
xx0ya8mtbMNg/lj4K6jI9rG+aL91L3OGfnNIP03PQaxKXMECqQFtRqcJBELwbesW
C9UMlxAJA/XmPegqAAXUWin9nszHVHBzuSMVnjwKY3ITHqk1Y/3VpMzLNC76wpE3
FaZbhVeiD/okKadYvkyYP0APPJK7weJEM+ZL9+ncl6HNzvfcK8+rpfAda8nNBnAo
wj1/IjcSDTy4B32EDStn4HnJsdOPkNCi9isZg3LuexrArictfEFW5D2NBRoJv1VG
LT6oTr2NO+Tc4kOirWSlL8vnq7XTJNuwKPq+pcu2g8Ys6BPISPaLyn+qOK+Wjq/T
oEa7tPQMRwiyInb2z3qSU3u9sRL2VsnxVoU6g+x/WkTTJAmHgTLnVS5W7QGxSaqz
mDhVZ+wD6msf4e0Es83jTmxzY1qeQo8Xz+lD5TtfEUmocllfBTJZvTHms1rB9vrN
VSutoJrtcReT9nJpe9kc+0saEp8OzelB/wyEwsriHd5oaRMQcqfta9cloXh4e1wY
qYp/lfKucEIiLoDaFULJeB7D0FAnXZYo0ub4NkZFaHB1RwyPtVFF3zFZgdJUjCcj
MX/DKc0Py3G9cx35RRL40jU2zSF9T2aML42gOKZYLErjlAayGRgj8KDI0bTvbknT
5nFo1bzDJ/t6toOK/zFnxZw8I1rPRmHNpTW4mvKmVIPmYMEEfuR7tDh7KfO5rxz8
VgDa6pU7WSEWNf9+oIhNwaIu1xNpgrlAYV3VfDK3Hkcpr3bGHdQ+MF8e7asDWVZY
KBmElXG40H9h0P1/tSf+hrjplOG+5AUbSHvoQb5knfDXwJBC4/hwjTVIn+ZCvjj0
/ZMAi+ZIO5tiUP7GW5m0PAyVbWaENuHkatoZWjcRWAR5BsqAvfxBTc0UhXY8EUle
dJPpMTuwZdm3nt8SnL7tNl59W6l4yUhm/zL9IzgttBZi9NIQVlvPuYLKXoEG8iJE
qWH5FFE9m4F1tuFAq/Tod8iehV51oKRUdeB7o/XeTGz5+rBzayKHzmpQA0wxphgk
HmDOSMCJTZt90xqjNomxKAR2354E2fXZ9yhJg9Gu9MqlndKBHvBO7Oi0FhAXmS/P
rGa1hSiM38Ej2yWxbbOa7FcBmw4uzD+9CxPAQbKGGhvNExCY3abDDWtZGGFjxknn
mtUNar04OYGS/YtFcNWsydcfqtEIhkXlBqnPHIoCtlU+FGnLh3QC9C81r/AN4RSi
P+vdBxBUL/aAJw9vCS4mfloEODAVdvSN5d6E+D//QbWsGKwqtScuiy9Tb9QtZKpO
nbyEFfB3nL3jq0FY2fF1lPkVGRYroFWiqTlHEGD4k70ZnjFseUWl0/klLv7O+neq
eaKmRozJPMKBa80BnHTFgsoOp5YSnBlaH3tRkPk/78rtXF/CicXMkOLzTJPv6/RX
D/0EUgPmK51d3ijK5RoIsawPFQEK677pDiujaAzWOu8PysKA2Hz4E/Sbtn4keZuC
UayWOEqND2kfkrC19SVEIIuyGNomzwOdG19i+6O/6dSPQ3cT7ZhEf5hy/LF3zKHn
nnaMQc1WN3FaXCoqBl4jFCVJLVtZ+u+oICSpWQRwONp15bh9zUdE85DcKITtHPde
E52J5MMqy46XMgLeUgE6YfStSVBGPPJ6VGYxQSx59qHxb5ELW/Ovm9WG2DtUR6s+
jSoXnxBF1IaMN4X8miZoFjzEbQUu/IKKRNp+7zrJKCMmfV1iRQbjZDt0e7v0pidz
AIMLfk0nE8LEgfz2tVbuAD/oeUS0w29WooQgalKXax+47TxxmfqvOU21AT5RAJxR
zoKkbvDQZCIBFT+IeqIOUJwpWcFSm4Hmfm3v0Yh0DChZyN3LoVYhVxjjdHHHIDG6
QLcmNlm5ar5hmr3MgNK44SL31Jw5VkSVfcJ3+bOZbJCOeapO6vQSj4LNz2QtTN5u
SUxuHGzrab+/lo1uIxpJxOJbwcFsOEmhYZKW27LV0tHFCUvdHh2szpDLNqX81y4H
oe5m69tJYoSDm/rigkWFXMWrRt0/jTgwrOTj11Rs6ucPlIN+Szb35L3qrGHapz8e
fArleiGAHOJowFfL/sc+Sox7uMiEbUSwzY/3XXJu8aNE1KRc/qbvbDcc/VZOL2Re
WvQVrqFKJ48v86RcDCoJHIYDH2k+QRTgOHCuO5/2rar6zQU/OeI3sPNYEExLJ0jy
S/fhv4zPB9skswCdF2q6CuPMzDIsGNcJJ9sbPLxReHMSCR9Dia0Tb/mTORZOHFyK
WWyBYr5ngdYuaeLv5oRXbtFrMOAhAEYrb7+YAv30BCgaJx7/z3ScXzcE9yXlz1i2
sN0/Xs8EkLK6Cx2NUkH/RbKfjsP1gFAiHyc94GSWl6Oe+2A37VtY9MzLW3+zLmVW
ylwwaTCF1QbGDrKN3lFDbulnflcLMD+qYM0VzLWpHGUoWoJBynEyLgm9Z9qv9uXe
VohZ61T4opTeFK70k7XNCHe7FGhgjevwH0fKx5KogXzXsnMZDB5DVEw+XKfi9jlz
xST3dkI/zFl/rfKNNZpxXxVgyporUV3kv/zB4jDu99Gy7Aw+Zu3v6agI8aWKatT8
PlDpS/k1pIyHm53h930WmJYqKMllOnMgzaSVEeLRwdHf4h8cdR934aEoU1nffB9T
eDAMax2g2uTjVjqYbriO1vBV44yMIypWINi663RBUfpViLhoq1TvVlZqbKH2hFti
fJKGZMZTERYkHx+UqOjyOTJFK5IKWGP9YjvIf2kpw1+3ADipv4+F5nhrfPivMUzc
yNFy8Rs7nBZophSWFd1cAeOc5Y4rxFMf4zp9fNrqI447AugcJCFra1x2RnO+gOjJ
wYHhnsmMyF9plOI9rQz332L5BgEYMtgADFR40Vof4LdnpoyxraadtIF5ae2S2tJb
8v86ebckYR3I+3+/+yEHmFuSejBwFl4krOmPhwpk2A2nt/ML8UForlLkzueP1zdy
kqCou4V2odRoCH0H1M+Kd+cNVziTxHer17mkpeSrnLNSu+u8vgG9e4JlVuqjKoXu
4lawobOnwtc3H/Uges4blelbxTRcSHwcADZsPMEkqZWAizs8aPdFD+pRev2GrZBs
NStXbuWZa7Lnme2CQwIwTO1uMNTm6fZFN3KcsUo1WfhCOudiNoJGOl38b+KaQp/y
uD5gZTvsSbLWJO/gnGMftC/cKrwZAJXFNSW3iE+Wc/Yg+4nW4pTdaE9tdfmIvU4T
AkFw/pb28BhEY8D15df7mfs7FdeznssV2tcHFZpnTRz1hRZcIKhj7dgQJMocS91K
NC3ksEDSioSTHtzyvrPvGuWBkkfbqC26rK5y2xxDosBcbmmOXIk2MOWu7mfNncdd
Zd06gcMcMyCTK0y9Y894grXD8/XewPWVlRz5UoncWzSZAzqfcsnQGhGSp+mPBj52
RBnKsdPe1Ve3l+rsIEvjANrYr2R/xRgj5tDCbGu2s1g6B2yk7YnI/rcrzLs+/Q3O
EOdhcWpr5WL0rBiUXAQOhdXaU2H+K90MEJKt5X8iS4w5HAISIuTU7HVCO4k6guOE
M8IONvcX8yK6FJhbWWutLhG2h5IxtW+Uh0ePIrd2BuEiRJ9c0gW/wDx/QsDmOz/x
oAyt2S8U8iMnKHKY07cdWRSAsUWkoWxq1ZiqrpcwU+j2WbJ1adqfwlczZNBlvwl0
QSJis8oTAVoM3Ogatv+2z2fm/s2NfvGGN8FREZgnTatlm/3Yd/VcGHeJNMXU3/4d
TBUk4MQ1aVnYvwjALOGrLEOYe3NuDIpo2sDdC0EqLb/fxQXxesBibrxIFDOGyHhX
619ngB0DCMOkTQEjsCJe5YdBh8NDMfU4NzLlFjC1fbunSOKiVWtWAfvFVOsM6oQG
kPl/6Hg3K9XcjIhXPj5p4ITOL9sZ4GNRlm6nPWPT1qznm+COSyRY5T8zPrWO2EjY
LFFEXaS7++aVTrw03DwFcgtPImYqv/2boqFKZBLMBr4Z9/cX2KVwp6RSZwPqUWvb
tRM+ZFrL4rfPfkjKeXEdq7fUNkW41nRB1058bNWCZNH9HM2N5waiEcmXdvTGkOu+
P+iFfZRpsmGqeoLhQvzRd3TPt0xN8D/Po6l5GhWWfyqKPwoG1ZBH7B6qvA5COpOy
lVjXUm/xV1eyK9MSp05/BACU8A8//JXw3heRQMyUFunnZkcl+7JvlmYR76fDVDtD
TlkSSROtopxqZLiX1/vVQGIGkkO121F/lMSVYF8tke/ACVnMCWweUjcqDSjA2f+x
FuDVn76EFn7qz7nbvC0OicwazCanLoZhEy0tlukXEvIM44326zE233KGobnYipH8
2yYaYCiPABzQ/m7iHfKWw43jAdoRsL2T0i+NNN+2sCSbdxqJoktT8ouVw76l4O0H
5xnM6WIHeEiw7D4OiytCpo58vaWkVUIO0ebmUjhReJ8iiGY4QqaR3S6XId14AEZh
L/O6vyQnQheOPHYfdvZbEaK3z8VMsXezPgJtZMI5sIlDw/chMhR4qdvygL08Qfuy
7NY+MIzQS5tegeoEsXPvqa/vW+54bMCt5tD3OfqLcHTIK9XyDkfcTzZTzg8Wzxdv
xYUlxT+1OfqSQs2j7i97S1GL9MtrR5bH3St6LyiNxixM1l0M9ee5ThRb7/Xygn2M
Zbj/9w+0FxfPCVaHP+G9dOj3/SGaBkVSsRSlgbna22wgk0tEzEQvq57qzXv2uO7g
oQS+mYe50UMwvpXFu+xJLUS8v3jEnbrOxmrhrqGNFxPp5GkWHue+MsBrAuEjNad+
/7wEGMh/QTiq9J/GbPu1f/Cz9Lm+BzqjVSvKYrGTqNZaJuhPUwOq7O6rwNhSCbR4
MIZRsPcbd1kqbNbw5CWsPlFhk4GyZXO6+DSNt9lY9lJ9zh0MGi5f1UDrzac/GBwl
tsAuiepD15VQ1+jbeZvsXkKmeF0D48tL18hoWSVbEuJPfpS8ZRRODJ+TFMoODWox
ItKc2mwbxG/RdM2fb+IodHK49cxSCTZrLM8rAsDph6o4am7hO0lCQI1Eja9m9UFi
W46sA5pWhST9pF33riPoK/Ud95aeHHOCCuy6UY/DzOq/pL6ThBdj9eUroJTraxbK
mWV+7Q42uKavhWP+fKEfL2qt6ZF5SuCk9zd/y24N2S7rwB21XIIxUluHgvfGtxrr
Pu7QZRI/YJX9i4WwjgKlxdvIfPCeVckms8HxzaZSWB1CPg2fJlyjznX5S0qxj5wP
iduD9I8YSW9zY8fSy8xYf0xSawLAgrYj87EzXKz+06J+XfBmYS9cGDbhgToOhMzd
Hbu1f4DAY38NwYjhIdM0J/YmnW5oPl1gdEU8b7hrCKlgu0qx+waH6WeH7ZkU7c+Z
Lx5bv6xc7Q8bp4i8gh5gkkKpK/4KLEgx4Yu9Vh9swHIeGw3X+wr9KFzD2dhs17Zn
jF2lzh23NdltajTwEktGar3EI6a61hI0ROXzQPlLpMwkU6CTNiIGEsU6aSV6IM7H
wcfb4dnjxL3OHEjRAkf6Dmr+HtEKnQuvej22kAHkhu5CELsKpbEiND2qoKIa8ALz
fcVmD+RZmUTBIvleTyQ7qSdKA8wq0Ojh6TBvp+lI8IkK/a49xhl2Hl9bSiwj2Mjo
9n0RTnSh5yDQ4l5Yy3Zr3I9wP3uZS8V9/1Yvg8xNhRitcug2/nTt4XooALX/ebmg
QBc4FD15joUgVcOlN/mZ+FgWQSJKfdsBqLfPDnuaOc0/4gl3ETGQhHoFwnXJPrxJ
Gsi1mtN3dp5g7TET8NWh9jGdF1eolASMGbZXeFLC49Kjr2BzV3XLAtmWCRmoFW5W
t+LE3PRbMEtnxld7/GmZcWyS3wpTbjbDPSCMqQkJEwbnEaVmY2c5g+SsgIbv5yih
Ogfm8KN2NZr4SZNt9CLKWkT6QSpH7YeQ5q73IZFwEYZVSLyHnPsz9SacPGz3JA5P
DZShpCZrkn/m/YxO0DfUoqZsDmcXKwTzc3K3zyrbEWQ8XvOxjnOiaJ5iDBcueuud
Q3Vnlx6ONrK5/dylrauEn3XnI4bfX8FPA+F/AhkCe+Q9Twbpwqryzz2OoIUn4KHT
wEWyjs4Z6GaJpZP01Uk46zD38m50PtXH2lD7SKLUC66KzpCnIzu5YylvHn5DRbMU
Y5M+I0Wvuvl3FtdLb/5gYF3m/xzGdHpcp8mWnRDkpjYL6WIbC9xvUSVo5C3KJus3
qn5kZon01frOfbEpSfp2CKiEvutthOvTppk38CGnIoW7/gA4HOcaaJucmxorth+F
gjr2bkhOPvqmy3BOaRToOHWIn3Cpy0algFteA3PnhrZxANhPq4y38B8C4tvJRIg2
+/YgoWWLmnSYqi3X6i+ar9c7NqHhNNfucl3cmqTpq19gQL3BhdkLbYikxkigIG8Y
84sp5M7Z2JS8hO/2/gGm1Msrvugk8q4e8pH1KOyNVkzp+xaH3gDfDCAk09ZRukIE
HaCSvy5vAjbsUIkWR/rTkOEZBBljkQ+4K8jOBb70hgkr3xomn7iVgQYYHdtf0m0a
gBHk6Uc0ztht/maazcMWyebwqllDkXKApnezGFRc+smCHSMaIfAjEKXBbCrG4GPI
J2Jq5ff3zgvluwWBHDpQsTDziGE6xlcSBg1bZRS/tpgfi823OC9eepeletSyAdFD
X/N5k4RYGuu92Xjt0r0b0uiaKRveyRQ+FJV7BoyDag6zGdLkYzh1lMYknL2g/JZa
fnIstDfKWqeBl864w0FNJpjdD11bMBCMWPAiqVAoz3tYBzZMdvMgsSuSQRTrOPBX
D/BVvPzu0UUQGK+5gKKEmKjqQgYlBnKtNbI96z1RTWQEUVJVWqoL4pJ1eTU7zRxY
pa37iSWEBFpFr/BQWfQV1hiSJVz3OfvUoYh+vf0QVNnfjHQ0Mf8mNHXyF3uwekBi
2WosaoY8GHY4xADo3U5yw0crlUWIS48BZMMQYnklP/VaQvrrENgVrB9evZV+YND0
EBoNkmKcWV09REyH0yd8iZiCfN2Mhd+DZPprjwmLanTfqB/7ITbAAqGA1k9ycnej
PUlIUJaC6p6wN0L6xnfnViLgnX7EwLO0vJFbmPbBNmCG83tXQhB9u2XLfBw2CtwP
COk8F5ehSQ3QKM88KnwuIngX7zpFIMwgSt9Ak9LU9bo3BsL/Bx9fbSbyTbsU04z6
qc2+5dvj91abFCFBlDkDQU80PQacb417IH9fRzHobRK5g2+0lgFMxNEH38q477u9
zG6+zKxCqQmFLAJrtR90Wz/qMJZBVj1fVdR7X82pdpLhg99R5LfwDuPtnQf1ki/K
y+f/BwGvvTsgebWGSaQ2w9KWL9S15Yr34tP7i5b8C6uquy38OLJq/C7bgDxz2qMD
Ydv61xPBecRoLQDD1s3agGN2ndOf+wz412NCdA7mINW0si4b9+1JPPHXvO6su+HK
v0hktW4iW+5LStczfJCYC8TqqDzzkqtie24fRLrpd4KneH0Z/gE+s7YvTFqEPEpP
ySLGnkAleeVrH4q3rcsWLX4oj8MASZ1hy3BX9jG7kr+lVAMjYe4YEIf638iCuUbP
fsMboi1Hr9QQDOLZ7vb/hvwnB5EbpQpf+H20Ao4qzVmXoyo4w2SE/4vaYtQc99GT
yzHtahzgH4+E28aBfSfgj4QGma9vercH2lKPCWO9/2no/weg4noDMC4P0ddVBbds
ER1vfrOoIImVfC9k0QkHjNgt48m7mkiUUqb+RdfHXyR/VOm36g2ip00uSqEBotgd
rGcospZ62kzj2E/kiuRfGXpigziRjVkP6kjQs5B8fD1vT0ByKR3ma7sbmOO8nC3a
jHO2LkLY2XIH+D7lISFttgpt5bkhNjjAy7OSycaY3CLGDCQecRcA5PKfa2inSDTJ
0aEbcNa4P4ukLus+ftThEKd+508gnuQjMyTyXAg5ymbLHjDDuJ5YbKO5QWb9J+1/
+Qp4mz/iiQtFIU0YgPz1xLW+vTWWJ1gkaE0yNmQBU2JZsF0GsthBTXoDDDacUZyZ
v8JpYbWKbBcE3muZqXFM2xHBohUdmygMAsp6Ga8B7RQJAYLmwGza1/Zlb4eeF/JT
l42X6gFb0GScbivnEey8Y3xnfOwWJpb8KBGLScwB8Slvr7yyE3IJ1E1wogeZ7u95
gDO3aAfBN/59s6nhJg+/cjzl7EAI3yttCh1DIvJOZQXQVmmKjkjrPK2C692rYZsS
RqVYoNe6TwIVZ/Big//N5XgNDVbuuVpvS2sun/tNlwr+nWgMcnjAgiVXSoKmiJur
h2XLdu8mCa8Ut6ZxCFE9wMVeJbXQLyWoxtMTgCehe0KF1EKvRml7p2SD6KI/vGWl
LmcfljbJmQBejL4sz5+Rq3Y/LFy9XtwYEFF/QA0Tw7K2sI/auvJ7NN84XUC/D6ae
ZFJSE0cSd4Yj7BuTSkbbM4eNcrCAbtmJxMyAJSO4pNcDRev/1FEwi6g9Qz4pqZmu
j1Bcev1dJQVtTltIc76l5o1vuTQBzjtQU1zlHTtpw3sNJoSVGdFqpGWdaVxJSHDM
/w170WtBg2qNcInZKUv8hqikkovv9MzNL1iVq1AvWqV4KtYTMR2F2uI9DujdHhfm
mDdHxpuHIz/xH5OrvlLcoobzM+jdcad3QDJr+Gk76hcT44hXJlcRSAIJrOXv0IIn
s8Ley73TruB5r5k7OTuuT0Jhe2TOhP32mkl+NmvOK0eGs/1cA1GI2Bv7Ei2dO3QI
1qZAXsiGNoJY+Gz5zGhf4JUE8fwM7DchLNAe0OvES6hCxXcGR7n0ojPzRCrZKoMW
fCHJpzO1rSJbxoa2SKdYDNRQRYC4rt+nCcYgVOLPKeYJt/aZ/k7FKxvbXOZ/HLOt
cnKy/AcSlh/01D0q8DkS5FcuDwHQSOYc76Ng688dzK5DSp2twNJfipGJnhTja1rS
UU+G8ydwTZpvIbJ+du+eJUG5nWBkKC5/2xgISVeLbR1Mjoe5dBTjavPuc7EJe/O/
8/LnwOvpLl3weMB5ooVZFTIDyo69Qf1+u79eebw5b7b+xTUV/R3cZxsk9RDHQM+/
FY2hctsnUCLWii/l+cFGfewtvqLGuInIbpnKFTAfQtW3IOCEwU9/uGBWOaAXDtOf
C45txDCkwxKlgqyom/TPeH/1UTfNumURQpB8NNSaJoM2e+9L0VCO9SHMHuhzLCfO
Nx+tuASrFsa/iXdSNhHB2bBKDTonAPJ1F4bK3i2ApLWsBhbZCzI9jhgDh6mUg557
B180p5haBfVLo05MtaT1LGu2bdCIeT1Q57csX3ikDrdgtdpe1dGS8m8eqybPEcB6
A76h6+bgJe/+Z+Svh9hrn40q2lMhyJHHAG/wdWObK2OAeeLiSeaaeLlyl02iEWfk
ryClUBu5amYZZ6Diii061khc7neTKNV0wFHWMzXPMGRAYIpIz4YSt8zYhT8FZbZo
Ho21wi+FWT3gw/QuFoZSIveoMahMyuEF8arYmN6nUwfFElSR4ZR4EEnxIWO3YqCs
8LRibZLLEdyRcxZqMSzgXUYv/mWaRP+ACrSIiJYJvCTX30qwkkJhWVE2KM/WAit1
/HAbjDeNRzAq9+7Hjp7lB60+Ac7udDsPm0uV0H2OQ+GRvJXOar6V+dc3CCj4OTwn
2I/njN/NsDIIuqN9+10cy8Eqi+w0L4xIoeFQ5fug8W+VnrWwMqplyWr6/1Z8vTot
JQznXAVvGcB6PvrEZ75aH+22JSIcjF9AYvSS8tpz6C98VKH5iZ/4EfP/AOPUpzt0
8y1me+eAVNFUGYalnboRlaeddYxvPCJ/0KfhU0Zxq8eWoZl1vH6B6km7WL1qr9WR
YjnsP1o21uWTzmB61WjyU3lCNl68csIfZY59zwWTAYd7irk1lffE9OdopIjpAWQ5
XGdQbo4Syy5Aup6M1wYAsom4YRvcEifXXr4m/TDBvMzRO+891dMxFHzvEj1aQELJ
vGs3nB9meYyBnTNwi3hS5CGU9bN8AVp5AcFM4vJKJSf/QUCPhsNSqURemjE8kfOu
aO1FnAknGC7cd0UnuoNrgEtA64DLR4k8ZtsvlwcFzUd4D9Wo/PMJdYfaOTUuWN97
B+G0sH0klTz1qoRWmqyIB5Bla/z7rFQ76GRBgKkiOG8WAGjYScoETPL53M603iz7
jGKDnyVrk9TqIZeZeeiSGp+rhrwxoUQYOiN7n/upjgueFsqyXg0J9DFShQvXkY3+
4oik2cueWkbX8aI9JMBrIeHK/Lph8E2iz9MeDOfLXEHT0X8xArzMiigM+pCDQtQ4
tP9H2lrYw81chi+rAPewKr0jKdWiA9d4XfiRheHEzLbhtKnBvMWNQJ8Cf5PpZKUW
RFQwIhUj6ydvib88tAh4KavuzgBwxm/hxSNQb7vw5kZBZ2Y4jNwboeXQH8osgwKR
gBPtPl09HPnjewyWDceKE/2QLbxcbNGPzpqXtx0ByzF7Jr94NjUYUza5P2fJCarF
B1yDssTSugxo8/o75Epte3Lhw5s38iBWt4/Zp67BlFu0s7dMLv1xzHnpY4+lT7Ik
QCAOgIZm/rh6at5h+6v7+MdUVGWNESz6C89z6O06Baxw4KThMdOHLCgnUuWbufh2
UYB78eUKlGz3/dVl/iltihWDQE0dCkx5nC1+VT20dfdTy2kxyhaBnBKMAohvlRgK
A2y+atjnBcYmsquq90FxNrwei5IMFd7Cc67NZVytl+vWP4sruOcWr71ZnFnBstQe
QSReejEA/aI2Xl/C4r1LYq+r14lJmzZrzRIy9FFyA+dK3anJMr36jg+NpwFybqwO
9LekQcKqkkiyrM0mAIu3wHJPwpoOOJJDqlBrz3Fym55NhfgiAkSwIf4jDFnx0GTI
rNGnVe1nngCmwmyGbtSMjDJgGQB7VYaAFp0o4wLyzYuHooxVS9TAvbYeZaYtKH2N
J0gCYLIgGpVjd9APOfV2g8jebK3gI0YbEOS17s7D73t2uB0GVeEdS758iHmOY3OL
2gVxY25OKUZqGGjpSpSkRH9dqYKkTT/78A/n064//fbWtH56LP1I0iOAHsCa/cz8
KrEUg4thVzHTtJlIH1Pbx/NJ78ipt4kKJ6UIVoYtmbrFq34xj6ZcQmsrRXrkKKGT
vvFGn180levAQVaMllShiY+M5+sxEb++XSZVJs0veaAiL6ARpeurf+1qCf4TXtZf
FNYjP8lvtz1K93BNjlOA698ZrPKPEnLjxvgcCy4cAu7EkALLI1vLwYmcgebIa09F
bjeYtVR5gGVw5zkcC9/yqyIJES0TXHVw4ZWClxnOK4mm/kYxK2rxmsCiMUgsBElp
6Z2XsUUuRs7DymJnq7t3qlfEzXVGzv2tWJkHeyKpkAazDVasg569WmzgWwUpzrI5
SkN7RiLSC0EiI7MY5vqBanp/QlSTB05G1W66Vf46BY6+uu0+XLvTH+AMMHWUh6We
sy3yI/va7Ndnnb8HqIXtHMAcroVQDoQRqjR0RRqJ60DCF0JRuRVErmdsJ6zZs8ge
tB4sgiF8U5LOElrJAd8pCAp3JjDwDmEhRoKeYwseUQstGPEOc1kScQIvJ4lVFd1H
8vqaZ0XLSQm9ezzo7a9K9QU07rdwG2DhyvsIELcd1tNMA4cTY5K156hSV/VELpUp
MBGixJULpVRLQ3zp3Bnzok96/Ak9bVrzS8Q0KOMfkeI2A5kUjLg9DNYYw5yPviHb
Nq7rUNF4KaqcWc8uztksWewEUJVLL8Qzj+vDCxPKJtYPyeRmCsBED/hPqzgcYMGH
gLr6GryRklvF6G9anUobk4T8xm1nvlU37JFg594JZTWKYTofs7jD5Omw0mRspyH1
7vGJVdVS4gEA/g5jbfBOdDegsByoL8a0qKGhTXI4gOXWl40mROwAQJ3CFMuywKPK
sluogh4t+6dX38Rdpn5TW80U+EoWmWao1VM6auAb9PmZKWHVAmDfhgKNxxpmhgOD
nKQyr5XRKodfawcUVZESsO1zYL62DjUFUYBlF4VpsDl8MiYQOZb97Xnfyr5YuAw0
NI77R0VgsFSrsLaZPZpOQOw6fyetlxWduAR5CW8BRFfXXAlgVmIDTP/pkiumSUAC
Y1twnMOQrxIH7vTWbnVyl22htS0MT52Gop+g5hsKJwa8IDbiZjY5x71GNeuyuSVp
TCIAHoTzdEdFUC53XES0hZP4VNTunfVz9NqfiXFF/vhVxB0GgQjtJNIrLFHHgKVr
QfgyG1SrLULVPhccPMpBNN1dYnXRtdkF31Mg8Fu56U5pFiVYITUyGxoaTb9oMEvM
TyCHUJFvN3ii5Q8HXK0BDlXyYJaCiU4vUvvJI/VOEZMVMbzaX1PyxyiEo99XgfMR
n5Y1DiZfQ9kclMdJxWOS5iZE/MAtdNFKKh+ye0/+P8UPkmr2KMB5Gerh4gtC5NdL
eKoZP87HURmD9q9+hiqHxUnYygf2L4b1tf2taR+ovfMifing7UhqsA3tW6VhhxP+
suJPpz5evn5J26/gWGol/lOy3uAr/65QyUVHWukQAx+6cYZ8DzfIAlQb3zp09jZp
0l7Z/SfVoSDYF34lQn+olqM5BD+XVzfWDbuNBT5z5f6ChMV+5wS/XaM1Yi5yC78/
+6LBpAM0bV8TPdTftj3jjS9iIuf10b/KwSY4xgLLaRmkju18CBigotEOTqs9dc8j
aUu73jF21vn+bv4dB5hKUauzxhhv+EfA7r48rT6E/sDlzdmijMZnEC8SV4sUYx5m
fDWlwqBTqPxMcdFTxbgfHJU8O1Bg4b4EKAiyAisZ3UeRaZ4WuTobm5PrYPus7ket
W4PYs9wxW2MoaRwxtbB3+dO+1A5wzLly4qM/vudvoxUYt7DeTYkaBvdEGZ8soZtY
hMRQnKM/HTa89QGlyN/sn5HAEbjM8M+h9RFdYRFAIAjhDccTt0674kmMmFLXod0A
`protect end_protected