`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
ddtXksX2+yylW5zu6QL2Lhnb2d1sD00763mmSITNX595NcHTEkwn0zB1Dry37fOW
FufOhVzEJp80NC5qZ/+F0Vk7Ik02dIR0elf3clrjeJRK85K4e3Hoo4xn7YbFUIms
l/8VZSb14+JVGURjfswrIyCUotIzlzVYZ6gzoZwDXIi5gQIBf/gI+KxNXPaKV+PQ
Ufys/12rjO6aI/pPlqSm0hCvftmBcnezN2hk1UeXgOIuKZnogjOsf0iJVX2aOOWE
6pD/psybjbnsNB6kH5uFTA5frkzIzkzl5d9+YDm9OyC+k84E83I/7/j+rk4L2dah
QJOvksSIzN867/4Qt8qYTQ==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="MvBXkzurAa5VTw+1JJ70nePUfoQXBvZOku/SMmg4TwQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
oRtzZL4VJ4iwysPsC8SXYCzXS8Fw2gtZTOskLcDV+1B9Nzn1zTyNtlo6lNICRmmK
ZRVu2BmCc2G+fmzynYlNTnSa7C0Cuel6FYpxCBlOuk3OF2tzAmLAuDyOH3Z1Yjzk
a0aHuoCdIRKv7BrZCdALt03JeUmXKPdOmIlkVGFl8yw=
`protect rights_digest_method = "sha256"
`protect end_toolblock="Jn9CQpRhJt4rnzZPRk+dOpzAubz7omckX1MrFd4p81o="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 13920 )
`protect data_block
gD6l00tciPUa6pDNTk/+t1gcgy1iCdpjTkA/bOvU9JA+cpFEv5u/7dp25hHk7lLT
6tYtR8HgwcLXTcx68BnPlzdPHkVIv0lwXo6yhFVkYlDWBcqD9ubowgKij0UjlXmV
p4anbpVt/gKvAYRDYe8Q5F2CQ8AIsxOuOcJ2vhCPchS4QF3n7+oG0MKU5ZyzxTu6
J69cyJfEk1dN1/jsYsyC20svlP5xak8V/U1mEDiLNggQjepkSg3xk8SI1qOHk1LT
pcrGilCzawUy2ao8BnEsjnhorIj6mv1JAG5MqBzFPoBBPZI6M1d8ZV1uZ9CovJDZ
lmun4WaHsw6XyXcf64nS8EiGN7N2syN9YDVHt+cqOvN5IvaCeypvkN8swYHsf9Kj
cDY+hO4uwEAcV+7l7DC+jAgI7K2JASHh/XCT3mlJhSJSsI3Gv6WdMKAp2wdxgwXO
vn/J48ntlqFay+a4a0YLtUi3owgtIz5BEBq4+zxxrebLEzHt4mfj6lHCuuMKbYvN
QBeBP9P7kiSaxPKhSLMWBG4PebohH3gC9+SFZtWZ2PEdugHS7otqwrjft8EENH9v
xQMaiknK7TgrHXJIH4F7qQXn7C4thdAvb/KGueYuz6K/4IAiOcGX5EYQZ8OSv1SC
qcLs8Nu3dEjAlavUbtFZEPH9DljxWZ3VfedWZUuGCfhXP3ZQ7Wjq5pMK86h3ghim
W/z73oAaBfT4rjtNuTMeCr3ZUIfHB89ACItjDisSr0LCvkgw3vxKMDcYgRpTiBqM
cgkKjh2mpcWEZD3EYbtSF5GxNZCHHzGUJ5XKPHoSlO2xTHBoT0dqZtuAid3FvhXo
JU2Sfom5Y+zC8TG/4wzC6/fiKpjHBaGr5RlqOu5t0dqirj8JhEVzJaoGH6rqJPAp
rGymJGtw6HXkeXv7RbubXo5wpCSVzF5NSQAxJzbnjHcDmY6dpoq55UgVfW9RZhLZ
0uRUDaonr0lCmIoTzJj0+KaEJjRnU2bllTmhgghn2Uduz2Qrk7oCz/0kYpaX7FRm
4i9346/KBEHdJB4r+6XOqVZXt332dsjRm2VEfVgpe4BItqJi5AY8/f7uFeYBLRou
z0Jtcp4rbEincx0aBpX5a6TvAdzfLagwucOlZI/OdWZQxB4aw8egOC2AYCZYAnwO
uThHZ0yKyPB8GNG9UIbaRqK5d71+TL1TjJtkLFpdDL8uCjJbJMfj9y+oGpYTJaEd
wqWt0dz5UfvzmStPLS+nK66j6HKvfI6OCvT7ugMMrGy9whBPKAMSFewdPod6KtHW
O6nwnY6eLqEnZ/UTDVPNngBlrJ1QV7+Ly5HkmhlUPy695Jdr3Q+Aea1O8FyfKm73
35iPKgCpUtYxfxddEkg9SzKEWIRhUelnGVetgrKvKgtsCZD90Gx7rexfDOxwsPgT
sZbRSiEWSibPwo5H528195zC3B+B5U/pRWmWMgvdSVhUjWFuma0/tj4RZDww7Q3e
yGnIhk3S2TpsEyvWDQssB/C4HxIVdWIkJ77YQGbmL9GNsCkN/9JEtOSQ/eUIARwr
EvhEls/vEpdgSZ/M29IpmrXAkrn4TWCGnN5RvpWQEsFLs05nt1QWtASYlkXvvqpi
/DjoMfoHcTHGaDVrTQrWRZttz1dQjQo/XQNxww6HQusTleuTyxdZnaQIt9RWIBsK
X5MoS6cKLDKegoRKORkFp8SySDx02wS1Yp2DFIp+anN9awRnKupjjXJAnxuxUn7k
rV8pGP0TXDnUOk+4PFKTud8QwM8begR/dOUer7YZruKOZK7or/S14ivGw+1X1lOm
9j/yxREEhB9rIGvkE+yjsVVXySs4CTevQ7OGhdSIbWOgwy0OoMlcIci+H5W/7+SS
v8ciIdx7DL0FBi0/7c+/2gowD+r9ymfWabXWdhUlO68iLXKQLxmXKJufHNwXboPG
i8TTvda/c5P21mu+C3wYorIS9vIGgt8Mu7+2dFxkOfuKc+FXrMt+YvMMQCH6I+/k
QuGBbAuDRC2NDs++q4MUDEh6MLGzSu2NaNTmd1DP/lDEUCcg+knGoDrpmb5SEgto
vcNC4JP18Q1Qxtp5G2g+cStf3gnw8uid7BQj69HAbZiYDenHUtapdCd01hEjdpgU
BZBuqCyXsIrAayi23S5HUPqWtyoPuzVgX5Kf3dVVWDozc2xnuzOrxNib92AuCJ0E
7e1cbcgCOTYDEjTeVZd/rvMAK3H3AEO7zzNYmxGPw92SWR5IStZP0Fe+Qpx3V07m
fGzii7N40eUNZohgGUHXAiTOy07LskVPc+dhJabR8VUJ8aHoXHGTssRbzSUq1EBG
rfw0oUZJt2cduugDi0JX3JUnByenhsJFwIr69j7mXdBPw3Q6NvN4jwDnY1YGvmPB
7Lg6X1T1XsNPTmL5OalSkzjjXwHh5HTY/mBe3BgAra8/hIaeC4MDBOBdESL2Y9yy
QJw3/lPNkyxXvJSMtciYM0a4mNXbhwzSKGQ7uKln6WIrX4KgkNFnCdFsXLURst/4
6fgR7ERW3pRoI+NJnVOyxxrr7D6Gah6KMhRhSjWWU8DqBtqHE0EHc6ou1h1WmwXc
Vu1QK7O1ziS0MxymDQaqpsnMwHLpsSnvjH4Gdtjyqs8smNK1vIynrexDv9qtCT4D
fWi0x1J5D3AGsfPyqyLjlkpA6etZ+HexM4Diz7Ov/Gv0IDIvngNa78su//wawWD6
+r0Em9k0zMSie/74remgScija9+FIEewYTD//Qv4aX7ClTCpqYVIi8jQpTB+CbAF
dbha4qCPb3JFWds+drAaDA3rlrXDYzssTLdiWD0RvbCLb5kN9JqiX0tYjwwMxxh1
3P+QexZDBVipezQeH/2KI5UPGeEvW9jpN0bKp4w36SW64glbJURxk2fZxU4RsgLR
EoE85XNH23HmY0wGUGV/h5NbHOl3EcSdEdNlTykuZ6Vx/gKJvbFELstw1As1Pa6G
g490Dqr6Bh7f9ndEbwmx90mG1BoZk4SAlcJ5nhNByAHMU6bBxs1m+EIbe8RzOkAN
VuhOLzbaNy3C1U+C5nRs3KMySwTbycpao/jD55BcJos3UyPJaahGCiORCI1rgb5i
ju/XaQfPGomEp+6mMdGUPkCDBfupsQdR87eI8FICvwWuD53cNNIBO5GWVe8mNvW4
flil6PJV0nsc8HQug39wY5hqF4JDMok9lMvJd9dYI2xxuPT+ihV3Ncqy5RNcNNAW
3JMrPddYlPrLoRQS/peM8r2onlvzJW4zBWPwa3hzCWhpJp2g4x76xyDZJ/4Fb9FQ
BpqO8TSga+XPnYuUAk/9crOWgAYP5t2ut4Ro2bThAQ3D0VpeLCSH7u13ACXR6oOo
1DKmzSx/BaIbmgSeXOL0ZBWf/BgP4zI985CNraJuaMG1eqwfgb+UZXNpp+Er8CoE
T176rx9QY+J5U45AAnMS7+0OgY1s9OGU4y/O8KQM0keuO4rJcb/rYw+LdZ3yCIXp
ijjeQrh0Mr6q0Nl37NdfkovIM44CRH6O5K7kDkjTgxsGfsYfjdbNoJhbPfglZ3NS
Zs74AZfwAnmGEoY2uqsE0LiFdqEgZhsrTIoX+QtmYQaAFEcGcN9eDmgKZB1gnT82
lh2dK/0a03qHiJAfWGPOMLm0Eq7shrjBtV3mB5zOi4Qx2kP8ql/T9JLxa3jXggGu
c71UbygOVRNpTRUvT4jjXDBezaFpzZhGKnXC39c/EesBfZ6zYqWVSLgpfHiNQhqX
Qe6pKmFT2sgxF6pH6wgtdobruOdlcEmdywAi6WI2kAUAhagTqEBi/rYfpPcfM4ws
3jQeesgFgrQDtN8UaEm/wNJKu1FWQ2PK29HyanqWh1xIj95ggkMkhuee2FiTygye
G6IhWtjfcdnc7GtEZ9o3LhLT5yYqU+U/8SevEZmpNVq6+OtLn574HwKOJwQUavQC
zkuEek53I41q/ebGA6Aj1oOZfr0T0lDJRyTb1JZgzA6yDLn5UotcsSc0BdZ71vAT
l1Hjaa4byiw3vp3mkY73HHLStbO84wvzNWLOgrvAih4RqXXsoCC3pcNANZzDdHVG
0VSY22QrAekPOn66g3o2uVwsL9FpBMuJ6EVe4X/wVvgjoa8WOt137zamMH2AY2De
2c5/IdEKhhoR+DC8r9lSUsLmOzX8KbWtkJag3kmnf0TdV7Yps3o7B0lb7Mk2dgiM
ksPlHf1FUqkareGPx/KAMzV/r4hCTVozdX33hSUR6idosqwKv8XR/gqGfdJq/8Lj
AQO2fP6ytMOAmybNSRdC+n2vqdJzHQJ0X5DcIbyc2uoc/BNnrHI9G65ugIB6QRub
S+LIS7rIwxENX+Vor4uwR/PpINd6/5JEdFNwTMJH6NlR51yHOYsOoTcvN5BwJyKP
rSZzs3R7bQPR3ubpwb7AtS6vonyjCMjWPQt5RZhdQbFvyc7z/E2drkW6UK5HNifp
Uzzzpt1QL0GfBo6x3v2k9vZEbyt4+xlMhFV+mNcNV34vYqbCc/vHd2uRUrC1YATH
9Z0BLzG/aG4YO4RAHen26Ahcj5xJWJ3FWqHi5d7gGArDXi4fMQSk2ckqarsBvS79
xtRonAXf5zM2Hn9mSaltgwXcG750LsQWFgR3wujoLK4eX3d4Tu9+XoMEBV6OWSRf
Ielsa5SzYE1FZUDQiJw0nxgK0DOgw2R22FcvzuMwukkNyczzGnQNyxVaY6yEianf
sKD8NyhJF9/6ncLRCzo3LLcGjcW4a+wVad3gd1q5K8iBJXEQHxnbYyk1UH03FxNr
oPWIO3MoxDRRMlMdRIJbJej3+tCh6i1eppRrItCT4b26qxMCgwGhA2C11JV0CYXL
KOjqV2+haWZYOfFtz6medXD0JAQhiXCCSY0vePBsIJT3bl0yfjtmzt13vmsBRKb8
u6TQ2vuS9ow+UNjr+1mnDzrPwz7xTiLHfjbnFUnw18Pxmdi7rc1hUcGTxpUbmUj9
BDKBwY+TkBAaPNuSc0rM1lBY/sKticB0rDtPULKWsxs6t0eEtYzVzo77WgPzNoq4
NyQi1KF5dkLWhGQJeOBAp6wm4luWnVH/k52of6j7gPPu16FI/xowMbfOFstKSoBo
OcET6vh00U5ArKtDmHNP+ztnTIpW484JjMmNbTerQRQaSCZ0IIQA5nHBLBq+CLwi
N1i7WBanZBsqa1r1PGGFmi7SkSjT3evh70lKQHAkFDzCxbkJYdxXCiyKE9nO8GZk
pnsiYtPNJW/crn9nYEcr4CV+oW807rNEkLBK1l4cngyukcWovA2Gq4S7SjqGWmUP
mCk5iT37ZUolY67zQkm0QX/Su18zdW48if/UW7iXPAbfuCpg71+8jiKim5Vi90Pq
8yO1Ec3/SQfMyAFFAd3MvJ6svGyWaQhrlATQQEPgTlZIFVMfSRRil1+Yu1kAGQaV
IuahPkdz3aJ4QelXDSM/Vo+HeTsp4wlGiZizW57l0kNx2NFcf9H7IMKCC9Z3pMy8
GmLxIpE2lL2UJ8DkJrnusSLRHezoTCukKGkCIEh9s3i42WX87amBU5XEZbtE8cA7
UXPrwHJmodBbr3sZ8c7lIoO4d9TVsmv/6pzLtwB9M1iXDh5M2w56Is1N7AqJCrGn
gmkazCId0WOHU3UrnKl49853QPL0NcaVm/kxFhwmm1D/Yh9MSftYSsS1+tAXUVax
oMyj9bmolb6NnUwSbFbVoXgeU4DKNY7zqX6EOFQIIt8//a36O0RNMzZ6xrx5TN71
XQvvlqCYhcGLZ7xskJ0E56xXKRKlh5MmYRMLOnSf+9O00MYSqcLKF9WqruDEcLqT
E5Pa24rQiBK4NHBmp6P70Tvg0ghhRkyYxZvPf53/Oj2nFUiKQ/s7UbRnG3B9G95g
twgYCU715kNKte/hXPEdGUvl1V8UURSS4qBE+6sJaou0d90oFMj6dbpD7TYwPodk
SKngeoccX1PGeAvLb4WLazHe3bcfd0XIhSfb/QfUX1NrDms0yqMauoJMEUJBETXE
aTRoOtTKWLLWDJSYm2ndb1+fsJQTIu6OCeBMXQnjUAMa4+Ycou1EiGC6//QoASxL
vmG54h6uSh9kM2TIZ5B/kFOvzjx6LRMNndC9nfoQxJKN5G2FQ+3SOWSl0NQOplJi
/Yb+pkFT8HBSOzHXULxtvDFpnhGLx/NHnZ3tudBU4QwPGDvOO60xWAxLgPXSGFcT
kTnKQJaYZoyACQSPyrHXodT4n97BYMaFqhD5Iu8A3gvr0+UwuidinyoXZdcHkpv2
rri4yZCBTZQobl6AMrZeiCuAz8vTn3GYDR7wsnzvz/AYtjmNosFKKKkaqWNzPZFK
O21BDsSslMpXEfT0KF8C3xFg8Rr55cNGUT88a37o+OTExTdTd9MZvDhn0dCBfOgD
Y1ciMslM/SLhpVCpaqIYbizOiNARgc1b3Vq0ZOI7n6DOh0dvnAbJofqRk7l6eY+c
Ka+krtBdAar24XbcqJbtyvQY21y2mctrTQnOM08n6tIHDJx7YhK4UWyqGSVlS+ZY
2EWQuhNV88BArmUOvoFgZtUcHVCyjW+mRF236TkWmciKy6ppr2CRpe/MrJq/Pu0m
JGh0ami+KCLIuBhVMsVoOqezbbsv8ZlRoRcgJBsuUmHC4grLWpAjRvl0UAEhfzCP
hFPvHY7Bq93b1orMZXooA1lW24m1YhwDlW2jLM+RmXj4MsUJybae1+YsCfyxnqXE
mDFFfj9u+S9A+KuAV+TT6c+Dw6LvuVX70EU7Wa/xOWt71Z3br3wxGboGDGiTpFGn
IqiylK8vZxkQolvXZVIwnyMbPeA/zMGWAI0GEUgta/6bzDxgfvbNz/XG7rV5dfLQ
zR1Fp6T8qbwDoTnTvqwMFF/TE4Vn7/t9hy6gUe1ehOjb7/kA1l/aa3GbYWDMsr2f
OgJ8Xh+ylCIzbkMX93oaiFqlntIig3w6Pzr6+pkpQssaDVh2rPrmz+9XnwrvTJ8s
GCAYebCuoyzqhgrazR6ob7Ck+vvznVQ2BpKEpMolOPMDiaBqRLsMnKitC7lQsQCa
/TBwkmRBtLNZbGLTHZ9D66JQ3AJq3mt6U5WutkAOuYzpt2bVPgcydovrJRc6uY9N
tyLj4l+PBVvMq5JmyoziFwYAmwyijLB5TxwarN2I/zwyMxjvz11j/o3yFyy1cSET
uZ3U9NZAstMHy7bd1qcfqHmpgLxz7DrRyNziZezFDGgBXRhaWcFJJTJN/A4nnYna
/t9H1wmslLwabmUJEsn6kYS41QZ8gLFTHmHGMrBMJu8ZAJ4n6H5VUpvQh8slLMCY
o+OP4H41+i80C9kpPOtIdHBw9l1OweckU6Lhs38BH/IrV8TtR66rPQl1/A+Ke4a6
ZpMDZI4DCfscK3GdnHeq38Oo7qWDpZM211G04rxboqluhekfLzuoh8sBhPUWfmHu
mYZU2YwnSVFR2rDLKIaiWIBH5xqZJRLepJ46qTASP66EhxJGHcg1lhMnNFggFp33
yxv/XQggfpwQ9AUIVjOZLugOPElOsF/iSGenvw1VXpBsPzkkzJmccO5XAT6pb5BX
pxHdf+OGUuADrEi4BBTKYOoMSef4EmgVCbBuhXWVnL7arc/O+TV71NrVMUYKLc0Q
ksctvQdNQai9+x9IbBFLNcKnzu19hj14sKYVN9f87orpV7oPDr5TFrdduSx3K2WN
iw5nMQLnYrbrfYyVquZc9c3ShxK8mr8Hq33DYibK8IQM4GL4NkFDi3rLaL1kAO/m
R8o5JDcPwGe9JBaH2Z5/8J9/ggEaJVWIRlD/OcT8bubasVE/st3uRQ7zbLBDPxFP
hjKKWSFzR3BcZ1i/dabQbnN6oJK+p+1Kmptz8sBKugqU+fmppN+nsyKDmMMl3OJu
akoFCXwdY4kJx7v0tZc/LBO2ZWM3ocpcGv/E1XbuWqLXji2OLGTUJvY1wMLJLxAS
WnOABWrnNkpK37kgG7BOeT2jwLXOWufMD//qrzXYS2oaoF9/lGZSQsydvHenxbgH
GUc/KaDylQsTyIHF0PPaAwVTdMrcMPvIpa9QcrWaYjdXwyZ2+NRcTCHMIOmptdXy
fKmtdwfGISPw4eAs5o8BhEa9axC8EA9Z5XrGmFhK51i79mrVqSA4ThmM0Pv7NKUh
ZwebBot9MUa2tYiPgdbV9kv+mBA0F71NVE3KNxPXx1uwXSdn/ralRFYR4bXOVY+p
hyZzVPRoYNZHiPPWn/stC0cnX40X3IpROeRt5J1G5PgG/rys7bVfljchqdN9j3cx
5pYJau1UWeasMcoqBYtgkkkn8RaYyfuxMsnKoQ0aLnzXDo1qGJ4Z8Wb31sTUVRPq
5ud/+Glrrl2S86889hpN2SpGyzoUVCPpiuSLX3jkeLRAWd8iuskdP0u8CkkT3C80
LC0ZIhlZ30SnSVi17DVVJUJIJu2ByVIjMRsKzJleqYzt1EebFo9ombvLXaaB5G4k
/ygsfXH00VmkMKhso6jPfiFPhlvS50mQmHdrN80x1QxBhEwukdvsGYiPsuhZQ2+Z
Qn2lQNM/xxNxbNKCl1771qtUmL/9+R2qkg/d31P2s8FtZ6rh04BVV9Ga0kPlFrBt
RbtIijZoHPV5KMWOD5GNhuxmUhJqbvP+dZaXZALtPKX0vKLLfGDMAs4jfnUh9qKI
2D/btSxswlE/Ve+uHfgfxTGLZHzdT7huF3LDt3AJE+9NtVbmkfHvnO0FxWiZIEZq
6C6ON79+rvY4q07kvZNefk0B13jm9QfWsxUJat1bQD39MbQRoBo+XUyEK3xOGFX+
/90iwfr8ouWPn0vMafekIfqIJvU5kvzlFy4MeAnFTAu6eRv7SpKCDSpSNBz2jbxM
Jw+LXLpYfgPMXJojyZs4315hWvD5e44VxAMtk62qRv6Wk7Wz+7JH9e72l09GqUTr
KcRmKzCwGwh3ANq38s9IdVlvnEDl93njnavUmPOwgFtz52X6utGflBB4zNexa8cJ
bFT19fBHqFLpiMwobP9oVDnHYAX4CQMavko5OY1Gf97UGQgGfX3hYJcZgBfv3Y5e
wjT24ETt/nm1L8SXKT7EtfsG15v2wV+0FS9Oas3yxjPEzBxnr66KlYCn4nmGeRJH
XsXSWKDIopS6+zsEKNSydZ1a+KrUnk0v3hO8i56kGTT3LEk2q4rE73kLzV0UVQJP
qju3xk8Kb21hSZxxu+mKSwi+yX7YDbGBilInxZKbL8n/gKuAq6fjeWgAi1nove5G
D7ox7+sCp6v+IU85HPlvwmFIiBYCTUNrIoD1BIaeSzopmXz7nu+RwJjxzqocqlGy
SBB4pSG8EwF6giyD4Krsuie4oX1iCPhMK81uZ8BKSRdBP4Hi56ayXvQMHZDMGefu
JR2yiQaSeOVN2293l2ISzr8zzDOfugwkuEtVKngFpp5VHkqEmj20AzvAN0nuGyz1
cyR9ewlLyc63OnrvxcYmkovy7oPn1xDFdBt0kUifpefHv7iUQwFGyTk9TVRBRuH3
hpqhU3JolHQAVLT8wBx2JZrz6FPnXgpMN1Pz7e4rxuF6Xojp4WKU9nKUC+LrCbYP
tu7f2XnhzW42WMaj6fQLrYx4MLwCCU5ft3z3b56kPnqHcai9AQw+qs5RT+bnN3+v
1YosKtUNzmuuihCtGyTpLFWTHRckv6kWHMgQDhyPoRxKbz3RsZO9HW/manzhKkDl
+q07BjAL0CNKx86kmU+wH11thJMOCfjJlkzfvp/f9YFDb17dlmKdSiMT0qIjc9Dl
YqDfu2R7JXgohvbZCgSbDQlYZl9n8bpCNj3FjadKngN+TZi9MLESnm60PomzmMw9
3aCtCoQFSs/zKHAGhoQbBm73diYXQyo4puqRqjyfpSI6pvVGAU9l4vBRP7oYoZ5i
vlQElZT4rhiMWAKqD1nDSIwtV7txIC0GBxnmI5uCQt7BduV2LPVvV8UgeUBBawbk
YlgwhA2+pc7B3q8TYbU/hawJhSRnVyzi9OIGEr82uTjafjKuE9tZfIBSMsBCWd6U
9eJ//j6E/XYOV1gy4olpXUMjZylLLFjH5yOn0NMOEzDAwxpCoZQY4S0bJz8RV/8X
mgjWw5BYBRDUUiPiwObRtA6Zuynn/oK8/DFvmDoTz4qjLbrXeWc2qOKSzduX3j0B
iWZYpE1kkU7EWXmPXXpeWG4+ydhArQjZ21QexGp249POZwIQUtZMX/yqGmO4Jtyr
+4djyNAwDuA0+j0j6+TK2T++8KhoIfYJ7G7H3EP8qN4dCH2KRehHpH4QKtu/99lE
9P6FaYBVYgc0xpiQQlRW+QlwddSSkKVlFXbg2IYQhYozUEr7EHigHFdCD/Km/BrB
S0qNN9mTMIIHV8awmvXBF2qBFhJuTo3M2Ymp8mRTJkabFEoEo3QmnEr62kZrCt+/
gsMmVAueiU10tUsnpehwl1RVhGN2koiW9jhIBHKO/RDH2zr8eVZk1Xk+y4L3nSjR
aKUNYMh0OUeTr4oyIe8TOh38pOQiheUyT8/v2V5yAHPd1gCi/1ud/QlEvAXYW12u
sWtWpHLG8GrcV/rUANeNIfOgHgUokTHFGNENcJDJjMJ95F48yxxR22wLDQxwTAI2
UBJ9fUWkUweJp1KJi5xodmU7Ai+PbKNh9pbEyQ1WDFB1BTaU67oxDAQkurF68kMj
zJ+ajQEujuenNTrrq1bYYYC6UMOVD2iUT8RKbt4jFLcir9eOtP2zwALu2mvM6tNe
dlHNluZ10hnHdczhgxGmL4D/7ntXd/PzC6wHL0gN/NzwLHONt40TTh2CLc+gB0xs
Dao17wgvLdAg+KDKYyfY6+VBUYfMpSUcNAK+PIo2dxAFY+jso6ssySi3THMNUrkH
cL8kefCYddGA4f1I+dSR9gotBw4ubAuaH/TKhQb0dFhsyNGABWiOB+j0bUlpoaUF
9SGs5RqytamWLQ07I3stIvO4kf58IK5bzrVeXtOWUg/lzLw5mW5K3A9SL3R1sptu
HwG1ND8+MBWcQInrp5buMP1Q2CSqX1nQ1dgWX3Kh7g57z+Y75L39yVo8BL7CcT63
wM7Wxavnw4H6OCEOq8rNJ0WyP9sUmd64IU7ypufjzHDn4+ezvXl4JVhIPBILqROZ
hX9KSpW9qIUuAcC306lyu2HWfdW+6Jh8KdvFy1quPqyBEWWhbpecOtfclWqe+Ebf
90UM3m/yYCfMzsOk9gZt73OC9nJ8X2/AXcTT8LMezLHKdBfKSj7dLHfhGd8Q7Uci
WU21dOdjlAgZkwf2tceYpozztwLIn75/PSJdK7lGfgGLHcWGaJr3Cgiuc5wLJp/F
hlSVmGxj9R1nkFT8bC6E5BDc3dgHi40uv5phHAIIVIneS9av0/gtFxHRKmijyBOJ
1jDuE3XoDMxe8HWjYRVIjfY4Hi/B0nPKdSXkjZq/qczwgxMrSelFopaB6e0Sh4Kz
wXKZwiycgGPk1f8Xhyf6T437UB10U8I4+WT1mKBj7Duyxs53YIBQyxMoKvbdYIaN
2ls4DbB9lGuyC8W5HfB+VYCku0Jbi9hDv8BnNe97+cOmv57cYc8uW95UFWY6fAql
V8nKMzGPEhFki+D6Z3mIDHC+VuZllj4I6mlLHTmXTFTZRriiG02FBORT/TqOB4Cy
lw9GqRGf3X2hu2bJk7K9sIRJVWYBDzzQkvkhNwhbU1ksqKDF0nbaG/9ZHU9sbtIa
lbGQwJjwVSuHq2KMdu340b7Q56E7jSKje0DX5a3/dAVnaVwJseJbl4c01UJiDl9y
OaOctHelEgUdMOg7etfTfpN53g4l//fjXfvKqES/zh4fPKDfTVHGvqxO8Ti52QtP
xVD5mzNUQNhrkTyzrH0gNlSWzYK9p+WDBYtHnzAkZTTO1YMdsOlKh9Z3GmcRTMB7
2Va9+grp3oBN7RBOQNzZs9W8OxIZAxqtXih3xeEbA4+DSJRWfBg4QIS2BzK9BQgL
eDLX7C8X+9icTJfB2rxkKUe8KGJCb8dNXR9dwbi2nL2elrY/TE/V423fh2IdcrWw
mroFgez4e5pAHXoqJBsMjYkkC2BsIPFODQZpJ97/tRkFhwHEe85TzWPIoVSR3lR4
5ByDNfGx4dygHP034U0MnPppqKFSN7jH81MfKm8uUEh1IMftzh638RKnHR3GGf5R
Enq0zJhkiVImXR+MMV9wwJFdkwjC5Tvc4DNXEPO92PK1pgjXDr3QsBwSCYzw1FF2
BrFujXftsmWey41FRF35uJBVI5ngCHKBl4Z4O/ZiXP1L4AfEzNGuA1A2iMpuPMml
80br5W3TYn0QYL4D/Cp/+ars0oXj31ECRjbF1q8y9HHtOzbEBtaBOSlKD6p+7Z89
SkwkE8ByNoCOv+Cf+dUoF/VHNFORp3Vl4dJ/7uy/eE4Nx17JMT0YMBxynalsytoq
tz2YI/2nqZ6qWxnZS0biMo65bFraiGwBg4HEAwiJjRjtX4x8k/J+EM67MS/Ijltx
dYgYC5JLkYxWOZnw1MgBIaYSsACg0OBIuJ93x8haDTMIG6GtZSbt53uyV2Ul0Zir
JPahY2+msTOOqvkN2FU2Iows3f6Ls2QWzJL4Az9PLWSgjKLFLygywMhixlQpJSQ7
QO7E8JLF7qYJlRYoFpoRTlm+HURxomjAJkgrei8c65SyxKELUgUcwy61w7Y0tiZc
zin68RLvg+gYb2nCWiG0j5LwXMJXf5Hwjz2azEJ++95GfjzEweK0DU9mZgFtYjwT
tOj/bQjzhRnALR9DfvwC6zmBVGOZ0W5oChAUCOMlcKe7u+2tW/vGfVj+dcAoVt2Q
JjT8bwp5gZJdRIQkCgdTLFUDVCh4yOiAUZb8ovSTtYp0Xs8AIwz7xzgDluTXJIAM
27iB4+qfQNjYoZvJ8xoRLfwGJO6WN3qc1IJ7tyPOBKBJ/Rzqt9t5JyVWd1UbuYQq
age0bGqRbvXsE1w0rZVjkwOUQkXdM3G9VwW6Urmn+xjJb2D4h7zRxRtkxECuWnKV
91ciNq0GD/CRC6t4Fld2NhOsskfNSSqWoKekMqKbPRUXSmMgq6y0FWZRPa5RsNwr
U3XL06E1Gonwmb7XNlc+XrYSg6VHXvikHh7ASMVyigtknJCjeh2Sx6Y6NUpMWIxs
tymrnehy9+k1THIGRUFg0Cxd4bRGoCbEHdlcLYpqx2eKV3YdWQEDCf/FniXMawPw
tY9OU9XNwxxooxNyITzuepKN79PpnH91wq8TWGojW+Dc2j1FlYkbLorCc+dQPWRZ
ZGASKWzpYRcgKe/TIcoq3G/mEN+5sEGdn1D++J8+Uk7AI/q56d4THmvfRqdPmKiJ
TndaFWGysB7iGUTaAaB2RbjpLagjHtoIUs8uaiBCPr9LABbydGMvpluMl/kWHaHn
TdaBC6zxC3L6P/wc0nM4k3/YIQZ9JNaswIMKltzFtK0uezjWq78qDK8+dFv9KMOs
mj61a0DEvgDq8GeR4YG/baIrIF52JiIrYUrIeMUwOiPFE+h66zyh6JuKHOX5CWki
zAqLHlhFOzbSOObKKPXWSRt0aKuIIASWDAF3BF0Ka1dlMOtR74uXYzk+4NNg2nYR
mlN3iloHQOOp+CBmJrH7Ib849hRX8qc79y3Ur71vrhsqZftnsh59hSZKKB6cGycq
PGT+qrQ0DF5K/u0+QIwF3qxlTwtUJ4sp2wsCEFqpu6ypxPl0Ym62jO9AxtB2xF7V
u10baxV3ZbjPm6MG4tJXKsDwn+o+tLRiozgfYXJUYP+gkEOBnX/nmCKzSLW1o6Wi
UXKrI9Mw2MeXku+cXP5bJXHQmJHk2zGrZF08B8WNqAGGsUuJKHlXv6eCOAoiTEt2
4SpNXJlIzVRmnoPJhg62geXQSMhdbUh/CHknshvegu/FbQUXcd7NfT//vG0iyt2f
Hlw+5NxHWczMu4ZwfX2CpsxpdR5N2kzML83fdYjFXLLcD4JXG/oI5uUg3XtDWg2R
0edTNgs7Xu/9LfMxW4HjJAoE8ak+gZLwhQl6A8W4nzmTgGkZvGQV8Ffox+kxs/pq
mtMWswZ44k3a0rcnelo8W903HI1YfOD02IE5mBKGk48IXzkmgUalyVD9Lu11piQn
DoEoVMl7yxN/uY5xKQ6K2THefYhZzUE4glb5T31HUZnBFO8DXeZxZafKUNc8t3ET
ItCFseG3Gwmm8h8DlMikJNj89J651YvVeUaBOiO+XwESj8GinXnkMKSzQfjOGLlJ
kNwUR9SDcFU3RcZSJLYYNJUG0eaGldCWXForTFTL2ZH7lx9oE3HGeeLgaWU1FeKd
Ak862RMvJvJrlL2ZjuyMXEUGIv35mo8+O1pmakNt23qbGCG3oElXI6pORLhvRmsx
LLRBJkeDcuRU4wHHhTFkbeKvibLcUZvhfYJuMH8gCGwMg1f16c2n8dxpcyLlEIcu
EqVKBzHD7SaFemhFGN0LckuyHSa6mPDn/7zoqFymvRguXqk6I7EQn3CvZkpgv4ec
Arw8WjuTVj1F/e1RqGQsL3kr40w6u3AoacDm85CimCXjGWX8aUr4iGOOgG9ilwaE
RavyxPwhaeIIhnGnhpRHcnnGX4LuVsmHwGSNs34PD/ZFE9lDwPZTSImoI7V9nEB/
cmn/6lWpcYqTODjFr2b6LAMgVbXQSFaH+FyYG8ytjXYQVjlZn8n6XANS3O/rBdhG
AiO3LOJWEzrh7NbHl+a5cK/arnzeXfAoYPByq/Td4dmMdMBEGiwy77IGMk5k96Hj
OlLu927Pl9Bc1e34na1zipZCMDWeNtTEDpe8HG60xYes0eX6nZGfmqHv3Wz4J+Kb
lFQIBj7TDs7GmkweIR4cPpMtIDVch0eOjmX9KRckMxbazeVJ49jC9rg4KNmBVSd/
OwLg10TmxEw5J9J6FohDkLWcvpiXvgiAmnnubC0zH5M9ClRrnj9YRr+1pyJCCZg+
LJ+5EZxUYvg+SDwf2pQlGwLgt3k5MTsSgynLJ0y6pptBPd9f5w61Ib32P5cE8qx8
rxWc7ppwhgi3kC3p82BOR6zesqJSFA81FCKvbDAVbDTOaHYB/3asZJoQBSpy9ScX
l2NZXT8vwmBtJS8U/m8OYRiceqYIrLlM5cg3XXRzzXnhbthD2Dx/XAvrLvnsdtPm
AM0+njAW/MkT0fVYbKcfSdPQ30aJns51hglmjieBDxQjtanGcRvYPf0pRbvH1OX+
e3A5aRzwuCbgnIk+UXYR2xfUG+bXpGvuLXwzOjmIDe1tQb9RY6hb/RheFPBo4PWA
9LgMjZyrk30ypo4QTOdrJNCqudCRQ5m0FnLk5CYWTCryVagW8VIRmuizJnDbtkZ/
qvwqF/t5cpxWPdz9P/TKvY11kp65Ak61dbcsh1mcNELtnu7TFdneU+7dax5xfFKN
CFo0M0iZr0sonbzNr7CppVpOHMtjbe5TRqFzU7mH6XIly/K/JVdgAfgFWUSfNCaH
n5dEWzF7mxFRMiJMCY9vHn+O8lSD9WQb29kJ1HhkYOGU/5ebUWUgCJZqFEbQO1LY
H46ahfexCnxl2zH/3m3k6SxOTm9KAf+5lmTfODHEsDnEi5V0qoT63liA3kjpOIBf
ZKf935YSpUgnUdQuKd3MTaWcAEfp69iJm0/pn4aXR6pGmhrM/S8+JAYjMHHJJ5Do
/3bLHYUXJbJD0FCf2ETn7AB/On8xy7C8ZM4gxcgeDu9BUijC82NvT3arcJEXFOgh
Cos0ZG58Eau2C0U3J2NFcTM21R7tXAZGQZ+Rwn3PvidE7TxXX43xyMLdO4y3+ekq
mDjJmYmNdYnnPLxyYHhl/yHGR9g/H8zoffUUhICIWfjQWTs4Mgy7CambRyA7lALl
F84v7uci5AJZNaeuc+qdBAM2n4ks3cceBPdShMxhDaWKbOUGI+QcVKSIi0wc1Uxw
ilVBN/cLWNpn4sVhpVvvR6egTmnhxLDZO0+ovibVrEtdnPs5Y0mR0BF46T4kqYIr
rBCi76s1FWQ9G41JJFFW2kNdLJ95Fe5Oy/UPdTfJlpXJOcE0j4xLf/HH30Q/KK7D
eadi4D39kEfqh92eOpToC5b0of58AGmp+BMUlAI+ZZMtCqsN0J3cuLxWPiGkCa5A
m/A8zw0cdE/Y0r2h02dQGg7WbVFavbaIIfzP3YzDxpI5G5W7i1yFUtTo+/fokoZA
dkwqRYlPCqRjhoZ6y+9RZGNqr2auV4gRqY6n/nG+8lF8HwJo5UHIZp7lmQSY4QWZ
ENz4xd6vMto8/2F9bTHVnbXPlZbLSV2hbNnMyY67k4R1hEuQR0OSTREP1uMI9GMD
mBrocL77YN/7rnDze4hoGXvker5WDTrhxyFUBVj6loFDXdE+TA8n4ZCLy56WUyMV
OenHr+gjP/LDJVqv++P8z4Dm8n13n1bNX3i/BNNI3iuG8tPkOendy5ySGcBBuvHE
i8nnogk+l+TqZ2qBiVOrE/hFFRo+69fJ6K6fPCI3YmENSgmCnZ3w1qLhOjc1wXx3
T8FYexGGzy3t6IearZKTwOBsvcDIvKq3xr+vnEJzPsO49izdpiCtDyP/XeBqsAVL
9ZsihR74RoRqLxdftEK6Se09XSntICWKQ7Fc00pAZ3VXOkmpJkaxp1DCO9yZArR1
nggaI51SMufszRepQ4k6gPG7mQSKGbp7R23THrTKOwAzfecgaAPrXAhGmGKpRHXu
RY1xKQqv09MW+zAAqOQRMBkHw2qX2AsErKUgIOypZplzv+VtRuBgbw4ZP+TJA2Du
dFFvrSq+ki1R9hsTHbiUE/sfJIOewn1/Wrdh+ooOkuuzElR2xYc03oEwSgNqDNpT
F6K8WclNDwxh6qFJUQJCXCSZoEIPwIVVOeUNHHpaUs6K0jScbXUK4rb1b8VJUKRv
p/qWzJQm3tovqbTVrgdJQIBDJGzH/MPCaXP/AohoStGv2s3jA+I4HHixjrqgU0Z2
xCBPSINH5YSQJyt4a7JHlJ3FeVEBkclu/hFLTV25GVWyZnkjqtsWNeUH9yqXO4+z
mFo9yjmEDHk9ZcAGiwJ1jAmPxbIjoJIbJPUIhCtB82sT5/c+4RXeXF2pvzVsrkwi
RSjPyilys/MO0v7iIX7v1c1bfJJIzEFNeNrzkDBxC46jfteJbjGii0BMpr3QqbYR
BrauPQcYIxQsFD7/vMuaXlDpz6+8S8glojb5mP1EzxhHz/FX/AJUxZccVDlF6Qal
ahznSsRbjx5mdWMW/pcvpvoMH0/zBRowUIu20V/gXVLuzBL+eaNZp9jRyS0a0iWn
uPt1tpwwu0kD9RxVvPldBTU/jYYj+htyxvGVMPJHA/K53Glg7z6g2VhjorYVz0vI
5dGMsFzArWSBC1LANA+6P9OtULNdQgPGpuWJy8e7VFmTm08K+pYkLtkp3/6YDNPu
amHGeptHL1fLuuAKAb2paqGrpfBjicDg8Hpl315wERx0NvEcDFAItnRSqgFp2xQR
bgge3/V0QQ3e4ncTAyZWcQVX2TOYtBuVBI7UJp42qBq28OoR9p6czNF37KgM9GmG
72vjWmg7m3HdNcMcuEL3kd9fQXpirTrRdlYq2fEfVLbLeEJxsmC6yRnlv+/TWDs0
dPB6tMt6l2RVC6fPCDxC2IVt3CYx18bQLVVX3dzozl0bcTSImztIQyYHlAKG0EnK
SV2dn9ngKtF5M3rbSFZU72LpWZ+52xNZz6nSlP632EDx8oEcu8pAoKs4SXBgJffz
2GnukbdF0gWHkkOyu8MiA/DSQ56hMo1NpGv6i3wCrAssqVDNFxZrxHDjuB74Wg6C
CU4oBBenbasfdwEz2vSAHA/3GxNpB9HsomVQQ5yPZlOmmiNetjftgOWsWJOu8+rH
60FlKe20yJ5OCHBpU1sOcqRaITaplESxDWnrTVw1jplnWexMMGUmILttv1Oa4k0A
B0ru0HCt+2uTfcSach1wqCpVqLa+DRheWrHl86Wl1Jc9Ccqo6LjC3KyoKO/Hc+k6
OPdg/YqRScLAWMhIzxuTQnWFApE24m/VLo6mZoUWfmSP0aeAEwwKJ3aunfz5QczU
/hGoF6NOrUMKQ9BEorbFXlk0JZ+p0O+VeWxua/Qk89yvWm0dqjujAMGz6iy5/SkY
YaVr56Viar86Jdo2mHnNL64QaRNPFZPwM1JdoHsFqx6VLummy/l2czZKTAyKyo0R
mrJel/CUv0sPTDGTOyj3gWvVZh/4czxQO4x/oWiSp7olfDzBgcGehj7WnqMOYNws
vxnLOWQIV41YZjXJZ6LfQxocrIpVFCeuws6X6dU2qNFEAPMuaoAtFGtnqAINQFvs
TtjLspPUsFx+3sO2WGzXhN4+jz68tEHcAb3lEumoGMMdwnwNk7zxAhkpzU+5Dth8
SZeCaBEmoOWeLcDuOohYAssXrJMFmHZTWoznOB0ed9la3aY5/1QW6o0c9dgLA+hA
E5OxUOD6j2aZhC8HaIqY5SBTeZs4S61OeDyYNEqw76ygeBK1B7sxUtP0nSWcU6uI
rN9cn6oBhZ3E+1wUZZbFmFP4KpYPlC9QZfHHAK0Xd/JkGrLdG6lyGNqvfaUHOenC
9hIjS4d0ZqTmGTD93gCGPfUS1Gu6ALBFFnN+8wrX0fWZtYLEbzguTZuozuINYK7j
GOAnBlQZhcK7o55N5fHPB1f1H9G/loQ4M35+bef/n9pZgsTnrP5U7c/dkhGQzzCe
ItZhPmUfSauho31yaEjGlGc7JJopfD9hOj3K5mLDuSMcn9qLHF9nY6geZB9Q+m90
`protect end_protected