`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
ddtXksX2+yylW5zu6QL2Lhnb2d1sD00763mmSITNX595NcHTEkwn0zB1Dry37fOW
FufOhVzEJp80NC5qZ/+F0Vk7Ik02dIR0elf3clrjeJRK85K4e3Hoo4xn7YbFUIms
l/8VZSb14+JVGURjfswrIyCUotIzlzVYZ6gzoZwDXIi5gQIBf/gI+KxNXPaKV+PQ
Ufys/12rjO6aI/pPlqSm0hCvftmBcnezN2hk1UeXgOIuKZnogjOsf0iJVX2aOOWE
6pD/psybjbnsNB6kH5uFTA5frkzIzkzl5d9+YDm9OyC+k84E83I/7/j+rk4L2dah
QJOvksSIzN867/4Qt8qYTQ==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="MvBXkzurAa5VTw+1JJ70nePUfoQXBvZOku/SMmg4TwQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
oRtzZL4VJ4iwysPsC8SXYCzXS8Fw2gtZTOskLcDV+1B9Nzn1zTyNtlo6lNICRmmK
ZRVu2BmCc2G+fmzynYlNTnSa7C0Cuel6FYpxCBlOuk3OF2tzAmLAuDyOH3Z1Yjzk
a0aHuoCdIRKv7BrZCdALt03JeUmXKPdOmIlkVGFl8yw=
`protect rights_digest_method = "sha256"
`protect end_toolblock="Jn9CQpRhJt4rnzZPRk+dOpzAubz7omckX1MrFd4p81o="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 1504 )
`protect data_block
gD6l00tciPUa6pDNTk/+t0OO0nC/UTtBwLB41d4inuAUA3i/ALrNyoJVcBnAmEQW
ptbcNp5fxEUJjnOxnedyZEuEBxWRieZFQnkRdF269oPaWE4NkwAxvT0tzgJGiGv9
Uz8ecN21pkkT+0BRq15L6JUxXxjP+KpGtQkR6fVOD6HkZa1sbBSlWnapUbJLiXpE
RFcYhib3dwIL2NO13P2IbiBuxupEJw9qivLPCJJL0oYDTMIsZeD6o72jCiVSw8lU
at7aosECcFsZm8boxWzBoNTctJcL//vekLXBmfWJH+THwLKCVa+Qn9+Zjp3Di/ig
UYd8L6VU8xhN6sgKrpmQ3pHPxL0JVwB+UxbPZp1X+ZimzCNVFb9wcJAtSE0AM2J3
4T3m/uZ9YGvVJL4Gkh2/vrqnMqzYD76gooexrtXdN7HXC+vNpI2D+AqJx/KKpZd9
4grHlm81f3DwYikD+TDUH1uCsiBY0IAwTTG9QeHWDeJl0IUSufx5lmoAgAyudZWG
KNGmRvOIZ7ZF6clc9BYfyiH3bp6mrCuD+Wl6Yn11itJMyOYMlTp1kStSAm0402Js
VKXoeyN7Vuwcrglu3e4aTD+9BHAaMu14XkR3Xe2xMmrY8+/csOND0vXLwapq60UR
h9YlwxhH3v2Cm9XARrS/bed2GH9/A7HNL3tEF5ER9cZ6klVFd6hKbqq7a5lr4oeV
0zy3vYztXSfw04LwRQE+cwirw/NO6tGxtd/0t9W24olLmvopp8rdTbEatpECtFdK
M7AdXQMfE0EzP3SZbOLh5AEBxv0liZEv4QO4pfDGKyruvCjDOuq1HLTSNuhuUENp
rPqw1LvRd8fH5PspIyvJ2Paln0fKqP2xUCvOV4VhDeUZ6UTUqCDzmsyyDo0sRQkX
Z/XIgAjfrtJ6Qs7uZI4+ELfN89VXiqyh+3+OqTe1RItIqOWzIl9XS0BSEAtnsj7T
ZdGfP5SWPSFEtCRkqJCh68syyY8J9Lta1t3+tfbIc35qJ+FazY8ah73lve8bnG/9
9AdfaTAt6DDL82jUNwkPbsmJm3vjOXp2v6u4xKCoUh6QfwBDrMIeXKNWEYWUYuqL
ryi/6ug5+W/oVqx8kbImUMogudv0AjPg++75ZETlLgtEtf8rs7qh3cLgJuG7JM9g
elygFbpMSGQCAunilBFYruJSKdH5RcVtWUAgE6NtmbgbJcGs72xeIo6Kgy4UoS5B
Ree5G0krfzkXQD3G67TQNW+A8RECYEq92JPz0a7yR089yIMHmNRwUL/cymDXdMlB
LT/keOkby7hPww80FPIJG+LD858hhVRzwHnOYZmLeMhjpu9jobo12P0kbWYiPMnX
A6M/v0NcodjmmNoFfr08rUnvUp5SXep+ftCpQ0dE8yZcT4xzpkOlY8GiagqrmTmS
3Z6QaLCv45yOfkhsl6wvhTFaSLnusjaA1QXayyhvwlrRUj5hb+VKGIu/MFUbxodr
a32OHfnBSLpzoMG32ta5409jO1rq8QPmafdC1nqSSrSYj5E5RX6lMVGKzOKYl67q
FJqOZNHRNsxJVW0J8nx6aKNjCMsskDfmkbSfG40MOvci2prEMvGIh768CksCSWo5
FM7O5+IqQ8lbvPk4UuGX540ypZlXF3syS4KDA9gl73hpBTZ4ozp9o1vn6eeDILkX
v6pr/H5zPcbw73bRLF5q1Cel2XYFYFZQvZvrsMQoGyaoLra9XhutNCzAVfLhVQR/
ZGRvA9Sf/ulgJ7FWKJyCqKUt9LAvjLz+MlJhV+3+10Op/KdcXaqwfcvGoeqsqIzG
EETHwsHDkz9P1olQtz4/UTEUuiiEjmSrkm4NZIMFJn/HxWnTHCmOKT4I+pcpuO8t
9vCtsKvY6/GUWUzZrQNjpbvvVfj6cDaHbi/t/2wVanhStk3pAx1gBPAqtDb5yLHG
3TtqRyDqzEE2BylkECtNrQOsewF1UgLwS/6ySsxHyznV0viZiSpd9M48BMb4rmz1
4fYvaUZHeYjy9HsI37bW3w==
`protect end_protected