`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
ddtXksX2+yylW5zu6QL2Lhnb2d1sD00763mmSITNX595NcHTEkwn0zB1Dry37fOW
FufOhVzEJp80NC5qZ/+F0Vk7Ik02dIR0elf3clrjeJRK85K4e3Hoo4xn7YbFUIms
l/8VZSb14+JVGURjfswrIyCUotIzlzVYZ6gzoZwDXIi5gQIBf/gI+KxNXPaKV+PQ
Ufys/12rjO6aI/pPlqSm0hCvftmBcnezN2hk1UeXgOIuKZnogjOsf0iJVX2aOOWE
6pD/psybjbnsNB6kH5uFTA5frkzIzkzl5d9+YDm9OyC+k84E83I/7/j+rk4L2dah
QJOvksSIzN867/4Qt8qYTQ==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="MvBXkzurAa5VTw+1JJ70nePUfoQXBvZOku/SMmg4TwQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
oRtzZL4VJ4iwysPsC8SXYCzXS8Fw2gtZTOskLcDV+1B9Nzn1zTyNtlo6lNICRmmK
ZRVu2BmCc2G+fmzynYlNTnSa7C0Cuel6FYpxCBlOuk3OF2tzAmLAuDyOH3Z1Yjzk
a0aHuoCdIRKv7BrZCdALt03JeUmXKPdOmIlkVGFl8yw=
`protect rights_digest_method = "sha256"
`protect end_toolblock="Jn9CQpRhJt4rnzZPRk+dOpzAubz7omckX1MrFd4p81o="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 6960 )
`protect data_block
gD6l00tciPUa6pDNTk/+t0OO0nC/UTtBwLB41d4inuAUA3i/ALrNyoJVcBnAmEQW
ptbcNp5fxEUJjnOxnedyZEuEBxWRieZFQnkRdF269oNY1rr2DcKwVbSJhj0g0MR3
3u+RYDydIxuzRI13YcPgwLXWPBivjzuhSWFFCZ3Fm6MM69AMS22nE5nbp6Ntm6mY
c8Vc+aG0XhqkRAQfL27kvAHeD0tvfWRDhg8FYQnougDJ7PDTcJGqa7y884lH5tDm
GG+wq3qOX2cI/b3bMhVZaS9A51ayQ/7ZYKk6btO66FmocgKBVPQ0Ff10+NrtK0bM
OMOy9IlHV12vuRYWlFJrmLWk8/DzNVkJjOD1aSHSVEOytVW6WPHYwDKcwUVTYHMJ
ZxcEDBJLhaE+9sAB07BvpW3KOOvR6QO9ycJ1w/HAE0p/nAij0oXQFuUB690Ww/H1
yQqxD6E9B7cfkKyaCC4kUMcnu6o7DeaCJPZ8kABvIf3jQ4z+CL3//T/swImaVabi
z6DWvjGNQzsJaMwCTiDdgqoLr/7cmovsDt+DTzQGUNK4hA7e1S4duYQPZ/8rl4ea
IOZOpoWC2eYPqm1d5J1hMCIf6EE2z/6E0Rb44R1c+Kj5VaUXCDcVyifroR6YKR1l
KKuDz1vS3Ffe9YsPSWwrioxIB0CUXBTsXRFFpHAbWdOO9Kfj5kUbpXcxeaRmV92z
3pW4ZMUIn5sgii8ipeddtqRcRALdHlQ+6kytzEWzc0SiJanPfHDfzhG1Hj5I8qf2
Z2LIviTiCu3Lsi0vlyWZWABnIbZt4B2AfB3bKHAjOkuAM8SRdgzhPrVqmh08mvcG
CO+nvQLgoenCqoWw5R51jtjRLc5n/YvXJLELJu2Ten5pzg4cZ5rybXwapufwT5uF
IcWdS+RkCxirdlw4sLh2MliS12IjvJJdAafyqemkUfngBYv2QZt3LpAjwTY0MWeQ
jZq37kbUEyBMEo4Tbfl44J26i88HcTXe3WP9kPYMxcoSJsZkW+dq9ZxQvysWS+N8
gEcKOq50EY39wAK1CaB/AayZTPg+SnPsc9b1XiGav1uGSIHHEArCGc3TGbBDD/b9
gvnnbSpEtc1lvz96SjMruFF1UxpwHktOx19/Tu37s5MS7JgFkSvXK+BDcjuWQcrt
RkNgdP4Squ2rz0QOunA6XhAhQmzzOB5GwYl/8TYPCkdJfKOyR+7nHkAWozVnGeTL
fc17GDse85Hn0V05ofXHk0HRaQaMyEN3ytcfLa7nUYmEP3E81VYpP9DD01zLAnZ9
vmErGk8sVpB0suPOJRRRLn1vSRJ3y64cq1vMF1MiR6Nc1NU7JRqII7AiGtnIHGJH
QX8gCdCrGtW4R5fkyxlLHvNQJb8+B0K6M8nKZx0mzEStJHJ5Kxl9pxRRCJswK8wr
udpS+THRieQNhXrM6wMZHmcA6giUGqcgxLVmywbpZwz7Ejsu1OX51oqCVFt935Tg
Iw0IToQuQsW3fzlce0Dlqr5i67filKUlzdfA3XZrzhfFze994yVW5lO+E0jSsO9N
cx3BHw6gaESeCRzGn9E8GY/GiDwTcY0Dl/PgxX7exXama84uHU8ihkdorZzypW8m
8cckMSZAfzCFKsldKc/92RnLHmO0Aci2ScTFpKXCrTIzDMNgdG57nwmk5PngyPj+
jpT6HD3I9DJNrGudtRZQRPzsZoBlH6MFJ1iN/8XfpnupN7euz1cwy4vnmLlZR/tp
rvJnPpRR5YzbOrE0Jq2suQVNdf4r1GNoib1MaGnWTnVK1Kgaw2So5tMp/0k8wuZL
CY5MMllrcJBl8iylYfPeZ1wIyhSg4PpYs+HSfvXvlRJa4mM+Sboy/zFYcBM1ZMYV
JxiVNl11Nsnp0j5JDK+e+aakK4gR9Qxrm2nZ90AMyy1UOIktZMRaupKNjj0TzRWm
3kZF1ftRWa6bG/XnLQj2aqHjA+saTqsu/iwDI8RYBZbwxodX55J/kGVkGRw/LUCF
Dr51mYrkvpLtWF6bzBKStq3fszl/AbZigmBJkp38aYKDgAfuOnqWw/6Egvmj4bWz
UyWWh5UYPhZDHsMBk7EFrD5qoeurKebwQW8jeBC82YQZFj6dBVRdTDo1X4hLmANA
+3e0yykrkYxRKOyv1T9yrufeMKqeT6CfaD2tuw8jTWroyCM46LG8ZGLDyyPVNna9
X6Dno8NVTmtf497WGj+CjjPHP2a/x7GGy1XWd/bb310rUEmDpdKB5xC0/qE4cNEW
uRO++k5X7mak4Nv37+LT4TXnMiGzicGM+6RPTYpfL9w+0nGLRTDZPnEnnc6bvbjW
4FmYV1gtUB73V+msppReVPqx00Gm52lmvXxP2SovzOUA0MkTZBz01ktIRLOUGd8C
mTeM5da8IBRLUuRnMTB0CMpsuwT2udBif94zSCXA7/1026av8PUEIi0/6CPOqXBZ
i/n49BStfBILN01K7uC03q1FPvQ8rlMde84MvEyeGlAIjGOYb6iLC2gcdebcIDHB
xp585apWuBOGte+g8ttos84Vnrkl1x0/uTFHxLetQ4nCiVzzmHABnPA2Rbn9stUS
uFrsV26iQTr9t7GIlGdb/FxoMj1+haIeoiCBOKp1wLZpR1IjRYVsETv32RR2rb6g
rvUw+0zExkwY9FXYG4s/ZLx6kMZb88uS8aUEPSSIrxnM9V4LLNxfw9lzRsDt29bo
ce1MT03ugNyhVtVOJjF1l8LSS9Wce4XuVdcn6WpRd7w/cZQsWvePLy47yXZ6+nIy
DkR7q0rH7JjQ1jluhkl/zJAHccf3lKLchi5pzkjmOcqC/CRgIGjwY5mP+/mDkVOJ
kLdmonePDYbXLcBPT1aIcvUxsDrNo/RYxrD2Y0oaRWJQ5F+U7B84+7b0zy2H+PKT
7H87C/pwtEUOrDKZmBXWTexnxtWkiAESsRxZGlzQwkeN971DEmBSpy4ZH3OYwpg0
ox15WsbtdaE02D/bTDgMIj6Ak+HbBavfXjlZWTjlkVU1F5NGQD426G9dortgEu+W
+/C1KY9ZayBNm/mE6xXWDxed1rgPMrLReuWipP4KKZ1pWuzBLXlX6DbkpMOscXXt
eufhB2JUh10gl3Ve9Tq9eThiUG8PZ+wsoX9XPcxvgnMVXzqaHUKUt+dZjIvw2DxE
NyelHtMCV2aTE0nrvroyV2hRjI2Xtt3iaC9yuRsfw9rWH3ylRTRcBZtRLT+S2Xaj
9zuRBYFauRkBdx8MVd+6HDD9rULldyuiAx1Q1/OCMOeJgavPxAzprclnvIrsR8zU
TwCAjMHftP/L/XM1C6oHfD8vfpWgeKlrzhA7zOBT3fUa8pJlWJaQX3RjjhUn3xj0
uktIJ2VVfdBe386cudUyT57LG1ry5Tdz7giJ9I859d1ClrSgAPaWSEm/E2fA87RF
MdNaDY5pioKKCJqWCplMRaxo37k4Jn/PBC1vBgZ/o529jTGfk2ig8mTacz+y51fT
WyGTfqSnrR9qUt30q9EuyYJ381LouAbifnSPUk9bKHX8i/ZwnQEFPZZnxUHVWWgv
WyCDpyKeIhx15aobpktNai+UZm25Gez4Vc4vFFpa7RfFW/V8UqbxPxKg4MqaKXjb
yKQSsRCUvPl27rHtwetxgNJv6gkHvJwLRbL4gp5iYtmEY8nN3iasrhjtPpQUXPoM
kref2GKOG7/gli4Kr0TJr0kSUNwRSPZ6B9wjrwpR7lL/UtXQawbovPCdoly4RvUl
HAMJ0AXF+5/1gj72yB92ciQKHzklxCPGnTmJxcge396BlKqIrS6hoGFBqlOC7cpO
QnIXZG6Sscpqe+gNdbxsk6gK0xMd9dlmucINQ+Yn96Y5sj3BPNdCwRkIy9GmLmuG
ezaiytnY3UVs7RBgcQ3GpuZw5/uJI2Xb+NoPi+8fpfVc6vQiiD2WeIoZvqWoacSw
wuSYTibIux+HS45aeDv5ScS7fl9+mHagTn3lvtLKg5MXGgSwkmoUaLU10i9jxYWM
Alkc6PWOavjH4rdpXJdVm7iactu8w4qTO0rshbUwwDw/qA6yQOGOCzF0k1Vexy4i
jjtQYtwMr0bE0f//btgZNyZ7XPMsb6ZqRHv2txZLLa4UBzZDNTH2fdjiMpFC7re6
U5fFlb8RRzignJisgaA/LiWsClNAZXcU4bxteu732pT1lLGWtXDtpEGLk6e3Suv7
kuI3VNTXYJiP3KPo2/dy4hVUkhJ86so6MietJL4bILAFz4YdlSKV844JHaHbWvaX
VcW+RNNKBmjv1o8qZGWy8Q0QQ6E3K6XgKGwI0tQo9GmBR7zEPlNRObVgEbRYXNdG
vvs1qaTqDSlyA9iSKxJuKX2926S89s8ELn2Op5D8IC1BhwVwdyCenRcKlRZ832kZ
6Pqu36rxVsT8CYI4Pyv2llrqYz1+8rcC0kMTLLK4NJvs+9O8CD5x4aBqQW+WgoFE
MDvAj1GeGZ04TEmIi++dQmQkszATSOcyjRmhuqnVJwec2GT2XwSW3u5NOyZyGYpz
51FyutMYqd6YX+AooVK6eUJj70XGQ/fohZJkQR2CCEV/FtPMyOlQfosg9XR4QzM4
0hq13uWi+5zNvpmKC1f6Ryw8C1rxjaFIIT8VvSUP4QfG4hZCrdLToImvyG9gX3dS
Zu+wAwDqarRINOynLCf4OvT3r7GHLcTv8SrQfGYsjulGZUD7M+mEValUy0P+1vSo
YxyisKy8kKLtaLOC3MIMQAkfYl2ZbuLFzJzH9Qs0W45WOy3JaZAbpXSX2by1JaeQ
41923nOoDNPrdbwL3xim20i6NyN5sRWIzkQhWvYFVh63oKgE/zaAV4P5dPrin+DU
xCYHhGW2ssIMOBTUyALZ3/qDNg/lFWG5M7kJfUhXwwAlNeOaIhCM2AmSKFOvuby8
Ux3JGazmgCzllzD6cwOadYS3x2wwE3FxAQuwwQf+C8u8xC3xMGX+aAJl3OL1lwPY
Y+mS6yD9L0qJbWJsjYHzUX7xq3DKzLCg29keOTZInPT+f4h2cqGTF/6OiiHMxdV0
jFk3SrAdS95mxQh/WohtV4UQ0r4AME//Q85vW7/LYjIT8qWVdOXSg8r+tje4xS2x
j3OobAsicKa4dfKNLEULvDrbPjqCpfK9ttBmez8uy9mOvhW4KfcBGTrI31CtGXqx
6PIBulCKMzsiWKCzguBEaaWAcLBUk/tjlgzXUxaOTjK/hJV27OMo4jxzYEabgSyq
wlzxN4JkqCVIO0wXczZbE3R05JAIdotOaXBZsJ/ySuiSPy7vDanWLuwGg0cpbei2
MtE0rDsHlF7vTnhLcXam7TMLMBUoJ2blYpg0ZkqKExf2PSy6udbdKnbylXQY4l7j
5d5aR2yRTz09u+Lne8wh2eq09i/0JGjXmgOZj8WcFrpiOoGcSLHJI5Gk4wrzB7ZZ
M5HeaVuzBTE8aJuDuGEc65BWHBAzOEbancixQDSnVQf4XjMcpgH54jknZMYulOJI
I/NzPEwr29Po452bM4DSBKfx3HkRSMJ5LdGQzBrIDp7Bc7z5ao/+zP4oB3SMKm40
poNNvndIqXNmDutAFvtdZqUHCJTncuiNF56HQwICzVfnMGn1hM6MKognThSKLfIo
tI9f7ssux4R5fKd9WybjtLz8m6CbYazJU4wmaUyR98NSVaQ1Ij2Giav2kA7Om5Wp
4wDsgiHPaZmsQZ7llalfRFNalyA0J/S5E/4fr5gfWMT8hNCwkLT0Ad7gwZ8YzQl3
5ZNM5lDg8p+/nJ/7skV5VbmptdAE0z+YbhbbnQDq/6aHltmzL9yUdHhun01g6+54
EGTJ9CVAi2uOStrkk4GqUldlt+Y8fGP6bdd85dCWXmWG9NiQP2QT3+VtPrAfGEFF
XAJtoYHPDQDqSm3obrUJbsbXupTJf7/DK0CIKv87+Z2tqQOC2MNsqgBZcfZG0VTP
yxmoCrBcgaoj2g+OWZbysC84WPQlqyyzt2HYNfR2SlZ7/H8cRZ3RRljq15/u3Lzx
wnZmQAfRua2Tpe4K8Am/JQ+S30vIrv8lUytdXzFtrxALsVyhn8UeoExs2INfdAzi
sWWCk/K9vEMPBSekRBgFh/a4vCNrj0yUYiTCt7AKcjrE4KS8GdtCg0VCasYLLJbW
qsppGa2jLJwJIiy7Ilj1NC6F3uPHSOLnlLa6LJtDNXSVRG1asxwNeBbuSphloqzn
vkU48rRjirO7AN1Oj9f8MXyKxHmUbM4OmcgXWTumMljd1pUI1P3AxX4S+Px97rNx
Aq1qq6koFIAoKmSUE8rcUjzKBlwRNkm5bux7pE/KFRWTeMC3Qt3aQm2hr4kp2u2g
3yIxg4SNMrQAjMXJKz0Rnuy5ApK4rQ+04DTA/kuoMsuo7OdMlnTBT2ESYPw5s/0e
y0BLLb0cTirQg8GUenam588YRV01kxs+G9uhiaqnL9apAndNXrrFMEsEZA8Wolh8
G7d7OWBJYKxeW4KVonFa6igOXNuOEqKEZa7JegzZ8ko2a6kdeNvIHTAPBG3ozIzu
PUr7tiUiyB1rfJmAIE9+V0PRrO0q5jU04d7F5MQui24k194ochw9SJbQDOQFuMv+
RtvoGEUCTRvDapEVe2/IOSxym7iH74Y+ac1IFMQGBpD4E9zzaUgkuba1xRnca+sA
8MZiQE0NypV8UcFo2jMcL6Gk6VaDdAbsLPsbv5oKxp2mFpcqQU1kbqa5U2ym9Vph
1VGeUjAVk6k0u0CQdG4Sax33GCQGUrTFu9oA2wluNuMQcGTH4nEX3mC3AOA05n9A
4QJMn+4sn7Qd0t552viOm7oGrw0JOHaGQ1JIw1Tbbkg6G1fVd3i49WRkDoXgImLr
ueI6lMM7A9C2SET0LnGyyUtUFxqkvSLE78TiYPZPT+HNHjpoV2g3YdkyXx9OxARf
d7M1s7CV6Dj132nsYrJACfj/kojwKH25xcZf9aGaSC0y30PiQEgBDJ5V9Old7/ap
U6XcD4XHbP3b51f4h3g3ekyp0H6lFUGgE0aXcRzAoMeC4b1CbyNPyuXjXCyEZdP5
ALkopGg7S3HRa+lODdMA45PMR/lgC00uLF2IeGugkSAbcWhYGWQwYfkUbw8u8RsM
VW+hoXMGeYmPTgeOck+OI/mc2ARgl58YSj9kJI1cLGY2067NnKWmZoyuy67qQUTP
Eez2WpGoVYXXE/z6VEtNrEmUpwGCIlcKWY0Q4WzaI0ATljBrNAqPD9e+UL8luWfS
iDmEB1hUsZRElWxJY9DLLs/G3dQ3mAUvx0yrW6GK5RQJTnHF0dUp+iBgN7Ht3uT9
+/EUXjtPZ83xfRPuPZW85HQ1jLNO159BKk/fMd81N3ZqdGd8j9qZCyehWW9QpQj1
QBY4WI4BbJWFddCS1Iu0UAFVUAJ1UL9x/Q2mUNXN+SucTt0fNAu2z4W2cH+RzJm5
gi0HbWfANW068iNp78upCPqfnVrAcQHFkdrhrvrnNIr+0A2pJm5Gn3Vfqiqt6xCI
rJ2nRGWHNyuNQ7f1HeByNZ5p8ZUmtQqRYcYRHp9n64XJEJL4Ji01I+RoH3ZlRd8w
hM6WaC4Nt2pC0ia3RKZuEMHZyTbVr/JjBZgmiEhBACmIQieDiba66/c4WB4itvGI
5+RZLZYlw+/iTRfKM+fjjKEeWQ239MWzDa7OGs+SCVFEt3nhqzgMFOKjLW90HaUb
aB35ac1tDMPeODsI6Q4G88Mk/jt8WsLbPmx15zKvNdlmdR5avgJq8hlJtJPgpLCn
x9XRSwBGqooC/wqqSbDxDUACBqnaVsHy9vjSR+aEaGvqLrwypH4G4unzRC8ohlX4
mPxEt+xPo90BlJdE93YAHi5Z0JOHwRu3MctrMkkeoDu+hrI4b7gJxjaPWnT4Bnjs
NBhFMnWV27ovSIPNbeFz+NfkIKHhwJj0FtvAPDCS2KM/WERd1eFoPUPV7UDAJobp
ueW1Nv99u5omvkQe8/SmN0f7yJbysOwo/okzaPgGRYZRgdl1kGetLwU6feIJW4gE
Xruhg269BNjJ+uy88eXPOJxSL0xNEkpPEjzhqjH/KpcaMU5qXgTXV73OzYmkHRat
7gkCIIjVCPVayk4qyL/8tZEGoe3kX9Ym4IjEBNNTX1UsGyNfVlx/AXuCb+glMv+6
sPdOdUCq2kNFrAV0xBJliApXMP+yCyj6xZ+4pUbDluDpLgTyACI8tEKjsSENeoN4
YpueNgR1n1YAMhXp3LeYG9vUh+hPOwvdcga9CRpvxIoOw87HZPR15qEs8uWXd94C
huke4E9MYihfh4lM75GnLzS+NuEeG9bCLQRSS4Wi6vu7FqD9SPe+ej9xuhc9rZfZ
reFUF7o/cLuQdkRoNTVvkZtbkIjB3h51scAip7NVLg3mMoOM7zViRdwU7T2Mudi8
/5BoQpLVCm8Etr1uXmBuE/mSrkfeEaeA5WFyKz033Dj+ZwKFYbfQn3bmZZhieHzF
0hI5w6P1D9R4qmvOXojF7iEGE9MVg4+DCRKJLXGYuL0ADNFvDHgRMwCL9Whr7s79
MEbYmtElt2BOQohdtf3xapkqTkTC7+TIOCLz1MBUuWWzBmZfJ0wTbZDXhKu2xDwn
SiME4jVfaQKXDCNI/+4IANyf051dHIJASmqhuF5KQQCX8zUlh5+IldM9GFMpAehK
Z3G9m5yLY8GP8OHa/EoynnlcbWO78aYf/GoNj7u1XnhRyhw5eXm744JxyLsJ1fPL
QSzllt8lltjIS0D/jyN99H4x68R1PCSXULVBz4blBPZsUIPh4maEXffTAw3kCjbP
6PAtgB2143/EaMtFph/Xk8E9n05ZBfCjLBlF5ni8MTHBdTqxAesP2lZ0ePwEKMHQ
qvuY+D5srvNVgwSq0GEoP5Lt2xZcczFQXQfQnzsjCGQvi1k/NsXcqloDqg2GgIux
hGXSXkp/2HRhWrDQdipP4oeBy+lgWAwSQiOfwVZK9PIk8INi4/Em96lFOQTPnRZ6
hUOUL4BVJ2eTkQs3XwGpPd+pQ4y+TxPK2Cuqq4iGjo++TgfUFANkImPTsxuhd8v+
oVyM/jYnjIInzBXkj2Inv7AMKi3QlAuLObo0rMEGeofxc0GU48jsgiLSx6yp1Oc1
4RV+7XW5YnsfM8cTeTc3gxi2tycVK0LQ6vX8C52QwbWt/p1m3ubJ0PHmq3HCFDMA
envcjrBaVRju4cTSSUz2GSQSsHaF2ehnnSXDoQnPYBs1p3SFKqUeIdhHa9UnCEKD
YDX20kKcnZHDFNpW5s9lEWik2cNLcHQ30pnSjoOYqezAlPyYJi7eYa7JRCjqKlvX
uuFM94aNicJXF6Mbh+c2xWxve2YKGv4v1VP5lI1uh57niqdTJIDm+kD0m4eNKDJh
`protect end_protected