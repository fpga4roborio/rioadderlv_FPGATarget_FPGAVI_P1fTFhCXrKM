`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
ddtXksX2+yylW5zu6QL2Lhnb2d1sD00763mmSITNX595NcHTEkwn0zB1Dry37fOW
FufOhVzEJp80NC5qZ/+F0Vk7Ik02dIR0elf3clrjeJRK85K4e3Hoo4xn7YbFUIms
l/8VZSb14+JVGURjfswrIyCUotIzlzVYZ6gzoZwDXIi5gQIBf/gI+KxNXPaKV+PQ
Ufys/12rjO6aI/pPlqSm0hCvftmBcnezN2hk1UeXgOIuKZnogjOsf0iJVX2aOOWE
6pD/psybjbnsNB6kH5uFTA5frkzIzkzl5d9+YDm9OyC+k84E83I/7/j+rk4L2dah
QJOvksSIzN867/4Qt8qYTQ==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="MvBXkzurAa5VTw+1JJ70nePUfoQXBvZOku/SMmg4TwQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
oRtzZL4VJ4iwysPsC8SXYCzXS8Fw2gtZTOskLcDV+1B9Nzn1zTyNtlo6lNICRmmK
ZRVu2BmCc2G+fmzynYlNTnSa7C0Cuel6FYpxCBlOuk3OF2tzAmLAuDyOH3Z1Yjzk
a0aHuoCdIRKv7BrZCdALt03JeUmXKPdOmIlkVGFl8yw=
`protect rights_digest_method = "sha256"
`protect end_toolblock="Jn9CQpRhJt4rnzZPRk+dOpzAubz7omckX1MrFd4p81o="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 7712 )
`protect data_block
gD6l00tciPUa6pDNTk/+t0OO0nC/UTtBwLB41d4inuAUA3i/ALrNyoJVcBnAmEQW
ptbcNp5fxEUJjnOxnedyZEuEBxWRieZFQnkRdF269oMYgbT+qxfCitmCMREFcG9n
d7OAWb6ZdQ7U1yCM2w50DSq+pJDNQADSvVGChEy+5lsBHHsAl3/WwA92Sk/aH8mW
LT3g2RdkD5jnbDyMo2I61JC24AToSqWiMyp6rspq0IY1wVhNO7aiZfYPMHBEVWt9
kl60JPLoFpBYzATYLYuMWAMjj97B6CkuIobHHpXb7Q1ApVrRGzrRdspadpeRXNaI
fgRpfHgzos/J7Daxsm8YikOWwIhaQmbRpVqUtHijUgwSCz/R6Oj/Q6ItCzijJMw4
D1+h2MZv6Pwua4iVy73GuNGDI2SM4xkPwV1ekP7KlNoybcVLtbSn2y//WXH+ii4i
kG2V4nfeI45CmTSxIXumLDp4g3zA5Qby9qQy6tV+rGdZL3u3VdS6SwjoG31qyHT0
sCqWz2Ma0cn3bYPfhYxd3vw8HlXzyQ2eanumbq7Pu+j2Mt0j08p/+YilLSh/H5bh
5yZb/OGRqudzJGLxTsyDaS+HidHi0v24XhVcMzxFdOo6NqgkpCBXcYTCS9TQYxeT
S7pOyBUSbCWMR7oNd7nVMbpMJdt0KN6JA2ZzYerZJ0yuyWYbCBdzAEeigGgju2nr
pqDDv1NTTVdweRbLE0AlwYyk7UNbY6ehZizg42RxYfFJHrDiNT813fafozczGjc/
Opy0qhUGBcN9/lb17fFbfcBk0uG07QtrK2UGAJvoBALJ1PQlDttRLKPYfLDNa164
97rolE3xVCmD/wuEmr4J5aXaYiNLMCeDrhdmdJjYOW4s5e3nJ56vqoccDVLivodT
JqnxAtayi1joYP2HyRN9vpP1KsW4xAxx8zj+ILzCU74JKilNW8hrilWXa+S+ZVn+
EAUQOygIKYx/d3id1lwNtoxbasOBs1B0AK4ADsQLknAmrfJrwOGBoIFBIiLQ4BBr
2Nlkry5NhlJ3TGDMZFW4P8kGf2ZIbK7kcBTiiGO18M2hxYg33y92z1YHx1HvSw31
+v/ge+p3rOdxRpZeUHkLnJ84uKGju7h37qkEELVWhxYgEbUn1H1TJIE4npoSH4Lx
sCzojppXTRiadkn9lspv1TPG7AwSO4tmJVMd1b6sGxJ496jq5r/ewqrk6K634/Ot
HdzaS4uO3Wu5X5JslVCyG2Ty2cSZjiUGw3FUmyNMRqg8czIwc8qQoXK4pgJL1OV6
jzh9eKjdlZi/48ERjPAX9ticBVOd0SsKeTQrI7ApEtylaPWqm4fMszxOT/QSQ7c+
2CxLabzsS8mouKTs5o84gkTuFM09zhPzZEdqT/S8NPPZGjDbVkNxUBWJYrMehTQ6
3+vlB95QMaCKMxZD8cHC0/kx9xSl9oVxs48kPhTCbnkwGo6VqN81KsS1kSxYTLnY
4j0dtv9wiRZD07oitOdQ/00TiN+zzESLRr8hXgYeYAlT1p9Ss4Cb704ybK+osmDC
xXSarb+q6xWwABm6Yn0WD64Wk/e8vsoXW3o96I4nyNHztfh8bB5pDi+5SHihmrsC
VVDWRV2bc5HDvw7OxAoEve7gzDbYvDYocGiQDuOvTpbl0mewc4MuVA4kkYIbGy9P
1sutcbX6+70pCEfCkONt30kqxu1I+IolPsQQGsS9f7mKA8NChc/pIu2Wyi/SIq1Y
jwfLKg6bRg9QM/Brz5DAwp06XHYhIsXbCV44kO1mzTxHiZZOV8Hg9rBPwHjcqINW
cZstNn6BHlst602ytXEgsA1pYFg5fNw0C5Sj2Ec351BZK1YISGi/9tvL39Ox534s
BQxP3jOIKfgfZ7VWyb7r78PbF3QMkv8FhI6tdTihCpn4VprOYJGKkQSrH1QRcxhd
ohtwM4CJkb7OebFX6eRkA6B71tgTRXq0QLY9DOyNKlrucleSZenHxVTdsOfNhQ88
mF1nQVR+fZOxQLRSvzjM3Kl+j1+X6rerUpJW8wNuHw0H+1gW4AAGD09FxXam1e8G
1BRA56TvcbTkdXTVMBRbTz0rfSD5LteVi4o/cXAYgyW4YqoqJxBa+VEbHr72ch/4
h3iDaJ8ESob/tq6tHFfGJH94XVO6WevZBR7XkAVlXGh0cR33QYC8uOdyGxcUF5iP
LegiUaJFZZ6ySO8BJhVynH6xSDVhC61pUVYI2qSMOO4k316mCAVaeUrAy+UrV1KU
tdGTuRzxNipzruP4G7jdcErj7k08r9oam6iysRfdNvCdTIN2xtUBR1Kbexh48SR1
e5fuLAH2z7qGcSWNjcUygfhemlpn8FJoKk7Kzct3hQbWB95iARAvXmjpwhIF7qKw
Erg6ijF2JvNztVARBfQOMMv+4cmA3BzIGKqfCLUXExhHLxmsB9AkdVnwLhTVWJJu
JvJ01mpJVuWaPGPDBQ7NZwMqkX5+zB63iMdXF2TiQmB75vfOD0AwRfbg2AaMDFDp
PFUfow42AZuCfb4JXfTLmwYhPxhksk1Nhwj98Qd8nyHiEn5BKD6IiLLwFl9kmSxX
0J1zXNdzDnafo8X/vUjABvy33QnI8d0dycTGX2cL91QvmKhf5Hpry4gUO2peA6hP
EBfbedeZDb7TvJWYnbX7rqAsTzOFZxXo7yNOTABq/jk/+hpawlxYqpVl5/dzyKhU
u0Q69Hg3+FgDOqEPFSPOBL5gGZtts+mLdeMZUCSk5TDnTsVgCUOPgJI8wfgGybsw
6X6tG4RxSvDUt6Db/01TWa1q+0f766Xy9M9gtM5RGjf4KVAg1/nrBjx3exgOeOO+
hOLXgcecHcBLFJu9fTqabkU+bDqAVt5SKGWnRC8evRYsO+hT1LuuTEIevvXTCvvC
0d/RYeV2aEdQMd2BkYAS853TDCp9QIKpJOqdJ8azX5rm7V8N6huDBWSD1AR6C9pV
MaJPgRBvBO+FU0LSCVIOisJS8J+6CWULTGE3wp92gYx0Y5xtg7f7a0nAxWufPO8s
mhAla+pbdrs72m+K768cLDMALkoopqLFNkMLYKTfTQWsNwUhprgzRzmnbqWtFehh
fZzA//4ag5XMECLybD9C++UmK3wfb1XHxF0sD6tgqLUsVfOtOMRHZ8CbymAri6VV
Ay46OZG4arx0viU+JT97rnu7zKU28sNblzFOLGTXEwJrxvU1t2OK/OHiAipEaXwq
xN7kYRMPORTWu0UvebfwOEUrQs1X8GithqORtJSiXgqpNDmL1bdyVivY0bt3guad
H6w8nrVWkroDkNtdpVt6+lLB4hZpyE+AFoqzoWT1eGCocVlEZzfQnpuXdKM4+RBv
+EcQkp//+q2gflbu5+RaSdXLVm4nlS8U/CwkjiwQoJXyH6Q9oLiRw5y9y+Mv1VrA
Hy3SS0xxk+/VCnrYohhjtCHGUbfKj5qKFR/9vYO8Dclq6KRHt09HymL46u5c3FDl
W73k33K3MFoXgCbNGAZDxDvcfNLg6LuqeDM+cYFk7N8YNhnaAAzTg5b4Am2teWmn
yJ2iepJqXjSy/kdSL39mHZXIBBuq7CORCLP/CTHHsNv2/RE/frCKp54bC/OcwmLm
8tdADopO0JPzYHJ2I6CU7oUkoBIBE22aNnKyfpRPA09510qhK9dMh/MQXUyU7dgY
tFEy7zG+kyS1qbbZMSBhlUw8Lh7YEjzlRJ/GIIlAPcCs4xO1gsZjlesqffP00182
ROmm4UI8qvgJh9ddMr4j2nrhitg1jxKW7kViaqEldn4QB7FlyiW9D7LoiLd6aWYC
3SEomgehEfhBTlKa0WVl2w/ydZKe4j59brSMJ2Dcvlhkv7STy8TEPgdAXTOG6P9s
QqVYK+ZUMqZScfNXXtjSL7+oo/9ijlg2mrsRwGp/OK1C2iWQeN/w6Pb2D8eUuCRK
ExPkTTysSPncmayT1yD5s6jzbvfc3tRlYM6RP8xaZ6/f1Qa6A7jIaxse5eDOvvEE
uEQAReuEoHtYcx8w0nAf6PyC1hKQJtIxv4/qI7GWxqLDj50bXUtgoA72rGxbhz6g
q9sIfdXEUHL+BE+TWzvYFhSN81IhzLUSHUdHO0otLVsupGAnNlvsKcN3icrz+Q3Z
uT8R39d3XbM5T7yTkFzFEqdpMMg4LfASwyaKMD4LkrtNmvwU2rXeeR8yfqpkM8k4
tRLAbiyHMGTrYAEiK5S4iBWaMEWouyt7qc2lwvQEeNF//AIcclIaWKWNwKxX2SWb
A18u39N3VRKVzeAhvddJQmD5oWF1CFsUgij/RtVVBd8XnWfZmN68lCm7wBIKkby3
7330RhzVnCAn8h/Q327nE5hC0uyTE+Dpf7SuMUB5Da0JyJlvEMTGVOO7mzBC22+W
4GrqqzDxrGAex2DRaUkCpFUWGatTJPv75g1TNBTREiAJ718x8PiuQsejM/8Ldr2S
MU5M/0DzBz2RaJmBJjWC6Mqf7taMMkJ3hbzp4cHln4B2gSh0xuRN8vz04MlRHFMa
kxvD3V7QoBVBdE2E6hsvYQCpxxmkObsGViuMADiI3vvUn3ed9bzuxF/etx6Tw+im
EU9fHkHjz+R9AIw8VtEhLOhQRI3+3PQrgBRsR/4R7eDG7v3m/+KakzXPTvI/D/OS
1o8v39K0WsfYnhiiavc60vIeiJh8jBNyE6uwqtOV8QwGYbFSc+CeZzIR4lpKnntv
Kc6usiPEKYqH+yrZsOdtSgBbfFpCJujTyLVoNoxbkaB0r2MNoGLdLrO2Hk1AslIa
KK5KUFfRIz2eNQJmAxO4zlmZOfEP279T7WWXGyW2n4NVpNH0b9Pfy1pinJHtu427
Q5YowkQvVM8Zt8WiF4iqhCNr8n1SGJua1IbPFR1qEom2zUukY0Ff3I8Qyu4Fg628
UY04uPihFo2JDWdj+4aUbY1YlmzNN4jdRwaMk2PXTSlS7K12knP2VQsX8udcZy3k
tXOuSUFY6axdgujhgkcbBk3CWda5HrdjSWFKtxXovpQCVQe3L+4XJbCP6sg9QNb5
NrPkgwAYV2oJFuW7Fmz5GpXpxJOPluVnGaKdS+55CK1gu4Nhtr1wQU04UT5W4tw+
4eJW89mrbit24Rc2gdvtEpNIFvCcXo6yKES314kV/bnvm9WNAi+6Il+Y3n4ftG1p
a2nX0HI/7hWfSA5A0kEGyElWTEuUAQ8LL1wFJu990WLw6aifEuN3BCWo8d6MNoIS
FcbCnfo2z7wIOdDxIoMjQS0r8NDR3w4Lg09YllHTlOM28lJ4fkLMxSVTH3FsEMfn
DC2uuLLqHqlhw4H3hn0aW5Qz5yHdr1py9lhR+fULi6qJ3CeBIrB1L4Sp96McvE0N
Dzbvtz2SQAve3yYP9yX+Mv19p+l0MTAY2ucbF+K9dssMtdYIpmdx4+yTCcd3AAir
edRDNbwNYIHVz9mPADKM/YO/qzXkXEWYYXwFTBjQwK1M2eaek+EtXePrx/nvaWXV
hZdIx5KnFfPlC+oTUCzv93utGKzsnc+4dgne+Qk+yx/p6Kfw/vWCl3luLQx26suw
d70ZTZ1p3ezRm5/e3I4yLs3iU8B1jzc+t/9z4Kv72v48U7+GvLuquD7mtgHrcQHp
IrWefkzaqP4/KKsgqzRdvjLZ79lF8gR5yJoYgqodjmdCGPTNx788n2PpE52UaVwb
+N2PVE2E68+Y0qs1Cpi7rwf4Rz4B0Etsiy4oxiUaZ33csboxPCfGTIq4WtSWM6wz
pIJAbeK5mkxCQ7qMWbC5p/VjvoBrffC4mTrxVpsMqw7ELOsxuScYh9tbvI3K0GnY
Wvc5EBpYTasJvoq/swBDMvczxSff1WIt+wWPzYAhm1s9CnqM57xOZGBI5EWYyPFA
i/c3DQpCmZEyUB4XkW1K8fu4ETm/J0WGV4r4xaibp9D4VJtP+8BsTgTdyTLUcH/C
NHYGyljB1BpHiL/KiBCuOhcustysIB2+EPBCs4TTldjgcWPegqHRYPv0SLc7T7J8
v25y+oFWcPrDefWEsX1pk46fynEPm8dWMK/l7rzHBxP7lyy4Pdrj6KMFIg3e5CRO
AqZPmtUrPTTOVTAQPL22s9V0bKAZfWDag7/G+tLw6+aQmswPKMRwe1SiZSGnyUer
Ch7hMY8rz6EGH/yFK0DbN5um1BLA/w1k9oVYvb/kFEa8GltMoX0ovSQz1pRPapfc
ffA773O04K54uky4ibrIwyPvKbTKQyCVdW+u4ixkC3y6Zwy1jn+wdD2dU7/7HoNA
cHuhlDlJxE3Vvq8VXglTTAGY/wqXoeAt/rsZIzHVgLbt+bdWnvk4K4HAcnupGTpK
jjUySwaXPlvXFW0H1UjRlCkxBSMYbq8gCvzHCoQeo3xOJlasDSSs4x2I2ZuG7kgQ
73Iw1uu64junkNd3raX5gsd/8i7vGU+nWbWbuhVzbyKTCn+VPX6KKQvMc7Ydnfyl
JIc0RMnvjlIJPcg/HGfj2RTYZ/nuOURiJQSvZSbXBw63cCN/HoSmQC+r1RIzMza1
viFTC3C1qpN9FVNS9XourCSIMP7Ydpt3oUQCIRs2oQtGAeLarBRXusF0hOfh/pji
PiLkFJm8OjqsiKwOvUVDt7LZYZrfdQauPBNktpUopjGLN9Ndg4cV1r+1IQP9gcek
xl6WJJHIbCF9PUvMoengmSNlTkkDYT4bWHzKdBtuG12ub49DoKmUBxOL/yDEZ7wf
kJbt6w7k2TSmaFlh2hGLGGrNXOLYF7+tyw7fmYCZLzi+ukcLGySuNGpM98HHIfzC
RyTW1zoXLaIqLlaTZFjTXRQXSdNDsDFLPyH7XRc1A60YyW0Mu0p6Y1ngFneq58tp
EHayF9ydqBxrZX6y2ec757vG6L4cke7Qe80jMwPzFcahmDKck7nPPvB2jEYdk5o/
X5Fv5/BIvjMdlSy3+00pHsVMkywrBX28WX1ADk3ddyw6OAQspskT8FLoNMHF1pgO
dkF1ra+3to9jyfk8TkBasQXjq52koDVce85l51pzPF9K1vVDIE50JEo6sgbMJXtP
OmLaO5YS/OjX9yosRCvFXRUZLz1jwaNsx6tCWBrhvKecFPka7s6WHWqYdUfsRJ99
+6klxpw/r19Kt0boEF2i5xT7WmvNePOIQ2Xlx51DKcTHXmbMNL8UY2IBtAKmHI05
K2f/EqQpvoG+9+3oxsKnw+NU8voPlD+iOXCMrP9XSae5gLC/Y0d3Eh+8cZk9Vjrb
A9GaWLT5Nlnovy34JDHx4qmZ54Ms/ZlMQPDyTS/lIYNddqFcVqsdVIADmp+Soj/y
U1mrX5EpPAoH0kpX3sR52G9slmPe6v2CHrHS0r0/hIEVq5SYnKiv4FFsOmOr4Gmo
Ja+Y0Wfdf4J8Wzd+GQ4jqPRnHb7S9Kf7VthE1jJy7HFL2OdS8+17q96/SVcLidYV
WomHRomdeZ1tanHsA3qxnAUPirpds5quhGejGgVACFsHp5r1tHicJ0W8nKHbUxcS
p5KCrbCa6RIRk75vTDNpV52+vKuMVxhxrOtmcyLj9s7E6aEys1QTcbb9hdZ+Muq/
+GbXpU0zE5u3hC9nmmxPLgw17pI6Y6notFWCtzezBvxOFRe8IKMftdIPjjznKsho
JkBlZbEKha8cdAEKZhWb5TvxzGw9+uKITT2MbK8E3bplBEzCOQOeoBBfkvS9P2/z
5OcLk593PbqLRfTCcREaiahqmzavWmEuYSqWXOflS16BM3JAEX4To/lNLkfw9SRr
fgOIhx1smtXuxgQ/BGTxKiL9lVkMYFN7j0ssOonWe0AyUhSSsha4l1BBwAUJf1D6
e7MI+RQBXsHeDUgM9Dg4RHYi2O+miPSYQ0jd9YVVqf512oymedYkurzQG7wfvMyR
LjgnadmxRJbd0tPZ++Sp4tY0t+VwnHAL140Nj/e5W8BmKLxSvTTi3039g5nHfMYk
IC9JpTOWnwbGDunC6h2f2rjM2bBrmhWgr/tPJj+CBgDkEoS45TKwXn1Wrrc9ahYD
aXdLYLrXGOwXLRwYH1tXR+bFPjddQW6sGun5kDjsmkwB+GJg7x/IZnF1ziUJlYxO
KloC4ThUxiY3G0uWXecE32kqSgAcmviMmMpS/9463m8BQWoLa2tJhYUMoAHtvP9J
KR/aHOdxbqQoLdG87Y2dT3odneqI+YZLUeFxHXZXEf6zQx7bfxm3O9w8RuThB6yO
Ck547/hLaQSVar1M/JhuHeTo4Vm/4YKniyINRH37oMY03vW68asulxACO3G8jp/X
NMV7kw+0/eBSqdoiNLaUBepQLCEHjKKf+Qr1V3mPFFjz2guvOhR+a59emwx9Ktuh
pk70krRjwr6q4RPHmyFmR2Qmszc90+wmbkRzh9lEv7OxihG8Vun1AR3PeTCQPbJe
9mBeFnITaampU6v6dgkMDUPoTH/01/pAYt+1n0fQwLSj9+Pzd/QuDX3cy55pnVOU
jLOGJPYBM0e+wPdU9Tu5k1I4ZRm2w5S6k422VDKcUkp87k1FCgkt9AAAkrgt+JI3
2HYYKbKvkd8IA6YHFyNWj8CZqhkPQ/+JVPJqs4l7fm0zrDlHTqnySVLyEKcKDfPx
LUsJrIW5Nc6zCndks8eSWLZ2lADNU9/J4rpgHUHs+HQ9Vwv0+MKn8pY2SY4hOHqC
yuql3PenCIYTmAeqmQ2Je9qEmypzO/mLXcmboYl16Y/FJHjOxTN5+Maglit4Ly35
cm6rhKjCQ5/ckzlipE3qyph6q5zZA5wI702pnoXFoDTPfVaLhOSEMo4tMt9F6ZIF
vKyjmrGr2NRE8gMYcxnh7m02LKJws/0uEiOcU0UP2SVI4f1jpdI4lASxMfUVg47r
jA0WSD4ad/AYZESmU1Aob/FisY+i0o4gWasaEUmfvkUlxr0z5xjXAsGDwKExRjgf
43VpzBzIx+vyNkmb2CADpFP1NcxInpl0MtwZdpFmi98NznzVcTVaVX0sQmmNXezu
HQ95nQhWiWLf0eLsuf/cKzC6gMo+a6ijEXlRdHuc61AL3kP2H/ZTrH2s9JwVDVUm
Gr6VdT6CyWzLqcI4/WmUzbdsS0ZvTBTVSF3zzjuzCmu4VJ7ce2AFbiIzGoidzSpO
85E3WjWg2BPLs08FN/xhevHtzUPv3eTyf7GgAkX6S2XJ3vSyLhkGKzl3+B1onDM9
iZxS2UaJeqSrXbSuef7yOlTke2fjbIivRWD0RERPIbXjtNPV/dYhRv67tlttS108
XhLJC+ywLZaBj393XtAwuU5V7Qnjc77qsi2VifxlroPd6PtmI6kV9ZbXHz9UKuK8
Rnv672kI/5hv748Kfnc+I6QGhiVgRPZb39yHzPuj1V47FG3CK5HHegPzw7opYbQi
atqtTc1dbbX7mqMQaD7efgdHV1Pu3IUMft0LiXMdS2+Rt9/Qcdyz3uTVI/OxCb0G
Liz1haGQJcNLfbq6vNvoPP3eMJ00E83MVUyc2/SsuqEBGTKM7SEIw5UeKOoNLMBb
yjdXOQj1xYar5mkxFzfls62x9WTjsokN1fYL2wz3WvqlyqWEdKFiQR6k8KH35K55
RIleggV68BywBfNU0PFw/F/hEBTc+1muX44baZtI9AA5oHoHW5Q5SVUFb9/QqZGk
xo1RibP1ARHipHW+iUTCe0Tx/ZJUIpJBj8qOFWKa8PMF8Y3F/w1JE5EbwGyLt71h
pKTDPlpqcVxMo5qaCSvzPCTTVNCQvZOdaimg0lIcZsB16rIrZf8HK5pNXTg/h96f
zV0QfQaBuxnB3kIBwKCsg2n2siz0NPHUxGS85sUQZcO8u8a9o0B7Rz5U22NVLOhy
e4d6Np6XUt9uKZwGdM6z6hRwfCWyzC2Y6fZffq5k/w7jfEqV7I0uIcLhc1QL7k5H
KznBYB6m9xDG9dfpi11Y9HtjuPvJnWnCnbFc6gmQq7hXvIHMc7K6nMuEawsFlhqQ
YtKNJ1mVRtWCPdGSNfhNw2VSsjSj+Nz0fcpQZbh5+slzxjVTbhfTXKZiOisMBL1D
pqdbWFxRD3NNVbsE/ls65JuVNpVKUnCT0Xv606P5P18+DXA7rtbv2WkfTprzf6b8
6+3nz1qs5+aCYAiMdNySk8RHXzkXnNrFx2OB4rUS1k8FMjXfHiEXEIcpzrnhIPq0
PNucLyZeJL3PYnNIxuo3wldmUga5ChEYP6caOM2EtMHNYRVqZoWlTtLvQsQdL52k
9x1U4PhSwFYPFVCsAGrxwX0echLBHR6nueF5OAmxZp28PFQ/dX5arIysQWfN8yO2
iLwDcV/TzrVmsbCSWmsOXc4Ngs9J4gEY6HAt9CiaE7hQvn/HXtlRAltsBCPxGfa2
KIejBR4x7jeBclJufHIjmt5hOHrr4NeoLR2avK7jGPk=
`protect end_protected