`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
ddtXksX2+yylW5zu6QL2Lhnb2d1sD00763mmSITNX595NcHTEkwn0zB1Dry37fOW
FufOhVzEJp80NC5qZ/+F0Vk7Ik02dIR0elf3clrjeJRK85K4e3Hoo4xn7YbFUIms
l/8VZSb14+JVGURjfswrIyCUotIzlzVYZ6gzoZwDXIi5gQIBf/gI+KxNXPaKV+PQ
Ufys/12rjO6aI/pPlqSm0hCvftmBcnezN2hk1UeXgOIuKZnogjOsf0iJVX2aOOWE
6pD/psybjbnsNB6kH5uFTA5frkzIzkzl5d9+YDm9OyC+k84E83I/7/j+rk4L2dah
QJOvksSIzN867/4Qt8qYTQ==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="MvBXkzurAa5VTw+1JJ70nePUfoQXBvZOku/SMmg4TwQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
oRtzZL4VJ4iwysPsC8SXYCzXS8Fw2gtZTOskLcDV+1B9Nzn1zTyNtlo6lNICRmmK
ZRVu2BmCc2G+fmzynYlNTnSa7C0Cuel6FYpxCBlOuk3OF2tzAmLAuDyOH3Z1Yjzk
a0aHuoCdIRKv7BrZCdALt03JeUmXKPdOmIlkVGFl8yw=
`protect rights_digest_method = "sha256"
`protect end_toolblock="Jn9CQpRhJt4rnzZPRk+dOpzAubz7omckX1MrFd4p81o="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 10240 )
`protect data_block
gD6l00tciPUa6pDNTk/+t0OO0nC/UTtBwLB41d4inuAUA3i/ALrNyoJVcBnAmEQW
ptbcNp5fxEUJjnOxnedyZEuEBxWRieZFQnkRdF269oOHRL1qA00mhb/ZYmD57tZk
fJ8mMb/EGKusw9/aJdaUm/72fWgn/fZE62204vvFNajA1YwgNLJryOJPfT0tsssX
9YgYSXlcSOEiDCpH8n0si8qhUPvos1jHv+FyGouP6rfhaz+1qt1MISJUY5wQ1XBc
WlDLqFVmM8gUfOUWy3qE3Y0u9zFbz3dpmrXbaEXhRE1iM5tlpgz6kYyThIBnXAVQ
pR0d2cXGakvIR5Cdu0TMeCmcK9Tzmqir4oJ2XgG5YWLjXeQYaQaABvJKur2UGfQf
wzItkLL/Uyu2g5BweubPNWxUa9O82+IuKq0Hf7RQwG3BtE2dZkMDsw2aS038wjly
zaBOUXsLD560fiop4iepRYGIaLPpNS3K52tWQkmCHlNIWDhfgqsHE4+nqlcyOlW3
ubJ5+giiZnrS6IOC2bAJSSAe0ZQYD0uiSW+hYzd1NQvREqQLS4mlbRvUFQ+ha8U+
RHC//a2FVDxqMt4EzWtojMV/sHqDvroWsK+dzl68BkAV0xoRDuGGTe68pA6cjFz+
oCYY3A/T8clUg8y0HuwCaAXpwvWabg8rCzhVa0QV4nx++48l20GvGcZUaxW4ZmoS
GJQh5fIP3qq8zPaK2r1k3LbLUEsTFoT8COFDJ7gqunyiNYjixjOGloFUyKp9iuIz
vbb6rfJbu40LjzjrLX9yLsq8z9w1PWFXNp0GtkA5Ad4kZjnDLamDIecGVZzhyrU8
AXgbnO/rVDHHFEiFe3qSjfq9RtSk31K+aaoK5iQh9xSPodu2MA1LdDCI0wwiblLZ
74ZOQDnA2y8KYk9lq2SW//rihjtB04665uee05J3cE9I5jG+ZaueAyskTXYGi4j5
YoiYKxsDKUJ6d7YEJGc6OIN/0aRKqBJ2Xo9/33YvzxAOtFdmNEeYnOnfmEj4B4GF
cnS3PfumdcrpuKwn2DCEoG9CW5GVOkxQwKtxLFZ37X8jSTw/5ktIMWtbC273YxXs
g4Brbw6XtEbS3OA1GiRUC2h9yHxTX+10XtYNq/lV835LKoGM323n/20LPtG9p0Gm
LKCfLi3ljexCaDTUiUDOVfSTpLBN8DtBaUICXuHLqkrCALTwc8x95viBqoiMKodp
NXmeyMgs8lJxowWijF2SZd//BFKuu0lUgYnE8rq9xL/6KIG6XhcHFuqpHXusgyqx
Fg7BNj/sKkFIbbWPxx3OzamKgbFudimQUgmCKYQnRrWCt+Auc1PL2eP02hrt7YwR
IXPkOnLlTfVjMR7NK7Z/rA+Jb0Umonhwhql1USN8Lv1hPL2G9f3B4uKheW9ec4vS
GNTOvJr7OozTBlCh2B2VmWJqhFa12Rbwn88LnS5Sz/JwlZVdNl5AfTZ2X4gaALs0
KIBVksL7PMetEkDrW8niDlDYjjIFsU3+kwu8qLwS990ThTrQkwxjpKW3//NB+47z
PLDS46iOsyalsZV1Ex2ad4zPUCxgHnGipn3jnRXZSlTnxhMOmzYOmh48xYwqWjlp
/zr6voKjGKsxKZdoNlCU49DR2WtMMeNOU7GoFPDdCe/S5xVOXgeRcNW3w7qI6S2J
jiOkgYx7Pn2GJm9kw7t+jNRbnQuvpBexTmFdbUwgzych35Fbky7INcqw3llRoHzs
8HxuxkQrmsdf09GOQDZ8Sv02QciykPUR3J/qrJdxdDwjPQYh/sOBkJ4r00cx27j/
F1f9wzoFDEpfGUo3Bi/o6Irzh6M4QsARhFNQ+Klex9852/LtiaOC5ImQ62StyRY8
vRmr8z1lMdE5V7AUsrKT0bftkWFq1+cUu2jiB+ml+Jtw8qaCiDTa/3y1O/Tixoyk
fxtghAdvF1vkllifErg3kPgiyGDx6N7nn5YERufOPJIxvuMvl7nvu0LldvgR/LNE
mV5AjCdl0JfdS5oDg6Xt/q4XB2dKZAE0T/HoF3HTFOM71yJsxnr9w4utZmkHgS97
nmLRMQcdyzTwnyTkpFB167DskyRRHQgCg4QrzPFPLkAOIjl+4j5Wcc6BPamKhOkv
KkECIKCNrAmlOCcJx+HtnB24q6PJG9Ml2NPZLvs66J08yWDBdX0G+qtvI6sW9QE1
TxgH7dJNOpHmqz3GmPeA/rlyVnC83IkAgjaKiZuh5BnXKvQGgh9xe7H27hKcdvc5
jXHBvfik3jEpuBRfXIaKa/+/+Whi3IQ4Bxq3Fx43UAqvN81wiqRkOVddB+BAfWZZ
TOpreP3Y4AYpAgM4YoRlEQsQ73PFGIHONsYfdbmjaE/UUfhxZACiNhnY6f+E6diD
vtlm/jZDkWaVGJD7AUaEWkdu0Ueck6f6QOp+lkhnyAlO2Nc28LNcT0ORJpmxEEsY
b6QkSi8Fp8L3l0GT+4293iT6Nzn79AiSW94NRr/HX1cnmBxTV9WLI3cO+UV+nw+p
aNIS6qNE2N2CzEs5tl4fJ+PSDGUDaqVvUxVfjJ2sCIurCWpQgNirPXQMXOMEbb3w
Y+umAhItyFaE/RRg1+X+3hz9MlVOPv/PbguwyGVk42VLCNmYTqDD8GHYkk5+1B33
QQPMhrPukKLCAMrY00FYHzurC8O8gwI1BhCW6mMCAFmCMmnRsN6qxnGw5AlTHrpr
tjCir6H5hykOpEwG1KjaIdQgcrbKsmNekAqdUkXw8OLXvgEbcKcY52Xs/2zd6x2q
xW6LUw39ynXBQLW5dksacYIMTHmyA0xvwVYti96JEIR/Vqbinwont34on6xf3M16
NodRF4pbvg5h35kFBeUy6wHFx4qSo3jzAi0C0ki0tRvtLwoa7pW8P5vAKyhVBY1I
AQSMVkw8+udyNVwK94y3mEZkDOLNlrsLYvqAY+K4doMD9yAI9OJ1tMG6wik+jKAH
tZNjb7w8HZp+J4sFX9+qQBe92Azzx1nfd2lSws5RvHTzn9tCHKO6tt/4VqM02qbL
m8UcZv2ugLrR1kyUqOB0FhKiDxmK312RiAdgkmyVU923gbKbSlRF9d+O8/IGfQ3X
x7DpGmg1H2pkNxfNTRdeLYYZqGBmZj1dDFaF1ipqPv8nDMmFB46wylvxglw6jerb
UBdUI34zZbisMaEhcyh9QyEXlVEk/Fc5hVk7bL4U7qO3fAW383YIBn1PW5zjdknX
cvj6phDOBMEADCi2dRV4O+LQLron/GbAkG65Z4Lsd/UCAdQYO4hdU+CA33/A903T
dpBUG7cL5CIw1t2+MLniHZK2A5TExFyP+LcETcB+QWIL3jjPAtvyp3ZR9v95OSIA
7ILW0oZkwR3Zv3nLKOaGaPiIxySMcIUgMlVZeTg4rpBen3BB45+wqCKnJ7kkVLM4
NFrttKUt0NXqNKegKaAGZePdo2lFI9rcC+TBTV9ekv2tDBq2UsLTdvdrEvkhiExS
UiZ57b38x7UOQbp/eBaa2c6jPTE2SZVF1XtP4Hyhe8wUa5fKgVuom/wnu6nmWe/q
q1ocxP5FIfxOdOlEue++ZhSyMG7c/vYh+4svWpJHi0tF7zks5/bAjRm9PtkVKTTO
ARVUFmFe2iqTpkXvXI243iZc70XVHBxOIESXhMWWYyVGBqajtykA/LpmwSy4iVS8
tJBnjFcz92HzJM2N2eUozSZTLvhwfnt3HO1v4opEjA18zT4+5n+SLLUVfoqFoPlk
x/KGuqbmjqzoOlNMkNP95t7gmqVLTmi4JrOE2f+SqLec2BJToZl8mf1d2Y9g3RC9
vYnvaHusUq3Vp0uIb1AsM4i4I/ram1DNHs+LLlijS8RZfhWSd7WMTsHkQy8sSZr8
FcKjw0YHygEn0BLnOY5rl/TtJe0p8DMXEf06HZz5mNS8lyKsJpxwSgxjCizcNHfn
O4lbW0OtiYoVtJ/xb5FVcQmJOTiF8I2pxzdFxsR6Ny2/kAAUi39vsJ8T9oZgGY2N
3H4R9wBFGVxNlRi0Hat2bXYkj0os1VUaJTQ/jZkBS3Np6jhsjdONaRJftm2hGXaw
RMePiotU6X3BVhEJ3sDhE7aCgBYniniwzSEHGzzaoQkTCbFTt0lymDYcByCzR0sa
QsJA7m4NnQo9kJJoGn9sAqO0UHBoMF1clmZpOSR0iD4nm90+9ygtgehRnsZrOVcA
k8Dw86qEJ7yXXj0PwvWnwsqyONyjd903NQ9fUG2KSTyj5k37J4zcKM8BAlzMcuJP
2hMhCyl4gB9IyvhrV2GEsXsqROo/T5ewbe7+Lm4UzMoDeMN1NAN1fjbDw1VVXdf+
XrzqayUqvr67HMCUGQuRxgqqRo9vWjDTJKVCC7uWmSDNK621Jp4OgQc7dTmFhSai
uwOejzpivdxczGncW/xn2IpYL3SabXdxC9PbvXlRfziUq94v2m3CO+S5t+paSuoQ
Mmql2dQQJXqJxv+Wje0LRcy72xXKoofV9hIYG8IZxzhEECSpLeOGHTM6pI33aqV/
BmYdxl3V2pu95VA63OkCuYD0eNrZZc/MmeMKU67sOrnvv2yGO1dcKC8LKIAN2S5c
ELaOtBOBGic7GC9zJLxk23Jq/usUljRsiOo1rGLdh7XN+78dCjRRiAM+bgpmTUjj
Zo+4cPonJmrmnwute+FOa1t7j7gjGSuiW57aiXrSLpcYPfPOaCWKOuQ3BrKa4CtG
028E7XhZ+iNQbBtbskFvldK/Rm/hFBIdVuF44X3mHdi7W1Z6pxFPF7KHLUiJ3UYu
pZMtAVjfAxlsrj7WZljogg3VMqSj+JoMLfxqWNql4wV4+w7hfhI+bst/Z6aCVDeh
vRF7+CXCLFIYaeK++n5qYv9TDpnZ7Vf887hD8QAJHKJyGIsGyeop9j0BtZP3GA7Y
6P3BaeiLyUfhhVznzrzly13DMQ4VGyfGczYkLdC0YPHnNxRZutjP2Doz6IThtAuV
8GcHzdFDtnszl/JMCQIJ3vjglmbPEyL0TJki1D96nTxduSr8dNajb3xz8otwjunf
Zdo7HtSxHm50daw/Tol3K/RvXaJpI0L+Gy9cVVWP8Z+aSRXzbDMpMFO9o/3k0jjt
GjJ8h9nBy7aqK7ISJ024hMFdx5KWwty12PfdDqG6yLqppw7spodHwiRV5U2MYCnz
yoek9JjTAOo1xMKijHjv1uwH2JMlQXSgt+tjwzC+Ocg/1VmVo+YZVHmnYc5cHtK0
NBUMy5sqDwSfsJBUnpbJHE6Uamtj5ZRgsd+o73oXUjkgOJtWT1aedAbpGwU/xezY
/wvyaveBpCaJcu5exV2YPgYXDiDwctgpdHSpii9YaNocPCHFVpcIbZAoOa8bazwH
HDJdCM395Qtkb9BD6R3n4hWrooP8ZGxfuxOzlRMirAdmfpSdwy7eTHgIVPWDddeh
qf97I+gix9mopXlvpEjWkC761NBkV2eE0BWTYxylvIjdpoXfzscsSAYxq/u2RHDX
5FXxZnoYhO63gW3L1PK05T4QR3AZuCDI372TUqTyUtqZ7lCHElZA8bHXNTLXmfRN
clcIYodRLCkLRFUjv/WKTuf48MOU9icS6j0sMqoDhzFq8r5doP+iw8/X2C7LEaRe
a5Wl6+KjATqxUnNIhtRoP+rHDBfkSVKk3VxiFQZ9D1e4Mwnpj5/xPazxGI8aJFwZ
Uyzr9yHfrhIq4+iS/typRwg2rViMMAC/F7DM4yhYzwUC9b7oo53uC5ZG3aIa8GIM
7edple4Mn/8lFpdQoEVV4Y5q4bNmQJGQVK++jzHaD5q3hRQjc/YdnsnCaG7r3/Em
Wj/twQ7ppOccHzjnM2edI46uKdNobPZzpa5UfOATkhuWMkt3aZwCg3MXgU7oYmEk
GoCXiID8rmj3EKh6OXSsyFGtrITk4vcnvD5muFNGNX/SJQvER+zE1rXvajruZfMO
DzTCTFRG6/ALqcrnTvfQ0ZwE5VWo2JQqLxmLTeddmd6gP23B5fL2udzUczkk2abA
iWPG2wWUFSVTHXU4sky9f/sIEqHf0cwVyYnPoaHLnv2PWo9Jjn1rlsKa+/5jTksD
HiXQACRdV4AwnXsfk6sOYJzkReK15Yqvwq5SpaZ+lUHHJn8H7yArRiawa819pjSO
q+cFocjXpKsFbCt62LS1v5VC7zJEcuRzkScYbhUKSQaYlg6VlvP8Hf8xxcu8hUz0
2GcMxKr5JmNIE1+EAymzBMHWbpipY+prWa8UC3gV3texgqW7NB54rkCILwD7lVxT
J/SltdF/DyoBwXQv2g7hrbQFNJSIk2lTW6jlXuuTuG3ml7g/4WiV5RSzpYPOENTd
wiUlwZ8kKZ8L4iECmIecLzdl2nioB36EH9yNaam+jZNdO9vFqtwgq0QXf2RLYYhk
tZtqL4hI+BeqnNLfh++xw6WVEwIlMT3/aFKx5qh9HtefW1W3yi4kgR5z4sfGIvPf
VN6faLqKQK27MGnjNE7KriCOxVoTsHlScC6gcQCNpuWE0PIrXJ/Lz/vV+1Y1Z0f2
Q1eRRzLUcgBHs1itSBaaOhx21WSBktBgC/zaSCVaiMk2MzNsB6OwFgAZwDi3w7rF
5gsDZL13ZUVrAUJOj6AnXnBqVaAF9shzj0PjXwn3bRdjTXx4zGqAaBdkdrz7FO5a
kIapBWhj8yKcHByPtXy1XZHYYbL1qlnUiR1u2YRtC3nuXokQX1wH0bFTVc8Q5Ftt
lTiL95/FBH6NkeFCykJjTsiylukIm5tpGSbvafnjOmT+eotu4Su00aUETfcr37bu
QIXIoYFvoyYcxl9pOVvKcyXmJwl97b+l2r9HSroutMXnhO/Cg4ise4PStCFMjsVK
F55uDqR5lvQXP9KcDbdKMyVdzsMb+/QNnLs92HLm4ClyA5RFJb+iV4yfoQvWjas1
pSLutVglvrCAQR3tSgyTqufJlvLuIxHBZyxh4L5cWZkcZAA7lmn6DMgFCYm+sxz+
wf/fn0UO6dJuh39pzGNMqs4HGt/OjRK6AKTWmG5xCejDyhIKs/S4aAXfZp53hjBe
Qso2WXts8IP+a1ke40yHjbEjvnYThNcMIW6h9UvA9frdEgKAjspAfea1rW24TsFk
FYOuUMpXlRuEwf6ERLjaD0Fenrtk1sOtTawcjgf/qJUDCiHTsYY6goEbxFSAVZ1L
WpQjrfJXsuNLyvF/lxbJxJLXUt1i5Xh8gzIap1CFLYxaVuSrqnQszledhIYazsGH
rRXRrjEc48TaBGgq3bl5ORKAnoxVOBp9h49oSzinZz3vD5MasdxuqZmYDMA8znRa
GY29+7tNy5BDua685AAXcFTRdPbVwxuC48VyqPJrD1HGg494ViXAuotyuBbZmNTg
DEG+nLh5Hz2iaPVtDQkBdcKgs3QXSzGJCX/VTJQIR7eDaz+GKYVtX1yMVkmSIkkZ
rtXVcuzh5iqzf8nBCZVlwL1uvpxjjL5DiZFFqCyHNbCdrOHDhWr5sjJXbYxiqSDU
qO9+4bGHIZdu7DtQFShUXrfRMP8/4C5Dmce1uiUCXl5hbkIWqQgMMzh2/BuqOU/m
VQGjd8uu0+e2bTalLD8i+090TogqPqcFchHgvOnIkf9nA923PbhXLNw1O0K0fhUc
jCxOFGT/KClTR8yYKEjbHLe2hju8bwlHZR6g84vAK2UwT6/ObL0JHOfIYEkeJd1z
kvJF0OwcfaWWy7B9jgGVaw6qWArdPLjSJloV8HlvCA9ShFSHqqkDf6acOAB6QxDs
nNl0fZr51TrZw2LgOJL4syG7J7XZMq6Z+0vY0zeCiz4W8TugK2akdXh/t/rxhRcr
JC6p9z/JhgJhxHPs2R1UxbwBR6xqmxtvcVp0Nrh09rQ0WDRlc58O1tkuVu+iht2b
f2TvXrsdBP+j2vVAy3B9yqapuJiAMVUrSoTj1mM+B2JX8317SXOV/GOjAGDPUnhV
znKjN4bDmbbRskBLdD7dL/kn5I8t+LlJJGbXZJkhKKWueQaRYETJVeils+UR/WNY
k1FFZ5AZpu6+2iTyBssh9w04bSWzSs2u7sJSO7KnjXWwYYOuhCoHW9gMK9Mo1b+L
JGbwjJfRk93Bh6XUk7CV7tnZZu0SXbBAeoCmnk4S+tZVOP0vDYzDgNkWsJ47ljVq
HEETUwNJE+5pyzMhCM34DvowDZwCaNLJiWbVUsWF+vY29a3DGF1jF4oMxKtK+KCU
u9DX6ybw0Ikqnmi7Q4TCnXXLp9oy+MyznOkMbagpf5OMJE5TaO9wShO9+dQM7YyQ
F5YTSlReQm5h4GoxA7dAIwB3CmgO7WjTknCM1/j5MqA6+TfZp+Y/c9HzQ/ihIRCU
dmLF3OWXdYx8+8Yl1lMYVewI4ZbacYVVF3DUsZ1pZmOydiOB2KxrtBlqUfE+UZOt
5daKsNQrWkAPHsfH71n5zhwLLqVJQ5VAxSQrfaag+VvogMlIZhUtkzcbbN6fiIpw
rPkPemjfosvQFXVFpOhHqfXSkgmVe27n4XIeAohetLdq/XhNc0cfHrZjDvGbH54V
GxAuL2JxicWhglPbzDwLIqNNwBvxy0XYTwfa/zxh0xWR2rcVJPAsizWLNFEv3IXP
NVqVkW/5ixdBH7ukUcQLHk5SOjGGPLLsh6nARubIOAB/2MYnndYh6Dan4kXuwczT
8nC8J0fW2liVoJ4InV3YEI0ON65cTvGEPpJn2rLNvjnTAFdcU1QHNWtPh62DY9we
w5w09CyKsJ+4wu15xExqu6Om/v6qbeQPJnLwc2lLHYTArepuOt9pZj9Sp1DEF7wE
kPRM8rgz7Ol3eNSpWduVTTYHkVcKSX4ScpakDKlgi7IbNfxx+SIY8WIxAen5GT/E
tvDrAz1A95wQ2crKggeC0MI0ghLEx4MqwU1L3RR0eecuvqp8wixxFgMG1MnB1meU
Yye2rj2QBGT63QWV2I2N2/j7M+M7STZ5EqDZXa2GMpnNuY/JExNkafxTxp43Mh5h
MDlZmOIrh4e0vDqOSWbwfZ4X/6zUTgCY1ChrDW9Pto3LhY8MwQKmP0sI3smOcVkw
32h7gLs2mn+WB1JPPtSbyLfEw+FkjoU2FiFEO/LfEmlZ6WOxFhuUmJOqNgedTDSE
K/aLhKuRs+VahVtxWapeOXQdLkSs2jltBO/AaS4+FuCEF/ztoMms14zzzDMyhRds
54daVTdSKjU0iXtQG+XX/q4l4i/9YaBDAdqNsSIeKvAQx5jLChYwcTGEiE6PBaRy
0M3U9EX5k0iYXGtdOtOtPtlNpbyEIiNFmgjE6Y7e0QahN5/HB4WSdUa63Let7BLK
2HWBhHiy+6sEdAid0dXH61aY54iw1TSa7BLRXLLzmnrtxeiQrNj7+LxtdXvmcV+Z
wYzqXRoHHIUhGZmnisOHFZ2e7/44pCrHNQ5nBYH945ZCExr9PqEmatDf7B4CNhq8
mGNlSzl4T0hs0Q+bjyzn/61k8hw8a3NR+UNBMWOiNtKGm7zSUq7DywCIGUhzC2Zq
U127Xfh+LotTfR0DqPuJVu2jJ30Zei4stOqjcBOJVY5eupzORwynVda4AbvpDeB5
274NaANyFds92JA2lx23QFlzMsZzOtLxw35N74UvIPvxztF4JCtZzBoRUVQyjqJb
PDO8IzXy5ODOd19AVZzJSOyLyEyf88dpjUt58ZOhHtXjEcK9O/2e/tpmedIpimwk
7h6qioLW95TaOpkoz9bFrunzuZyhVK0Z3IqJUAdm+lwSET3z3WBzMI5Z+gwXClHw
FLl7bz9LhtvJFbr6wd154vWXIRBQruczcWL3eg7h5LJtdk2e5Im0F0mqkJ5fzd2+
fG8aUW6wSJH/DHvi1ospzz44oSdMMllmSHNyQou/fv/G5O4Pv4BA4c2CUvFNtgCR
5PYk2Ch/LU1V+e5HkE2Sa5aFHrOiVNOX1+ep7pFkVzRwgB3Fu2W99JjSrCpeT6H1
MzVK/NTAO13ixaRnP/fSG4YgNGGPTerCSV2FjAECIWbp9WvjdSJxDke6fMitEY7R
suidwQYtIcDOo4otk87RgaBeA5SHkzJX65/1rM5Xz/QIhc8CgrgyG3l9/z9TyaKS
QxSUPnDNO/9v+Hr7xbPIhzYR6DiWmfaYstN4df7mq+wGK0JpEU11W856ZOEY0J4m
sgwBYL2sJUB5R4Yrhb/rx0ePLO+Qmy8qkKavI8vnEeJbXpnT8nQy+pyju4TrNUGO
v6pqUg1chKjad902GYOSHl9oEbiDkZCSAVxrhPFz+RxMqk0mbAX97PbWw0usiTQw
F/YnHStkS7WMeb05hE2eg0VkKICRjQga3VRjhmXSYj3FprL1Zh4u3zVkrwLmlQZn
PM30UzEzd95B43RSqxL47QZGVU+4HNsR7Iz7VxlR9bPpipo9NAkZmws8O+lUtmDz
FNLum8ikBZWC7FwiBfItG9fYz2eeS/MWnEw1tGHG3VYVIWTo71TaisNtqVB1+cAd
XzkEVD08AWciawxds0wm5yoiD/baWJ5EzA8wun8lKz0NEYPF8dywU8S2JFqS15Rm
fRQMUfecQWUEUsKCcY05wXZx/vwM6lOISL2o3K/ropffwlZUbnQ8zJPFjeukG/pX
jebyus43aKXqKyBbMaVOyzxnaPdfNATl6NCOTt2TmsCZFpn+JlMDlpR/WBbcm2l8
BWT7woLNyM4ETAKDdwkmLHRKQQSlUAjnJAMliOGckkj0EEmP2MpbQjmw/af0pKJa
Co/kewUgZRGqxPcC9rhu7hQ1xKGUlmlwc4QPtuL5u5aTkOvDAlWtZGaaSRnt60Pe
M/hP4l6hKWScM2PJLrgx7iTb2ETV3+3zoX1MZ2OpneflYgZftpOnZSnqJX3ScmEq
tnNPRJEsEb1j/VAzZT7IflPNxxT6gtlnv6kquuioGbgLUN3tVKmGKPGzlua6wFJ8
0hdiDhw+9hTfqLsQnQIJefBZuJu+7rFblGODSG6ifVs8Tllob8sPee7FGymHWX5p
K0C208wrfGwK/50JPmh2K3jUdk2yBhzmXjtVoY6h0KLWfcQ/Agjyr48ObpQBV0HT
jXmSFKb9QUlFhFJElT+bAiKKgmYm4jtXETUCsK9WOe0yBGmjEp8dnf7iVOhoIHpY
rDgXc4FQlFPMgXNWOs+ShfOwJSf6kTNiXwL4fUSLJWV4jjLOOCDugbITrx6vUxHW
CdY+MDV21YNGhPVWnZ+bC6DhxYj8CAK8p9UPCsR4Yp1YMF1i7PG1Yp5s1DNNpvD7
CE5utx6O51lW925dgUcb/JMIWC4pi3FBedLiEGsC7yEIlO1Vjm4WLcL8raQl64QN
y9IPX0sTItU4DF+m/PLAQdkuK94Cj9PLp1ycTaZ4dfBGx+Tt5fdiJXGR77mdQpAr
87xClG3YF9FWIplTBIHJvObj0uQbXwD3Js/8qyA/6cieet93lKJohYad6vHL7A3/
CaOWRUPEOJZcNAmb7jIKp3XOrXGLkTi4FFlsdInniywdo1u1qQvaMHO08Gn1nk+w
5T3vYqyncJ8EeS+xRCWlArjB0X63fwzqLdo53o7VWXa6yuR+au03aLcF0aty8iOZ
2a/rAQ63r0Y84tQhuUyrsS+Rrdex5zWsV7VL2gSAeZ4tfyioCdB4kCt09czbWisD
W/+jw+5ojgqt1PLOf4Nrarq/plxvp2BiHO+7+I24Jy7QwAOQYRYcZkf1R9eP9jDK
8YNtqro1deGXlsMBgNVyJstajcCDdlTRsZxMIEa7cNzby5XrHX6rE1fFXLyF9Pnv
hcrGt7Fu47w/J9geTW/f4TMvpkAQHb47w/Pjm6PGlWiqN4wmPEMZYtSFYrmYLrtD
1L+1JX7oI40YBVvQrfqqdfa6U16czlqbOEB03UnFDetIkXMU+2fp4gdFQMBDKfZy
6bOSHHNI4XWP8S4rJSfUTqry/wx458pR+tix8Lt9/oRshtG8w05552Boi9+KxdU8
tAxDC2nxkh2X7cDQFXeJOmI3mD/6M74CB4w6kAIiLzz+SZnWRW56CnwftBDll44R
J1ug1r6S29wbjr3IS7xVSVpG2HCAnPA2pbhGyJ+XFQh0xxSI8VDLyAFdXgIO0MeD
Dyny+B8Zx31b/kS6RLlocAq9AIAFmZtJN2irBhNGwBIcFu//UMKYbTRT1OWqfknD
gngdT6GrJQvdbtV2conLOK3NEu/l4g3J52jIEHzmw6s5rl0nKrvNLr+7ElljQSVT
LnosbLtNYzswWlV430UpCxOINy6vRcuGPnC5wJ/Tyg2mxVOQVh/JQjg8zaqnNFwI
Q3rejXek7nIRPtFHvH3ZQ745VG5ud4d9UNWoWXljuRKt/lyMmtUVIVAlHNk+Wp/m
t8vuaStEB/ARtc9qSqBH+98YAUth5bxv7SlzV5/DhABw+ZSRjU7arxrv2zvEQ9CP
zwAn6WB8HVyaVwocakiyDShGKDkChyz2hISUoug5CCc5FbDKvFZjKqMnP+oYK6uE
f/KWniKZ/yTRM6BI9GrxYVtgzWk0/SUm0rtCC4BXuyHrFvmiQeUlwiVBqBIZsrgL
R1fUYytdqu/B1KSYA6EoJfchb3SxnopueZXn1WQwrLMSwqvSxjqZm0P3zVRkW8/O
mkX5smr9o3u0aG+6ntcPN7506vicm53ypxNq+9Ccjo1VHKW6SZv2pB7X8bFfXSX3
Il8Plc8JJiFO4B1mh6fpKRSiHy4hPTuFzijgkHw4yUdxcH5dI8c/kLJvTHEimilV
0GZoshEy5xnFixkVy1PnCYKor/gTghGzQel1gPLI1qrdm0lI4YHaQos5Vr2g1HXn
Ah2KCUr9hu+Jim0cZTJLaHxDKBKyi8Q672w2TZz1u4SUiXoHeWghbZgxvul7AwQ9
d7iHMUq+nrF+JBPolFVb8USxxyOg5PiVWa2aUlKJhxeDaaso8lTlcBftQKdU1V9V
TAT9cvQcd22nlFbmKDqXk76cQQgrKToXly6Y3SYzSmQXcmx10Yo44P2YJwwrOlTq
q4fP7lVJCQ/SZx5TNNIch1F4BdhfUBtAUKYap4z823VIA8MOQUXa96Mw9SA9xWn5
IME+USG0B+f9xzxvws+KQflKUV4edWBJGlynkt14o6RH0O7R2n1C7olRtNOzpL4l
iqyjwrCy4hRKa8Wl/AElY6Et8mq9eK/V5a6pPrY0Yzzrl6f/7n2eYEPvMJepQv/X
TmAtHIgbkGdPnrv8scNHY0RlrS3bdxxP0zz6W5JlwDcP+IL6ifssn3wBdrLASahr
Adfq1Psh3KNCnrgxWrvnzf9OTCOcdl5PzjczZN4zwM6VTfd4LuCvAEEG/KmdaXBc
ylyQkGFZaBmdvh3N2voGJ2Ku2nPF/GjnjJL3VCWEUZk+t88AQwNWFwKuRSjRLAWW
UldzK7395NXnNTHWm6YYrYtEKET8qq9KbuObm3xbvAD4rfZ/EdLCf1Vv2i/68mYN
lr1nCfhucCRyFUCgpb5M88mVbPRf9j5ytXhm5qYhyYeUkbZ22NSc0LaF1lpqT/m6
nC/c3QYOMTT/u7LEgkbA/EtDO/MAZElHzb9oVOHJWNdjoSpzLW3sVKnrqNAAZ9pB
yUlHv8ktTbOGoEat2/UfnfcCD7+Vib1Gqyj+XL/Mo7Kh9emLyTNMwv73BFDBXYdF
2D+ru33/O+gOJeMugXnMcV2kBDAPx61rgRNGF8WfDHYpvEWkS7K1BNU8AFy+Ouhk
Jgw8PJMlxsEX7iTH6V/9+IkKBpF+5D6lS9Jq415Jk/o06RVlm0t3IvJoXU8qkW7+
z3b3bokTRmBfr4hzY8o6CQ==
`protect end_protected