`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
ddtXksX2+yylW5zu6QL2Lhnb2d1sD00763mmSITNX595NcHTEkwn0zB1Dry37fOW
FufOhVzEJp80NC5qZ/+F0Vk7Ik02dIR0elf3clrjeJRK85K4e3Hoo4xn7YbFUIms
l/8VZSb14+JVGURjfswrIyCUotIzlzVYZ6gzoZwDXIi5gQIBf/gI+KxNXPaKV+PQ
Ufys/12rjO6aI/pPlqSm0hCvftmBcnezN2hk1UeXgOIuKZnogjOsf0iJVX2aOOWE
6pD/psybjbnsNB6kH5uFTA5frkzIzkzl5d9+YDm9OyC+k84E83I/7/j+rk4L2dah
QJOvksSIzN867/4Qt8qYTQ==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="MvBXkzurAa5VTw+1JJ70nePUfoQXBvZOku/SMmg4TwQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
oRtzZL4VJ4iwysPsC8SXYCzXS8Fw2gtZTOskLcDV+1B9Nzn1zTyNtlo6lNICRmmK
ZRVu2BmCc2G+fmzynYlNTnSa7C0Cuel6FYpxCBlOuk3OF2tzAmLAuDyOH3Z1Yjzk
a0aHuoCdIRKv7BrZCdALt03JeUmXKPdOmIlkVGFl8yw=
`protect rights_digest_method = "sha256"
`protect end_toolblock="Jn9CQpRhJt4rnzZPRk+dOpzAubz7omckX1MrFd4p81o="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 5216 )
`protect data_block
gD6l00tciPUa6pDNTk/+t0OO0nC/UTtBwLB41d4inuAUA3i/ALrNyoJVcBnAmEQW
ptbcNp5fxEUJjnOxnedyZEuEBxWRieZFQnkRdF269oPW7y2WEPIN+gLUfl11ksvs
UjDAYUmcxlftuI4xXIM1HaFZtFNudxmCQo+iX6QpDz5h2niX8EdfY8PMc373uDVu
E62A1BN4OV8ycEPxaYW3dF6mQd9IYmxdjhXvUXWuMr9RNVGyNDk52N1GwTgReY8b
YRjuoMkQJE7EbhHIdA2A3nkIIysD9y4hqepGc52f2HK205Gk1NJnBLIduORIoiES
xTQ1cekh6QlSXLhBKwE+0qEn8OT1Vcz6aoKbQeJkPZQxAf4jqot2vF53teZGvxny
qVsC+//73CHDDQcXgJSitMonJbTCe713Xit6++7qgRS5hFBQBDff8okd4d9wCLze
9TS9rYqRTNsU1mcDI3v2tgasaxfte9oo+CmE7esm7mRPQfu+5QBQwgB8HR6yGUsc
yNHkoUROZtwj6ZcKWv4BPC5MrYnRB+jxP1/Eaqjk7nYRPEiHDHn8S02BCPevQcf6
/MZrhWfuqxQvMUU1+KaoArDXOzFOMAghG/0u19nvAy1tknYzbTMKy8ges06n1Wxg
qrRVmx5IYpaZ9PcF87L0Zy5atpopVVvWSgNGG1uhDfWQvuOK6iH0ZunfHPN+d6+L
3aNV+32sm8owVtQ1Mbq9YrSrtmD5SvaJr9Yw+lgS+Je9HWPcOYAiDKQEpZz+zway
XLaTK87ZlBSij5k3TP7vCbZ4tX/bMJBHci8R4hB2UYP6QcsmnHoFgFf5BI3qQq2H
gWouIKSz7O5QKbvg7adizfOEKqk8UrlxtvD5J+P1z3vi7FkE9ZCI6ydnIw6xO1Et
tKrj6xeZS90M7VuuQdYigzSDfeeKyNL7+lcHPGWWte5KTelNI+0L6GXhnv9AZGyq
cfLM4748GOBjGt+L+SyLddyDGUU9NWtCZXbQGr5jWxrKa+HTQTdkWrrxo9YwdkLo
bySbRarPOMm1nukqzt4WgnUR8Bijxqxtq9PI+kZoHi+IXdOnRofnqQaN39zpipi0
+H8pfMIyaX9cVc7RPZA33XEkeKCC/U7OOUqVZjv3KvC4IgG0M31NhyxUB18Fvg89
NHxY4ENn2lJfP+84pQZ7MsCHjsPCFNunWPfH42tC5b5l31UKptd4t2gT/gubg+g3
OLw8NSND9yVBYOE/ylqNsCiH8Yra1R72lAUDIum1ArsQj70FkfduIG+6h9KWTS+V
SVL0adf6QS2svCEZ/XxiQVoQu+udTO7Ua+mtfIaAJEyCdJlv6uDLxdb9X1Jcnnne
GLFgUPzeHX3lVz1RQxXsmx7mendDWls1kLT7UKDGp795NMG1biuXcvWrh8SEzoJ/
qZKhsPd2Kd9nFp7WVP3TFXIxrPCUl9gJ4lg+CnjRSgvbCFYMnijlWdU3csgs+nxC
MDsqhrcCW3Nl74t6DrdYwF3GdoVdwCDzYsa5/TzEg9KnjVOO69WByyk3j8IyvLxQ
QmkqrQ5vRfZaxyrjh9jxhhi2Vahq4EpRBXO/c39FKr3i5vl1Eg6/yBqtlBAJNOhx
q786W64ZGkRLsiS2/1qdLtJs1wIVQm+qK6S2urTPmGahrJgcMWy0rrTkEJ/baHhH
RvyObJiOj+QJk/2IKyjiUEPcKumcSvk+q2yl+HPVWAonSUrL5i5SLYNs/VwVh2G0
iGj9w6xWewzJLyGr61rwBdRe9BkyP+mYIcK7u5bTXp0frCzKJwyyTfcsFauIrMdB
t4TUJRbAsf/J7c4+Anc4TIpP+gSP5PZmFPj14Pwr2duPIbkFV0tJIdqnVJE/UGcL
jQyrswqACMCceO3IKy58PpZdJfwdSyEngj2+Woi7kyUMQahG2C7nnFrUwf3Kmsjo
vXRO3VHjvjDNYSl6spIyYf9zmfK6Hy4glDHID8RaGc7/BsVpkEAoksqSQmxPIYrG
uGdVpKX1lEhlHvbBJekgrqpt20ViHUtejwO9oHPWA9WeKg5lgi6YqUYtsDdlOS4B
jVm7+kDeqFZF837Ifeqve3MDEQi9zGKndV+xxmZDZFgyYmqsBVZiWFcf2TUOYfkz
KQ9JVWfxwL9CBG+f7+xTNZPkFMG94H8zHR2qd+/5W0Ad3wsb0RrTnxfQcJTuNvv/
DSsXY3nTc5/SvHEPrwhH68VepDtMdkW+VMGNeKoLC0gFjxcMeBJpO9QmG1O/Uy1p
xsJQilnUVJlwqznMZrTVyGSXrGLfICGteV6jn4js1R4EE10Q4uJzkwBM8AIcipWc
3u8dQxosmrQuECYXxymEYFq7FklWrk1OtyiJY6Sp/sx3FWmq51DT+6gi4iDrgvyC
eYMDhgU/yNdTnV1EBsP79foPSN53w0Q5s5BIxSnJl6R63olBvhl2XDrl/rJfFNP8
dCzSJj6Zh5M7LJ57c1EuD3zWeE25YJ7n6CW+6/z9s26B954g9T+Hnc5AR7dWdHx/
XiBV+EsNnHvGYtNY6+2mXaLoHq5jgmVrhbXXnxgldjHLHCbBEsHI3IUBFiX4xGOU
ZSCfhxqzwVCoew6z+Ve8AfdtzEGgHl0wBAy/cKYINxlPoV96zIuT3cnlvg1+b/vG
s8GudKrjONW0jkWlGkcgWIdglxg/dp/LQTSXcFj8/1iPjlyS+iT9bqLydm0Hpc7j
T7bS/268L5zSBwrYQ/h6I/Y69NcpaqEqHpq0O21u0yOJ1KZY4TjKMWq2rLzwxHPS
f0azxPLZdgZx1wKkil8575KRJhU3Wn8t15Fi2/y7YHbSZ6cIYRb05CJWErTlGggd
4dm7kTzkORkpFMQaN7DUjaz0i+LJXvEYqGM01n5CQuH0U0eWmqkFs5eGM5CvDzmx
K1PsY3NgytJQ1pFwxaLypV8OMsu2a1/w6FTWVEHeaTNxQE9pezVurO1z1S0pGNNb
ESk2umw2gD5ZcGGyVD2xGR9yJ//YLqfHVWIOMEoqiItykRfODgRYapZAJah+COl7
sb+velMQ7Xv3t0g+AWdo0eBQjyOIk9uVy7rJvlUCzX9fPVfWuYWA1qGIZUjsvADk
/d3dUxQmAEuhQuTDubpeY7nCFh0ze1qnoh4vCcpbsqjeJb/jSNhVv9cDNHHl21F3
oAA0RoxHM3lylsGlH2VDPWr2eI3wdqM44pIeV0+wJJqg7kgyxCvYeMBFJIy8i2XU
ZF6uvAIdrd5XyhN6zeZWXF8vw8imGUKJn/YHoKsUuPD/aOgCtBcaDFC13seV7o31
kqlAwIjxK3PHS4bYQ8BhLzB2qlyYcED2+RE00+uBumPlVw5QJfTQ2uoZsTgpvPcA
H8PZOJq0VtUJv6ExI4Idg7dtq+Ood0nA8qL/Ymx9y650ogP0ps0ijJ6mI6RmT1x3
mDNw5sl3Scs6AIvMJfiiDnzkjdKCm8R0xcuj34f8+mjSt9iyOBLQJ/ZXM9g7LklJ
hTewZwy/M3Jldp9KJojEINm8pIZwNTLzW0iY6ZvcdmzyRIC4DJnfs70TZrEU1Y0u
jAYl7pWKxUhX2kB0FrNrC4dKbObgVTsLp2RIhWTW08k6ANLGzsCqQHpimGjp10H8
sTMOGQ55viNDuM7B/vvDuJomwTGERuGPhG3LXJk199NaPwfBChbcqbve5VgcZBrt
n0pmPP2riMnF/jxm5Wmou41LoYWw8aOqvY49dGe0CKRU2DXC06QVs8Fw5Qf0+FlN
XPSWS/4HlpiwvZZsfOnUyVB4EtoOBtvEuXfEN9XE/HTUjNyfK0RhQA4MiA+A+AZZ
fJp7AFAm3uDhUpQmYgIOj4JwS5vIcUKQPwt4rx/tkCS1rSfbk70HWIOPFhnUTDqk
U2kb+IZeWTn9x136yq3uOFi0XbRIuFbrstOIIxV9OCFgdemRVvFmI+k/l3A7pXQD
3YNhWn4/mW/wVn6DfD3+Ylb9yej7fvvDqivXyx8WSihN5Uv7MgTZWctadLxXptOG
DfhJY1eVu9Mp8BzwaXACgZRapSv06A2EUlwS+DzHVFU1utbLTsAYn2AIqdpxqHv3
JUFiYp1GNWwCJHDnNLjakDTnthCWzFkiXTw3JUf2ft54mFDZreqw/0WFPDp3p+lU
yq5eSO5S3TTAkxjNO46RgTczx6BWqxTg/OVV+/ZtPRgJpoU0kt2kAsk5KxJVIwtd
c6OUJAIEEy+aJJt1Pyz0dckebrQjVAefZ3V8LKDLaUvqYPXTIlF5DtSRQT7DJWrl
H3K46QpNCfCx7m8wfO/lgN3ZR/imetKLmtkELFFibAnkb4vjviySGgk5Dg9Tg2a9
MQYgzahObmT5So9MLR6ZdyV2uswXG1WjZwz1O/Dhzi1yUtj2KBmwnDwFKz3T2yOB
MMaa4Y93dyZk84k/kVpVjpjge6yerHk+KSdkTB8WUSCAfMXdllEYMmneHik2327M
GZpSh6YmsnvaA6km+upxZ5Az9Q6W0mWfGNxETTMd7spifSht34NTsrw1xICDr6ep
Ma2XX1ned8tMLWhwMGOftVjcZcS7MNBjrfGaFtudHeZd81gm238XaRfzZ34xcDdS
P806Z0O0jeocLl5n6L4aUABkobFKjhCg2rCTVMB41R8WjMA1+5LlnR74UzOhIbXH
Zn3gv6WiFrSM2RcqyjLHpjS6E1iFi3p2POXmNsm+YreQGQ20J0q3f9RvEi8JC5H3
KcfRGrHCAb51rvZrwZ1ufdW7XwpgACZqNdrDZ7yB9gEYlg4dnSTW/INGThF2cpTP
oxpMNxE7wtTQhjxfiRyxZ2h+RCz7lIwowYUqY0erNZcGuFWCKMpwgska3GEyTf2A
sODWwHpeNJKjiX/0nXezTTZRkUra8I3LMYhJqJM8QwTeuY0ymkfAxU1uY4+Sx+ez
j233cOlqagk25a5CHrvDxcLAop+7XGVSBdeK4xrbhDqzdcC9jiV9sv/4Qy31M0jD
3oDUDuWP2iORJJVsJ9UfOYYd0cxUhf+yjryb1hDf5yGeK9C2WgCeXCecBT7qmkzg
B8Iy/C0YO4+c3jiyvcelO5Cojsj8X0Dwa0OIKgzaO+V9ruQny8DIgTGsjlu5yNHO
idmFp4x1JspoAFqdvjTxGHjQuf+P7d0gIJ/CXhmkm9uBqX6uDbE2b248ywDUaQdw
Nbm5AvhXVG6l0m/jC94ykD/7YuAHGWcFYhfYbL9aDwahNg7Izi8LnrzExF8Q/70Z
jxE+4xT5fhvNQtgjYIbpxfBaW0utzBHBmmWUrTC6Os9JAjNcNkiIcFZeOhsDsU7f
CLKilMIcUo1RuH0P5uYXEHsVjKPQlVmwzMolEsY2vxiZm1UZAwnr6S7Tv5XO7otM
BvjEs1lr8nh11A2aAUsXoK0vVMV3yhGik6AlYkjDrFlpLXJQ7bVwyTFRr/FzBWAW
MmtpSQnep0DVJAlK5Zxr2ztVqDSZNPXZgDzggbsJZgcPLshSjtWy6WZZ2Hx7g2yZ
w5jxv7+JjkhbTjzd4YbBHWjprrQ8Il/Khk4XlUvSIzDimuDyHAlkYXqTkLggKXxL
1jZwPf148DEQn3rqyFh4le9UQhItHSHJ10MBCTq+1cL1d5NGf/245IdvaAzrQxM8
Zh/5Hod58jhLEyCv3G8azzrFY9HlW9WK4Jk26UcP8dXJrzdHTuOqUJ8gs/ahIGtb
iybbhJYb5VO4nmeB1KWUKTVjcHlOjmssQQvsDq4A/rGsRVmK3fgMQEYu125s5Lt5
TDcOLWC90yaO2LPV7sdbLWHSrdHhWDmIWObBF7qEBD9EOxZ7WsIYV0XKCbpoe8rH
4I2VpkTn6bx1o178zc5FnyCZ1+QeXBADNEb9NzENp+ifYBB/TnJtWzWFkSl7m/rG
tiKuHHxmq9xGIvlZEn7fl/t6PSCJMxnPqKQUyqZ8ZvCpxoO+BP249nYIk3FltMYz
D0tTPjGco37l9jDZ5XfzoLQ5LDyj8fjI/qEdAOcThWVYexzuMwFewPb5qjeUXYko
yJL/pY3HF5cs/TRcU8LcBf/H5QjAm+6jHDmnk+n6QOa2USFnhk2/YQeWtvSflffz
gTnGUyMl0k82YCVchEqpIUlquAWiaBhBPo8jdMd7gC8ppy5xaWalfUcT3P2s0Z3o
bN7cMqyDRzRqrzGEiV1/ETttJlqibf3YTMduOTIHcNYO0uI52dYp6qQpygIVor1D
6NWYCSKhLCdVsPGARW7fSr5PpdyprC3pTN+uD0u/CXhCV3tAevabeygE1JhsNfOH
Z/GApONb5E8m95qr3ATfetKM8z85gceesh5y8lcXNaYdbhcSBaMbddXP/fCYJbtE
H2S1Vy9w8YY19lJ1Huf6U8KJLDAVmTM4vqAlS4fuejauu6yH9Lzw3pzvuKUmb2ST
vujSrW25Fkt8b6Mq1GmM5WyDheOTcCMXcQxORZDhL1WLKnK3714oGEI/lSWf59TW
xjJKYqLNCDm0m+jPIOv8s5iBHdRMN3NlUbqqkYFYk17ANgIeRC0B8Loqs9qhxFDO
wgCYMdnFMAsks4Y1A3ouWlGpObtHUkz4qUBhVkwoLMTfi6aLyELJ76o91oqSu6A0
hCVuPmB3d2TS3z5+B6rJPRQIraVYh7a28S8dM9GBxmHLCOwSCVm78B9kGjQmfjp/
hggQ1qwrY88D8g2f66NRIVkC3cpMMQqLnQHp2UyseNI7FM8HBDujAW7fwIukhsjF
IC6kLwq7Gvy+G2uW2F4CMfP5KesvTZmZkqn25oJtdxVbB/h1EZV5pzGVu2nPBQen
/eWm/mzT15HkUFax1p5HmwIWdf8OclUWd/gW/T3OKxIvk63QcYOmt1pAX++n3ZIO
vQNVnbb97iazRnmi+xaEufdB6OIPkaAJQ/HlhG8UzM3NvuR88i87UGZZV88K9OVG
Vjdle+lCFwBiatiTVIczrxx5oAenao/7T/J6Qq/xeXTYVLKlIrpuQnaIzQvdOdZO
Ioy9n2/aA9ZThk0ioT+yFWWJBCuSX3LmZHDU6TORO1A=
`protect end_protected