`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
ddtXksX2+yylW5zu6QL2Lhnb2d1sD00763mmSITNX595NcHTEkwn0zB1Dry37fOW
FufOhVzEJp80NC5qZ/+F0Vk7Ik02dIR0elf3clrjeJRK85K4e3Hoo4xn7YbFUIms
l/8VZSb14+JVGURjfswrIyCUotIzlzVYZ6gzoZwDXIi5gQIBf/gI+KxNXPaKV+PQ
Ufys/12rjO6aI/pPlqSm0hCvftmBcnezN2hk1UeXgOIuKZnogjOsf0iJVX2aOOWE
6pD/psybjbnsNB6kH5uFTA5frkzIzkzl5d9+YDm9OyC+k84E83I/7/j+rk4L2dah
QJOvksSIzN867/4Qt8qYTQ==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="MvBXkzurAa5VTw+1JJ70nePUfoQXBvZOku/SMmg4TwQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
oRtzZL4VJ4iwysPsC8SXYCzXS8Fw2gtZTOskLcDV+1B9Nzn1zTyNtlo6lNICRmmK
ZRVu2BmCc2G+fmzynYlNTnSa7C0Cuel6FYpxCBlOuk3OF2tzAmLAuDyOH3Z1Yjzk
a0aHuoCdIRKv7BrZCdALt03JeUmXKPdOmIlkVGFl8yw=
`protect rights_digest_method = "sha256"
`protect end_toolblock="Jn9CQpRhJt4rnzZPRk+dOpzAubz7omckX1MrFd4p81o="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 9648 )
`protect data_block
gD6l00tciPUa6pDNTk/+t0OO0nC/UTtBwLB41d4inuAUA3i/ALrNyoJVcBnAmEQW
ptbcNp5fxEUJjnOxnedyZEuEBxWRieZFQnkRdF269oMNNFGQrlArf+0RxD78mH5K
FNqdPRdFucyEY9p5N5FNPloMXdRoLsv4lcUs0h3bawzrk5d6cqfklrbrBGpjr64X
vUZhHz2BFTjDrxJcNeaVZlCUEZdGsnHZtVIWyvpuSYkaz6SZsmJetp1H/52jBU6i
xqgip7Nq/L5nulaBzz8RxolXexMKJ360/gg2Y+tPzJlQE8zz8DSl4Rs2zPIHTt5J
4nBDlrujp4cYDVtznBztUZpiAWNiHzXvb09atx5FsvXMoxwLXSrtv251LBYflRPD
QPVbukBHKWeI63tI3lNLl+qTO0mu6hSDytIiegl80uj1hCHj/kvf/Wp0BVR3zT0W
zyIuBmIflywViNuPM6HIIorVTb+o5Zz+NmcW4Gi8xZ4KWivtyCG9SEjkggO7M9RH
wjhy/AxuvvTaHxsyu2uEhb2VWtX14jYS/8SUyQGfhWSsx9aYIGrYYIWta30IKBNw
vzl+yo1oDOIdYMFtqfKGjm3NZxmFLAs27EG4zziqjzXe1WudwcseCO7yiie3u+Mu
SpksMJ0tLsYLD2MAUP5JTjN9sE7/NkHqzhRez6Nx/2znKDEI6cc2yL7XdpEoC4dt
O+acTxO2XDOqNdMaNZ2P/Fltunn1BSuelVy3OTu9oSPAGzjXfrmTS7hOfb+sdvno
qWPTki0V0KKjWr/4vDk++J7xsT6FMtMSWVnWIZ166wpmJjvImGJGt9yPnfr0ICVV
2W0DJZDg2hXnTXoiKjMYAThvRCIvwhXhi6tiKa1CIIuJzuGqH2P/wGSsSDj0IxEC
s0yXDwBaW39xsb4GKYOEoT12nsGx2Y8Xb83VrTrd1ew//6sXfvtP/Kiqh2qykSYv
ISTm0WQrwcOYZL/jDSdjEVk9uArs3234ucWIrjn8scb2P0FWVvpzn0dTXX/DjPZ4
lOv5gNzXA16hYSN7++dJfNDhT66zBzeldDkzw3puUQt5pezX/Mg9epimtidRrLlN
k0mcHCWOgtEharr2khKnnlUOMnAMyVk8Kk3yDJLqOkDgkMfV8lnC/Jq2zzV/JaDh
Pf+Op/MQjYsEuZxAGsG/9Jb7iARNcIcmzGkBrG9MrHbkqgJF9F5X1Fc7W3mF+JZe
hAyfR7MTJy8cwW5/dsU604yIhFa27sSKBtUwnpddBRNzbeK7Q6wmQZ/X5HcvRp4u
mINvj9teNPApxjd/AD2+0XNfmd5W24ZfObuLT/Xy1Y07ysg+8oRv/iIai8Sf6W9t
ahkMWgy21IvXl15VOJRN5fwJuklJGIe+TS45kt30ZxYVr03AfvykztS0hP61TfJk
swWtBNhaMZwWNcsC374ymfNF87s/uhz91yYGGZd1x3cVln/aa2UExQK2t+XbNJD5
a2yhkcRrYn1PbsDxriUoP2L0mKRcEhsF4/O3zdVP7vcGnZ5DNzXW5rHTv6zgSULc
MbU84XPicDwxsz3s4FkWjcGw6nKxa2svCOlCaOW00D5U2noSm483/2FCF7vzjE6a
tzoKqFFdUrTB15s3oBrPFTpU14qTx6zFw+/b4NeXzWnpjowvCWjcd5Adso/MbiWk
P3UzJQh6Tq0K5Ixe8o+JdeeDi5rJyxWc9a8c+mZCzPueXKVO2O+FvuXGp68OY0Yq
+pX+RXp/PwS2vENz+pzHrayzl9cj7obmxijRXissdL6gsbFJLS0fe88TtFyapENy
SuhSnFQMEyaM3wBkG2cT9hpKqWjWmWXF4026nuhufY64x9qzKvIWEF7ZdMLitVC3
vIi2WLsa+mkf/YQ5SLDzDSJOyrO5xg5KHHXmCMRqI7bJyrQ0vuLrF6VoEZxslpPN
+gSEo+7+etx6fg7K+KFIk7iuAimO647VJUtA3i4rJVCfe98na62oKd71efj+BC1A
CVY0JtawcNqwb3nEnkS68cSrzPRx58qfNgWArA68lIY+Wo7x4E5qUiEiyUUvBsBM
IqGeb97eltSYWGuR8FOqwPtqEjXWNOHS+WqpUr2yZ+8riXpAdKOPs1auUWG89O+8
2HmraPVcAWLydUq8kGMzF/TY3gJtX8k6f16/nB7Q4u32NcJhKkE17H8ZnowN31oQ
BDc3GAgmvX3nXfus+edi6+SB/7LNobTZTA46ug7Done1yH6CGIT/ayX+k77MaqOw
HiYhMTmkAjmS65qU6XBDVL5w/WpF7Dy62ngKNW46Q/iaodDph2VJu0rSfn00t1AY
46f8DGOnMzH8KEsNc83MXduyTtb83dzLU4+67U3GQUMr0+rITaEoQ3YhXN6Kmh2v
KqzZ2HrJieT2WN4B1sJwbCICYhye39vTdcbplfUpnlY/alRfVKPpkb7++FCSZUgO
FolxWzzhHa0yAQOHdScj2m519bIiPiO5J4mdRlYiVI2wyE3EIGs4HATd8DAG6V6Z
GkR+HR4hb1QC7vmZDPSWceuZ7cAO8/FwEl2y0uIdC++ePMlVxGDxCnZ684WixHh5
fYib6QB69dFulzHxLyIsi9dOtcQcpnLuXYNbGg+dug1UztyGpW8c6ZPvDwwT0EPH
PnCLo3jb3Hho2A2zF+i7kdNPNK1TdTBMZnWD17nkoBF5Ar2ZNZo782vjShhBssaX
3U898xjtQUKh2/kj8ViMsaSmmZ2W/K9lfUHkmNuUhGi/RmDWYxI+IX7zrhZj72b+
Pu/Vkk/sPSsVd5t3Z3nllGXHnpPyXvHsWCVlJ2f22FW1TAqv2JXf1QVQr3H9dNaX
G3k5NFQSNwyQLMOSvXHOTGaRFlRuNVXNis1WYL9HC3PI/4t0sIcSM60LDIiF+3Od
MDn7jvDb1cQlh40CT82d4ARc4vKMWKC07m6ABtUDv5I+8NF16OtOZgf6jftfpUY2
pm4Qu0s8r/PCiKePetPzA9T6blZVto3k0sKKpWsuKohcdNtSDRmNY61iXTto62L7
RsZpU+dBmgFFUsO5BVkvS83WxJmt3zjVMyjUpMCQoyD/ll9K1t1p+/j2SP8Sa8iI
uHr6zT9eZ6APaf9PLbiQ2Bp8D2arciwnE9xvca/vjG4NFPO7H+ivpK1hhmguiYwu
c6HbNH2UHmAt0SCowyXFCHN2NAC/tipri7v6URVMnvQ1bKl6yKpfxLCDpfo5YpzY
uy1S0V7HAANdzaSkRyqxu0drtsLJ8y0XfquInCGRMNpMLflUri1DA4Aymy4b0tqB
sWfpSMX5JM54lJXMqJBUD8H5LRMePYNKYc7ARRpLYeNThrgy5aXHMGGTefDZy9Ar
VKMJmAL07zd0OSsiWtjIQfcjszOvhTyDJA7Pcup+ynYLF3x/7iqqLVt8ozpbDdt7
EaziC+8wnlkgT7WA3EfOxgLnwsYuK5cNZX6FG++YYZncxIRfZquamxJ5O8Jb22CP
TQheHlMus8NY+A/xX/AkgztA+nruwO5Ezri75/ibaLvKwLT6hCU+nR0QHc5Z9y7L
l2lTHs5tVWIfmZj5J/mKehtpT0nA3Bcvc88A5oCrmlm92ZVgZoE5eYhD+Y3P0BSm
gGBCW1B0hjN9xdeq/+TQfkFu3wQL5IemwbWnBX3YIZnkIZ79go94too0tRNfRAV0
+86dq/NQX4PlhXVz0xlwpm/Ouhp+pIsAJhVltawRs5eixLA0NxhiKdBtEe+fhhYk
p6JLkgDvWo4qCc1HSCSv2FJCx2OnZqQagirzeNEnwEBX8ZxV3wcWdVLIVxGQ+yqu
j9QLySpFFeyMuyuv8LxeWfOuMIdR5mxgAZnZmjl9FFhjuXCQjH2586tGQZeSsN1/
IuPmNAaFs7sitmzW7UNTT4Tzwi+LOLcVkHUNpb+TSwxqmYfyL23hBFtTLNhtxljJ
PHKztCZi83zRDGkFjL6CPScL2CALqCeLu32gcfvzUYVTBsL2taGJQ0ZdM0ggcYEi
tEGK4ybpchkQ1+6PHeQPgQD3aXeUUBe5fLIMGSOL7cBdUfnm03eW1DidXOzLbQdq
kYrJxyuXDhQj/3dT5rU/5HUBaw1pdnlxXdGI+meHIoWL+8otDbYU3UVHCAIV2fKV
3DaY6usrxk2xO53fjVclX0iz4TSjNfd1E5rRuQp5PtAJCsrptLsytb0/glq9bM04
5zDMdUVfc1hFr3xqhqGY21eM0FHKJMSEFSZO2qoL8JV7rJ6VBCbQ6t9hLWn1AkKX
nEyMeSxEO9z7G5gR+l1RnN5qUe8psRad0gY51i2JIUibuGz0zYrEXgElo4HW0AHU
Op6CWb5rP4ku8C2X10caGtCPMggSokM8uh/U/PJh36KxJ4HYT2uw6G0qc9+Loc2Z
0D6ZMi6tWJ6XwffNFP8hXSsDysSo2+OsqWitkq4IsYh2n29kmvnIH3D0md8XK4V/
ggfI2oewIbsPI8iJfgNSsuhwv++5coEb0lOqEhIDd2ZAfFbApGOQSO6poIGOlncU
L+uPH04B7USuJLB1BupGJSJrAQTfNn2T77X/uDVKu+4ZLeZnMB+Eph+dnR5iVxp4
Yq4HPnTGp5G7qucSqqEypaeKAHcCMyMUpxTQcxcVATFgEwRWt8+fC1Z8xY60Une6
JFqrznDFvcEBrhJeUNexzOJlaR3E6AC2lee/U6WbELIMfhUwz3JQO1gzbDcW8jFe
m7ZqCF5/ySK7RBsj1kUG67ukXOD5UVpcU+GAXGVPQYvHaJu9faQFFtZhFSix3s/b
59bCnyTD7mFQ0mVa11DDrKJO5dnyZhXc5UsoKMRUuBvGc+sc78H2fkn9GF3sF1iR
OnbLfChiFhTx/SJEqPGJOhgZ9V//J1cizVyrdgGq+31ngHHDSinOxJauejjO/gIX
8vGj7A+NXUypN7wJVW/4q+0T/bt95yuu+m0OTrLCYU/zI0HKXgucvEQBNk4dhiiF
kNCpvLmUP+CEQH216lIE6v3pV3jp/lmBXhDpyWIUp/CWw6XawwvpOHVhLG2ZJVcl
M1sF0k31MK8XHvxZH6DSOHm4+gdyYOG5QaFQVuqqyuJyX4hZc5XpYBA7IMXJ848/
ljS2MLR4VXAtWcHuknpTdyPeJ3tq2FRxWJO7FmClCxiLGXelbYevv2aar+Csy82/
B5F4Q6dZSxVjJtjCxXra2NtSngNNzpPt5JD/draqW1+f7u4I+GaGHmuzyWxKA7NR
YjEwqJ3z9HgsF32f6ebymdenWXbtEi551HLI+5cbfaMxmgU5JnkuR08u33o+C7zk
loevcGT7US6zj3JLfKNeJM4YDPeJ1tMzgAiTqd0I426g9aD00SVt6/j57kv1nI2F
6YeqkQQ7t6pEpBqypGH3VP6gTKX+UVi357EHIpOklFUnxCLo3KKTCgESszZxU95j
oKbN27GoXCjGSJtkI+chGjSHsZZRMi53/Tsi8r+Ig3nGxXsXQ1PX5vSyM4zIkOtz
BIPk2lwTgd5BGaSYXP/j4DlcWwIVENzg8DWeu0VAbPGvk91Qw1IX7MeISW9zU/OF
YO+GfEbOz5XUtoO2reiq7/YG9taBwmC7r3/8B717kA585tSq7Dwy8VebdimFQM6B
QMumFOP0HihbtxSPxF+K/N1JpbfTKGAazk3lq/tTUU4cvzSc/VQ6eDFrL56v07R9
P1mMsgk3R/ucCeWoBfgrCEKrIV727cYUnre5ZkUuWzQ/abAzH8JOsQ5LXs66vHvS
YUVPgoHVXIY+hCqrEaLvM0ftO+gEsoQP2khSMiYGWtOf8U9c/DyBsF39DD8gLE2t
8vMEyCz6XfLRl6XK8nnfN5p6RpYN2rkZO9iEn1eIug9JsoIWZ8RZ9OPbAO/nu0O6
NOcqoNl1cwfOR3pgTjqZwmTnEPBJO0srtiNEIfCSAKvICGBpq4lBIRR3YHDfkohb
EZtYTT8m9O7LlsNXzV81DnerygXgjx+gVoaE8QkmyWZtRqOyr6F4MSNXdHYEVcRJ
4IZ1wCvoP1x4UtdxIs6POQDxd4iDMZ0Y3/fQvl3y1F7QZb6YvDr4u8FdHnYDxDRg
rxtexix0BSuWjwUc7LBJ41UmSKr49mhbyYG1RaYJH9RYHG5tSSxgo6kvRMLe073F
K5lLmNAds6X8mkgXmqEvYof2DgZXH58KRKJwqHpDYQhq9tsKye3eLqBD6XZX7aBt
OpRKvU/iWHxyLI1nsN6uvZZnhN8M2gACrjNTceUokTHHNwBa+PLm/3QyRvlExwFk
BMPjnfw3CueDeyEgRp5dVFSRXfk699eVUHjsmF+unC0alf7msQaZImzxcM8s7+v0
mQv+BX/XIjSUrwjltGJCLc6xLrEy3SkwsAT451ae8cL0HL3wITY9zakDvPOHXNBJ
Uzs4wbEhJDUROoABJx1Eq3BDMvYYkpB0qnLrWWlfuNd5UnRr72O1K9XsuxHJw3Sz
FaKC13puyOJIfqK7KiKIraS6/hXJWRhzVLlmGHh7HqGy5pgvxXwVK9V89rYFhZqW
V4pAIcTHH/Ayrvq/9ewgHObeGqhufJ5eeF2ey0lvTIgO8gboJbbMHKTVz+stvD8P
724U7jYiIuFcKkT1naedzLW9LGCu5WDQJgPcFq4ppUVBuWOOuupGMvkNLg01Nork
qQrAIggjXx60aohxIsn4r01RPPZULgC92VOTIy+/cHonEHVZdQOSj4Ugk+mCrgHP
+YWCoM+51rbsYOTEx4qRpUrPOUjCA5zYHTDkyLe+At1dvO3u6cApUhqDAdCLMlnK
LAXgy0yA3cqa5osgmW6lU+npBERhDpCq8Vpjq3489ify3NCd9AJfeOPlf76J1Mz6
OI+57/iGLrlWKMqVNlQJDAD68Pv+jNNOuPBq52YZPMWvQA3sHK6OtDNZR9HcHram
+Nxutv7xJaUiH9A2xDX/Wt+j+HXOUs5UsEIofUjVvAgz0vDmz3NFNxywQUPFIA29
EiRVBskxyfPmXsESEu3aQ821eccTcIXT0nW3AmznQ4tajPwXU8Jp2F0qS4JDFhr+
eazMflIc3h+uC+sSsWwXjvpJcp7moCeefXPtYoaC8hSGLbZzeSXR4cT9JvXU0ck9
Ct5b8H0QVJZ0yqEGbBGR05AErzD7c27UOROZEAeR0zfv4antHvirqgN7TBxyrK+d
QJltU9pgSzSI8GKT7nKhDGbEaji0zJ1e3D58cuyXvLYbCSFXu0UAENVDvXVQ6VXE
9NYmcq3b91yZkX4qFiuM6mIQN6ZXqCiuSoyyus0+QGEPM9DWdXNH6+PLvFKlzfCG
ZSO+6hQ9UQg6kMR/r9Ojt8TvVtfmVinhcK58UROrlJ54dH54aqLsQNMh1CVLEf/k
6xb8LH0giSe1sNxUV3aIvstejq6phS7VwVxE5xtIoL+5+SSbNGlEnMW21VbEQ66c
mpoiY54zelZssMVWyBVWbb/pf2I18HL1YvtP2bfp2uG0bYkLtQRAwFkBuEL/TFtZ
YkEltACcSdKw0t86lyvxtKNYdePwjPVrOUt3xHbsKA/GujoOlrHflrBVg45wtYvP
Dznd/AzpZ4FWKAg796P0/vuI1ZorIrgKvtfSUURrb11q+oq3jSFa+kr5BKtgpp1Q
FcrwQzf3X2EhV8AQOwpRTLpS7/r4xryGBKz2dLu8YEvlJXrdUXpmu969U11w0m1r
bPeoYiPyJfXlig1O4uylxkGxNSJAt4atiBesv8Stcn0rfbc0sXamCDKj5L/aJu3k
eLooBC6uYj4C6v77DzBFEeFytx73RUPUflKwKeGH3GOYfxsxiPoXK1rd87xByUkg
LwYkbm6S83esAyPBvsxcbbaZp/mp5++ftjFlqloz6iPe3yp27YhzmL67ElFcYfZ4
OK65tPi0G++n/JjRQPimL5Qm2n+L7c1jmWOIaKATCGBcfdOC7pJrx6qxmv+NJvp8
3kiDcsngmpSsUo3JRY5oOwEDBkQnkBwnzyiZH2KoMRlDwIhCYERPM1iRU3CXfikC
z8J3VxK9onStfmTNjjRWzGtMLxNTrqgzOihUQOA/1p7sIl8Xx2h6lqQnyWRg9l32
Dwm7Tf2OCN1RZjgHxi5lac7AQn6LLPMYejZsbZnTMm6d3/atR5bFJu48W39hIWum
LyIGroFwecMSIOx+8StWaYrruHxAGk6BFeUQ7Ymp1xGUOoTRKPWF9V6d7efKgo9P
/7gD2/0AqPsQS7bmREPgXUzSYzlvBYSg3a97ZyrtSbL6jQsqe3L/Cb4A21MWSgbE
XAQFgViqb6wqI+4oN+lo71VAIW50JNNbuqBrZLca5BC3yEb8x+lsm3WPbs4LwPjV
aqm+BSDOXatauspdWIWuyn9E+TjCh4s065gqePMpUp/Sxrm2IMglLwF/QJELguQE
Rxb/7Png8+4lqdz/lySbOQVpAoTQLuqWb3WZzcT0jiJL1jVyIMFhU5uELF+hH62r
Cjg9sArjSy5Rroe9rSw9pt6ZAkyhxvYktJi7qOjcS8NWdHkY5PdnX31gI1q4rUuL
wtw6852w+8ory2CzhTWsabQ9o/G7/zWBQA9IAv0h+grGk+yx+Pu8z3WIoWEx+AOf
xRGzn1zw4hX6tv4KmJPSpcNzQ1UIg/TvG5tDy2CsmxZo9Kc4n6eYhyqBafSC+Ffj
8LcDeNkdBtrPonp0P7OGgttvy9ckSlNgAuP/DRlFl5x+GMO8Kp1GRlUyoiuK736L
cCElKwZDx0dBDCr6ys6EL5xcVCglehg0iAM79ljjH8RZIyrUT9uqsiYXH3GACrTo
DkqWd6omMtFCB0me56bYn5Z/OT5N3khh9R8mv7NvqY0u1PUxy2gvf9wDa+iWPcOQ
dzgmbq6DucQX9DcJoWRvj6p10PBlOmraqedTDVfgMx0Cs5uW5LuaiXMzdamRCE2v
9G8yT1fLVqKHSZj1WRAStCiDbA0/ddxlFmFjL0jRj7BRuuehOjV3ZCEqojnj6aLs
aqjZ5waK7JltHu6AXHEXpUykdlXHzsrC07TsfedwTR285gBFG/oSU3EJLJZe4ZHz
WRMZ1JsYwKh3R10GqhV1to30B132R/pqGsNZK3RnGsH+lpngoABOVJkF/gqMPdq7
eF74m/6IExQafHcGoM5oUE/K0P5FNfU1/suClsY1lHLkS/TolrNbgJhqCaFZzih0
cNQVziwmulmXq9KstZVyBjmQM7fX72Z4GGcOtvN8/eXDVSK6Bn0mtw26utndZyl2
Wt1TJND5xUvuKclFdOb85BQ0c4X29Dlzg2t1H4BwNME6QD51WzzFNUfxd/zALvtZ
mlmaeXZ2HaY9cIfY7b9V38kvjtxftlmTedBjBh8yBXpsCFgKlmbKDs5FqudQCDLr
7+MNXP7fumgxqcUQ3PEv+WhUinvG/2DAxE4YF0HoTfy8OlC+VN1BV37JYeelISen
w/VFZFVyJaRSFnosD23TVqW4fzZLTBLElyqVZ+J99e9Vd2PxRu4Pj6SWZOi33fHE
gG6gqCTGa3fe/rgJEiEqke2Abxsjd7Q2LZiH006O2DBr9jmSlvRispMA6Qg+CWDb
q+83df3P8e2c14de0inINJs5472sLHUNG3b3dPna7NbltsVzB7p9gO5etCGXQPLm
0ko8q24NJfHMwBwe8FSRCip5SU8BPvOZFTIWaayei33fXGElfrRWu/4BGtuk4okf
KYDr3/1Oo2AEvBtKJCF2e9+EYPs5Gn/Rj1mASluW1Dh3HXvQhM4L0ewxa55l0HGJ
INouweXd0p6LiKyAQ6GJ74Hx1srw7J7HHg46EOZ1j8Azs/Sjgb9+I9cYfQepCdeI
utrTSLHpHav0eh3zqSwF/Gba8VLKdC0bFnfvn86Q5FsSvaDE4oipaR0GuUv1B+Ol
s6/qJIboTeHgtHPjp/KCip9uuCxyPb5r/42TLjj3fvVne1w0zwagXK8WUhGkKMni
P6i2SpwqcXPWMuE6LyUvomWcW2lM3/4k3KCnF8CZWhggHcQH8/3YaP2tkKngL+4X
QH1B8Y3e6+6l5VjO13qcpjl90aGSo+y6D3dsxJoCrnbwMco8wEKSJcaxfWLh3AQW
DQvaaVUs8AGd9W//LctF1MWDVUYa7IVS4bDdsaGU5WFEnDV4EKsWzfgUkEEEg4tO
pajiH6SRqgLVYY0ZMBU0f598jgB2LYLPD2xm51rKnJgP9igVirY6vxwHOAizp/cO
mH4qQzTGRR+TyEr2xEFCLPgK38YPVbGDGvfJ+DAgl8S59qIulYdHHDhk8CoSTyug
dix53thVIahZJlI7w1W8IPVMkGb7YYKq+U0ooqKSVT8jvs0tIMs7w/hzAlH7zOaj
/jhSb3Ipf4bHf7JIPwEcdeuFx9XAQqz6zeaDL2ohmp4SnyW8XDcNpzevOpbyWcdD
rH7Urn32hWglIq5RAxvp6uUHOeqt/u1da7v6IihA36j85mPWQHel+tx+ELYXjLBp
2BIVJR1YjHJmjbcARLWCg1CMtBgLE8/8MBl1K4yk6Bqwi0bm+HfzpPGK2z6OkX9t
DLBAbx8A8wyBMXWq0ad+7CZ51vVacAWdqorBERYbRx+CeoxjQCJDoJd87Cgok8l0
aJYFkYVy7ez7C8d3HD8iBR7uLIXGprKlEYyQaGoGGg0/2ztAb340d1WAEMDpwPxV
MfOdqMR2W35Yxs7Z7hwVvGsBKfahIRQVrKUDj0dt6xxhG2oKg6kel7exUYjDa+4C
H8wWFhkjse7xKmGMaW9BL53hcfYQluk/LNw932Xg1Ssh23qePyazBNoYwh9NO5o9
Ok9lDYO2TSt4g3qyxHGJ7vDY4YwH9nz/QYLkh3OWvZ6YZr0hSxBzPcy0bBtKyVb1
Es/DgC6fnj4TNmen1NfsmhMZqfLeB30fIdrqmjndaVda0nuFuggZHwgo7EH24lAe
Q0/d6Ehi4ZMHFcJ6OXA52wzpP3DQNuOQeTTl1cEUzopK81J0/htou+OFaWUGUoTI
VhSXAxk6CRgr8aJOEXgCnhR7l7WsxY968l06VG/QxUwj/nJIT3RnOtCo0ynzbVNi
SlhckcgEn6QzE5N+taMtZt8arycSpvlrSCH28Jedur0BNmfytbeUc9iBAjlCUTbv
1OJ3xkkjYY4R+uTP76EwSS+Sl3CKzYhAj6w8lfGCEtkvzNqh7spkN3t9bhuR5Jfo
R+V8lwLIZOAZPqlBlvDkPz8jRIZE+6Vk9+2Ho3FwgC3i+ib1AVyZZx/H4sN8kAPj
yhvDxrddv0DUqdcsp7qDt1vhFU4NNizUQijrHwUEUwqkfxGihTGl1XaGPyZ7SLl6
ON3Mv+3qGg8Si99ktkvN5R3IP5VmSFhZads9gErI1Dgt3K7i7gtQb29ZIZAj4F80
FT1QAhitVFRJ1itKG1voYwd/aZb7uIlVue828YVVH3m8yWjuhBX82wjZHXaQp2Vs
jwLhC0muDOIoFwSrQsy+/hAXcXLiMkryPSZZq4hg2xCwiJvZVzG46bFnf/wNYdQX
MLE1PVBXPaMwgnZqdnta0GgJ3Phj3PMpO9WkwWi0/cMJDSqNuP3uPm0ba5A1uHvJ
UQXwgkJOawAvR7ytff9FJkakp5I/nD2hO0PcM4BYjPRrJ4YkkxCBv/38PhIWYUvb
58RJbAvSUKninTQjL0VY3IVrNaEkT+5GmRyfVnjgcnqOUsEkjlFk24LHzZA27mTv
P80+xiG3XMCc+oSfFNAD3hPq4JXtszIJUv+2fG10mjBM4LSsP2enmZ2D7wNrDmBZ
y0MFBEJwNrGQUJXu04EzUSt8/Fs4su2FMBKibk6WjtuISwxnuFNlkvRts8lu02IJ
UzAGM8cHYugkCYJLB3xRnaqwUN60++IY2ZEiNHQxb43Zi4OMMlCMCB586v0UgCbl
UlYrQK6yewHrTw03bRCLcP1ougMLpVO84buA31A62FcILFwE5758TzjpmVAss5AG
yJH4zKhDsngs5KXUDrR7yMOqKPzkoLg+qVHzNMJb/Z0EXzSCsFZECbUjDg+DVabR
FGSvPmlFIHXgw7C7r4v91St+6YFzTHSrteY9eelQTlmn0z3LAoPawyDRq1T02DtZ
aAAWDpZRT69FC7Wrg6qApadsL7eO9hcN2c5vJkgxxMg4wPcXfQE4GYAMeHKZdzOB
vfLVWc5oYtgr1bh47+eNy+w3crY+tbgfl3XAzs6n7fyTSYVOJ/CeQnBTmPdzlNQv
13FVBsTnSLX0NNqwDKaDdS3GOkQe240P/M3nzRS2CNm0IgEHR9S2IwCW1GVdPaaU
KKOCJK0eFS/dtot6S+uhKWvR0qYCLAgfB3b+vASKudc7hgmKPt2KDzPdD6rYOqL6
sNyc76jHhabGRWU62y+BgJ3eyiibGGngad9Q/5qE3tpgbzJRNBFMphSL6s4FBe9O
q6dvN2LcLkZ8avi8pO3Da+6Q5vI1nxGNT93XejtUfr/om8awpYPVgajHmzBq0SKy
zArCqsPcEHGuvkMnKccMjPWm1NPIYWc+l/Okci7W+2dJ0S3uH3E3ptbUItMHR6O/
GxEIrfFy2MfDknwi5h+aID58eGfJEl/GBpJDoWqWwd1i0ZRfOZkPygSSVqoAf+Ey
gSauD7Ekd2JSSjJH7Qfbr++o9/spIKk/L2BRafR1j/nNcA2I35IPQa/KRXZ2Vd5u
FxJKJvyTsJbJwY1cFL3n/ndKaYxexyNblogFA4QFYGafJUMFxUi0zi550XpL+wTM
zwa6YuFXhVgxlnXrlwTz2tQt+sGAjbVu/zv6aw4BV7Yhzr5DA6L9plwcv/VGHf5T
7vvh5hn+g+4Un5CTgAOaQB+R85VbktbDNO1/at9I7x+gjQ5fvKX+ND8J0MsvwkbU
HKcfqYuBjROj9dgMZkapWVO/c+R2/2FFjrz2zoPK7GC5uYKIKNrBIRKUzAXp/Rl3
SkqQyEQj0MDToBp+elLzjYAEs1g/HQJite1Xohx7pu9oDTxvUau7iNd91HDkofoV
`protect end_protected