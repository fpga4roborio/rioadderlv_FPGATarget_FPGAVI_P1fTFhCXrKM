`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
ddtXksX2+yylW5zu6QL2Lhnb2d1sD00763mmSITNX595NcHTEkwn0zB1Dry37fOW
FufOhVzEJp80NC5qZ/+F0Vk7Ik02dIR0elf3clrjeJRK85K4e3Hoo4xn7YbFUIms
l/8VZSb14+JVGURjfswrIyCUotIzlzVYZ6gzoZwDXIi5gQIBf/gI+KxNXPaKV+PQ
Ufys/12rjO6aI/pPlqSm0hCvftmBcnezN2hk1UeXgOIuKZnogjOsf0iJVX2aOOWE
6pD/psybjbnsNB6kH5uFTA5frkzIzkzl5d9+YDm9OyC+k84E83I/7/j+rk4L2dah
QJOvksSIzN867/4Qt8qYTQ==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="MvBXkzurAa5VTw+1JJ70nePUfoQXBvZOku/SMmg4TwQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
oRtzZL4VJ4iwysPsC8SXYCzXS8Fw2gtZTOskLcDV+1B9Nzn1zTyNtlo6lNICRmmK
ZRVu2BmCc2G+fmzynYlNTnSa7C0Cuel6FYpxCBlOuk3OF2tzAmLAuDyOH3Z1Yjzk
a0aHuoCdIRKv7BrZCdALt03JeUmXKPdOmIlkVGFl8yw=
`protect rights_digest_method = "sha256"
`protect end_toolblock="Jn9CQpRhJt4rnzZPRk+dOpzAubz7omckX1MrFd4p81o="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 44896 )
`protect data_block
gD6l00tciPUa6pDNTk/+t0OO0nC/UTtBwLB41d4inuAUA3i/ALrNyoJVcBnAmEQW
ptbcNp5fxEUJjnOxnedyZEuEBxWRieZFQnkRdF269oNJzSvXzmnZqv6wyi06Io19
Uhp4Ed04PUc3yjLdbocnFkcEP6iyRKj0zZVIx6UHmQ8RaDZhNKIg8rh7kB8tBjIv
dVqHb5fG/lAauj8R7B1xt+LrGctf/TLJdoAGbTXy/RWiVwAy+zqm6ldr1/kWoVLx
wcJocbO8iBXStWdj3eYgFF1sgCn3o1bbL0B0Iqg3665SbTUbwl+pZs41wwfXqR1i
si9ebQ+PZSDFgNprngDM8l1LEJq9d8KEB8E9bAQ94WRiXih2rv5mXIOj3vG+Cw7e
B5yq65MKNJzaOlDA6T4jlpZiqnNyQ1m7eKlnxVc0d/uAyqRmopHleuQoHvAKr/UT
7tD4IQcG0WuNrMza+4dt/Y5w9hzHWOKIIWtgmSKneJQyKySn+3to7xqSIhKMV7Y9
wpBzr5TDdmhfuHnP9SIcEDXxDhJvsAdAKA8rsMwatiB8n28H1HHhwg0Bv3Qv6ldY
wjdEd4y0JasMUrlIneWFxu+6ZtXKAFZdgM1KSNY0cQJZjmabvLO7WYm/J6GtGEzW
Urc28bmYlsxuOOg2ZEWLoXpGEB7QW9tCSodJF1hyiJH7lPqBwQ2q7lYeJa2iV38B
QHBAliu/OeKMumZ4IPNHhC6FpjfGzu2HbutHJMpDd0cXPXnn6yX3Kzhnj+6IFuEB
FzMLPxy3aqBlrdI2LiN8rRie5pr5xuvjDORLMTjLn3KkMu7Zc10/Y/PIuzxM/7nr
+4O1LrhmlyVJpgaqzFtWVLfDm5XeDYAEgVi4ISn45R1Ext9VFevUV8W0Zl2uY1Rz
8MwQS7aqpQ+tdwxlezxzMLgI0o0odjtwNFLM2MylmjacdiR/ju+2+lNjFZrb9exr
WfVcteSGN1344ONVDEsieEGGwAIXuRn1jdzfEs81ubKhpXA4q9ZZL2jTUTOiP189
yBdsVDafnfauCF2di6VH5jw/JYGwf6HO19Kg+0olY50qG4lAXDruh6Im9u82uTH5
WSZg2Gim22WnLmEb1N7UM9adIykoQ3FKWPpT50oAvM1AsZytrc6LEAjAmWzDfGry
Vr7nn6uSTkwsZ4yokqzfm0dX94yraOjEuyuISRYGj0LHchbW1s21FiiO9PTLbO/b
NcLH1/cKx+fNQp+MiB/US+UY1ctemU4Gw35lAYDEMQFYSgQMcglqYfG57Eo33EIy
LT9Ji3Z7EpOsH1ltsGO6oAIyTKD0XDovLxHOUInrTUxHUlr7J6gTtzD44S1re0SZ
QEczniZzj+Y5dOOaQGsuna8/IG+hH8X5hqTyqCCSgf35zAvP+8MXw5tr08OXb1Y2
0yttDzDya4M0WUN9x5ZDA3sD2v64dcb5FlzIeD5ATzHKDKr/RZSCPHovC9SZWWVC
SMwPrst7kbfl3PuuxgFYYmKGjapQIraPIAJRSU60q55a7IcozSeTLkEfX6owAetw
yXOsf8M4jk22HyJy/lF82GqBaxutk4w1WkXO5aABgXBRnh2C6eiLk9TwP9ADTy2p
hmO9bnibxZfMGo5k485SI0WaxeNnUs29JIaDD978XT6Z08y4aV4AE+mz1fRc4oP+
ZY4lf2myQfXwaujLFTkEfIv9y90XIH4tkEm6WJLqIn5EoN4t5VycduTpk6ULGDKy
eZz5+Bfn5qRqpRueVPng71asOBU9QBdBf9m591jJubGODXcAgiH/SvvSOth3XBep
8Y/wEBatiBcIv8LFj256MZkIrv6f34Y2/L3I8sg6K7PPi3nEo+ANhnYDgetnepvR
GQWSlLgGPZxTCnoTplHE9a2lYZh+t6NiWWmT9W2dWRYkoGqzld+0LldwCk09+iKr
29to3lI+AR7W6DW1xZbaewMsgZAANDXAxGQiNI/E+Nx3tR7/R83N0SrNbyPFXaMW
cS5pTX4Al3u3npoDbNYdzxOI6TWN19CBH6GbIeoTh90txxD9UxX+WcUDau1u9bZo
T10FimZYTF8xpoKaMWy2xH+Oy68kXFg2Ad4VzZlVBAQUfWJMmGNE3dZvOrjw2vJE
91JNzdx9mE0ZPsHZH0h947roSJOmKOZ4sKrSdF351XHINj8MYIPDrhc2yoj5RMwx
ri+WIaQ0EoKlHLTMH6HYh6q+w/goTK13KOGEJh59mOyO2AmqvwBAYjsqewK+0lly
rrLgKEaJP/x2XYtONgNnNUffAw49bUbRV7Vvvin2+FdK3e1eTDoW6fvspRAaSxf2
EpGuX0NB+aK0IotJFYw8/0OzDl97JANFwRDjG+D1cyU1BHI+jg9HRZCFsPAy9nYm
NKlClaOwLxcZotc0bGvQh0dC3jeWLnRWJYAa66Q9osqf4pXrq4R5WBzddHa+7Cvs
MF9RMQTpDZS3+O40f18JGT9oL26RgHrwFuLa9nM7kncBznlSwGH+Nr4O1TAyHJwQ
Vo5fT9x1I3z5iP30rsscFHpJYzuMJsoN+rX33GsRsArFIY71DkmHpyS0Q6gGvh1m
u3NHJ+uCUmWGH2MEycHEwlJ7rBrLxNvomSkWKcDzMc9uZBls4ixhho1YJ+qP3bpW
hrDSZaOydyYMEpQ3CfTXbmJKkn+yH8QioezN8BflogOHyE//R1HaAyoncdh1QJ9w
tdwb23ATuqlpznQypSf13Q30os1dCX+tSX3SDP6DVtGJDo6nDgWa1c2R5wBr6gog
W7HyYRDWxLjTC4FtWVISo5DUMEPhpZ0FpNtdoNp2rs73zuk10BHta+ANV3pZy831
yiOCYDVV2a/Z7WpOzvmwzatA2BkMX+5hbbN7cNH/aBBZVaapNtjZ+MSTojNxs/aU
dkN3zZWeOEOc3JVH08rwkUvVFWzHA5dv9l3VfW2ZeRDy1QcMnf6q4rV8i6bvvDF6
Nv5nyMq9HNMYdX+MDhkw5Av/1FsSoQ9gjQTLP7HFyzoUw5+Vvl2tGhaC2786jkjC
JBUMe4cRUd3dA/cTgccvg3IvwMOVQHou4/DrIdbp4MPB5mqVfR47rWtJ5m/5L4r7
ebsFmFTNsV7U89tIry6ySyADFqXdYjGchH5TdK+SliIKYM/Rnl3VT0Sorfq57zmG
itZyTKyGgJ94vjdEsg/VtljUdW+K28paI35/iWbTfvWSFi3+H8NIwSFLKtpErXzX
J7MwAXZf57yO+44BAfVtn1ZjHJKWvgp3li14gwP2VdsUGq66GqZLLGJf/lNUJhpf
N2PIJGv6mQ0330/vXv6hF2nlOTlX3GB95vb51X8NyQ3jKsdB27GDtzQeTZmhyulo
vZByJTzqbXPitgsm/H9nlI7jWwh1kFPcRxOJNZZvOgVd0JFpEbDk7mZsGQy+BF6/
unZ21cY8iusBlv8rAwgwm89UiZDhlSKXSl5BgPFCdz7L/WqxEpZtErGooFeggMAJ
dKDmAukfqS6t1o8Nru7amXuaxxVhLL9hXyhW1qt+0C00A5KqQPVsfcUk3l4SHg+U
HdQrAhMz3wVUvKWkWTGihMqpMOXeF3tQeaICOWzD7HSzVEiAJwC1+RUPPF79iMBv
0ZjUUZUg51gcbFSeirFNhkIowFkjpyUSSWZSeHT4uSviof//5XtLVLFP18E7yEl6
dN4sQJiOfBRbX3N3G5ShAKbfmmdpAlyrXnx7rGk5JHCNA/MbWMhJNsm13befBFyF
3j/tPmSG1nQb0QJXoKhpxNKe4lVOqN+ra9qD4p6WqSfJj4+ETjlgwEPCBaogOHpf
UFQTQ3TK1qM5maXrmgpLxY9txtox75U3MXXNiIJd6ryJIhv8dshtRm7T+k5K9ogi
mZH6lvxlMLaHxQ9tzs5nsR/2DzmsMDns0y9BWuOWfP1AsawBKkzkBy3Qpf6U/g7w
NFVF+8IptdUU+XL/59Hf02D8thFKf6QdmHpA3Wt9UYhKtfG1ZEOHhakGqqsRdSOJ
I4XwX28/e1dypDYV/j6Pq7D1Cx7RoRbP+iBY06aRs8S/Kcs5D85Eg9urZfFTJNhz
fZUnRFP2hbyxpUo1k0yXvMW+PGy+Al6q/dP5De++Ycvn380nqQJyr8nnv6/C8Cqv
BdPu68+8HeLkENaelm6dGCOMJRAu2B/fWWX9WjWUbYoqU2GO2uX3Zn9y6+UdVgbR
DSl24BgzCMkWLSQ8h34XRsYJy+AYsxFYj1v6PA495U6BIQESs+9ShIi/g9QHSELO
Ss+bthhkM6jTIwP8WoB4m1bQs5+Uirsh8GyaxS7lqdfnCYa07knujjU5dENTZwsY
EV176b7XR4cPEutBRAzENzJxVdFDBpeZg6oPoW4sc3M/fTiY2XT6erWkDs3rEc2R
vuy1htP2UgZPgAM/fR/mcgq/jUlqS3w1b9wkJqbm+O0YEqJXJOQOTCMuUBGHplkI
7y9+OwcFyv2y+ZGXe74JHMm9s0xQma/JJvVCIKBfLKU734KRdoJhqdLT/Xh1caDy
ipnlaEYF+iOmAIBpjV10CPurq5K+ye7Rem5Z0NexhYRaCfgvgC0W3QtpSm5PGaXH
XGnuTyn+K2Pmlca5+gui/W9UC0JQtxDAJNrQheS2VUWeNewtZTYl0paq05CKsfcs
1p9RHVzqC+FD/wJAYns0NDWgBtQ2Q5poi8uEOKvF1XXwtgWe8nIR5g6EX5GBPbga
TCNJ/BYGMjaqCQ8tzPLjYPOSIIETV8C63Eg+HQS0D3yRDww7RI3nfUxNKWubWt7w
sPDt5fhZ6DhMoIFJiS4evpypA3E7q7k560M2h0rd1g/UFQzeKTLaxzYEYEZGAQk9
pXAEwLKI1WdA3DPNoUcbNsvMFzROwLlQ/A6p0vSOmklB6gvm++VtMztaiyBzSEcB
amc0SSwxDitG8i+YGMpkQXi0zusWm8I8JpQm2vmFPiAFRlNxIf52CgH5oEPtZc2J
RiTOAXN8vSwjEYOVP1a2uV53LIoUhXO/JQ3/uxlRGGt2yEIi9+XwuMEi4fJ2IA6F
cVo3wVB5WiZd/NGf7xOLOfhxY/Xob7jlqXMlB65U5Re1m7uXba75+19jFccOjL20
OS5lNim4292E1t0BeznxgwHR3vvEdHfmNxGbCYkJt7hPdj5B7OsSz06SsKK+7Klj
ng8gUOuDjLLnkXDoa7kgGnRGp0pSBTSkIr1KA/D1QGFp3A2olENm0aPhssSJlmh4
5hq6LozfpAvbh3t12vTtoRErtQ9kjmREaURHND7BnWBphTaZ3m6PWUUIliHb9uXI
NFGEqOkTmh4ipT5OLlnAfVwtYx/Aw6rf8tp693POSlxpUjvEovIb4zYtrFrB4Xo1
vUpZ7/AChYtysybcF0jfOf2q8af0r1VJinQHpWh+vkNEBoFbgxHahnpVbFDyPx1a
eK70Gd7I1zpTWXUbEIJZQ5xN2O5n4/kset3pBcVrAzBTilzwkcj61Sl4GKcqEeZE
u6wvm9A8eifdwPC7u9BnlYd03bXMJgfP7Jh2zrwwcnzYEoI2LOiuGKF7LctZQgL2
O9ezUpc90N2mttuER2OT9JWXs13N/OjQYyO+H1sUR3o6tCYl9QPZXZVm38YmCc6j
oyRepV3JBJ765W/HIypkCz/gKM76ZFO5MW0j1dhO3o5xx8oAAZ1Zz6WKZjZjIiiA
M55ckyXlBT6405D2g5NL4yBrKcsBmhZWfCpubw4P2jH/QbOFIhtjdJKwecIYtqj0
VGhdrGTNH9VRRcRocBPckZzbKqWACLf6xvJWba6pbCHNc4WwPVHnbirOYD+Uf/Aw
GTIFPUf840Z8cENhqIwumld3qSI7ePN0m/OG/HgmPxVW8FV8cqN/vvFs+BE6mSE3
I4vBmCrNqB9djLR290dwoODhX7u5FyU+kHbXP6Bspfmlr/PRnHPUZYFGWtLscEiO
HTIEV4QyiqN4B/x1aZOL5tayABlFxIebPnARkjYAyQ8Ctt3BiVwmV0b8ZCge00o2
Uz9e21hJKScPDkklNdXLRrvRwhjxODlu/CQHsL4rpkdFaExWjcuKtnCQv/+oIfEb
vdJbS7ZzgxfG4CvoCro0wLX3AF88q3isUtm/lO6lglNAG3figQpQWClD0KIzSGl8
n2rexBfsq6gBTqBH5E49c8jDehT34om6OmOAc4OPMqJaJqMF2WhlD9H4fWZByLnP
OqFukDJ3Z7wvaJ08deC6DUWlCfuO/vAdlyVbYLnZdTBelZyX9nTX/TbTLjWhDv4j
4Cthkc/c+EoIraZ1XUgt+OktTN10Qc5JT5fdLRDgZbb7G23p+C8azbOL79ye2l77
6bGR9QbOWphksAEf0o0D8pit5HjXkReVoRGgInyOZWMBOBUzAViPRi62TxfRWjBM
VXB+6FVF9EWYNiz/SzOAXL14G7BNGn7H0HYzn9lY0ycYhB187Gyt8ZjcykaBY/as
JxTOF2YaMFBIxuGFZXiE5DeHwYif9geFCLF+KNanzR/M0+b++Gv/o9e0vYrnWYtz
xEcfcg4i8QuLYDy6raJZb7cT3S2OHymfD6hm3JQroViz9fudB9GIhsPzlseOHkXt
VlOlfrqsXU2kyHwXpVYPaQNZM10+gdDdkB2+/aTjZXYz/fPjNj51MH0v1PEXc3ZV
flJf7rObRO3dcX6V+h4LLtFRakjjHtaLTVC4EL2WwFtZsoCMbNcESCNINBerEvk4
s4+a2Zhyy9zpBkgUcl6uNqciqj6z04gcFIsDPHEZBBn8wXEq0TZVi5jfHD/q5HPV
r7FBIVovBHnxN30b7vNuSUe/rZxR7NGAaQpOU3sU1C2MuB1cjppZ96paa6GzbGM1
cF+KA6zeOKeNpF6xKSD3RNTObK+53/x+vHZ/4TsEUUmLsE1sob9hBM37thkXNFh9
WO80WcH1OQM6EhKRTC3FZ7b1ZD77nI65F4hGvOo9X04SSi+xAdeelcU/gW00HDH0
T98xUZo8uEAOE9BT+pSprjL2IrXQK8MetNQbsAb+x586I3TcV/vGQHcL7l73tzrc
S90CgfsTaAdozPNamYUluSyo7p/mbJWvMvzg60aRHNSXBV9s19aoo3Njhmz3mM3S
Y7ntFPJKf0j2jbcVf1UC8NzjcHEb+ODuIcWKcK6g1WbajK4kqbK9VMVf3bK0ypcK
3kgLV9C1iJhyus/M3sBZfhTuDoywUyaQjmdnrhVgbrtAuFkFZxQF/1VeTLTCvEdW
gTG6J4rjTRlHNYIOavLJ6O/5xoGWQx/mnR358HTaXXHfbR4IwKfW8cpq89yhoDll
GEztua7YsHeWtbcdLKRDFNIUxBOTWbi/+rf8ljof7NDQbWCAfyrG6QIF4GKWLlb1
13UkVhfB46MizzersXOAVt36KNU+HvA6yoz1ovw2NfjNIUWjxL+adhQRZW+rZF+b
BuTHYhrX5BB2YAmzkgDGoEucGcsaym7AZAEqYmVcHGPm1VRWAWZqK07bslIjhrEF
lihRFJSDZOPDkfE/J+GnTEL+z/THfhc/eCjJyaMjHRaRcy/CcC5can+jRL938OXU
KDTzHuxtVtFa24WVj+e0W4l/T1KDD7MAPkIF+B9r1kDftU5iPaqlJXt2q1l4DHKX
/xSl4HVBRECd9z6rR11r5jWUGSp890cKGEWUHINCr8tdIdX64+CfteJ/f1Cquvuh
GM6HTHpfqdI49ChF0PJAClkLcEjMTlnBuaPUREb6QYRNCp34bkG70MrEf2SVRAsI
Sq0ucc9My7eoK0s6YIhGDBt9oxgh+Jvc3WizKngf6gjLQSficFyzGWblNnnDmlIn
1hbmFd6WxCx50DE3okJTqsbspBfE2B/+KUSv6kR/4pbReex8+XmR0RhA5Drh1GgT
JmxKIPLABXe2RR6g+TVOyCUfz5A408fHXsa71a/doQPAhBAhYQjZDobGnh3YGHeA
CZHiGF+lKqZiPsr1YnPGGqlHUtGfbB1mqDUwM7EPRX2KdvcPfPHwF5QtfoX5QCcs
9LSV3P2iqjI8ocwDZk+CGUqi39p1Q3R+Y9PNkkK50bkUkqulogaRE7xCLRl9VvYO
+2KDPCYNUB5N+1irXcbB6Eu2iYyPeN/jBRpu9AyZZVoxUSrW0Lw7KFPe6FCF79bO
rIkWrnUggFj8BjthkI3CwAp100axjASRLIXpw8TDEZVXuhSxXal7A6UVwbQ9tvos
TSKzpzwADUuEsLjf6rOL6CTG7x0xUwEHVL1jZHPlFKpjlthxriwNgTLriitiFImm
eh/TLadM+SC4WDZrssftGQj+4OMlXs3Y7X2LVmp8IRzHxEXY3Uw++Sv60KUf4mGA
GhTsV32b/66sPrd8Xhq36JrqVNUaTiJ8Q5RpYTIY1Dt8mBvttKmH0GMc9+J9nTCC
5BOvSYE8IuhJ4dQ8ThEjvSQcZy8H6ysh1fhSeUupw6m3CUavtlseXo9G+YpLYJlp
x/JJiPUHhy9rlb2tcZBmMqQrVSu010h9y8aG1PjLqkwb9jyLs4laLtTtDYwTmeit
h2OYrXfVWZEhcXXwmHQtfEK4w4O5xxVuu2hv1e4MyHV9Bj/81Zl0JvqXLwImiPwT
Tl6sePhdMMW5MwIuHOkW5j6bEkhsMKf5bY2OQQc7VF/ddD8VwWDShsWD+FAnIuKw
VAqFeX8ssjWORzdkmDDWxUj2flI/FWrgFzQ69KHV6j3MNJ1gYF10T3i1pOuFohma
KfuN2comly3dgzQDGCPqR5FNPY6x0XQbyPi9mJsf3FvJ7LuhSHk1e0V4qxVhZT1k
8eVsXt8PXOs5T/nxihCXtJ5EbEgCdMWD14csxsZTx0p8uo1YWfZSR9KochaNfZ6a
dVLoLA3SfPbLWx/1RbSwey7vhxscZyirwWgC9SKIswzy9rlI/nOUyI8uMkudi/b+
/Elws8qolP4bgyVdYHOTjWnoaZBn27xLc985gBodJ/xIDnWdzh786lVvULmOnfBf
9l4qj/U+XKJxTFyL97+UPotLKFdj22xwCaWt2s2plTEqcWCqXJuSYWvA2UcGg+i1
8Q6JpqlGcYs030Mc5JOL9tkTp4a+5gWw1STBIOdmaB8l+LMA7PmKBxt0rTMmaK9u
rLQG6GiNxATj3TSWDbqDJSukNi2mjy+o65SvOcltGOj4Xs1OtqTCeqRVQCCvqcZG
u5NhRIPLy6atbf9GltcX4uwhXXQcWNHE14+anzpJhLyPah0hhsXdhtah4MQ8s6Fj
GFWCwABgdyZ6tmwclvnRublk1GOZE+6g0B46vGnmzRs7OUt9R7wC9+qgJ3umtKiV
IUkvTQ1fxtMsGLvyxPolTxETJwEhWg+Jdsr39Kd4B4p8vP0x11YlhL5tFHuE1hip
ZqtvncqZssQa2Jqpz5hDtKH2SfNQPwJillep2oBn06rpV034APevN+wadG7xcdMB
ODcwn9t7KsjNLxT8zx3G2Qp5mMBCRpKV4YVydFNSwskey2a7k7h1CE2+bVq9Xt0Q
m/VoBEMVRV2nR0O6K09HhgCCN5qSjruZXzluKpVLzF8kYetFxCtHVg3cbUoW80BW
R2+32rqLOyV0xL3Lz99upmJfyGNMRqyV5CEXOmjmlimOq8AkzVJdNtwnmt06OBEa
3JDIeG4nrI+ieOkJhJ88ByPQ7lP1o23aadpzNREKIDO567kQ79VZotanbLY1e97h
i15y1oiSvW894GwwO6QY+qXWK6+hU1GYMTiTVAOff/L6MM6XYxOgFuOebacs7tut
9zsZeL758+SYyjtwj0zwWJSxWxaCFA454/jMq/JHKFHMdoNECcxTzuDAlLb9mJs6
fA9De3IMLQBAE2wpQaTtvx52hXxzld0xMVSKzTW9MNSMm0PLegxUcBZuLKhpAe3x
BnuYEshkShnfEphuyiTwjxYuNqCj7wXyD8KlwiWwT10k4IfQxIoHH7H+UCcvO0YQ
u5VtaYMU6MY+WRjgWwj7Cm2fbqVG4/ir/150fb1I0ccWhHb1/vNhHkDhF7U7dbyA
KC4KWdXAqWANAxZJ/YR4+aV7Mf3ZYFxV/Ywio05FMWEPgUi0DunVXlO8hpnBJEaj
DW9nOVsuRIcbaSlnVeq4RhqabE/Kwz66sdtzufvrScwuK/nrpUo1knGQbkQlmhTB
GECPSn+tzBPwjKWgP3hFX1Hzt+CsBwdly9PQ7OJ7KvibRCY9qEiPCg3s11RQ1svy
FMGzSOwqM3vGd8ahvn6whvtG0EKe/a4UGvELtdFWnTA79BtDzrSDyPPT3/MARSdH
hzji1UAgG9s0hAcp0TtW4EbbBqaZ1Glvn+HjEDw3ePmCI4kQn91yWl1UibydwwY8
dLIgglTkqFkPL5/BfWBF/MqEU05wy5Y+6obiYV9fiKszauTHjnI7F5xmzFzd6Ypm
Vdc0ZVcuFhg5Umfg7TCXIO1sIKrVTmchkjEKfjd5VpA7eJIPKPt1+EenS660fkZp
udDDifC4CMFkcI2cPlNxZu1DkHE9g502KkpdUL771eQyOVOex73VqBTwuxXwA17k
hkvd3RSyAvZ3X+FyI8uQgefMpZswEutK4UYGhYcwkLuWmZ/i3y5JTYWmn1LMUPr6
3oO4kHzMbaslCg2DbESPhxhlWjlpyUxWELcQoFkR9B7XpuPJWLHFNnXKNCpq1yl7
oQUcyZhlP8c5BlTKjmOpEz+F1PgCqRqOdS0qb7B5ErwuBcH4f9ixosa9MM057FVm
obnj5XzMABmhcmhkypwk+5c5IfFeke0pzDZRMoiDSfFNFClHFI6MuUkpt8VhbSYs
ZSN7/VyBLvwIj+o3VKvN1E86YzgE87Dds2L5kUSw3bt1VUTHbgfp9W9CLfAQ7mtr
8SAUxzlzqqXedDX/uX78K6iZ2MnMedXyIg6bcGYn8joAMecO6uLnTqoZkCq5pzUJ
ucnoW/WCVmXe3R03GqZAKz7EZiMdLfuJPtxvPIAqljnmJfN7kAVi4v4pzgfD1Hqw
Ca8yYKUn0XHwwhtmIbxTjCGDM5zENQV1nretPOme74pjfytUoDD3llTYvbaZeGTv
9yKIN2GOa8Qq+OVTCkPqp/lKucsbpOtTQgY1YOClayQHTWKE+Vg78Bz54k5ZzMGG
JY/vcUgYLVN1wIcFEQkBQ1KUdbWuHMLlsBOeRClcT1Z14/eTQsTtesskephRnLLU
uqj4eHJO9KtAdoKE8HKQ5lRt6iabao+JgqSvnweHvfpERCkAuHWjOWibzLKxgDBc
LDU4RO52CL2KHYbAHaCgacbjTRG9LdWbFa35qhuQ1Uwoa5527A6+Nt5XSah/SdxT
ffa2cYv6xwbnK172h8e1zjHrVxi83Jp0Mb5A1zCHuoaymLbxIHe+TCjt8Jb6mEqG
pipn3MHJWmZvMiEhJt29gpLGWs6uOVYVz3j+j7kjaqqqJJeUUke7H/JQUhaumXLp
Z58Lx3XHbjC/8TlPI52JW7kpqysMmD5W4DGYuxqN0vFoaEqV64QX7BwMcr1GIs75
oUiGcHgFQNKRZCy2d5yVC0+RjJFtfepdOOyl6JfgMXjQGNqoQHMbZ3I6NXuzASjW
7jIcoGNIvxNCXD7gE9ndnZGBy9yY1npcUSDOrr87bVe/p4qMyXRsOG7/IBiKHkRF
E7bHAMQEGB+PXVZdt3iEY/chB2iTClULwyOkaJXIDUbXAeWJvul4Q4qUUoLWmfzI
1DzdmPf5VwjVYkWUS8rZ9WjSaQLNdXBldKpQW5aQ3kqVFehZkRVEz++GYahf3E0i
72IaJ0QS1jIjyyahNUuBC77nIAz5aZegwpTtSyyjqdD9UesaMs2CGVLB7YYycdyK
/WjswdFKqzBjHWcLwseMaPlTjhDNbHK9FXevcCF7U9agSHw6s5imFqCVFzgJtIOB
11PaPquebqQbAl+kiNZNPyMnyyQVC6dVioJbhAmqOLo/4ae80Za6FObfqp9lNvJA
t35uzF+PlGZIdGgi8FShqiNQg8Wppqb5YvJDwwResHP/hQml8CEqkgj7jjZWezv3
ewJ6MFFWkjOCUc9e26BSxfdGvG19Kd+K4sBsxCYBA/n9sajzF57BBTtWpakME0yx
zCfMPF7K6EAQ0dFyqK8Yp5OGv7UXPFpGfwk7ZtTAZ4A0yMg3PBb/Zxut99DsjYQx
eCiBcj4NbiXOxzdkkODyGN12M9nTBVAl7QUXyijOm7F1ehuwfHwd0LbGlPBO57Ox
JNPQOby2G+8pE7/1Dx/EO7FRW+wGJqRFl+C4G2VPxL9A1YY+LJubyVyMwza5s63K
aw3UKwBCegPKUHA6L9rH2xspzHBKnQkWIl7z9V52QTIpczOPJ7r78iC5MSRqzD4D
A0H13TZiHBqwangrVcFWncj595HPgm5H2VrdG6i2zJ0myJnWE6LNS8cLKCU3Gi/X
B2alrHJo8wBp7ooisT5ukpqSG070y2cUDPyLwCYf5zVNeYdQeewNJnjPxce8RR8C
SPaBEKvcKaVKeOduUvOjpCtHhhqE7oRy2J19QzfFPWKxmTS8ar8VqP0c/G3QeMDj
QuHDSpnGv+AuWuVgYwlyW4GUxz3lQetKQnfQLl5p5kK7SFyfAHQ+C8IsjTsqXa7z
iU246wx0wyLZ/GYmpSanVN+WlbIdk6l4u71qY6+ut9ogzVYMwdH6oRTk2MLXI/MI
xZ25hYtLmM9z8iLDFT3v4biMFCA6NIQe4sSCCPEo3XlrgrO+MRT6p9DhiF45rfq1
7rnWDPxzvLB0oltGtMnlMFe3wWBr5uWsC6uRruvJEenYRcH56JJqy3EQXeDDDjn2
USOafQzK17KoJpbPR2NvjGaWG9t85SR6FP0fHPp8ib+NTnflZDwroHMVhz6XWnmr
9U+L8nm+JNVKYwoJFqgDC32dPlTYcKudryA1gXWcClSou+8zKVmov9JSEmjJ3Nnx
qqQvxmaTlVUFmtatwCPPfUYuN0xq2h8I5kPXRgpyIlGTHmxaxDGAsvKob74IlEEc
8RI/hqQXbllBnIcHPJyjEML1o+aEMkoJlVvmTl+CrX786EbtiIV7R8l+TAhFfakV
4O9WIZTpg+mNYhn5XAGaHqHwHoYvnAbHgr2oMBqwmBHkcF6eByGy4kBz4LSqbKxG
j1ygrAGScKwbL3CMR2T8zPsiZVbawu3EFuIC0oTchTHeT4Y2FJyC/H4EN5vsVPlQ
FGcJemwMpuhYN9vOE37Am4ZgN1nNyAOX/QRhYJKXJnnypAPbCFpgecC5GnNDdrSP
sw60Hk2lu4GPAq7RKA9xjCEjhQI56y7jsq6MevK+yng7YbXDvSEAkkBY4GNGwOs7
xktzPKulu5DUIxrTx36N1xxuCupP46/5MIYmcl2lHFRtsdIRmaB2PaspLIHFjpB+
+XsBGn/k64Vog9PRhRMsPUqj6fNVIaMksQsJ2UR2jVeJ7GNuWwegfUwPkv0IlzIE
/ZjSAxqlBEV7qggS6PkyVV4pQluVIlpx8AIZdmrtlgPAp6XP+ipOB9Jg3TS6FnH4
aZD0uKzNrFBG3InDmaX+hNNMIe+sZQcmLRlKNoapiCbKL55AhiTmh4PplUMoV0MR
SvVCqwb2pIkhSoJdm6YZmfjLggUjsZteMMrGJElZUqSYU7amQVaDYn3IW4kq4nBt
YFCzk08XLoeE/LPqWL0IiwTIxyQPyroTB0IcR7YzQ4PGKR+XLlYAN03hl8r8y3Pb
pm3HSru7+rYvs3eEyhzyQOIMPoFVAAONaCbpFhcnj/SQnz3wAECWtJX5MXjvWZ+p
w4M0J0mT/WJRNDyc2y2VjRm/+EKd5MMo1I0QKbKafrmoXrqyLO8M+8WQ/pZIbaKs
fh7LeX+HY7e3knH9jM/AZxk5mDG8wUlmNLkqzDtfggv4ucbg+3eYoAgi+xcNpvED
qBRldwk8NUZcrxPIaAz+VPW/WvndwJR5QOE6zhvfLSVPa5sK1Gqewc74SxqXrXeX
b4TaworpR6tPcFGjuG9tMP4WNxk4wrhcmxTdPlviugxEMRpb2u+x+6hdY5aqgkov
HTsvnYSEjvetQoHXGDdg/XeIrz8cPOHp3SpuVDVWFQVvai1IwU8b3aX4EMsM9PL/
qZsku5ZM1YGqKeahyNyCCQxUdJwN4TTDZKME2sd4WarGTuqf2VEzaGu0Ae1SJL0I
oxnvJHrW9R2qU245lYIB3smjEADxZeVS91yNgRCMJgIww2TCS59rgoF0h7t98UfG
7oGmsG2QISxvG6Ro0mTuAJ7x52OnvitPHPW5OFzn8Q6/shx6Kqws3mco1HEZZ8cc
5bn2/GgPDUgAbJTRFjJEd/Pq6QlJYOYV1uIq5yh0zsh7h39FVMq+YbshfflMbdjk
CBGQ/2fvAD61tOAr3I9eC6olOxMPIGHwV8WBKKbO5UZh3DemZMYhsPDqi0Utulr9
OaswPIOOrhcVfBIKHW0rK1EPEPnbjX8xlejD5aT96P3pFWi2a01HqeeTYn6LyJFT
Y9tiMF2X7Ezi2LLetUNKW1/IKC25ToIDvDvocfdG2KehbzBtDFwQ3GiXzkvqF6tR
Lci5rgWkUbyZuE0CYStXkPpoUP7Ri1FwEouospAUhIF/qqEzi6y/O1yYOJALTVrk
Ndn+IBgefnFS4pJ8ZiHSvsq4ROCsa257jaD92BfJX9FzOv0uDPTH4iUpyYZUhFrW
WrAae0Q1+Wc0cwGd/EHI4ZM1PtHh9NoGnGaZ3GccpjGE3xve2kvuvibKXg1tTc+E
xgPCpWTlC1mnzpreIJ+7bxaH2mOP3/d1pq/QI0l+hm6eUAfAmMrlfWU/Kp/1kckO
OeiWGHdtk3ipab7aH10pbBoao4ULa90+i1B+sMZTeFs3MFHU0oydkwwfxEze74Oq
jNzj0F5Sdr0WtjvEssuKudjOlW2c9cLzuDfRDz7PYH6WhD08IdGZ6A9avTWFyIJy
/BjWpPKol8R3tQwa5gKX73YvHmzN12VLSEtAp9jE97CGycj5iUFro5QZbOiqxz2a
5EEdprggAOnCr4iX50DE3Ise/YBRqLDCDDy9/qY+pNEi64QnZJtPI1YbfUa9lRmL
0xIYwP/dFLQLVBvvvNIpjuobkCNw64EEZO6v/7TeC+p5GMlTIYIp4/v5BDkaIxPd
bPummObwKJ4KPiusKyp8FK3R/pSNpFZvVTAQPEjDdal8vTshHNFD2QrRNh7rL8aE
/r+8D8KlLN6GADttEh+05n4JE6SMJLbczZnf55rnAQUYIBjWki3rYyu5pyXLWbJ4
nfPLXWBI3Nm2D3lCo/FlOZ7zEvohoqCn8W7FUTuPn3UpLE/TIhLtrh354XYdQPkj
0atDtMrvxwv1zRi7s1+DuGKXyIaCaV4y1yKxuOAfYfdtKUIbGGCuqufVTdsfxXHS
javc5iGV5eTZ9qnspPDWSoMMk4TQn+bQNuDme7zHGNoyja1MeXnwV7naphErlObc
Or2wi5PqyzQfh17XwC2Ax0KmR30/krvesqg20StaVwxS5D4NotO7fVj4QdtmckqW
LEqquQWLE0ghhPkuXEmjfuJzdj69lWW3kam9XmsVRQ1tJMhVXiBrKnCjgdz9ZJII
fhUDr0kbxm9/PPEapc1hLs6L8iE07NchU4hsCYEcynfaeA6iTaAjSSxyxFWq1zqg
4tLzOeSlCx/qexsljjpYapmsskzmyZY+qhPilMfizrkcgYL4PrJFoSVfR9UeYWlI
6FAFYW/AWQWiyX89UFPtq702U1ccqqvnSxigaTi6HRNW4ZuEFK3Be6uysKUUqYYJ
3yyXWISn6N+1jWw+KO44CNgW2oxSf5mNL0vONs3+i5dCYPhfUsleB9TfdbyrZQ+P
23O6R7kCXAkCJDJFmglCT8i5krq88P51/73vbRTG21TodEHFyOugO8oc+Qu9RVKl
UotQhKCu3uB4LhfJg1oHnE5ZRtYTmW4/EKQaul6sORv1L7rCKojX3P/4rCM6K0u8
SM9u0xAkpLaJ8YTewulc/GbwDcKEjujDPBmJhMdqle4+Y5o9hgyIi44sgVeVfENk
cyRodmDv24+x/bZJBVuqQv/GJE+NSCn+lwG6mlaW1Q+jj6EE/cAX7P2EK5cSc+ZJ
oq7oqDd2t2vUrywpjtq27jGz0dHBn3mhYvYlDd97NE0CHCVIrxv5iOSFS5xQD71l
AZ7TOfPacIvBdRQjaIOe9BQ9UXUsbu4QcgU04h5kBJrkvQa52uptTJrVfP/nYejM
Da0lxcgDVzpQASV5VDlR4DUz1eje9Hy8UPXanGUNevC25x5zkalr6hGao2eY4zuy
bXtaYaZlBgofp6CbWjU8v0boPu+tB0vR64iIryncSi9jlK/p16hW+CwYAKXeC9aD
cyx6QZrdb4331t5hnaVfwyqzgKJzSWfh9KzTP43iCKhDiXNCI382rW9gRxcLG4kG
58btkWYGlDsOkFr/8OyfX59QlnWi58jjUkBUpg3LIgGyhraloNkOfDhCbQvi09wh
ha9WQfmIY43BBylj1qNKBFj1DLJ/LaaSHDGKnIaSPV1M7jfFxq/+glpKm3HT5uWi
692yHfKiMAjBlTi0wzAJUtIsEuVfrn8Jzu/J1Kx44pOJo40pQmNXDhLqZWrc+w+B
ZeYcWS3jR6zTZaTTEuA8Ea+qswRoTzFi9Uf8qpSvMlXi35xJnxrGSNKAhEmO5ZFq
yW8PFMx1hL+UeMIQXqGEi20sKvRe4BJ6nd+/V9rdHczymPxSOJilC85R1MxsZj9E
Kr8m0tdOLO6+yN03WYGrkm2+ofFkskPT58Ek02ExRsA3g7OMUBHz7/n63EnJHgNz
iKyhtl0fmUoim3BP+AYUvoTFNnUaoT6iD6+cC5qDDfm4fqJPFe6hYwtfnSnRaedP
fg6gno/grYQMqlGs1gQBxx0o5u7b+0PshWlTf0fnkcKFC5nv4yHZ0z8OyzunAs61
GkD+Spkrgrn63Lih5HvpoEY+V9RygtfZcTCLijKaDtwu2izzj7PmcwTeWsseE82q
hPCkIarcpvajQo0JVegFLyWUYLNooIEKFB+99m2NOTwVwtQASTcoq9zguDPWnkbi
SBjKuc3HZ1LP80n8UOR9hspr0IDl2iRPI7LQFk5Jx2/AFGkocOAf1hcE4vhqS5bU
GPzr3GVKZL8QQ3OA7RJgHPKMOoIyNK+XwSMkQSYYJPNdG8n/G6h74LNiYPSwdzKI
qUbf0I3xmrEJAtCckZcXqvb7PXXyGxonXD0cEUMxLIv7dwgBpu2ZXtpWRMrF3RT5
iCU1Snpfv0mew2eZLiHfJSvo1V/pMUq599j781rAw9Tuc9VD7GsDDC1H4/uMvpie
IUQNu4TqkvbYIlus+A4Hf3OF9xiR8KlRLCVbLqYImoKgoXP2KrwW0o/ENGTgXDSv
OZqOm+Wtsiq5FOyp7nIN0yZpKLYdDac7uBIzcFLuHVJG5IdGsC6ed+9ljSyCy/rU
YVIine39iLVsZ7Vkn8r0tDEe2wOloFXHmugjy8O/FoW3prua43j1X0yszB+07PrQ
9UBAKiYoE/bjrAWJG3JsP57P6d3MPtPvJXg4910DIUWHFpw4VigMoz8dZG7gXc+M
llwf3/AZQ1PUt6+geFZEfTAAL8lEUP4aDo8WqkTpa7SDm0JtYyXkLkEpaAzabHFe
LIFtObFaprAKDkegnLzxbZHHCwf+6e/kLkTCg0G/oVtpuDUGeKP0YGWOcKxCw2FJ
Bsxf1vlbhP92SiIrpQLDdBLIQr/8YwBQcqysrt0iudPnLfec3BLMQcNLczuUt+hQ
z1GUl1b5CHZgXzqIyUc2CyvSiwAwUcEb2CTVXEYfkczY93ViY2++8J/o7Xyvit9z
EV+YC9Pk4pq0lARi7JpjZk+yj/My/QyFkkwfPjfM/nmuuvZxJqB5R/gr+ZRz/kZf
JCLken46tQONKEvVQTxzgyu7rsCe7VqU1T6aSLtritjE7F4Hud+bjOvs7aYELCr2
os21Fi2gY2PFvtgxUNYh9PlzWP+W7CydZsYo5zqmY6HDVVVyIwo9qAkHWj2+SLDX
9QoKFXeH1lboM8D1RhZRHmK9VLWbHAzy4vjiiY6mB9YLZY71WkHsWUdz5Zf7c7wy
KUfxjCU3iWwj1AXQ+gW5I0uzdJsI2L///CCqvla5ZGJDpv5lNs3Y5zcKK3tXpDEi
OCH1MbgJlmRF95zfplF/fU+ckS+kGqE3SB8X/oHJcNtqlhDcdK3OxIXZ1+d+z0N7
IJHjYuE9/1dcSvunGbeSWuw2klibVYIhCSxQXyfM8Nn2I6H32yBnk+cMUq4MaXvq
edrdWf/IM7WKbOBHKw4ZNBd59qc9RkkJk1lmllT6v7adhNY96O9rvJB+FyvIINBe
EuhGcJ57QB8E7qiFLqyaK9e+ktpHumolrau5TK6lDmVj2iR0YJWDVKW3L2ACKl/K
vCD5yEW13pvuLp5DKrM1kTP8dkVEGPoWr+wvhVx7snDUDbKAm6Y3lay/ZAMD/FLP
PJB9dKhHe3JjFPcORxNn1R3dU/SLDbvT5WeIDNyFmmz6H1rXmyOgrrgAy3GD0SCy
ZVLNEVQ3S8j4rZOuTztxAiogiKbtFaJY+693g5eBkHAe2HSEvi1siw/TsUI0tPfA
j6ucouiyMi3JmRyIVfj0sgg7sDajjoQG0qqlmyDExccLlGxPQzHmHyVESHRL84HC
Cv0dHzLrRKo09mY7pFNCLGLasjz+oQFVqM6FGjrOd6bABU8wiRYTE8sxojd5eRd5
5BNUZ7ZJ8e5XQynQsRUHIjUnrMOfj2Cu/UCLQQDu0YTtHRJTbFVxv7qLMQZuOGe3
LcAGBpVp3hJosoxd/YwGmdEXmEPLhbkxmLVv1EZS2Xj5oKCs+/wfyQ3cvqU3hhMl
dau04QhMY+wHUDaLMXI/qgVH4/95RU5OM2o2/nYK8/UUbxewxPi/6w5lWiHOO/iA
+Tgu5mCICThaLr9tmlH+hKwnIo+MKT8k6Dw/FTrwUIBHfVZODZBnkD4JikoiVgLW
9bWD/wV1ZBNP7v9N9+V8accpNx9gkIdAxmND/HomsJmfiK0FT6tvI18lfm93oYh+
bx3Cb1KMG+XDizFa/rmWgFGw3/lRJwjv8kB64Mhm7of4tFIjG3SMktlvmzqeu+Yh
nPdklPK/Fp7ir6J/xdGJgRaqVkF7de8gtMcqB0qiWGM+84znHf39eenjADpYvX6C
lOS0uB2VdENCN98tMvMsumRrECxLGCnIpQCLCVimzX3iMtYycFjBzhjDYCJv7lMX
grpufFNNu+ncNHhcUZfM2An2fZC837PbMSsyXO8BP1IlVQviIRVJCHhj1E6N6pXG
6JUpc5HVrk7JZ2PLaql4LaB0rApCUV9AnsJ67RhVfKls8u6+AGF2J7UTs9eCEeMT
f0mknSMZrQYtrg+UtXSN2lLushmo/o1unEAlSSQJU4DSHF784GablNtOPtMgVQJP
m48QG331dhwA77pY6tv63mZGZZyWVKD6u90EqKVgZGXM1IN+/XcilLh2Jouhwr+k
Z2GVQUo6k5Rw7SeXLNSUsRBStIRDI7/62/gSBEq35GiwtN8rfFlOjK0AyY3NKqMt
NKGN3BmRC7kZ//zTw0Pnw/VJcm9c4zztiQ4ZOnvBvxmJh57MG+Aw9NarNGZqLQqn
sjRoW7uh5qdZknySxcUX7s7dUbXLm5uUpbt6BiVCbcgFCSMhCDKbCJvFTnz9Cy7g
hanrAblYZkQ1v45qqXMiUXcX7S0itKwZsuI9VYkWmEoeWHvF9qG+MtTgmIWKq05q
SOBGPLajXikXZ7N/L2IheA+zu7HqM1ie2ULLbRsgNDj0u+EsPC93PkzBFJ/1eb2n
7Tyo7NRY3kW2L5rWqOpVI14nu02Hed1clrxDWdzzo51wfDAM85r9/DDt3Iyguw5v
mxm8TZAyWdLKWYnApgaZmgWr9mL05av8rmsiAuj/ZuzZdZx8JZAFuly5FEqZdzhK
iWLOQGL/GgEHP3onsR2uxaZEUROjh7l5yPV1gRVh1g91Ncy3s1zFq0XVk/yZ0Fs5
ZV6K2IMGlaLOKCB8M0eN5F3cNYa7n7OrZX/N8AENmYl3lcu3evMwVnTkyE0E87fH
Vc2DW9XFOoBT6rDI3F21+p/hnCJh4Xly9nw7cmzzcmgMWkqsVImERBRsadCQQ91N
tgAJLdT9ejf9b9610HvMimfl4EiDJw8Zs+Gswnyr0BbB4kzCW40EvuO8kpbEkL7f
JmQ2fvHlbbNuyC/CdJelOrwKvLXAayQ/cGRGgv+TYaFLPt75sCsfv9i4Ml34Kkpq
lHnBUwKvwaOxfnEIEh47I5iVI2nWLC/7CtbgXc1YeoLgYLjLYlpM9dxV/55qiivq
/jlai53df4BhAA5S8b6Et+OyWvyt8sdLi4p9IoIKRIaXacYBoBCJfZ+QCMvtGau0
vSbrNvb1TwALI9D06nwlHaqGOUKUWaCGrStNDek8BHZdepnXcgwPtr2X5/rvneZc
2LHS4Q7idQUa1VO63RYQfDP8na2RiAcoDe2lTr/p5OA9KP0y/c1XPoR73JTCdjXw
gmu1s2g2208JmiO0FRVybC7cZrCcQQpLNX35gHej17tjlAyHa9HoQGpvqW9woLYP
DUWEYDS0YHPENbg8IXVdBaQP1lo5LY4HHCQQDIj0iBnrgDwd6NX5NuMZiLnE2qOW
25mbDaPxts8WPIlUy1lUr7nHUuu5P4TA6jNfwdRrY9YPhnH8OcaubMx5ufalAf7V
Q9IdBnH0eUKVzwLCQzqMDOfW4bsRYjqmUORuRH9W5PLyY0c5kSXegw+3AKYYM49k
NCXA9mYDbmquxqKE25GcvAuTd1QDgZPlQDPBefPvjSGhbfvBT05KNDQrJml8oei8
Uhu11K4gmPRlFLI2pW+lWuBUVFWzVtyxKNmJ/1UqShfUPilOH1Jv5KcNu9lxuecJ
hgoE9aP5bIMjk4G1a4RDdimM/sgxXdLyueuYpanhv52haLi0xJhLtvZG87xVZua9
NA10rX0/KI6yoSH5P94+WS/cZtQIsNx5fxbeC2IKUZ4fKrEiuN8ZqTmbFOqufqNl
QLLAYYMzWyJRgj3G8RnvS95aQnUuZLMSF/WQL4tYcdzuKvcwFAB9OUuALFWKh8+S
MzurstHYjclbkeZSlkj1uUw1F4WJv4/NvqYBc8DMqebkD6sr8+lyn3ZywoBrLRVb
y/AFov/VNx3Gu7VlT3r3EkVETFJDyMV1QAmmXYz6dvCWHvA426fnnfoD4phln9hp
qbeUpmdH+J/46fKUww/NC7e8mVUG34WnjTqBzcaIUKXfYXIAEI63nJHMZi24AH1I
xigmGIXJGHnfpM16jy2Rc/3NX/p9L4U0kOKXF9NcQ7u0CF8/kbvjEbMJJciwR2M3
TSOe0OeezuRWtLVzU9eAZ1zUFF2KMp1B/efMj9pomIdRptK5nAXSMGzua8nqkOKe
fZqoxdst7cql9E6AgCUH1/KGTIl+6iIPjAZHBrIeDZ3fcz8px+NByLVaoHYu4htg
4y7LhmJ8G4GwsKha3FA8CWtHSMuCq/7dsJjpubuPmIGSZr6lKBuaFfNd5txRJln/
irhuOwes5x3mC/Gh1qWTYtJEm3aRdZfz2W2B7GWj4L4o8IOBKqVnSqtK5LYYQ/Th
w/UFuu4lqy6cW3PAfL78OaLej+yc05j3//PmhA4l2ztc52gs95UkrtEn/MHvRDW5
oe5NPATEkGVb46KAqVrKlfSMB+S2k+07+Ed+c1llVmJZeN/MzySK9KAEZg0e8cEm
a4j2IEgtUtxqjv7pJtrZfVg7I4HLuPjc0F02FazUimHY7nByJ1sckk/5zqDz8JTK
fb+pNK+pkGk8BMx7sY/I2nl5Y2h0uQ+dfcNiG9hzO1Dxr2CwcY/LiprDrz96INIz
psxZ8iRSA80WD6y0j3HT/T1jp6U8F/qA0vgXO0k9gSbkkTgQxF4hbyRWRlB8TAGQ
ZDeBwXFS3TylRedTFZ6gelFEE6pmPA/og5fxP+im51lT2y9qxNBRNjK/ZjJ6LEtU
uicCDmTzUPpcMnZK7uQ6jAqkAOIV+0N15egpkup3DxgsnuuY3RHfu5dzPIkAfpzS
qpxABRn+04YKxAKHRfiACIrUXfxW97Br2XYFAN2cU7uU4dVr/N5OlPBYyWqmoiUR
2m0S1NtGnuqFUaystvUvO09uL6ih4MWPtyh9UyuZAnQygq35hArV9kZeK9wWtsXq
SltWTqnycvuG9NBjZ7Sk6oj/pfe3JQsawY0T0fZtNvT3QqRs3G2o+Co7S8apUMfc
OwVs/XAi2cpAdPYN6YPRTpe6oen1hqoblFE+1gZURZQPs5Pl92j4OQmbfY8iBgPG
vKXIc1AajEMlhhrxUVLm9xtvl0/qofgGL7buO3yMeHHdAHUxdVeqb+Nn1d9QHVYL
TrLauM17Gbkend/PKM3ZEL7sxfD9ERBVhJWI8pAVMLiL6sYkFpLSYXcQRt2HGE+P
7bgzRPDVch0jjG4NVdOtr5nfP0ZC/PMZ9KFweXijzhGFEMgWtAi4MngrpbuXvSCT
Mvy1RvTIzbmi7Fa1Y4jBPFCEHXPvL4PWK5kyZJPAhsrkPogImCQcT9ySMtHVA+fO
B46Uexd9SjGYXh61C7r9g/8S7a9MWrzg7G7Hi879F8c2CSWZWo30qGlcmt8AH8qh
lCHlaWtDB5pMCOZxbVGTmolZDTk5JyatMALszhgOkXRKT4ntPyKdi5Z2TRVVsg2T
9yFPb3WjolIf2fwz+Zp2I609xs9v2DX81RypYBgbMm7TvC9F1SimUtyTJPgyEiIv
Y7TKkI99PQMskrUIRhTJ1U5mjPI6ogQTITPHOXhnYsNsDRFShwdmaBixI2eMmcU4
faMY44H0Qx6/3iTPaH55OjqrjnOogEV9LhvUz7hiPt6yEbhF72MiMB6ZqIeeX5zo
Zo8Ouruf7EwV1aPC5f47LK4LgFdNXmRJ72uFBFiPmF1KjDEMFma7Tm10Cm2rOW1D
ia2Jgu0pv6+dqEt8BA06UwWjuKwVXnjTUspL0ywm9V8l1jproVqVCsiaJ/mfnDqa
2GEJeiC158+KMeHSW9sTW4tqfa1WcGUPqJPCZ/FMR4dRD4QY+GKT2vOHTmQVYiv2
dsT5cRpGYJbJCpJPJxpS3aA9MrweRBQOYGS6VJvykv2FSAyrbzSNuS6om9QR+t0L
mgo56kahJEdwswBOmTB0SEhW+Acv0B6GQqy1AzdAtPOMND++mnZy+irAW1+BQB6y
nrjgNI/+8C7o9AKx3EjgilsjQ6UvMiYKYIWPTPASzrFfwfNgK2Ym5wQi2hhcB4hx
dDJ6oI5C/IneArY3NsLA3mCS6NUQ/JtgFqc2FWMSYjjCvuRlXLq/y9fkjVOLeE3C
6mE+dggu1EKxaWCuEebq+jYHz6LjnAdLtC0yiJeY2ar/omhliidwjwjBVrfyfpii
1i22T/WIrv8SrxKM5l9Fn9JhqZV07ZJWh4FPU8BwVUhAneNpOu5jM4D8gArLayNT
4R8MYkyX5HKJFow6t3CeYaBgbe/ktERpEIhK2XFZHJtOYWScKDsSL25MPqMl0FTB
4RxAwT0vw3tDzsNi/+1WoL559rjukJMXVaIVjrbiMeg65BnIi9qUM/YdbGkFCB4j
z1WslcQDxqmfxWyqITnWXX6QDiW7p4Ev94kbvzLSIXscczxoRibMGyLRJ0BxBigN
6l0ZKVvKTo1/XZdvCem2zOu/LNhG/BvVfGykn1ApBZNRc6gBFbTrXvfHc32Vxq7w
glimq93bxxJODw1LdZj3oh3nwgUp1jGPGFngDyNmFqY9mpQGywUQjai00G3jC46I
4OxoxcXMDDQ0bkEJpPYdYHQBmWTmH6lGTPzlj3PVpAZCIOFvqQiBg6LZjqwJVEuq
7xSNT6CEtzuU2e0KwUaLks1DOgnyggv/Bo/bzIjPnugI4q2JeSH2pDiCihJC4Paa
gc+5l9HUSS8DJVyVR6ciquCoU85SZSyVh1wihllZt7/ccrI5l5EZf69UEJcd3lqG
XqAlxsredA5Bj8bjO/pGrGg2JwRFEKC06UHiDyRl59ENaaCQBGt9CugJdntzLxpo
oDVMb6XQ3C6lDqE7r1xBGanSVSPp/i1ocr99khTHnrtll2hZkWnl9G5o9VaEks9i
jvIwOOJ0m3fu484F+YBHadV9W7ebrVFNTR5rQoGnpdHBKUs8kLHOTnrQOiUPl5SU
+7nLuTvap/AK6w6AomGyGlNLTfj+k35zkJ7m8/IA24WxuXeTQYL7Ds4z8L+fAudQ
wRsw0JYW/gpOTUno7o3djVyb34HqHT2YZOHLPmYpHO02vcN6N2IOApZ/cC0ZowLe
BA7rHqyQ4odaPT28c2RFsBNV+IUROapj386qdQD0NA7hHhxc4CGCOuIaqmAaKlCa
anuMKjXxFAg18UWgNBCiUwOPfotqzPfSsMJVVv7xEzkJ90BzCCF/Vb2hYybY5r3n
b62SXfNiw5+qI3uy6+MyAKxkqasQD7KAFiK9DA3sW7TictktaceLAQt0ie0lPkI/
dETYVdXGS+TFZrVhjsYztGuIjMwNkdwlxUwXG/Re4MqLwhDyvnDUC4lwkRjV+rev
cUAhtw4FjvEV9L6tNIYffrmuk1uj0B+vwid0MuR7VYRJmG97EDXozWthlDnRQV6N
GcN7A2dD30jzcDNeYDMNLZxuWBvL00wFA5oTs+txateeB9gEE6ZQZhY4diFxw5+n
IvDCMcr0sObWpxrri8B4ShMiAx1LjzRErdbc47qpErhyPQ7TiWoJBvuoyPUzLT3Z
GbOuVDWSfy1JxuCOsRDR+M915mkuNzs+MMFeGZA0xtq4y7Kw//8yD7VCKx+/H0DN
U3MtB16ag1FKYRVx13V9y/5IB8XQKr/y/FAgakSFlHe2J9CGZImGHMXb1boyG6CK
x2M59UdJp4SPNdSrCbAYrszXHRbpaSQN3a+4D745/wspFCuLq5pyZbJugoChs+zO
T/+nd8ekS5Gp1kcJM6tXgBh+RjZz/3qo7MaaKJXjRvFmyPvb0BY/PNF6hsXt2cTU
ShGyXrozJ59cziEU3d6TNtDzmeL4CsyEH/QhCvejqX+XZmjG1104lW2Vo32quu7W
FtQZZ21TFg1eGdivmjHkusz2uMXlZIM7WT+T8lhVJJfFQTDLS9hCa24j5S3OqzrU
E7BxbD9DWOYp2M8+hI5T2sbbTnp27ExTEyAuARTTFy6xJgRHE4BjO1/bUKMWeEF3
DCpZG7PcPOyhFUHFJ+u/AUqYU2q+rgwWFUfY+KdOPv9uKLfGxaqNHpDl88Okk2Ah
M4XI0zEAtnxKP5HcKb/UDEIwjCDK8PHucrRYC+eUOUtHjyV2VbxMKLb8InmhP07z
HUnIaeW7gKG29kTYTy8izOD9Y1muAMHfIkQkYd4afYRrhTgPaSYEanrmPQOVpjKF
BE89wTpR2rHYLSEWBVPntDQ3jGTt+R7lUYMR9nvYRhjuPH5fxfvTQfMbHTp0Sy9E
Tb6EyOEi4ZhjKJv5UH0Z1aCxmSwMcO0g1l19eiE1z1yDaH6cFvxwFrFBeK4xYO2N
lnjpCs/s6v/cASuWzZR4D3lQPD6aCkES4tYXsMopyzQFFQK9PTGsldjJH3tqfXda
zslbF2bEDdJMcaEAOj5DOnvkEdYdTJFz39XU1DjooEsnCm/opJErVCfGBPi9bp/j
tXicrjxGcFJLPhOP6yHytC89mKQVNZpq3SaD7eOg5PKyd+z+SDtdX3/zcz2bn8i2
G9sMWMKDjuEkkEpPNJWLwU91pyIVAjZP8HpJ8U+IVB4k7l9shGzkfxh4Jky7V/Sc
9QRZRoX2QR9KIS5jNbS5ctPKQwqvHgni4PqvlxhFRwxN5WgKVCngu334dSBi4tKr
b0KsJur0jStv6mX/Xf5Mz9hS/+p1vukJwxdiC9DSo6Jt2YcXvqlWwHfuXebTBKjc
Xn7PkR0HGIeT0xGOQq1bvHbHD1mpJdxWUBKebCwyCKtdmNpDgUWrQ4VDLHIG0b9Y
C8JnQWwB/TQzmYypFLKmWvY079VoknUbEOe0w3Lr6EASvF6l3a17oBsyO+Qr35DF
71HoTsdW2rYmZ1g3Z5IuoAuxFElCOE3ptRklfPTEBtZpuT3YvbSjaarMQxvE6/xk
wGOcgitwAbmf+XYVUtastH8dZ6lsewasQN5s7YJ1w64R61RQRR9o7KtARzgSVuzI
rQkQ6/fWdGJ8N5H55SRUpmKhyL4DqcdSmILFZFPu+XGEkk9zkjDapsiGG0A/cZWu
J3Fl6Z/OtVw7IdXxCEzT192Vv+fuhGwl6JzNNSlbqaSSeysegCv1hkWAcvSAizAn
dhD0UDjJ0PYdykXKkX8DWodsLCmp+e+Bs5Y/Ewbk5yStSnm7DvMi1eeXFfdJtFSR
Is37hHsfMbWx1Cw4zh7Kx2OaH2YSOC8oBtZXQYXox+sPnxfNf+uOEkZQS83XgzQB
O507lig5fBYCesqYYz8L7f8EXNjgmfLEbWju3EW3qB0Mp+L3eBP1Cac23vLbIT06
PzRPIwiFTOFoWE1hj61XbaZWrNJ+iZe8B7EJ6AEy6C9SCkncME/Vn+dPSoKigiuT
zB4pZ9ApdFR4Cx4jYbrp1jlVXGvnKahDSfpMtyv4n5g3GkcKhV8iV7b/A2dI6kny
RWHj9Vq52inMmD8U5W8s3Kq9QgKH6/ZfcMUuDU819aFXPX+OKhuEElvM/zm72b3g
PElipwNqjzdtWuNp8XwLU0ZQiFaQPHNI3CMANGE8h0ydOxwkeAXAYIfeAAuhEJT4
OVbNcrbScoDfieiuIkIpHFUHI0xRG68V361zJxPzWwRZiRM+1+1uj9xloUIqsLeI
zZ46xvIade4/E+eAGIagL8NIA8OJvlaCbnMO6NJeuuuKowXsXa0nWgHcvUy0tlK+
qjGVM+IDT/00fE1IiN7BLyLX8E782gMqN+AcLa83vZYb8PBUchTZH1ccDK8W4oQi
6kcpZZyo/u+Xg4ifv83QONKyqW3CXF1oK3VuVIvRQAQPS7kuWpj1h8IYidzH5YWv
Rs78tME7Erj25tnO5SqLbyFanaWBXqeB/FbnsJRDck7DZCaKcSTAcs4E6wprrkbd
QOc698dblgSzPPaA5FZOsEq/HroRznJKxxIaST0JuFbPoGaBUEZzc/HpU0PBWcCx
broj/yyr+B6cIz1CHmf+r+ltJ5bKeR/HhhJPThDk3PrtokxWFoQjexo2C+DpzNu6
fWULVzE8RjkLAfP7Z+bhPpjZ/23EgM9GS3beIiOrnQvMFch2HHo3KL9CLe8HBYV8
K9XEf0GzKY3YhbpyYwTkZHTTYC/FGG9zCJ1/Te/+vDEjtDTNgvL284/IDsQdwIFf
Yih2nu/ihs7iLsAVeI8MjvszDS1ZmXFzV/YG/4DK0DUhSz8vv18KBgkg3MJNv1WV
KMAVZ9MppVyMYM+8s6skPKq++g66MEN1ustV/OiA9i/ksycuR/imq7bQUNEP3wVY
RyqNOU2ZqnpkwIuQFLfhOI1JUxg3A7FXr3KZ+N1Yv+jcTxu/rfuqDKFrgL6/oRX6
GdKQApgxo5BHaztnjg3cGZf4bApQc6H3tBRi9zrMepFgV5wycncnlmztvmE/tezG
zlcK0+FatrGc22xglIivFOPZEGGTvZQthW0Se/x0bXlr0vma58MGApNkccgK2EnO
v7HuhJmLqRjzpKT1zbcheoV8a/V9kwlgBl7sX77RYR+MBxRCDbXJRBdv7lIjXuQk
xzKK5+iFyVP6FBeNXV5ZSYvqtSSEM2cyzZI+PuDrLTiyTf5NOtJCrJ6h4ToOSFtD
ROD1IvS8dm6627ogJ56FLlpoB2H+HehbYZaBkOZsJXx6MU45lvrpi1Ug/mxrGs9S
0VHbhFfNFlYY+VqROBGpsdbZCQamaSNd9Y2gne35GBe1+hGE616N+bjEUvGQ+ZZF
MBd87SG+cfTkzHD7z0cHQ8vO+fHTcvp9Q7oIzq2ZeNtN2MZIgwgoWV3FCTJc9g35
EmINxDCJOL29chvGDtMDSJQFxb2muh8FfMxJa1oZ/+nO8iAJruB9AF2uueAVSl8q
uqYLQlLcRbCxiW4p0wouFtuuEhkm8enxC9r2MchdNjm7wtVpVJ+P4HCOF4aSFZL6
LULzbBJ3vIKFgnm3n6QF/qYBovzFouX/Asw/NYjpbW0womoAl/ND/8g8sg70WIsJ
yHX9KILWwJjBOfWeby9FEnk4Tx+nbNWsCPS8Z9GSWmKBlBEP9BMXsCvEpjZhuOGE
bxeR4pqk0uq41N6QgStPygwVbGoJRLGyf965mEWkvyKXxPxpci/Fyx5mcXJ5rxNu
KSljf64gNtCe5M53o2bmDfLWXDhm+xVHcwcYwCsTEiw1IyHgd5IlrpVxLSgwkmM5
Snrd5blcVtwYAdz9vn1iaUoOcUeK79Ct7ebblHV9F9egtd+LTfonwOEHayErvTa+
MaH1PLOg4kiPjyKGF/ZhEjgwRX4vpFyXEpyO6oXeXcR+Ou5CUa95qU8zGGtCHNyn
wP0BighTL+tRF3fYfB0ewUzJ9rv16UtN0gU2xAkFhuV04n4c8IgrWWnvx78RRlCj
OOkAV+Lyk17SS2Nlqz5dbUUj/GWMck6YN09i5nYjFhQBp+yKXsky8jfTrbFv4nh2
8XaSphRplGkNOw79VgMf1bNOAh6dH/OCU/zcwOobS0pxthMYUEgRbI+2l/8BGyRp
ZsOtyCx5UaUpVjXXlu0DSD5BqLq5FT4HgRQeMVsN3qtacwWRgm+RfA/EmXRl5c9F
v2I7naBHq2xj30LcxmChqO5Vjt5bc9YJVmSsjJBX+uPqn8qqnXE0mn6d//E7WKiP
opcAq1UOAESF/bxOiQOcHVGm4zkr/kVOf3JOFGJRUP0cdmeuv+z2OsP0AiMh9Hvg
DheBrr5/gcSQdLvSc6FbCSx8MLvPUZNo93KrwBASmEnQv0Li0/fnVO05DeQxOdIe
VrF0GmkP6r2BUAHUG9kdDwnpLUbY6U7NVnfFL575B94QTumeQrJjB2f/Dq8rC3td
iDu9BMWQPc3kFvhMbGpFFnW3EASleyEwABhzLk2KGHYuYSEgvAE3WAc+0Z9lYCR4
NRRFLUEBVKiAv1EGpKT3iSrfZ76ofbiJtiJav28oHByvbaqT9iY9cTWFqryXYUH1
WWacYpW9EqFJjjBY6NSrc+tvTgDzI1xhBSBJ8xNm7c0VlLoGiGpqmDXjsvx9rEoZ
wG5WBooop6Nu6Zn9/y6uW4JZe5rApKvvd3KQvF29RnQuXdjrPEKGtiwsDRV37f6c
OOeK3sQLxJV44XodxZKu13Ysyr1EITXvQC6vqKBvlo6el+3R/k0tqWxzdqVmlMlF
JzU3WqP3/wSLA64xV/YPWO4Yg09X/DRA1Opn+ezUEu/vVuIMmtWTPQVDVqp0WpQi
IJlU5kaH7Gi9GJz9/i1Wwigo+rP21jgdF+icjOh1lGqDuiEsGqyb8yetU1GgGJ0x
z3oTRLuKo9wvhaL2uCgj3cpU6uaO+4gOwztyTrePQHf97iE5B6OPm6Vk1FXxTwiD
MJH5vKNMDPXG1K+tRbkyp8lPGMZOM4tGYvXUMilZJbDOWa6fTvhyB7Z8pTbeRlIT
DrbQbT8gQX7gDZGkR3X18Hmbg0A1Zsq5GnZ/CVOcIkzTbaScTBN7LApdYsBYVXBN
Rqsb2Kjo13Y8nv8lUviKevzYCcVZo9bFxvReBnQLcj3bdrdWd8iH6dH16R9HzRpx
YttAuKOy/SiEGE8ytFrd4MszH4mYxG4kfIMcfDp8R4j4I9bzt/HJ0jpAY+OgFcUK
4au2OMYcr9Y0l7nQp0//llTQ2086PjmQjMtj2P7PrszJmGAOcrQVvFHq/J7jSufj
bBdbhmrPq9ZGca0zxdQz7pDL0f8femXQLcvERekLYNJNLq7CsfJM01Y+H2XMZaL0
mR2GcGzyyhkgW759A7rCuyaZsPZODny+9QV1pzj0UEqA2nI50NbQabQdveLnNzBx
H7+istTgzvP0qxppMsWf6yHRgc94eUI4xLzgcDGYuFgNiHK64rRwlQZdzpcQobxG
cGFiJy8kVpBaRixuqoUddfDP90LAOQhk9PL7Ercn3L0MaPZDPyKajI9XwtdqfyqO
YKG9zU7QHR9aQze0nplUrLhK0tMxpPX6pZYLt9vWmMNhfoV3m10YVmCrbGNpUVlz
2SSrcSRtYEYNiZpQwHAqHYDIACH+V4JdvK+GQBmP+tzt+YmaB7nJJLyEXO03rVyI
hvUtRMtQle2m9zWk107ve8/9m+HvkQxYFN8p/Wv4jmwJsgt+HYf3u5z5oZJgL7gK
Y0OyapP/hHtusZikX80eUz/PdP2p6mGk8g9rNqULY/BzIEOteU/rEFfC2emmOxQC
+0D6D5c1V57Mz1mdG3OWMe4yG06gYLF92YUKN8WzWAKM7k+A3nG00Clx8bqPUSxO
0YtVFcYHEsuUW0OcgS7jDG4dgnDGpvwT3Gk4f1oPGETj+ny1XwmJtSrHzfklOKO4
7az+Acc2LxItDMbekl5sfeT3AQyNuv5TgNrCMoVzQwdmbKPmtcVhT3D9iUFnMLri
y7ywU9AZXRgEWh2Ws/+eByY/epOLDUEm9d7cXWQCY3uEjnsn2shk0fVHuR/DHr7Z
NUxZsXB550DVFX6AlLcmMtILU3QFpb8P5VUFX/ySmEGJCTsdCQU+k4OH0F/UVtVr
XXtUE1PtdbeSDr48jB6o8Xo/39sTtQanLo1ufA8lwNrnw0lHJaDCOhmh9o96nSlm
CUIB2fAPQs3eTrmGNUb1JTjCuf9k3b9ut4Zo4kXBDfXXh/rqHyYGNQDk4jAxkjIQ
FQOfqk2We56J6X3arHj4uBU/cwDvbHgoj3rdzbUbJdytRqY+guJCIL3G6uVm/H1P
zNBu0sVahSZ7X7bu4Kj+ZeUa6t4gzShx42gYXGz2gLHHM3CqKiO1IWa5vSNxbOVf
+zYmh2BYrzY3SLcWhDSjCBjUdtG3YJhgBL2PtUN+ZIdAlaR7DYX67OMI8h7DaX4D
FJh8KmYqs2A3VMqit96t4/DGEN7pOmFr0TZS67GvIoxdvLHHoyPM9fw/SWvfzIQw
o/2RfpNbMGZarJLfy1KZytasdc1KjJZ/RGZBNc8dI4+xcBT0i1QuoaJ08fDtcxbo
skHg9SDjoV1ripaq+ZZ4BL6lRA917/thY3GtVk5Db79wmTGOVlNul24ZiwDWk+JS
UjtxIt3ViCderOQKmRf0DrKzPb/AyMZ8Fiuga2pvRv500S5SnG4BZNIQI66YnwT7
2Lu0l55p5v2c7XLB2ss0h7z3TOhhK6ncvis2o3wy+wbSZ/SioHch56C3WevUSf0P
yoEVFVEohlsVnWHJuYgd1LINzi33kllupJcEhMkridoW/+JZYhkxnJyh4ncYyku8
gOek2VE4kmAOeea+c1TUTrV2K6m/PNwfTN3IlUhYIq7FrooZh6JfWi9i1cHWTtsC
u+M1ZY6oaH2xuX60SmqZtNpDAgxUSkK0hmeC4QUVuAP46yGZ+TioBygGGm9t7c5h
QLbprI2IwDaEfA5iBszWWS95ruL/Zan3/dPamRHAYxluYXNr95vEYNVZiCNvu0g3
QFwXEIYvhlTvX201oSLqODZCvZXyuxwHcs5+X3MFTDl4hXWcAYak3e90lDZVxjKZ
ex89EwSw3a8rJSgxjc6CPH3IzVdAgk4yJ75vNHo9Kp5SZqGE4fvY7pRGcriSBGfH
DP5A14oWLM/rjnh2sQIXyPyX69VagDZ1VdF+Yp4IE1oR8IwfSjLnI74jm/3298ia
6AXA0CXDYsj9YM9hdlIP6NmTegq2rpZTe2nv7c3TQsPgvzK0YxyDwj8mXd9WU9ui
VUEf4rPsqPrsT5Xb5OQzxXxmSf3PzZ14YQWxoFgBoUisOU1FQt1b4IuMv6a9B8ps
cDYGLOT/ODXYv61q1EDWUI/jjm8U8ZqBKwNBGY8Na+Zhu0lEJ0ayA4AUdAT+6YWH
Itr6D6wlG/g9EhOmcLaclo16EyfupEIk9cTu1Sz7o/WTIyfeMrOQcTIwLH4xQ6DH
rcXjf3nK9rve2ucRfCuApnUeZEQsirvnq3qGSFsfRWEGG7oXVTJwjZXLEjTv8dSO
T0BrFzG6k/wMYT1eu354d7BxZFb2Tb9SyYLPabShrjrIjIcDbVXwuF6Oae41X/Wi
OwNtGjLNmVHzr0wAv5CNmGhPxGXFfPgNEeqOVwCOxxXfeyWPPotl7ut2y4QlkLeF
xSelaOQ8ubz3iMvSguM8BRcep8v3BxrSNwuKP4HbjK1M7RJnzDARxcIENR3YV9b+
24SSd+XU/Q5v5aVby64KcglvQwUkFFQy7uDpLcZjyDc90oWmC/XzALoxlIMr9iAH
fQ/kZBwNUik9CTDxPUSFm2t266LPvhfe33rcjL/X2Uv3u3jAQ8+LiXtmxOTpLQtE
sECBNpV5GIuIw7xDbgkB6XL/cvGkDkCBSOlIpAU6mzsKjK/H8hSkwm5Cngb++eSD
18zhHbO1OzS7f69sN1ZZiEkvAoqIEUD0asf1PL6De76r7xVtZWdN98molpLqBOzX
fa0J5uDPowcV55jNRKUQVsSzzEa/RJ0hpMhw7GKuCYnLM2de0Sns6pmwrtEc8rUw
XTt8y4dYC/j5g3wLh6h29cy/44mZ3J+n84CMsDQ6ZA2oNzA1CrDuEeJPxSJ5Sk5m
uAImJImrVBXawfFCuiIbCocPA+AuxU6e40pZG2IxXxg0wo4ZeQsUMhotg4YQS4Hw
jH/JikojdORDidf9RfEWWsLc4wvIH2VkaoLclU1e1B3NXm1gKZUmlXciMDe3LuDN
hF+G5E3tzWf+loe+WTmcY3X/6tsjdV9igOljdADJo4G9NKlzfeTAy9kwG8Jll4BC
Csb43Q7varPwQcLTZCapdz/aN0TjZNfH8jf0Bo6Mdz3lYgUaN+qp6AVTi+cr28mK
4D6vqxWJUDLMok834LDetLaDmCBVCZ+6P4j/+09plUApkPtuW5ZAg1WnVjNQpYZh
VHwSfPcv4Z5+DBA1go+KUrR9pxmyOHydQcQwlMag2d6MuY8lEt/2bub8cjndnjj1
pPdbjqfs6+HoHciuMBKsoATmDf4xWV+y7bVAHsrSnbCEofDG31OBc9BnIh9Y05Vz
2RUnFF1u91GvgpoU6d6T4Mc+FJhZ4xaZaxuW4j5kgPwM1osVuyaqym8K2gnulFYX
6DkYZ4E+/x+eXxYjKh7hEWeXXL9YQJvke93tN0J7LUBd7xIUDOFhoAe5kQ5mAFtX
M4FXJ3JSm9y1nuNxfSxCJH+i+UhMRlyh2NMPB7ymC89PcPEcs323Bebb4/aKb11e
7XQcUgfvRkO/8Lz2Hz/GSyUN13o+ZMLhfEjjB73lpH1XFf/KOUby6ZVM0r9FXy1U
KYC3nwVj1i9CNnf5WvQvKfmehs4fOhiaGrYSIXtutPxdW4UOgOl6q3pBgokRjKmp
TmwXDx6yRfXCFKxN3CRdTl8K1EPeDRuvJDGpaEp4x1yPgWqxH3qTo0lkTPFcKqCp
hrtkAjhHyhNbJ8RxlT+RXllma75dFkUTCgDbwqqxuqEh5F+YNHDE5t0FHfvvB00B
hwESpxcpmh/BQgcartGjEF08dhEOeANEygf6xCJAk89jt+va673qrgPhMEbQzbMa
iZMjqfe2kPJz+IGkhUjEZSLlEdXj62Uy+6I+JA3lbD6ckchSbbcnuoZxie602LFg
r7q/pz8JoiGHbBeeqviwP2dbtflvcsTpf9aPg2ckY2y1gJkcMD1AApwxYTeL0vAI
KzDF2F46Ec5JpX6rrzA82g655l0K1Uxdl9uSnJefmPiviLTYhHQyMLimL/nU8H87
k+x//vndlRRBzioUkKqlpBD5t5tKC0aR9yedblHulXnQ5POaaEgKZ03ZyNMyHtDH
07C8uYWXvHSnJnJUNvYt24+DRXImZXyZSnSQbtYhPHzZQJU2buWMHvqSeELXOQtU
UnB9ZJu7rmfIXahOhceUnxk6PSE7H0NkKiO9tcCuJDcAUhDApv8u8iXWkNwVY9Zz
w8UK2KQQKGk7JqUbVHHONXxADlOkswoQ+zeA7BJlCXkTb3Iqv+VxdFm+QFxK0mPp
DVdMrwhAeUDvalIbEXiEaFFOy9WbmF3Zb9HaSyWiGcf/oRRYcJPG0K6kDLtVKjRJ
mauA8qvIHXPkeyo2WIqeEh1z6Kp/amYTq6NA7/4QUrjVE8ZMHw2q4So3FZzvqDrr
4wxfa6DVpmT2neNVW1+9FQFo3XBoJzR9LzTTTfqfBgfFfBhRZp6J5vzHe0ns+SaU
zPyWbe8FfKmv0XchrAkD3IuxfB28Rj5fXqHAU1q6RupkUI4rk+/oJpOQ7eGGXjjB
1ugRs7fAOsrlr2GI7MUuRg9KFTSH9ZW8aN9dePx0STyVjp7uXb1SgwINO3MQRsdM
4npCK7mbllVRdvVucTQU+1qLxn7LmMg55mwbyoSewK0+fWcUR8RrJ6/AaEpIcXwr
9LuZVLwvlH0y1J/nx5VEnCU5U9IYKJD2oWg+8AI8397w7HkXsZ/XwsOvGFzkLEVv
stwHYYOAN8l5q57uc4zZyEs4RHdajzssPSA3bAJaj4/bbnT+RKaCJHBbROZF51+J
OnPOEXir7PfHV08Hhs3UmLSm7cvS0uHIqHrU1gEkAPXkJdwGxCS+Tl6JEUUKVo+J
qBZBvSTf07YhTqAnbBioQF8dYrVsqchjLmKw5WWF2HvI6ZnT4SUc9mel3nJ9tDAy
MKqhqSIDIQoTqhbq9ZLiznmIDNLFYCxTvrpF+GXdROEScpqEBIt4js0nCx6wfj3j
bKPfVwJcYmso2WzuhZDReLLl6zATq12iEOnC+42EtdJ0tSN/5vyy962l2aW1KZ9c
6udnZNlsl2VGh5T5G/uxiUM9YRvqEZrlkI80MXQOPidE4FqfeV6ppeIbx7xJQ/OM
c86ufY/83zfS3wCsjb8+aMUPuBJnXgDYTcbN9YqeDs99mQ8vsX7rZkFO7Opi04dr
apmfrCs+rkf26341U23i6RMngpODco89jySERvbFsThFJ9g82rj5Y+dBnCXpEUIe
pX4cZeGYkH5OfUcC/a1rPWimA14RIAD47ddzLRYF14TNNr9lzJ10m2FuaRPK4R8f
hsBEcv4fV4gbCVlnEtsqnE3Vt3nzV+j4WZh6sOBWVD6Mhb4uy3YlJaDQbynEFaIx
/ZZXZiMK8B1bOjs9PI3ldhC+UXNpsxBXJz6bk7yGa9tqokQIzVfAcYmuG47g10wd
TfymuVOJxH10l5/RZrPeUl00P5+2M03yHP6/Jgt03sQuKscza1eBxOi9jPh38Pg7
KsL4+qf6PHJGlnmqY16QwQpncdjCTiiGX+RGDj45wnuOPskbL0hb/JnVdef2e8bc
w+l1TmLJCMQFM/f+inL3SwMDUJ8rClVNrBUXQHX/IBx1kyQG3fgoXoOuwe98ozWX
jlPsWuC2xGFlZfA2E6i/Nx41pjvHw/ktDVjDK6mt+WG+zbxZ+sJCtb/n0aFVF8gg
yGkG2PHIlZbUP9TAdz53gViXdis21MZtLAy3MWYNTxBqdW9AqifLuIncDTLZKjnU
mzVIjUD4xG2TsxTOck4Axl+wwIuFox38tcgVJp/NKHwWC+v6z2kQH/lAXtJRySnH
06zLNT5lotA+lPK2tsr14U607pvxwqvm/WswZ1WzUt5PRRBYFM4D06s5EOHf7yzC
ZLy3oAG7DJ3UuC0+Oax8RTuRbvuvtdOk9qeY+OkpGKS2zDnnOIM2fSQr+Kxtw2xS
Cb/MqnoTE7/t9AFGt+E1Ek8LSQyE+4rdOGTi6EZREtNpmrDglst00hnq3zfppeya
Y+HE2Kd3B+kQBGaHW5ppizcWtcfyRGJXT5Hfn1ratNDQNrb2fYr05qGX9h2Y0iXi
4DucrDL8pvfqEF7Ht7oWSYrhlp82LFZBLla8LRALZ6xpJ6Gh24t0I+wzaNks6Jl4
rQqjC+XfjQPjPVK9uuhad4nC/NNUFreWeGqBkHjM+cwzfoYM0Z2Qt085dqI/kwBb
MfLtYzkpsYU6/2Tat1Oz5q2PBM3hAnSrcaxtRxhQeWGV7Rl92xOb2RK/QFoVB4FK
ORzlgSuiuPBlOEgC+HlaIHdbOhNuyNnupAbHaAVtSHkip6wQFsuYwx669XtJDZlm
U+fc6RVkp4GQpkNMRmyd3HSwH43/1gSltwOuYsSyTAshTmYUH5/4YM/2iXnHLYLN
4yUuhYjUXM2Tld4yauTHAFwE6qZR6y0ZrTg1t2ZsPVsJvAo5P40HTlOmWGkooZ1r
w0j41Pt45tBZ/+ZVlTlt4aO+K8Xykso+BvpCpstjw8gHSC9nVKxkJLiIqUnOKqOA
625SxItBqbDudpxiUWKcgznjN7LRl+TH3sEJ3E8lCZe5Mo0yCL+Wv5OylqU8xdSo
XPVCAQ8Wr4mT0lFAG+zqVjHJ383kYiAzD45NNllYQKIVr0zA1AgkVZvnlPCtnBo+
BFvkzG72iv0JlHcGoGw1/0JGrn0FJ/uHPAYM+tGmF2VL2S8CFpz506oxCQrStApz
uPpyDwyBvTyEjgC1ciCqPEEzMtRV9jSwHWqQ5hgrQgzkxO1Hf2HC0JiOvdZ32RJl
QAi7ouvjnO5kFvxLXgqFOHvK5l7A/m2R/ikGFFhCsw/siX26T+iuZcbTURMtEWrg
iasBORSy8HBkuQ2OkDEcwyOGlNzLqrKpZuLvOsBHihFaE8DXgWYBVxlLGNrfAVKx
+GRRvOHr/U8+vFsep3Zgb3XD/XhFMgmhocK8TirlQwXycYu8qC2/KTt4bL5Ls2vh
uCvWt71T7oqfPcNl2K04YD+Jv+fsgqAqTILVzNi+NSJ/wPtDz0nrtD4V+88R1/sA
GFH+A+6mUUTJIZjjBTRCJ9n4QjZbq77OphMbpKbwYOxJPtudcujOpuHHDoSrY+PY
W9mxU3NKjCmXZeok6h49F9LPlA0fL6xjJLjIass4t/91wA1IX9n4w5HyQs91xM8W
vVknDzWiHVzjWBozgIT3/9k1MC1VjAHcdL6s8jFY+BCM3YJV8GV+RlshbPjNwXGA
k2ZPVgNhieOcGGX6VzXzb4S7GqC/7SWSThyTpwlMJnjpLh+6fgxHZOIXGLJYj3QN
Ri3BzTlTdMi9O/OHQP2fZbJGYm9weAudZ9y6kTq7CuNXAos0FKQpdij48Xdp6fAR
ww/2w+KHlYN8Hu2fqwTb0qjqhNNER+HdThXNwGY9EGR9/LwWibqBmYOv6qDBu+rs
9IVGw6n+hbretUZI5bRffbGCeDC7DbM8+6vAPDJ5uaOTeiFc+fWsDrw3O1EvcSzA
XPfiqVGP8jQLE1iF9P9/ZIZoYuBQqQVlntkJEb8RHu4omathuJJZsyzA6Pqz57XQ
wKycASePriZKKgz5HNyQOe+FL2bZzyXoOmO52en7UTTJAxSV+7z/j/evsA6viTbQ
pfrjzoRAraHz1PkIerdcFzCW9cxtCVCvGDYXTF758I9l2S/XMz4vJP1fHW+GOQt0
VPvOqt8HIYhLDZR3IhByTY4ihK01OBfblhqXE9ubxfQw7uwogALE6oHYWJAKqFUe
bcvKSkM4a3mE/k77MuzPxpEaVYBPZA0l0uBLilVArsm3YEZyPDaI7Id9EARiDcnd
uH2nnJUzfTHrIUX/M2uryM6RDemk+qvCZDGCFI2H9i7OwbbUWeMQCt2H1M0S3uat
IYzG9oCy/7ppfnRaJzdww+jZnjVfFJX2OLprGiUAvHXU1k10QjZKVykcGkhJ4HYW
NJuqoCCfggROxohUZS1Sr80ZdIVndnzn1gBxjBdqr5q5tsyX9IZqlsy7Mp7rKqsJ
p3b9ypYjrMDFYMsLiZWbLKEImvOnrKgcPwYZJnU2ZjKh4ckRsjMGbbZHZ82qxeaX
drC04IEFo9/19Vo4UMs8o0RSo343RYpMw0cJlPIvpZqaiYBOM41gqoXzchuowI9Z
ixq9JUBPxCX8uCE75E7Lux+TAL4eW7ymAWNw+NW+gwbaEDvZZcfqKZPPIEZHvK9r
ixcXQ4R5HxHSnnSVS1Oi0EcqQbQ81SXwJwKaXim6EeTATSMnWBuvKXPK/3EiaZFF
BNHQGbWBAwcHqUbhLji+hO6dOdFAqQHzIyvABLcRQ2XsR8zV6NMd74XEB7d6st2l
Ob9OCDQq/yNPvFK7uC+7TwvP51S4PFUFi4G5UqoaxqPlEKUCUm7skZ3eL8TZAfih
ms+IRnvQlC+ba3L49musczyWO2jtt68pw0BNg0uSY6TqaAjkyoIFh7DyqPYdkB68
hhgT8YpIK7isOpQVzn+f4I5sxwYcNYLZx/r4uJ78JN7a03GQdNSNq+GpoYyiOZpV
W8luzUOrMS5LYpPAgSGqX5vwGFajlmNdzuE3XwM+yU/9jCXkmudjYseLyTkkAb4T
cQGXWaEdm5e9Qw+HYPeyvT7XOEbQCPqUm37Mqg3VVpgRCJAG4q6JW8sGdwqzwXLk
dHl+ALchQG557ISY7Y6N01hmlYlJhljEaeH1gIO6YcDwYDo/MS4LrpCaIerT57VX
2q9sbNcxjOL2gpKXDTM5lL10pO0kOd5porG8+ngyHs7Dylt00ABqfMktD9ckzOFc
pLg44xT4OEXp9SI4f1vrHCnspmqGO3iDRu83IytruU8uBzNLToA0UgqKHBqs1+c4
yUsDdgDaUbjOCQ5Q2UnBiVtXVbDnE86KzTBS5tpDN0UPoolFHABqkH1yZiN9AzdJ
7LAEYY4oi+AYCEVAUH2TKYHZ5nmfyuJvV6GaEh9m2PqysRA0QeDU+LRVEDNrfqG8
aygObH+rVaeP2w4wiCK03nTqU5ZgoJpu54j+ePZ9hjU/TtQf+l44fN/vGp/ZzvCT
zV094I4uonwZ5/1fkSyDEgq6bpX37DYaA5qr1RbNWvG+25J+01Kq5Jqao7xYy6OP
hT+9HiqJuOZypug/SMSw7c9i4gjX0UnQ+gUm72hCoSvBq3KLu+F2uk4t/CALj4jR
lzp3ZNSON/5Vd2CPiME2z+J+sBrKXVb1F64S9+VUCR5IUg6mk6ZAlLqPZD042WmN
ES8zhefKEB5NN8qo8C4j3OCD/GMADXPS0mLRk5srDn/DD4fqk5OhdiureTv8MFwV
n2K3AlOF0ku82ymnmx7yd/AF2CValQBasoDWRFx9jNTr9C1zafEqMa/F43EVam/J
yGXggJpbe1sc3OJ5u6hU7AEWIKEDQ5wnBJ+KzUTZ0nIAYkLwFJi1Ge03YVvPBSj2
vo5eaexpxCvQUIg9GZFjxEvzQeAMH8jKq/oGRflGnKKrvr4HljeVcEw1X57bjrWr
9gKYcoKDXnsVbo6CGfoy3nNUAJ5aftWxecuQUATrgAvHFJMz2w05QhRvkHDSOMdg
W1146arVpJIJ3Mp9whxT3zrTHgyEVP2cx2CZk+nhHqEA98uhMxdukLjHjr6Ut/pF
cm4+kMeBPbtD2JW2twKeLQ/+hSfmPHFidf6BCL6BPr2vSING2IiRRmUIGIybSPjr
PRjAM2sFNzbnXKyAnMCSahXYe+SWCXmhTRH/7OPvHstqSwhl1mnF50EFH6DfrpMK
YQrZwMicZT3frVBeIOz5qhJ17gur2ABeFBaadQu4vmbopt2M3YGELma4PZisL26j
3DZ3kjAst58KHaR+qKfh0SYuBy7Rr1BwbrHXkcHGWutiy+pUY/BQPbT+tX9Uj/d4
nMyEgt47Gpm6rXjhNDt2sR/A6WDm4Bz5h03kNjQ0dG0ehsaVbGbvhgu/sGCpbPD9
g62PFRX5lxVJBLimX76jIRnJlNCrwFKXXuGWlLUhhuJP9AEhPB3rAVgKofnINROg
VOVdnMZoLDprhYjwdATLNJQbYY6VBhHmFoBkVXirMkxPMIwKTNyT2C2P9vgft5V+
AVVVuxfFBw8oL+3KYqO4qcQFBBKgT/lRI/It4Dc2HZcZJ9O2jc1Fbe3jqPYnN9Gi
i9Gi//9L1RT8S7hf959QUfSntcNSgSDlAWuP4gBTpOmHhivEPEUTZxen2VW3L2kI
OJLlg7s/xznmUpV5SQfuWtrrHqQbBAmMgnV7w08PoBng3cq+S7HoRsjQi8IyKhEc
Bm/RA1fUJvRqF0c5R2K4KVFf39oBwpY4GSBDxa9l75YajmgnUkNmO/dmpthvqqE3
ybX9KW3vYc1ZuzkMOAhsQbVV/MgpZzIgR+pB9pJxiL75fzD3cwzUkRMZQvW2lPIY
YneEf/Cz+rZmcsxHLm6eXfmRfMXQwkIdM/70YGCuZJj2SFtxfFQjEcTjLwsVA6H3
rZHZNT2QzSb4aC7/agK5+IV8MFFT9ohLtZPicf3HnAzFlwPws0DttAnWgEY5tr0i
9ks5NqjtNUol9VXgxHO6Q7ETzf+7go+Vkcw4lPLpqNmDXBpdwXqlaFYFF6csQRLb
ZXolHHGEz771Hq+TmbPPfX8govM+h/p5Q1FA6M3WxV/Suu06PvipfUZs4THjxfzI
iQfDQkpt4YyffVhEE1/ZoWKtNPRr8bEOMAHG+Ely4CNIGR4Q3GmSynSy2EIGVuYf
7xSrR9lWif7g44Kr8lx9abroPVPsGYE9EbNb4La4NIOkcQqhsn5fqdamGWgXRj0N
FKPH4WrTylGEa+96HlCG0fHo6G1V1RxVS2N8d2AfO7I6aeQIaNkqNPm6+MpnvZmT
FGJ9kLWsI0ZbtMQFP+ZLQAcme9YCCgaswPpBk4kJ+4y8BVyX20+EF7KUjrzlzSYE
q0joyuu1RZ3OzKY7dvDcTSeCoufavY/8Mfj+UV8lkpJFaUahItuPQUmzNZ/Fgxfc
cnIs0nfcAyO3y4+3ZflPC+yHL4RZzZFemulCTSEgCEYugrxWphbSx6SprH6zLqgb
yWticH4J0GT1PauFGYGojc7XHuG4i2q69BvYpvnhO6+P7jW0q543Efgd00iO+R/q
4dOUiTVcQMn/dq/a0GicTzj/u42HBc+++SzA58wREXkm01o5SPbl+Gz8zTH+kyEO
BPyBdxeLfeDdrsvdg7JXn33WNP+i6aVCAXCbu1pTUvdD8LCHib4e0cr6eMU8CydJ
SR3FCMPzugTjsfV/GltgdP9UYVeTmLka8yCW4XNFn6MdSUNop88FMTeva8c92Avb
4ZFst4voPTb1gt9LtHedhX2Yvo7x3I+xx0d4qD+MvYFx/hGASC2BsF+yZpIqM+C0
V+GTWo1LFLiLuh3eYC3D5tmev0N7H3d+UtMOVXnSi4TDvyZBe4e2EUDV7Wx9ioUn
lnvGdm0R6KcRKQTj7L8c8nS2Ami3Cfk6okUCV/B9qVjgrWcy+JZM4eeZxpE+Vx6P
Me2OfOCX7p+otqYkct+pDtU8FJuD6mJPAsNlB0D1GM14ME5cK4gnGKkY06ZVrOAl
9EBXk2sMBjVOnE9QE5l61czOUfi29Vi9QbP3Ld+Zm9YCfkP9J2J2Y7CiXw9wEab6
gILF1tteZQ9T3ELhWE7ssh6efO2y4kcJvIoEF+f6McMahx5GrW9OYpewuuKnzIT5
UrBflrSAgJ6FfdIhbFeAO/XAaNTMzy3mU/b/EKH2xK9EcIpqbQPmrH9c9zGaxA2X
p9y2uDKaioyRD66hZJFuT3ypVV1TuAEZ4Ca4Zzt3PaVUNKocmKvBLTb/hCQR4p1j
/ZjIETWDvYUgtuyFFL4p/tEUEWaTWkjXZJJTpJ+gg5U45vAhlGm/rHnKHxffT7ny
we1X0ok1iCKD9t11/nlMa+AIUHq8DCY9reSL0JCHin2THn440J+tfyLTyY1A3us1
7W9pkbruM/i9ihnCw5MSbyEH8tS+KN2znfR5q8uvBqDYKBIut97pGTlOzoE0fFj3
AFnC15pbdv1ny3gY9s6MEIQMx6qh6u4Mof0Cz2YxpY+YlnVjx4Z6ZxZ5lydkjF/Q
w9v9EvD0ZCBoRM9pJnOf7UiZvukLJeCSnnyjbqB3kAExUiHr1/CQR9OEl0QeVF4+
3NmrkAT/fNEZ4UYALuDZeM2/UIHSUAPe9jEzxukDDcAZA6TcQg6dCJxNR/DJgfbD
RvN8Piaf+kvCN0SDv2JhBOqqfI4kU01CySp+9qqVPhH+Wjk470/837nr8FPfGgRJ
TGS7PDeGR6xNKmpOM5a87TmNquVc8hppKhtE7ZWVUu7X1iNlyDDHimkYVubHvC/D
PQkGBU8d1mnqs2LZZQHEdHbVF/gwfnGV1JnVzRqbL6qOlTgo7au+dNJP7cVkq/vb
nVvZk4+7iXiAFj5znM9XWH3MN7sACBqrn0+2BstVlTsR5517qCwkz/YU9hebu2sP
4ZXn4/f2yDQ1gOCRAbitq99zEa9Zmu/f+corWT88npcpx14rOn2RxSGcntUrMKxx
MBh18Q+cQAUyxT9NnZiiNE2gnitEXuhV1olaJ/ZCtHc60HgH8zQS6uGjvtgjAUnp
N65s9Rn57bM5zEP6R/YJSGDowHp+NOclb4EoqHQRIVjqbMcMrs6BF1XbZUv2430Y
HtABoWvVGm/ahgCfAsZlL/hm4SomFwly2IEX43SmEnlFayhw2ZNdcD2rh8/qb0wT
uj67+CLSHunZqcXmcJxSEPHV3K98Za3z69/T2BbdcNfWjHttR91MNq6Wz9sg09jf
60yO0ESBF+16Kv6wIXPsV1rOrHAHLtPhMTBikJ/Q5+COA0ejmxUo5BgkqS6TXhtc
3aTuE+KQjl7OMGsMG4Kp6wK66d+CUSHEohBnFzix8JuaRlNpMfawCSFwLrZIz4bb
PAULzQCjauTLLHPBp/1UWUvoTudaoxuzAQllzjO63rAQ9If7mnhXq1aBBn1Fen2E
12XRmNV/jG3FZWH9/2PmOANAmr8ZDolQXT26EN+GulyCJxEBtGOo0MVnOj4KnyvH
daluGCzOsOi/J4hJLeZVdNPVqW058+fpoeaMo8fC5ewa7NGvOHLKWeFOwr9q6obE
gPBtcsLP+n6+YHj2n5N5y4U/Re747NyWlvvBp36LRfCwSlF8zeLJJQnQ4O9ZFuhg
0kz334zDm9KfO0df3R6LD5X0lDfLU+w49hzG62kR7++E0IQBd4neSUpNun9eAhx3
MSydXf0jRsltU9VAya6X9sYReSIKOMMCMUOMF17dq/FSdEXrAAPfMcXX9rVS4qLX
t5RXwPdBiJXIP0r3LKa9HztiDVKJMIqaKixDsvVw4SkU2/QquBGgVaPgzW9nQatD
j8f/w4z28wnzyB6Xebx8JSvgT3nK7esjNRWLCpmUzrn9qUUaToshCPnOa2gaBIYx
GZLK/D/C2c4MlCulMKUqinfNaZSFmWYXGj94FQmoKjOMn8fbQ671Q5Q6NP5Ctrav
0D9s5E7W9davY8mQTZk4GvOZZf2bpwdlw99J5eMA6rpAEm7exZ7ACNmQhfXaqB3d
sd2ddRaD9ZJAkW6W/AN1mRhM/EJqCKSHN2pJgRYm9qRoBwctO03rpoMXOpUH4PP0
D+BX+OTexEIsqKOBfFiZ+Ua/cQ9SaLtA8PPqVIEKCliTnv4urCElHQNLGh7CmumP
WWPPQENpjWTU00DgpwYcB40kcSfE9CSqoeVS7u0CLgPVqtpkurArsCHA3gLAR6Yc
XpgzI7PRjZkQm0pQ9Byp/wvLnr91+1PFxj6mC6JPu7N9BgUcBvm8UH1WNaOqb/YQ
BAKyazW9a8/RerGPskinJrNZ1fki/t/5H/BDL0ZiMQSugQwUOa1cDN/BJohju8Ct
eKehdvbPM3FZgybpLAcePG7yhQXPT+DR5HA/Guk8t65kQXzQ2VUqvPT82ABgpk7C
rPA/nwD/YKZZiSncfGdHuMoKh+fjarTJ33IDQY8zAxmg9p61+PuVe1KV3RkBAQ+v
bmt2dhm8fRS/8+/BWPEpEOEnr1Zi0TAHMFNsvxIN5bJyKBJAco2MeBZg2qfNFiD+
X5x2MMUvkOCubvz+FRgJrSZjD5Xxuv5Yu/gIOYkDDp6pDDSUKICbTOP68uk4eNvM
S1m5wwLbhJBfmXP55sQdjlHNKlAPtuGj16soG7a4AzOCiD4wKuEjbXhy5qa2iSHF
CYqhqdrdInLxrUA9sJ1Ad7EaIorCmBaldi3mj/L8x2vr20RomuLlSrAwX1ki/2I4
obpvpGaI9oj/FVkbRKL1SaVC+lUsa4+rIH7zNQ/iMO+5KJ8QQ13IAsrPpuM5DD9Z
aimCOWxt9q7lVgzWSHex6YAf39DAHeupRxTuIy4PQIIB4hFvXRCii/FZFhS37ISP
1rIFau+sKzEEtK39Q9aOchzZFguexG6eJh4gcGndJwxMYH3TFTOZrqQ3xFnnuisz
qMc0Ac4EeKjoxgcc0UVHZJQdq8wycVTbtbK0EQonk4LU/VY2Nix7daIwmrI91iuN
h3Qe6DHkcyf4apLy2YCMGrVY1teX2tBYShMOUT4jW1TVmlhPOOe7vHLBAdGunvnx
pBMJsaFWtU1o9gRWE39p9q1Vv0fI0M4+J4iSkXi4mQ+aOoozTFuScUzlgMeef1TE
kGkVsqh8NGBJ3rVJ28NipCPgpUS70XgqnEW+QH/mT2CFw++evhEysgsjTVEHexON
l4L2CLXswvH5Q3aFmQqRwc1nJ1mzuH01yOFjA2PDKrdpEgmysfiMpoosBOVnvz2p
afiUnkEIDx9vclSdYCkkx8NmX4eQmjNMPRHgGdNNDDofiQKXcH1kWawMGXInhZwE
oF7/DlYMH5Uqlr+O2XORI5q+medQjdJwxXwdPwOAWpaBr/68gh1iS9PJT+2iIwg+
rfgmwMv2NCsLMmybG20HhjBB0oCLblTOzqQvdwwRRWW0uyMknj0GwYilhP4Ou3Fs
SZrNT1VrmN0SDLVgJh9+qFHD/TfpKLr8lVsCoXYSTwS6ZfCLRz+fZ84Y8MwZ4i9H
AmOqUBQ4cjXpKAy2X+QTuR134yk8XWI4Vnwka/v5AkxoffmTk6Hvb3TYc7mDhk8j
bVrtKv6c7FHLuUfCq2EZmq7BRs1E/6TCjBFVsitRUSblyv1zpOpfg0Y8WHM6Oyt9
8OHg6+70kIRm/y99lQI0BiZEQ9J5Y1y879ZG0K6KAAh6S0QZabLl2k6DLOE1snZR
Wwp0oRiDxRErgff7BYXoQj5Dx19iV4LbyWELhJ5o1iERt5jytwMEwKipWyHGuG5x
/FyHwzBcMdmkwT7xu+wiehSCJG0MMUbc8XC/FXMGe3wk7gMg8bkRhwhVCMszknD1
PDIuZQU9ns/NO/4+OX0KedyLC+4PA4BEMJS4vUFAV46dAUr6YB/dfBW7IGh9Qf0Q
D4HCrLkoHXr0FE9EEAo7ELExZdxDt9B11KOWjOdV+2wus2ExqRqUxgLHwnTdlA1K
vZHfb7JclwfMGKAkdTr0+iWAdeLH6vpGMeT2vODMIb1qhR4PFmplzkGKY1J8+BYL
v8vjjDxNkaRYd3BFNQMjs1U741nyVATC0pKnUmu1rWKPU2uvVwyfu4cOKrTzuZH9
OOPmePwZx1O3Ubie/yC1iW6rv280zReV0c/OV07QNm342DUM3mmXsUEouuVUHh1j
eC4kfF/uXQglnOali2Lli9YyIAP089ROCQQAKdN8SBAvg9nMm54lISLDP9sBw1Lm
d/IDq8DSv7BTPfqSVnHa0D0mHf6dr5MRWA/XNB16xfsHkb87TXV9VjbfX4Fr7GWG
VmkddJ7YEE6Re4tAG3zUuN30ejlBGGhYrURItYHpqbZDoJO2SKbsxaVRIpIdzwv9
9nIZgnPwqvdxHGgUEHE2TL7jwbz3DtySiJaC5kdgTvlQ4peEtq7jQzmnyuovTRJM
a32qxv3qKhvFPfazSfYr++jA65JeIRXdaySgyl7E0xJl/adLXS7P+IyGv05tOtu/
H3ktAWJRdCe5yxWsN6z2Y6MrN8uuR0s/cRRlQAImS1HmBiPKreOv+Zn8Pn13wYh/
oA62DmN3j9rJtUF7aOrMnL+kLfDj6SHVDyukoPp4y0RslkLxSx5jV+6AImM+PMC0
4np8P4T73eJmP1SQ6zllmEpfRLmRRkAbI5lxpGXXuw1CTR9oR7D9O0eL1E/XDDg5
J6nWg69IFjY3Hq6303TFJEH2I+AbtFiBaQ8Id9p1c4HuapYQUb8VROryw2x8c6sK
Drp5FCbhI7/aWYnW68sC8N27RkHgGyiIUfTvaApRLpL9Jiy9XlXq6is+ZT3fIcpW
1wh2BKLKOfw13/fMJWAnHhAg4IRHk09VjdbhU/BKXfOWt5LYpiozAm8rJ/MncE1Y
uMsVmLdBzdwx4ZNIWYwjA9ieCQWRRZJrwYYgRY7VfFntIWATgxYA18J/DnU4c4wN
U5x/sUfEfqsissBiY5KjvJBqDVQtjx3F3DdYwzo66Oh28BnUQTeVNEdgyt+uE1rT
B+4vxrc16vCecOuZZlW3zuC1YFAt5Tw5zXpONl5/yGQ/xFd/57uP5tt4e9F8blwI
T2Fxri8PPZ7pLWfOwkR+20tBscq2U441Vi/1M+CG65cKT5JMg2RBZ6lsz3EE554C
lbDShUzUMJTqXHcuCOre+Je3djX1gjRSzAM8x3HGGB6Z3tZydufrpfAbbR8WtTU+
S72tHu+Sa4U8A8tiY1+mLUlgGgZX1WL5ecWGXTolw3KbWi5TrIjp4EECYEc+8Sze
3CZpzaKy8gopW8QKhdh6HL3Kfz+OpRhHqI5obVoTCSV3dd6IbbEVu1znT/tTRZ5R
waSeTsBkj3MKni8vwtjCKGDUaYh5OuIfqnYrBv8fgWrybrc+QhGw8NjZ7GkGtLlG
/SlzhUSdkcjZj4J+WKZtFFdGhgdRdPfdQIJQQNr59Wd2hrn3ZDsxLXXuN5G5eEDU
/5/DkGD+SrcRt/20Q6ky0H+O0hE1v0VBhS8WJe2sdYLTUVZndfbCw6OPv2OVnHYZ
bvRqyqwE0rL8uzGIphfrRXp74XAXFMm7kNPhbsjHycMftons+DyumMkwLFtT7cB6
D1ZVMjyJcftyl0JHm7vK4i0cAsO/U7FsI87W56yLaN5yg1zw0GZRFCEJeqx6n8OD
y5oXBuWEPiAkVu8tsCopAJS+zIm4eVMZ3x2RKy/lSOxbIbMaYXwOkph9xGAudHv2
jCL3kPWQdIov2sqUAeIEbnBmGAsc4iI+Se2K2rbNzJDazX1/fd11vUc61N0HX/Zz
PPUEnsVNRLkiTu7zpEu/nYpIF/o0LIDMQoJQ8tcBCrnlHUFxJ7670EzMgfL8vMkH
wztn3FWuKUZASguF710y4Lp2YxPkJKRg3EdzAGN/QdfrxQ4rU0Itba49y/X0Me00
bh53eySMk9eV3uiKucNSF8A8/K1NuEcqwJPtZNKDxza6IVbY26+O7WZicw51J6cj
wS3x9U5YIv4SA1zKNHmKXwsrEg6IqRTTTolbK0/85CBuV73IZu2vFEiw8gJcIXzQ
EF3vdYRuI3kyRcwI55kLRie+acWPcgiOxyYJmBBFxwe6ZEM7lDYoIHvDenunb9FH
WHmepMoPdJqQQAhZWSbjcF/tunV84Jl5nhOAgemVizDh6q2FphjLC+zJVvElnU2W
2CKjFfIowxy6wTdjO0c5ZECERCatt2LFj3FInoN++dSBI2Fo9hECs+VuUVBhDZzO
Kkatw7KYJl28aKoM4/qCOETU9NJAH8Q+M7dCWED/+SzOb00s6gtDMPvNXbgkDzGF
BWkiZcjN+5mNUsPuzr9nuFyyQvdjShxDaPYIRTN+xq2B/4aF6VGrGyM1JGPdnuap
f4sSvzTAahU65VPyaLvANvMoEnaYOaXb6I5eD6U5BNwqnlELx2IYlJbpj9CiwXSq
rZ9Jg2veTZZBLeMj5XUVFH33pMG8wnSSQ+TzmEtWlzkxg/nLRYEE6rdZL4pzwqZD
KN9SyyzCgBYsgCpF8HMEmAmsPh9EUlFGR3LQQfrgl8WxMTx6aLPcglc7nc+2v717
TZarYkVu2PkRHWd/7MV4ybVviYxP1kdbiyp1fElZ8vka5uBWc+Lv0iJyI/3+Xnjg
VvwyMfd4HtE7AYQdP60UfCp99zbUzav9Hnw94LLBKSjqq5XeRrTnzX28OtNKJny5
rInRvXcJH5a5/lgzKFSPB0+iIxFvDXCKFEd/WP1nlfQaKhLMi3nPFaCf5A7442+r
OP+TTMJiwo8SIkhWtLSOuhDnuJs2Dj2Rll5TTh6Q8GUHP3oNgvfCaFt1nGazwx9G
95FSxKqusoQciX9ejC7NupF3vQfUq5+S0xHpnzGHoqXNxu02eSp6kvbFDueY/a98
7YuG8S1tmWWnt2NIfHKYAR46NRvT7e/VaXUbWCRYIjmBFX6PA+MMoW5Y2/zGgC41
Zna+cWdPPO6IlPEywY/u4TiPUmM7v1fbWYmzgM2eJsM5DKf9CnEw0810iovu1BKc
goOg8VCA8V9EygWD7eSml0bfZsdvd+xRIWfF/8wcGDDn24IAi+f6yxk1g++IxSmX
8ilc03zkiXCcJtla7dUlDbb+q3yZT+V/mjaLweNayKOuwi7MIZoeGc5FttgIlWaa
iSVikyFzHT/z06N9V+RKmdUtp6QdU53EfrfNvRBAKKWqIYB04ie4CbdV7nIYheeB
8AFWFSPKuWnpoyE2sSVInOn3m9taznJxcGnRxRcj5iZI56AhomQMesT/7cyySJAk
M4F+lI2ZWVYbJpF8L1h4aLoJFkvLAblQt2J8YeUqds4fUgBFnc1PCORJ5eTtIeuj
cCpNwHqWZQLQrFcdbmTNpGoZcJXM3LLMdK8Nf7qNeArcOGoTaay0pyfbinMgS87O
WaBulFhPxidD63J2kKJUz93yXO/cvuaac507Z0KoxGwi1uC3amrPqBEjz0ejGFti
DwcrlpFbT2HUFJjtIR+O5xM2pgCurZxZ3wEXFNAFApnutQi7Qhc8cJh6NdsjiScJ
ZC51F2njTgyvcpCrrl8vi64N5MWdx2jeBOz8XtWYkDX64+7zbGvB6a1XIGrMhvMW
bMuQFpd8bw+XTNg5nulpR4G3d7K5p09WMfOOJo6ngbC6RTzPTsySJaW6gdr0h78X
PN8MvYrDBjPmmTsUQ/tNdAVu8pBLcYUlG0OEJj6ivUPoTYEhc1JymyZZN2jmbNb3
F+4FOFDTiJtXyDFf1Y6UEDDbpG6IX/gdg4yJFFKlipr8eObBwFxjs5KeRdA8hVp3
FkVcEoYi2UXOuf67Wtwbw6PmjMvJwS76sKVFDNOnDEMPPTMFZH8OF//yc3A/G8eH
53Am6joD4399AO3BBjAxJcVAzhnDecpFd5j/VqKHJF8DTyOH7suF8gozmd7jOeNl
RH6xOUh0pElAW2BE1ai6qQFI78cBEF0O7anmrjUqDCn4PCma2hz1xpj+h7IKwsNB
Luuqyf28MX2vN/R8Gx/wMwJ7J63lZ/8ToAOiGtzLSK4Iutt8siinEUsGLANrCacp
RFiJfdU9faCEFzhe42zTLFWsE3SwAcgEdFHoUcBedxw33DGzSlfejv5+4JxlPph7
RemUA95FMf3Bm3c67r5gq8hd/K9NPmV4IuBUpMeV41/e6UOco0qz3dIG/SGVWRan
TJCt2tkCNCRWHvxlU9tlcRNrDKtdGRdx9PagLDLKWy6JDJSkNy2JxCrwpmZ2Ootv
aAvdRKB0z3bSjB58GNoS0oBtgZuRG4YiHhJr4HZPGsCgu9f/ZNaJACdE8z/ubE0v
I/yg/Ip+Cni+D+AusHf/7a4V791KjNzs+BAfkgVo/u4geLCn0q3BZsyVVwCG77VT
HuUaT+l9aiTXV6GSyLwrVWP5vMp6Tx7tFhwWtTos+/DQkWWdzqSbxDmJL0iB18Sg
WdhdpS0MpzYvd/jDM3NrEv0YL1wEoYn2IP81vBk5jBCt8TUVF65P4IxQdt1tRgjO
qeGrvdrdOv7x4+ek9UDnRvCu8q/Zqe+CyXt+OPofWy2yfMdXA6HeIxnrsVHdE0cJ
Upq6QtSGLQjoaxB2xLp74SHi9ZPKPVp4WQnoV9+XolvTV6rbpboex+5TlgUXTM4A
p1kBbFoy98I3mpVJu/KxaDy0189a00mjHYMTvrWyDnbheVETsKLycLCnSKsvIn6K
OzAo13UhR+S8hjX7/yNsky/+H/ro2/jBXHYNdfzI3gbAVCKe7C6nLrB2lKkTXadb
j9wHlkvjUrn6yKgdddA4uiJJyicv/fs9HEHkCm/AuIfTgSwxMmdBfwU+B3s5+02z
ykz7GfGa+vVmxXT8Rf/Wpn+5H2nhf31kXF5SBqFS+mUp/hFWEVHi892TYdZ2+pmZ
XOtZk77rtTiptS8fVHYaaEjrdh0ox3FQTu13Nj6m4ReN7IeXaA+COEcXIWm5FwXK
vuRCPeROCoV1Xm4aEkAcI7ZpG30cky43kWzd9ocO63+PDZpHwyHvSHr2GzBdR2pE
7xM0NnUhpDLjEsTi+xnABUYdM+cBDODcXzkVlTnVSOU/ESUCNz8UI9ZJ+FCHfwYW
MdivrruNmP+Z+cAaj9TMIie+wFIBzQoG1SE/G3dHxgmz1dBA24hBkancxYLS63Xw
cPu9vyUlAexEaSsMpN15QO9GYkf0VFwiqkqPApvMBM6T4Yj23Ltw6hJouM685yDb
mSYEr+jgvQDKTn56d5Sq0BJSlV881yRREAbFYn1Zcit8Fl7LRTWvpzGAWk/sgjky
LSYo4c4gcnYt9qrFJSaoX2UtXzG1os9dShNQCAB17UkX7p0lK8DgkbmtAqt8niWc
SzFDRW9XkuNlDDnXHK3A63H2Pu5vM0+jqf/BEIn5NbJbZ72sczaSmMSn2oBOljC+
fe7RK0Zhl72MJj/BNth2CNAywTGk5JzPVq71Mh71hykenw2VUuY/Y73sGU1OqBrv
j0LghLccz4AEtaH8hJBN4fAd7T0gU9tHl2kRYRJDXidYblLd/tONmhBMR54aZpJC
ycflSDYkRAyhnbrAz58zqSByum9wvy7D7t/jO+U8QsMgDJJS+1fMw0palWn5hpEI
82PZwREFxNUXmD9OTymmibcEQ3kDCY/sWT3gA25ZYFz9Uo7tecaQHNdSenKVb2Ez
EsxlS56c0yTO3kubsr9hGsRKHHjUzwNgfNXYmJbGTF67ZPmdiOQWXiBuISBX1Cgy
hGecAjCgzPLauuGppyohFP85sCkfKS6Ktyi2F+v4oB2u1AXJn00QdSRkds55BZi6
awTOw8VLDwacZa1FteUMG2nysdis62BXxu+JYBOnP2srXQGHlhT/kRrIGW0X/0G1
6uGX+vZAvdAO+I+ag2SEJTMO7ZOuIgGyfEyKH5iP7OnkBGUawMvPD2rHiaPmA3rd
rR4hDkKkaJXMlo+5u/D7+VXv9vmiSVftNJJLIb7qYjGLeNRQ5MoFcwQfhklBy6yU
bltlj979+VVxpAp/WnhwZuJpDtjEvAF1KLSfic57YGQn7MTOuMDTzkMDGErKYOBt
epbpV3odLu9dhSjxpzzeZef6difrLQlilWtr4IzaKqWbK6/K7tVCbhw8rXmlztqr
kbIcF0kbkKRp3fUFVokOjT8V0UwDHeSq0uRtqg8FOlPWRce62IMq02UGtzBvi1/I
1ZQYZPbDYFlJM8V0kVRQTU6FbG+r7A/fHPUCNKIBgaIvfZTB3AdjRchqB9K/rt62
XCPEaBsD/JURRFkQ7IXJ5/5RBVSDConqtkEi/m9WUs/PQQglXPLkNdffWNmG9eGy
i5gn+F/ElkdJuMw6lPHO8wn1fLzXgATmHyiko7kfGWrE7AUhBWzUWNHrilzwZKCE
3uwQZAdEdR/cBGsFGBkjwIo9lIqFds75YKaoKaOvxsqHS8bnrEx0rIvyOKDN33Hn
nCkjFLovPwrttkhzwBYcbXZqR+UBGVz1VU4cz5j/7rWUVvypp9+OncQKdfoadP+m
iXP35cnFH6x6k+IfziFMeYQfqUyqMblky+5lN2U20/B8FYZu8fgjdSxC2TXPb9sS
Ds5vp8ZjTucMIt/KE1yLwl89pI17GVITKFgs3LkvA5IW2o0+4aPsuGOIxeLv97sY
tkHGDurOI8n/1GuKSkigGqxl500D1EP4qz3DqHG68XcN8XNEYACk2K2QKkF7C1oN
1zCsdUyVkseFRAkQm8TZfy+g8VVCnWsr/kS9EDnJDUZgllfhsSGf0eCyU0feWHYd
T2z/HsfJIQdYnWq7GDArj2ukxlvgWIi9FzPuqLbT3yzIEKOFEwJKgledksCuja6I
4ARcQUPUetd8Lr3yvd0AMCXIsnnJPzFIHNM1UFkkvx3JCBo+l6rsekauRIUarnF+
BLoxpm/AxUJEj2smSMX8QzR7sFnWzh74wIxz5TfewAl6t2+hpDfQRl7/lmWj6/wJ
hzGXCzNgpOuyUGx14/bD/4vANwv+wlifvUq/rH7dK/tRz/txNYi3YeF+YF/MQ/i6
75n4FDwKhEID0KhR9ZQQVMrlqiVxzA1xflfIt96fJAX6OrbTc8FDiP8af+GPcP4o
lk/P7LD4eX0wUo88MNZO40lsunMWvTpFxtRXlmy+BBeIoOJ/lxKgCq9xn1TgMou2
tWObhlVlcKdUJPgUIMonW+Au9VVSt8Q7i55bqj76eMiZOgryGGw9n7gm1EYZ+SL7
0xPTX8qn4+NIowe7VIGJffHtazIAE/nBU+CxJVY2i2hq5WAHTfiatwVI/2pTiqka
3Gwkbly2l+aAddMiG0gJQzElKEUGw4bfDVHfZeMejBCwPPsuxR7cTOtG4OswsTb6
1ogKLDKmBlmtDPi5uza8Wi9eIW4Hcka3V/rK37pJaqHEyUaTuQbAMTHSWI0g4HDx
Ol5OvmphGYoVKASnAZeAOTFzQniY81GyMMnIZ2KSwu3gC2N3CoQRv6uoJqHeLaJF
lze6N8uhpuNt1SsBV8zhwNZm2eemTfmJeTlB46m69q0O2bWEdUoJAFVDkYa683Hs
CRdu73H7FIW2F052rW/E6LGOqnbdm+KGlKQq7Dwdl4wRBCYQbOgzN9DqjG1TTSRY
dZqhJtTCe+Pp6Fl7JZdE0Guq9I8gBHCRHRbDSObyw5kqkGZEqGU6HNoEsLiwcGEe
e7uzNSi8r2n4hAuy3IbUcLHlh3mNYcEkB94Gho9Od/fwFxDOVYat1KfLL7UPRgNi
5dNyZtTTJJBsOK66tUINWxL1uQFut0vo3D3+iqYGGQXkH0OhkerqjLQoVlW85QTK
Vt3uQt5ysnCLSNTCPh9wS1VSlfQRmT/obqoaaAuKiNbBZvyIuzXAivOzap1J9ZBp
mw3NTTrTXr+nDzAD32n2AUAL0h3T3kJaoQkqGRJcN2N/MSE9Jx1DvTFzEN3yyzKU
TpSruZB1YWxOrhA0Wxw5aCmPm9IT2iPy7/fdt9WsO5LbyLIDjNuRhaeMILNnrXER
xunUrf0qazkTrliio2UnyfI/KYy51pePYCcnJbTEIz0O+iPBbS6WaY00CbV+oJYy
p0NDI1800RssJIuFEj5hpH6ozmIFTdLa+1+vQkYZ5FmSZV6SwYImjXAMMrcLHdOn
C9xhvFvQRIZn/ujiaTovlVTdFdyqF0Uqh3AaLtlkFMENKCSba615M6TiFlrJFudA
opf1htszeeyI9D0lkYAPuj5szhDSh+NxXsvet/xDW24Yq9aoFZbHEF0Kz5PDBS0V
MBAx1D1JutHD6D4bhcN71fX7/kxSvUWsCtpsTH1gHn+TUYKlUbrpNs+u+OTAvRSY
N2sTl4cE3wTFWYbA2W3bbnhEb5dLD8U0sqVkWgQtCtBC/xlMd5mLK+EUpAGRJahD
a+IA/PdHclPA+D5WcAL7WMEdhnv47n9CM8ue+vUI9NHeqrLi5urlN+iVTuVP2uqe
Xm/w+Kr8sGykaC5mtjf/osfskfeYXT7f97zDoVH1RNRgVJ3B5PT62NbrG756crCO
z/8x0sLBiCwVVyUB27O8doVsslH7EehEpbish31K2biPt2YNCctuQBnQEohp3cP9
xu00Urw7GHh0/rEThE3wTRyhkzZpzBNAw0l+AOkkLzvb0cugxfaj4q+DItMDkU+a
TVkoQmOGlvlxfC8RvVKLQENWvIO180RY+3By04yPganoPzMqxAs5gaIyT7to3pxf
0Hgxz/nk4Xbv3EdBUI1tUXTTssGy/+nf96JcWECcBGYusd1xAQYMQX2JoV1cEGzK
tMH2KQ2Va3k5fb9P7Qapx0l54riExpBX+iD/hhiv535daZiJYfKsHxEG6LvJ+zz6
2ZBqGi+WUwDr1n9acqVk+2mJAZR0jxxZYHCmWK2HlMTEnTusZlma6Jf3Zxz+/Z2j
wdVmhqvx83FlW1sFhdU66KZXFBzWPaORHfEDjk958mT1vii0/SRXzdeU/XsMn+rO
NKvi+iLpjAQbFUl6yqwmNBsDVWu2CT/69OabXRXBboOs/A3eOBIJ1zVVfgWeSmyM
fv1tR+TdVjIkAtf6edxFgxtQFW4MNKpjQXjPrVx54uj/h7WRhXlEy7ubuCPi6vac
4afBqUPPKUHadmzdglCPjAtML94cKRoHnZIShZrxdR1Bs/5K6mvi00bH/hYgVoSa
nk2yBxvv/i8yhvBQ//kEwb80Okgr8P6iSgDvHU7YSlyYzdvFQMlqyLXRYDWDpvbG
a0tFc6xOPhAcoohrAZ01hZofIA5HVvzQY6nUUt/BjiZSbIrROVTdMr0i3usuf7lh
DdzhiLNZa0JayVGbRzoSpcUgeDUhCUbhxjoeUpIUxN5Mfp/6DoC9ifrxtITpysqN
uMI2VSaQfGFlXaXuIJC+S0gDmJABandNVa1wFi1LE9g9WqxpXiaD3pzxUdBIpL4r
w2zV/I6TClFz0ZmH5CueweyUUYnLUMAXBWnUrRwqb0pcJTyeyvGwchBxu8NS2LGU
HaUetdm/QzHDifb26QQ+Kiy0gNPBLO8UTdyS7vYwzUDUNmkwJpTZ2+t1fV7AjZMh
fzhEsF9JZgAbpYAWK+b7SMCr+35k4FCYkTnvD0mMIOVJbWvdn/gYW6FfhRrOvUj/
1pukAkTRd3iXA05w3wX9oD4R/ypl3f/9flUn2Q6EvKzFl1PVptF6nqOW48bQ+rbI
75dO6KRU+AW3ompxmJ/Cwlu/SgtXDwmvzaZK/GZRnYMs+xMYZGbcXBK2XdpBo2R/
PtPN+pBiXtIP53bDGm6Sy4Wa386AxdbxL9q+m07kdc6AOr6eB4FdheLbz8joPfuP
l37+P1mRwf3YwVxf01+e7FsptmGs3hXEr1a4N2w1DkgaFXHNL1lycm7XT7R29oY/
IoXx6QSfYRaRll3s4Tvjgr12eciByQWNBoDBxCiD1JW7QF87eJgx0RwckhdtxQA2
tSNV8YwJXEwNOvqCF0c3Lqs+0lUWhzsNNoqD/llUAnB/T76v0zkuU+8YVaciWlzC
Tc1gfw51erZG0LoGgO5Gf4mbuWUmUZp7k8KMdFTIdAt2cPd0xaA1VNh+GVcPAyf2
DFjBIlXvnm5iaMEhxxyJxHq5sZ+5FemgoO4pwSvlM++Ie1NGErEHRsvwTnwjtMSg
BApEAejSodduU/x209aFjvmbN6rxRvIkqDqtYuiJ87VO5g7K2+bGRM55NtNEd+9X
83yjDMLh64pSD2CVO1uOT2B0ThaBJgKfldgLmSc8dRRSQOJFGofqbnZzZZRpg8fI
69/rTS+8y2/jCEmGf7Sjlb+VR1VM8JJ+3xv8ukGaYsaddBknviSCgnOBsfmOxN7P
0caXEhCim2IoMevoAM3fjQ5smC9ebvIpkqyRCfPtGsszKnIshkAir5OYmGa6jsdv
r7nSgY8hoSeBHqUh2MjkgJfUvNgIxF7WP84vkhnGfcDAH1/bqBJEOwXLXC9rJuHk
BCJd6rkWdOeo+ze4sw88uDwybt55pCV3FzrwSoEmuvF7FqoB5XXvXhXlKOdw3ea9
c1p5qWnRz2v+8l6V71cATTSR7cmqNQGkTw5gQ1Qrs3N1wMhTMEAuiVVq8Y7QXF6c
OxhcZZbgdr9Arg22jJtXoOu1s9zAcS7eeGZDUbN3m1TFYgrHeYKVGPEzTtSyGbRZ
bhXJa+hzvBxogpTTCr0fq6UKghujoiuw5gwM6G5FUfd70JDwJG8VqkPq6F9Ywnof
tZDIE+SfIecw2pV1Vr2e1xYALZTiDCPMrdC7zxIS/73wHpkE7L8MFo+sFtJQoxOV
MAE2Hcf8RUCv9bWm4Up2EZq1t3X0f22xFkp28DEHxhsGrdCEy9SDNPC2r6EjQlG4
jCO+h0nRvY5zqDVVmcpdeLjldxHGICwmJFmnFqbZe0xVCx5v9b6/JipHsp1kXcrr
+GSuerdlIepAfcy1yX8MXyXs9vGEynh1KRuO4b41kweF5N/U0c6E9rt6WYJ9LVd0
7WLyBvx5/0BVtPinyphH4c/kQ/YuIA/OsShLu6dnRsay4YEh2rTAUP3vkzfHqEcs
7+uw6sAjWJiq8FtY+1Skw4PJ6L4QAWohsZwlVIy6RrpqhK1m80xh1SUqaxv5FYFe
iy2ei2CTsBDQajMKaxFvu40kpBO7DsRbz92nQVO0+pIl7kKOdCAw5ZgFFa2Zxh1S
56nUBdOwNk/6bBgTB2at+/xGp8AjLEzXyjnsJUqT2vDrKI12QnccDTaYreFHlBBl
eR+mBMx+0yjYq3TXomDHUSIL1dHTGQTG1zhSqfBMvd/Wa7aw09RotaB9AEK6jbhw
3OYGJQUgMD9PZrPwM9MEZoUxUVzrBu1bxIBZaJDtHCrChENHmbNhrLihgfqbFW+I
NJmVe8+fKgJhog2THgAjIbfMRiKcWA57Wxf7ayFvFAMt52grFvHu/gA3c2bJT38A
ccUddA0HH7eKghZNf98ouQUnEWwxcCb7lE2eh4tOVkzCX23/9fRzcKcmTg/tWKcj
7vzHo7mQ8FjgdwKXVBZ/SUGWw/GG7P96GvWPHMfXmxv/R1a/Yqf4XgP0RJgYfEYg
0+mDAf4Gw5r0VGo47MtaZ/gh6NwNaysOl2+zbJjyyaEVM5ac1U4RdNzJesiBbjpf
99Ait3vFd6H5ROE2UAUi7CKtNFrkqg7FhQ2IWW4tiBv4dUCiq3t0NgUucB0A1ySi
GJvwa3nJtDtNqoa+I1Cwp6ZZXQF/RP6Oo9u0zJTIgR1WvO6rz0UbBtS3q6q3TTSU
QXxvxmyrX+tkDUfODOpNS2k2BJUK3CH67QuL2S6/+xR3245HeuVPu4aktpxWi4tB
O96Hq1Bt/iYDu6J0E08hfQZJO9IU07DL4qIgVrKvJlqEzr587I5iJBWdjmHwkJ2c
H2AGJtPsdjY4hFJ9bnG5A/c/xF/T9HDGFjpJAC+OWVC90E7feqhWZarh3jjH+OUg
z/4UxotVQeU88ukTftMFg/1BQrS6h2rGTvQOCU8dz+3ovh4eQgMqA1HRIof7Oj2n
BwTgqYXyKWlkTap4vEv/lUm/lnSR+W6W4KjlRDq7icsG/x2AFtBv334724/DUKpg
tT7oC/AA3yS2NFEvS6n699hgaLBtYcFUDPOE1+mcxtTl/cQcf7tVsFOgzWT0124z
DTttBfPYtwhdVyKo6o/acvHlT+3rO+vRebsgIYUcNY1bT0k66GM72acfM+ljC5sM
F2p/T4XP4974f/FwmfCsfFniC5mBnnaEY5HFsBJDuYkXzBV0WT8dAMxj6qzLj1/n
NKn2q1F37j69Q2v04f8Tv0LtT4Tt20qis8UxspzNe7ytwey/CiXmCHD5/6K+nSiP
dxt3yMBbZQPJsYaLpRwx+1gakxynYk2iHIr8odf9wcSUtXuzS0Twm1cLh9zl0aTT
qNSDehb2V5z47koSLkSnI+G8RFo44QG958UvrSDBFqIO/2yG49vgyzWw4Np2AYpZ
Lfb6O3d4XmS7GR/riTEJ3ruUxLeUQHqu6Mu4Tcp+WZP8Jn6kkQbhG70QnRgy6wEZ
er6lm2+AFaaeoEefyh8oAGP8r2M+tzadPgAfypSVZGeJ4oUwtdKKD8hr52Ha2K/F
aLqWvZNMDTQf7qAAj62UqzqF7BbJaBxMbjvG+iJtjJTuQzlAv0f/CcH9xx1IyXBZ
lkRJNSEQnW0q6m+IvPjnLwTRH2o1rtWPEASE7/yDM9xHeeyQwHTAn6i0zN2B/OGe
6qg+E3pv5xM496Dyx9gwopTf15TBdKGvz9ybab6nRgsiWiS5zU8O0up/2zOAtoI5
6v/D3jp5mrrU15emmDbmPlWGTllgjWyBMNf8evXAD91hVRTdeMob4xlZkY+HMKvb
B+RMaXpjVwfxqYj2kAu8Utxw9fUFmqsG+tE+/XAKtKblUD9q5fRdovKzfhW/KP6o
rAYx+v5OQ/WYf0gE34AIZmD82caqdJpHoO9Xo5jG7RYYhTrG5YUid+tsFkJHUOyr
Z7h/V8hEVFFXVsUGY3r4BnoFUn5Aq+CrX7WeN3R0kDy1tzUE+00d42HenWw2R0sB
1UWnyczex6ryS73KBZXrkSnb7FhKKAOlt9zNsqVs7J/HHILuotHF03mryLL0eShD
5eaYWbyowYxVeM/6U4R7wTOl+P3n43D53AjbQNnu50FmcSNGjSCkgTJwT5+v94tE
BBoALfhFlTYLH6735S9XOdKhJcLsQ7XG88pqTsya1+7yxoYWPYCkfP85+h37t6VW
k0O/qRR219D0NqLnFYo6YaAndrjghmHMqu08KGVvLDYbPd8WHm3oaVAat4Cy5SKv
mEez/oRHLfoav0jE26Cmeglsi1ds+m4cp1GFq3/I06vIYMUkl8I0wSRoVG5utU/P
kLs6lfIEoe1m1Fe2fDDWpWk+ZdB4eeF50xB9wVJFXFhn/hHyjfnf90CE6fW55lf5
kpGdWylo7uQLW8mfExVRtzRhBALUgY5tf+qF9FLfwtodDISkQaMQbgK8Krv14lkD
vcErUrAG/mWxyu/Yu++kSP5ErnswkeTa+EmfSwifCMjSDUgpQSwoJX7T7SJaU7YX
/0yXoF3AxFSC9GlQiNepKzF2tXs6Iygyb7u4bRYFOxQjrARMatJbnur6X8zlGrTT
nqha2JQF3yo/etstjW2LMqtXvXBYJRqzURo9+9U2I8K2cZD64MN54wdrN6+nZrdb
PeEOp2D4282YPEZmKB/JRze1b6duq8t4H1qLhkKQbAjOwqJ7LPjyjIjz2DnUMx9j
sYMeNHpcTJdO/SDUF6CkhZ3Hzg5EJ9ChIjvLqudcwWxAdrvqFiP60pcJBKPYJFp4
gpjg15cNLGg1t54QLfVcBxLJoa4o7TZyP6rsorXBE/04zKEqzHiTzULrNTtYLWLp
wHfpxnWqHM47DgFTy7HLkdr1jLwmdPT9AcuVtzcUC9yOG9VIPzE1pzoTnkCGIXtd
nvW2DpcbTeVcfDTs/asHqdf9MbzUr4DYs9WB80Gwr/AnBhv9puqj/6mD68FA+T1F
vQVfc5dgniJ9gAdDwB1cJYik95rS7nbQggOJqQ1Io9fSZGILBf4hbkJQCkM7eD5A
jFAgfgiQnWIseZvEFupaFSpabxGh5yOJNPfcxuQw02/0PCcd6qcysSyT6NofPT5n
04dwPCI5x8z1o9l9SXbur18+T0ZHD28wIhTUMKpdH3EUqTGn7eDAAKkXITRKVLSD
9AA3KIw2Ltosf0EH7SbjEYNlKJw+XIAEikLManTaDk+9lnt1G1RhrppER9V1zE4q
C1AiIXTaoa956uQ7g0gLa+az6lQfsNOfuDjnyZtuq94eUV5qiPL6UL2dbXLbn8KT
TW11bHAUHe6q8/gpQ19B5CEbwLfpzXWj2VApmqXVrlQbFynEMUazo6bemHcWATQc
vq5eC7BPItubkGNDfY624mJ9Bnk8/MrgXTnQ6yw5fIWk4dkOrdKleI+35dfosqJ5
SPpyU8cBPjQXra70AZu3UB1xKqb71YwPDiHgZrDeMgE70CJHALRINpwpxoLShSvN
YCDE+5TD6+oLbnnlEvCw+XLlKRkRZNZX0G2HLmM0mT9DGidIJ3ugXMEx66iseYd0
rU/dX1/C2ie6LM+ZRElXBuKB5rxNerpHCUeMEtXGVRj6mgPcRZy7DVB7Ng4cbMWv
RFZ41xKBtRILRRSgO2DwcyJwg+UJu/7/Fb5o/9VZ5wqNyZvmz10Gc91Jr92zg5nb
TZ9bPvl4ta9NRSq7+wf8U+kam5nh/3/j4gMROPDprxYDM/q08VyZXK7HBdVtz/UR
7hbArpHqMhq/2sENBkMk24P0phQ46570qLGqpGDpP9BXHkr9u+pagMq8k5RNTcbi
/0xVa2r/HgOT+ZEvjpeHHzRT1JwfHpI+cf0+i/dpQ9PU+D8tYzVDs7wLkGZ9aEI+
QG+kr3hKN5o7SziPnh1ho7uhsCeKZpw2BSy+XSqTy6wAZPFz50oo3OLp93FVtUJj
JnU/V1Df9+PUATEkYUfpeg==
`protect end_protected