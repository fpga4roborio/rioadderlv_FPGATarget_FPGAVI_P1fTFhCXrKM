`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
ddtXksX2+yylW5zu6QL2Lhnb2d1sD00763mmSITNX595NcHTEkwn0zB1Dry37fOW
FufOhVzEJp80NC5qZ/+F0Vk7Ik02dIR0elf3clrjeJRK85K4e3Hoo4xn7YbFUIms
l/8VZSb14+JVGURjfswrIyCUotIzlzVYZ6gzoZwDXIi5gQIBf/gI+KxNXPaKV+PQ
Ufys/12rjO6aI/pPlqSm0hCvftmBcnezN2hk1UeXgOIuKZnogjOsf0iJVX2aOOWE
6pD/psybjbnsNB6kH5uFTA5frkzIzkzl5d9+YDm9OyC+k84E83I/7/j+rk4L2dah
QJOvksSIzN867/4Qt8qYTQ==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="MvBXkzurAa5VTw+1JJ70nePUfoQXBvZOku/SMmg4TwQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
oRtzZL4VJ4iwysPsC8SXYCzXS8Fw2gtZTOskLcDV+1B9Nzn1zTyNtlo6lNICRmmK
ZRVu2BmCc2G+fmzynYlNTnSa7C0Cuel6FYpxCBlOuk3OF2tzAmLAuDyOH3Z1Yjzk
a0aHuoCdIRKv7BrZCdALt03JeUmXKPdOmIlkVGFl8yw=
`protect rights_digest_method = "sha256"
`protect end_toolblock="Jn9CQpRhJt4rnzZPRk+dOpzAubz7omckX1MrFd4p81o="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 9584 )
`protect data_block
gD6l00tciPUa6pDNTk/+t0OO0nC/UTtBwLB41d4inuAUA3i/ALrNyoJVcBnAmEQW
ptbcNp5fxEUJjnOxnedyZEuEBxWRieZFQnkRdF269oNMNuiRq1YLFrZlVa7pSSym
SkFykF+HG6HZs23UZmpivRhi0foDjoiaTqboof9HT/145nlwiIpRzV9YBmfZEVvn
D2t0uhcMAyWk+5NlDs0F8nPnQ9o64KOCiabSv/NKc6mXogkopwV5AOqAoU33csC7
tiva1y4CIASdQPURVYMUcYIcLOxfJ24LwSQVpdzSqz2tWiqoE4s+40NnqzUk8Tkq
Ig+bqbrOyr60UrrNErgk/F0DBaWYWKMrrfFtiY9WIUx1qgz24RnNAnkzeuJj2EIT
5E4DzfGaSkIyWyWXlw/V1lSK92ftIykrs9nLg6JQCYibT9cgGjWFekumqY6Llj4i
cd28RXn1yvuumcNHYSPTPT9+j5O6MG6WSNCBSV9Vm4G9etGScjb7rGXYozZRyovn
0sNhxWA5uPXWZG2jDNk8UmUAc7LYhT9j4L/GiDW24vVVqhdjRVDjuzWUtpUZiCMb
l1IxgR/7mavMPVg7e5O1DKfESAAWS9qPzYnLQPb7jo288HX9+51B/iJ4xL+h3YB2
bKCWMcThrrrENk67PtufvDveauFJgffaV2Ht8YTgVpyxEErje2dhaKXQ1MUtTs5b
7Re5FGILBWlXQbgVmCG+VFgzQFO0Lqxyrm+L9rn8xTLOtyY/CNznbGrDppPXnSqo
tYFJFy2RvvXuagJ1rc508cKecGUr7xQYK9SvuoPfXqFfSEX7pnlcKi9kmsuACtIp
ddHBjyw+YDJsR2g7TsIP5t03qLL6L0Hbl6uRGimIsrve5XnetDmeZEQ0c67XVY3q
DvMST58zh3TrJxPHftYUvgC8ZZvPvMebopiaBNJYcQXe5qOCJjB+JwScUr0PMZg6
vJfOY+fCo7vknCrulW+S+ZAVKbwYlxhBH1BuVdqR50ued7kSo8jZGdXsNrf7NS4V
tkTPPsOl3AewsF3/t+O0dFGvljdAM1LLndFWyPzNe0fBq3LqnuIz4RO1BQQ7s7YW
RcyUHQY36x4ES45sv3iih3v1Nsgz83e8Cy+PpW6oi6C7fmI+qgbIBvdoppWJ11Wx
Q+uo420doifU/JjHykqC6iErrCULBAJYEG7Acb+5222NRsatqyOzOus/aF6jCtB4
1BUOG+tNovbWqbQoMzIUKg01aYX84vt3oPmLLmlxtUQFH8Dwg5Qc+NhVBTkpuvux
QMTla7Ql11KCYNTRSjblqk+4/vU9+vSVkmMQO94b8P1gs/Q6luzj5rNjo3nRFDVk
hFPhVuO+wo3tq/pCnOI4Nh7J0+fCEwZQWSji9yI6uky+7V4Cwc7Nq+4851+HzTzf
tqjk1sJONVEA/onPB5GPKCgfzkPbNE+Eq2Si2243/O5qGTrjGCOq26SrSIgGH1oS
EftnKUFli+FJk6bxTudvJUkeL9zEq4Z0pru9hbPFdvFkiZVvBtMazsvK7XLreyiQ
n5ODy7nFZuSooE1DuRt8cBXJUvroDhV35l+DehJF576QPEsJKbPNGiYTiiBgODaF
Dps4hMnPw1tjtvVyc5U7WwDbvRsFleyx2kAwNGME6p8Bnnljbbww/wuC6q4ouduI
UcynMM2cWrCkOvYNPE7NR05F6FNefMxLZLJdOTHn5oycKqcCc9MqlXAOzDK3GBWG
UgrUCG5tgNEckYctZ5m9XyqpYeJOk7pL64yAYe4zk8VNs7ztuwlPiNd5oiWpo5hf
XJo6S+OaaA2rHu5LOBrgu3ze7apm0QCbJS+3XU5qJ5TBDPqTUXiABNqEa9j4iYA5
Rqogi+ljEjwpObURoqpOHkCRVCVVb/k9kv2l0qRA/1t7A8vPf92OQ9Wf8LyL1qqH
J5MEGGQBWpgYR8s2WNpsecfgU3SFjyAwKxE8iCqXMUIGWiVGQc+8CIRINONkaCiO
VdgYd0faqlAsQG6D1zmx2YkDzzsCCOkEkCC9iO7nbBr2sz8arBezhKi9stwcaJMK
HQs1+4KEI49FNLGNzKB5JBRGRfuP6KeJ7fxlc4YxSUZzEFcm9wBwAGwGVxwFzATE
0lU8iKcvn46q2vSz5RMmCLkDrWBglLpfYhxlXKizJ1PrmoS6JQcfu4RnZmfYAB7w
9fh5t1R7MOP+Lfga6c7ht4LZFc4cT8vxzb0bpdpclzCzxUr1HEP7cYpLMW8SFWfW
9Yl94MA/q+EdY9YzSk5O8PpS66/CasTlSferOiYfgD9cdT3rDpBbf1PAc1KtHDAs
nVKRL3ouHvYiRdTqrlyrp5FEDm50PPgVQIqKW7qBzwREMD+BnG71cnu3FdZQNpQs
0R1T8XT/thH2IxHPDzrQkd+es20R6B6CdL7AO6xnBsI515ZSOSrpC5GH+LUpCrXJ
GFR9qprhwLGzI7v4Th2ls4cr4zpFXyNOHEF6xj4Eh1yIR4LkCiBtK7Wh4cyqbIdX
fYPyRFbF9m8CFKlujGYoO56nBWq7AoCVkWWEyfxHGutW/k1NiAHpUIEOhTFBvXCA
KFqo6kVi2cL8qklEuN0pKuxIEfBh6Pj5i00d5ooXPbjs0K+UYhOlFVlKtg80FKOx
4xewnKW88JqfF3WCGRCPBaYfxMJv+x4pgkWRd0mAXxmmdQ039CtF6nowo8NCLTPj
0W4hD3y5g7emX/RSXigbdVFiqplbROuqSD/01+ZteBdXB4EjZZfPRy0YCe5x4mH8
DvwvtdT8wi460kjd2FRX4+STuhk/ayaW0JWJtp3cj8fzeS1T1UkPNRDRYxB3EBMh
unEIEkdChOg1O+G0iiRq0TnsLZDwvOCYwRubK1P7Cem6HR2MoTLdkUegP6DKstEl
qKqzn1RfsSDVxU2WU1nN71oJJUPjNOzbJ3tb+bUv4cP+hS0EWan640g6AhXP4U1B
GOBClRLPWKnWmtPu8PaYZGTD22RqCrVM80UK/kNC38Jfm7vG2jbYmk4lkkksDs5f
62dIVj3BS8GPPu2MIGbjBTG6V3PddwnlmcPYuROHAq0ddAAP09es2A/snZCMf1fH
qdyNVLCehXHTRwQuu+6HpJwXbkhR2HI1i5juaZAQbIbplZbjpr2sEfhtscuMAJ0L
B9h4Aaxdz0MVFqwQXiR150JPH048xH11MEwGpWG8iZTtvW3WD/V6jnVPYwo+a715
0XPM78IVTY/MyTaQ3/aY0nTrU8V4p9bQ0syQrLMnuFDywi9W8gUiTyY65oNEO2P9
o+XCbsVTbb8FJCL2eNhAlguPlIXNH9rbZcgXMX9/sZ5bWzgHuC3wVe2lDVYZQdXj
oyKeUwR4rjkz2+HngXNkEYU8a1mPEEC3vbMQ+h/5JTNfaf8thhQrAu/ILzAkD4+t
0/GtuAnt/9Jm03OTCklYISxdfnkxuoXLKLCQ0sPEL6OWUpsSOxzMEBZoHJHSaLqz
GbefSJ7RUZ7IES8ia9U8bHWVmohH3tRo6s16FBtSLgVk+oKorN355J5z7tRzV6pd
oAyN4HsvYiSv/tSi+U2HTAxiAfHIuWtNAazx3WISFV7W1IEP8TOpiaDMPTBIxhkf
oKw+dmCPCrQWT2XDRBkjKBOMgw9xnOEI4rKmGbVTBD1aMkwkenAywUib0O+XpzTq
qF7nWn0yO6+rsRuCs4g6RNZYhs2OxChT3GZgO0OW8WdPwdrGXZke3d91y4pvSl10
FjO7PdNNUxfScspxurMdRqTZ8aTPTn5iwugM9SiKRbgDvQl6W1Lpmj6XateAgGID
BuoLaT8zBGjIlrgiDqEXfO+lF4+U6Uev4mNhGClH8H85jtd8fApPwsuDkmb4Sp+O
eoiVhiYIQNtuh4WcBkaOqCvqsyKcHD6VJKIV9Y4jINTjeZ3SPVLJeucgQJYJJn4R
sewMjPdFvfBXfwECuQF2HDfvFgpli1MXi2302bo3TeS+oAHXaJZdMWBP1nKmVDVN
FoBzJ87Ho8g5E/U6sFnNok0bxhGDCme7hi6FTBnoQKgBiwrB3tW5rMKui6sBZS1/
H7zqd8iVnEI1cRiBBAsnn6ws7iB3X3qZqyM9VgNcA48hA86Cw3DNbDf3HxMZvWt+
WrqOKUYnABu7oQH99jreUYc3YIAvzcN6zJQz6aq4RReIWQQS0JYbRlC8/LLOa6xz
F+KNw0T5ecQhXfz2CMZj9qmU1OZ55bJdl+HRU/xol/iEw3Hl8in14vNldSlsIeFF
ZhNL41rjQzl2Xfbh+eBdqtw1oxwiGQ0huGyqiETg31M5ewwmgUgMkGFZNrcnww6t
irMNfI0qmCQX7lYfjlXOKx0WTpGBM13aodFeOayPNHszjpCLC13jfPHdo7tSjApw
qvGcKNOfq+vK4HNkIa4QtwknSv30TGm6hjRTN0hFoaTbA+ww36jeRAd7oO70ooyg
CFbM2ggOmStlJxazw755uBF2JE/qftwzznrbhVLTtv0X7J+wXp/oLEarX0hsFlYp
+cbMXvUgWk8jAsz238IchCqi2WuI270dbzgkBvsut39qCONCglgTATyVvdFq9QCB
yMO9+Wr8cS7bbfDCotULO6/qh/T86/NAG0lhBU5S/pxNY4ymfk8HMXDbwD7sK7kb
DJY9itO9Ti2YxahKfazwsOoWiW8dlSBnPTfVd7mDRWVpJSQKSfe1Sn8r0NcfO3IW
/zc2sGdfCJHxYzVY5VVqsTryPSdM93IvAmaxJ7JF0EpPP8O5O0rwHidV7sOe79hV
Gi7JIM5kEU5AzfshBVUI4+U38RIEoLJ5oXgvAc/G+SdVLwpMOG+zlQrXoUYTAvXx
98sGuLtqTg3ffB1MryQw7nzDaut/OajaP9/G/ERPkbDLuYUUmUWcBwF72hpTqFBR
L0RzcJb1zkJu0UwFiIUCBOj2Mg+l2XuRy4nUUWjWN0lPD46W+CAewu2Bs6z9F//X
AF923drCC3emqqQMwUAVVQNrH70gOjS/dzTp8NDdTtlU06u2YH7cMG8SM4EyV6bA
c9/y5Gmk7N1nfZ0Y5OOyoRlimCRNmdthZMEIPddPSKMvHeP7xoBl+VfANhty9V1m
oup/v8ZddCrWUWxz9NWxmyZHns+2ovOIGasKZCqOt5R7ejgkEFXhahoMkxfGZ4Iw
oONxmcDbkRajx/S1XV+bo4/xlDZkHcKnzr9c3Blw7ab8kA/r8lEvUtZD52hPPw+5
j/f5CSvrmlwSqJe204yegvKUAujzVjHRQq1bynARkktAsR/2gjmuiZJX6aKTp082
BXsQPH+v1I1J3uUSRtw7TBTpDX7D1nAP2N9F6skoi6ix8AkkVV2lvRWxGP7yf2Uw
dRhZMc2MLbv7SROadGwRQGchim05SKnwtn+bqZeg7/eOtraQthmT30a0vTTPPHIQ
fNkypOS5vnMWVm45rM3MHiRExmAOL5K/eTRJ6kW4D16FZzAcr2dBLGl8n/E7E1kf
ZR65+CUq8flD+/ZlB2jlweNZ0eq8Jhg1rICaN3ZBhchNoQ7fmk5u56G/70Hm8bzU
9HxVNRhBF+895AzdZHcbnsDjttyBrm9sPRGESltXGzWrxYe1YA7Lph2avA/8orXR
hsULNGpCATAZg6Dno2WJJzLiY5PZmwlDw073gNYQrmdJFslxz1cVXfe95EtKTAx6
PtS7wWhXucO1W2Kn8if+pAuNuCweYtecw4k0/P1Spr0IRfWR9mzUyHhGPI38K94c
Iq/h24ahXML4F7XR+zIDhn5zeuXM8pqKJ0aZYiL5VsfpIVQURr3HvI7lk4aN6O+z
iYcfZ/Ph7bS+OAxaRXjebjsIwhTIToLOsbUn0vHNsL1/l05KsdgJQBreKVWFAbCn
sOS77OewnIqw3nCB2X/rdR1FagdTWoUa2q1FZ/XiD7xbwp6PPmA9bXfm9tkJb/OU
KxQnuUQHWmgujde3red8z5fDhm1FeE2mPMJroh//fCAQnk/ez3uqogfvOZ0/LM/t
DBDEw77nLec2IqQ71i78S3SD4ouSDWRHRuda0Yr1glpq8MoYNTwnJXBhxiV2oYdb
UUmrc96Em56qUaYBDzBNKOdSoW7qcBkEN6Qv041/evEA31aiut0grNxdJmSUG4zF
X6MCNVxM0vYC9xz3ua7vowX6zdzP0shpoRNqL7/9kTElFq5HH15b2oxeb7Q7A8CC
NiJv52dZqTPNARPz5XixEmZ1JqJEmZ1sTYfOLOSkxM4Hg4goHyYWfYQ6uE4dEPsL
V43i3z5XqEcpKEf1/8/OMvne8RFzadIa/IWVCaGEoHpwfA7a4pLkR7eN3X6dtMSc
ASTb4xVuoFUqiRERDeUueWeBn4+GY6GUQeqHm3I7vtqxd7X6fwkrDFnCObig/E+Z
FXPV45nWQcgqnGsQcMm7P2FZ6jG/a+ODI78c8Y0Zw2/vFEgXwZchuz3Y7CoX2jjG
5FymXo1pfOcxvy7tcMCMtZqC/6GG2q9m/CvKN90bmAH340xCs4ucpZQR2pDoDqJM
8gfkdxTU7xuxgjvqqbjqnuHkHVPFHPW3zcf+hzF4ggLCroJDLp8tLWgprkzsibcB
EdTyHcEmNDxAlj0C8p7ZPwUv5/wzRAnlyb1JeWRFrSu+gEG57MhkuiGjLs76zja2
Pl+DADiplSHH5PfLvw+x8j1fvP6OdyeNC8tGIFq4CZotAnCulNLBJTbwoXeLBDTG
nNOAe4U6oaGmL4AdWh8Zne1nHu2Qi9wvpqObUHPSiV1lpWw8wVBLZ0b0Qr8UMPtf
n4IXq0YIl6QZs/DvPbu9DNqRfOkzuuEBxULIBujcm47pmId84KdX19F8i7KtyWFT
4XslhQdfxrE8MYtfzt4rI8aB1/FDlJb2yjuWYIJFr666/hdiov0OOuOoI6SVnciT
rVFN0oEd0nLxE9MIsyj9z/UbyUU/+hlv1BB/y1LEjXbJahMtbow48LaJUoSLZXtq
6R+x+u1DrzYfKjkcxjIRFHi49PDyd6kA3R5qPJaPzlk9jMBa4Xb275KrnReLH9r2
fyhCCptt6BMqkyCWXPZjr8F4O2gmkwUFj59EvftGc9Lb0XDSlBLXRs21K78G2s4p
FmKDL0fMs+8MuKkMTHhl27+XGy5iIZF8SWV5yntQrnvfqa305lDMmcDXCLuYGZFP
HFZ/AearmMWBvpz+RrH2WmUxoa4tezeNsHEzGZU+vlJqxFx/I0sYsdXH0zISJfyF
V5+OhulA3mEHI2mDefTMs+sW/OjTazSeRWp/J9fnLKtzYcfzFxubC+gt4JDI3EhY
y37EgUvPdQMJ/19QuLKxeAwXDEorrzvJOju/mYEqhN0f5VaR//Tg2cSvvmfO9mRw
3hBkPCdmdYSPc7wvwXjDxLluLOaSMaUhWmKqsFABz4LiwQ54VQR0h/s0mehub9QO
4IyrFK9uYhxoL1APeygwWC5EkMFaMcIzq99dX5waKlhnTqGM/6WsJH+HVDpSGfWn
xfiXOw3zY09tZSMGrtZa/6BA4joBQy5joWfOG7IVEkHfvd6tiPxXotg9mtLPorI4
TH1vb9XUtmLQV/1pybwePInW9gDQbKrglssQCeQIeJuh9KiETK71DIsC1iWrhmUB
YKJ9dCRFwhDRNHRu7l9Hca3EqIApZ/WLkODHjR5i8Wc3cDyylcMIljkGli/B9/eW
vqWYJiIxlO6f5cutpf8b60R9Dn3AMsGd8+yx+DECofneNf4IfPfTmPPwaZvSQL5v
enXnkp6tJab+hYj+bO9lB0a8Qeee1NovCkTwQ1AyRd4Nfswy10z0xmkcvlV0XK4i
T61XI4AyUdX9z8Pvyxxectd9o2oRrAu3lQQJt14p1JWmzu8GOxJQZtR7oEuAFmcW
vcyjQcBZ7+/2N+I6Ah73FO1mNp9D827mkCyX5Vh/bGjSvIcsR/XVJlzjOYjH6c61
5UQVhO1Fotie+Nk+uEK5hgj9fJ8wPAUmjZoc/ymGgULGdn9LpLTrVm8J+4maHPxe
PugFLuXeu9hElSP2qsk38BLUdhtKlctDHb6SW4FjUa7clNkIgMvrT1KCIPKHs8la
pPAT1XCKEoGDowwSPDqjCCmeqWPwPXeW643kne7f/5jkiW0k89j5+Ly0sxt+uOmv
2DC1hCKDkoo8M2DcFeXMVjN7bwQrKD3sJ/QsQ2lpJSKZW2AeeIme9zpC5Kca8hn4
op5sUQMQPzkwPLzdOwqeM/RL4g3PkiOqDhnLonzGFypqs+5k0XeFB+A/Jaaya7Xp
ezJBd1qeMri/wCr9jVGBkGLEUhr//Jb/yHT/eIYI1EsuQ3cBpsHDeee1nhljNe6R
OL7dijBiYUZsue8aAu1OvNENGyAjue3NQfiaYLgz9MXujg1BHXw56WthyeKS06AI
ZG/jj3NCmGDqu3I7c1STSO0x3oh4il2BOOxfVUocqnbJH5Oby+gmBI1oGOUIBaCr
Nai9D4vdBGf58Z2SG4qUO7TZiXbn4eSbssltlikkFFl5vEGnaK2c6MQ4StugGcij
OpXijr9ZC7lNXJC9EaLUljlrXTsD6kZ1E3wFWg6yB8aLmeL+xmKOnwuOh8f1/Hun
2gmsNWztkiEQalxrvoRrryWLKC1DrafSgKgkGNbxvQBjzh64nnTQaIEOfLUiUFt3
pPK02pGU9KCs3Fsn2rgxp7DK5X7IqPO2+jg6oVhujiIkAnSdUBq3uGqX4sY7vYkH
K7tAk2LMOYDgde4qZlGymg8dadXkdw22IpRBsEsU1PxDCmg5ZupC/fN9vB37nZs5
x/eZhdhxT/Vj0z0ZyoBgXz4X9JseEAVnt9l+LZqn9W9Muwefj7knxqPu2TmNQ1nV
6UpdR/eTEnoVGQtCH+PyfUuK8igXhbiY/UX2csQJuc6pGTxLxGo/QXNjz0E/ytmu
oCsDp2tafV0wc8prqdM3NamUshHKMD1QHpwVyTiNQe72HKXJ9JTH2yr1SNFImBFN
CFH8SfND04Cp4aEKxZ+C9JYGqpbBpDk9msmyBB2Jo3vmtIPB7jyohGkbM0fUxdlA
e4V7jFmxb0FuwVg7jxASC56ttOxdzLKWDFSbHlavDs5egz11LxvpTvMB4NGtM0X5
8JPG45gItSiFGCcuC9+qRFyMiI4AhagCVNJWGauQoiDk18sSxc419C+JmGSVOHI7
gVtLwt5FoDf82aXPXvKZOh4Ma+fdZdjwCNDfaCzZRnoi039PyGE4TEg9dh0uYOGQ
TgEjZrk7OU5dQupQsQOj7IPli5KyyMbZqbEUhMdncfrYvocrH1pkqAyq7Inb/HsP
27tAVO5/87tRmkFEL6FW5kJe14cPMfmgBexWuzvHmF4E7j1m2s/2Jk38kaHUCFju
XxJ3Z9gCZLysN4kmYNylHZFtxJnDxzEAPXXYUezLqy/SesXt/xwkZ2tyEqCgkoME
Q8Nw97EMp063lBjYXNVhDLK+u7fb8HrT5LJ7R1TlBmuwGcFyKKTJmfnI8QnCLtTr
KIeLtqH0moxQL4Lm0yYZhdW+OGY38pQsF/5/FfVLMJvO1SU2ElvS1ksuKOwDnXFf
QpYR2r4gKTHKEmwd0PzDHKpuCAeaDK+HgO1WGQ+8+n27mWDlsY/kx69yZwCW47H4
uN4MIscFrjAr5KaVBIQ05MIOVh2/kk1gVxzgXsE7fgLMAQNz9o1qV2qq4XAOjR6X
PO/3HD71v1+yT71qqFi3dfbKePHkDdrKV3EXGy4fb8bA3WUzGHNoL7pwm7v5KEIy
sHHsGAJUuwAcDRChE3NNNAqCy+Wio1qVFWHhkq3zfKwSvH1F4G5RjxmuSfwK/f3M
Tk0/PllLDgxC/4WWmT+IcsX3afY/sd7h8GelIvcpj+uNyrA2UyPokuBxPO/qjPUo
u/vypyIhsLJp2OK8dTZdBHbS3uvPMcxdraaRGHfBmQcV6yWh1bV3y2a0dRvxsBH+
JCr+rLDWxCaOMisTRTdEKFEmRFmITqq9CtTG801TnHhnB2N1oPuEm9cPjNjAQwpV
4xMMSsz2p14nmz4jyA3eL72u9BRrmd/hRw603rr+trOAdgNJc/lf3o3Y0ahP9l8M
5R6pOomDyyYCoT9BlOdMHfHT4DlbY4ufdJ4ONcHcKqrviwRLKyXTrB/b9c4uTXEo
X+GTOI1ZUz9AdnyAn//mdfAGuYNZFIfLX2AezMvCKE5DjFibYlqrgPsmhfYjdfxJ
hFcPYYJhOHXjS3Hh/NDHL/ieU5SNvNI+Ea8GdAAVzc2rnVawjpFn7+ndGHqQQ/AV
LZkhJzKSQ0qbwjSXKldr0tSSUX5eDtO4XYvXuKoKu93KNu8SWXgx/98ugarUtWLC
YTOR5slf7S+IkEwVaq1yPCiRYuMaQZM4/SbIqN9RhInq4GmIgbneESaAV6S2hWvn
maiJGdOBjto3HZd3DQFroC6rOIhzeVaNqvx4duhU0bwxgAF74VMePK7eaTXIFvGw
FkwJrickKFUE4AvDrpw4sYTVa2VA8fvLAH2DdjikC93sdp/5hMC2TABrI5FJ9KkS
Tbu7VJAtKndimsrWuucHrYoNBEnZqR7maWW86PpUB5iBaI6rtPH/J56VgYHXFb5b
5QZ8zUZneSwHAgV5LSh9N6hEp6o0BR4UVSaDTrMsb3hYzXANe7p94hgX4DIayqlh
LRcE3lAlRgKbgQE9N4PvPp8ZAu50Tr/WRKNc1ELvh9J94C6gVO2jDaJB2DZ5sSCI
bFvovE78t1PfFnr4Y0i8K7hI6/WmYEDdRXfkU3y10aXb0PWJ+pAUKAi530KTIJtc
03Du1AF2OLoBxOuyDX44FofXACtCVywjmVhVjlOTakajP8ZytXM0ITXmXk/VjZfT
i+cpfyhzcuxIjOEj8Qi4u/Bn5iCR1B0LnK9vv1p1Bh+tadDWs1s4pLok32eaNASY
9QOUpyiZtLDihzayenqxLLfmbqbvDeoyI4CJU65OnemEJETABUghkj6fvWNwtXsK
Dt4OhP5frB/x5vHCOHsPlh1OROPQYgJ5Sum5cLvckBaL9SDnVhUrIhuJMJVrkk2+
NA9jdAifIv8eDwTBk4ERMWvFBKeeugxnhT8xolz2F3i/KFpPHVQUYwM+yoR0wYBf
P0LON8jBNlvRB+lLkEFHl5rvSAoq/V1YeiGwEdFUvb8+mFMwDVawYQKk1tt54wtW
m1FDlGH3BD2JLasrPWmQ46yChIEZw0Q5dU4xZL9+8pSXzsg6C8Q5nowuRIl+NTv/
3gthOXkiS0Jv+IDWkoJbfc2uGNE18b68MbaeKZSF9bnA8OqcG0nrc1nvo54oA8ez
OF5DQPHoEbFmt5Vp7HSJGFDfcBGFxPEErVezkvE1NSFfd0ona9zlM9cZ8q2R+FgV
EP17jQw4mKbNgckiSFkvPJTkKs17OFe0aAkl1FwVvPXXdv7z04aW5ewAPaidK441
DbWWUys/MuvLhcNZ4PGNNyjIv1ehNf6CoPROMsa91Y/0ynFM+8psF0dEF/p1HB0M
1LlI+UXcChQPK/rk+RkoprqB/wPz31i+tkCTMuIWR2YBLpw7BOGdHE3FinhtNlji
jO3KdmyzaVtQO6wGxVac4Fo48Vw/0Jy0G8eTlkrpX8DztlV7AIO4XfdqL71pZXVr
zF9F1ZA4dQ7h+h6JS32CEM3xSEAy7Qlv3y8olH5/J2TUcqIJAxIm8A+I20FsVVI7
fsGXwHOyGyPFP9SeQwnL4yLWOdAvom+qA4UKkccj2KYP0VwJfCIai2HEoTrFU8EW
wPGrsX9+cqvH4YdKO59fRYDmvaCcX2HYn4n3jV7jE6z0fHGS0tuYCiTV3mutG4zw
mgOJjcm6SThmS3ZMFRNM0a1LtWhHiKmRvYTLXrlVRB1hwuZJm14Kwl23227WzYcM
1T8aVfq7TDvsEOLYz7fcXgEK3HZ5JlfOGTvGiep7TqvS33fnEKLC7pwBoobNUSoz
CigaMTu2OsbBefu9Cb8rTh3rN64D6oZGgGg3TvTWohwEXD6ev9cI63B/KWTwTp7J
WIHtplW4c4Tkv81VchyGDHvzFWhVzEGewnnAtMWiJPxsQXuOHPFVVJ8v0C05107y
QyWbQeTyoj0yBcgcYlT9SKbS0mW/ZV4UFaNLSSbANnfs9vyw7VMF/liVimVJjRsn
yYay5MknrjXBW2jbQwV/kGEXSpoKuCU5A6aLPdWGKr6LuTSXv5OXs78s/1+JvqC0
H7hxDRVkfzjsjHYilgMsHnPOHaA78Re0n+GIOI2Y0u4CoMpWqvnMLD4fqHXkrvSy
MfJhmfHgqGLO7YV2PqHckG1r1S2LIEL9uzZf2R3feXm4tldC5JyngHpv6UmneRX+
/s/pqJRRRsV03vkYiFYs7jDV3r8hMdx8J4fJveovZrpuhWxnbEdU4ANV5YzA6iUq
8AFNT7g8dX489FRXcwTN0q/c58kjFudYumLJy4WDeHlAccoS88E820Zn+UTKEN/6
f1LgWX+vP0ht1c1vVgGpXl9TYPOCyJP7jpmWBjQ7FL6mwVHO4MbffTS9AnFXymxG
mtFp/rvRcvZc9/govqvyaWb2RL9H/0MUMWhv4UQMKC5O8DSlwBQlVKYzb6hC+qWD
f+Hj40AhfDf8Wa5uPzou24KNbnU/orVNM1JH4/DmtlvGscNGOel7qvhG/AGduXq0
G1GY5RtyEc2jWwgRIMKiQYG125Rb4MZE0QU+a/mQ1jdKyP+JPPdbNkAUwH+CVkn2
ttJQLRR17H5vSWwH9WaJd38zsrTyoLH0GAhs/eUMaW9/S0P9ZAvRp9geudyjxpJF
NtcvWBXrwUUPnYFkL2fge98anAspO6tcvUNqcdbqngfIxHZjZrEYbqJBWZXUgcTn
kcUNctdQu5njFwOUoNeXeRALmiYiK8YCKHjYy5dPbog=
`protect end_protected