`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
ddtXksX2+yylW5zu6QL2Lhnb2d1sD00763mmSITNX595NcHTEkwn0zB1Dry37fOW
FufOhVzEJp80NC5qZ/+F0Vk7Ik02dIR0elf3clrjeJRK85K4e3Hoo4xn7YbFUIms
l/8VZSb14+JVGURjfswrIyCUotIzlzVYZ6gzoZwDXIi5gQIBf/gI+KxNXPaKV+PQ
Ufys/12rjO6aI/pPlqSm0hCvftmBcnezN2hk1UeXgOIuKZnogjOsf0iJVX2aOOWE
6pD/psybjbnsNB6kH5uFTA5frkzIzkzl5d9+YDm9OyC+k84E83I/7/j+rk4L2dah
QJOvksSIzN867/4Qt8qYTQ==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="MvBXkzurAa5VTw+1JJ70nePUfoQXBvZOku/SMmg4TwQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
oRtzZL4VJ4iwysPsC8SXYCzXS8Fw2gtZTOskLcDV+1B9Nzn1zTyNtlo6lNICRmmK
ZRVu2BmCc2G+fmzynYlNTnSa7C0Cuel6FYpxCBlOuk3OF2tzAmLAuDyOH3Z1Yjzk
a0aHuoCdIRKv7BrZCdALt03JeUmXKPdOmIlkVGFl8yw=
`protect rights_digest_method = "sha256"
`protect end_toolblock="Jn9CQpRhJt4rnzZPRk+dOpzAubz7omckX1MrFd4p81o="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 13376 )
`protect data_block
gD6l00tciPUa6pDNTk/+t0OO0nC/UTtBwLB41d4inuAUA3i/ALrNyoJVcBnAmEQW
ptbcNp5fxEUJjnOxnedyZEuEBxWRieZFQnkRdF269oNhwJX1uWBa/PVIjj9snLqr
bUH3wDYWdo7LSIKgNv3osOxD90soNzQX3T+KF7lO2dbC/TdLXmCew9BTUNDKjUJn
cr0EiaDLPKhAvB7ANSLbDE4z5CAmR1nrpa8CXFjNJkv2m0o9jRCgqAD7h5wP/G58
Y6Tg9nkxrvMKC7X8woUhcWkXsnD/FMwb1wboxX2NuQAy5g7oBQmoRvTDnwLPGv48
7xgVo5ZhJWOhSDXywr+QfZUutoX0NPPLcsHMP0+tlZG2nhPWrYNqNAR6X2YE9MZ9
nyjwkadaq0FgFfa6lyDrMlbX7U68Wd+yMr/EHnG+J44Aq43QwB8ZyVXiwgcaYnhu
hm20ObnkwERq0x4eLCuRX80Ff9U63K4L9GOTehCQqgYBwOuZe/XO7Phwvgz/l+vk
Jtx1ZMKvjp/gUFfjZ2RAzopG8PEaDttUiK7sZ3j36mktvDDkW/7+ApTj8V1+pupU
So3qfr7ISAHnnEY4WCIow1FSsh0BxhXqmJGv2MAJDXf2ujD++iu1rbj4smYfSC+Y
jOWWw7s+W+PZ6zoQj7Tmy4fFfr8RrAdLk/frF/154UqB1M6B39u58z7aHQnsL/Jd
QUYoDbh2CqtMQ7zJ4C9i2ER2pTNQL/jfMG5t1NfTG9iFEOTAbXKUwLN77q/CxaJF
SXWe1o3b1OxWGJjNXpp8RdDnSlQeHDbj8KcVPsswMqa2PsenBrqa1p1XIA7ZOrlI
EVPRb9/BFNe4gi9wnw6LUeGmui06U1vPIFNkdo/hIJIAkCsdnIF3W0VHGu5uHGWN
MZXj9o6JbsZQ7OVpw12xG5zhKRNy90w/tM8I3htomhUCAp+oaM18xQlwjEZb/L5g
Os8lsBwgba8RWI1ahXeUIui79W50EFvKr315XhOcH2qZeqqJs+9qVLt9ejml82sJ
B0QsXAixK/IukVNRBcF/1ZnnLbkwRACjDh+l86qpgK5UHGl51Jooia++Hp/St+qo
AqV3yhmmSf9chbG6Fydend7EAnZSpF09m55Oh8qnHaEvA/WEdZUKfkTYZ4vWVjKp
xwxXHuNBrYHYWfw2lUyh0EpeydNML0EFKTNEEW7ID0S+nRnwi0FNy9GAIQ9WEUUU
dfQJLCRKZ3c6MyarF7HHjRUDVdeHEKzHPH3nc3aB/SJgdVT0Llx77IiU9kedylsD
j9x78jlTjdgkwAHW98on9oALZK7vLLOzbIwUWHqyUzTaMxfXaP9kbNzdNMqbU2HA
7F+3ROz/rbEdQPKx32W5TwXW+/jzoqhSENY93ya7fLV4FVlyrWbS6kPu6gXHyZ60
+PmSEtCM+++vUHCjW3ffGG9wOLhnrAybRSBwUAjjoic5ueBHYstRoh1Ky4wXKibg
iAA7Q7JEp6cQ5qXzM/z3yRDmrDB0dG68bzaxWKg20UfC8HpMI9bdJcDZ6BDnEq0L
a6xl6D4gAtJW+F2aqH20n3Kk/ey6x1XN9i2BZ3TConlAPnWJkBxsKWdS6avY85tV
AEuvkjj9EwGVnxhkaAgUCfw2uJVj9Q3UQUxshb9ezaHVV7+Kk4IG1aw3GnlkLyxF
O3d3x6aGEN5auxKZtMKqNTxCmoem3jypw7ioB6+mhByQE6BMyKrr3tt99Zb1MJIx
zYm8aA9homcC9ZQcwgss5sj2lGjStVqUGaokrZrNky7FEAwIhIwS/h/7YnX/NQrW
UgdKd6RkZJ6k6SwDj4YXH2W2uaW2JZC0Ez0wAu2N+HZb8E69xFmmnatj6SShkwSE
Ez4mBc86RV/ShO7TSiL0MqOxf68Z7coXmUippOaFqilsfAJUqMTb0Phz313zMHxw
BowtJ9AN1BwwQ1gzUT6vAtLbmRVozuFr+PS0qH1rsTNv9iqX4ayIGRVvrHWFy46H
csxCPdlSARonp74PItJF5zQS5GKZuGIHUDia1Jz4sW29BhzOcXiT85hOfxlKcONM
/cEVMcShMIv9SmZ0dGJgGY8f7xi47iKi1aZZCb83/fAwlaGKicAvOfn8Q7r7/Ftr
3Ga0xBYE7fBTxIhMxmDUVLInDvEcRofsY0u+rYtWQvEE2yVb3IUeI1fkpnzv7Uqp
nFdZ1sv/9Wb1KH1v4fOlevtVaRGp/h+/ly07hfEpXwo8OesrvJtCCime7+Klfw56
DyV8/TTOfFejEXhGl5j1tp2pqGTQn581KSELV+huXpb/4ekwrdvh6FqA3kqW322l
J6UNqF8J3MmZINk+1iSK/G3VIJ0KZoRVDXDevd8ucEeOkeOgmUNgDRqs9q3fA3M7
lEEz55MtN10PPvBjm5KZ5jgOs+kvMOHiBgc1oV3NLmkSORxpENUO9suYKZyGFx4J
q3fGsJQhikktwXoXLJ0qrln2z+NnnHXRB0qAcOzxQA/rpd2jxYkeIbBtLorSKLYQ
q3/5KXfBijDVZnpNRnyOe62lLRgh3cu8lioTJMpdAIP0Q8yemXS4OrnD0hAIXzXN
1H33krdSpg7gMNkLPPHbrS3MZqEThkTdpD0OtH+h0+xBwCpti8WZTk+IaWGQwLuX
HbbAlO1zL8o0oQrPqwgTXMLT12NkPmedKD94X/HTIwLtY7vSNYPymJAOhgsFtvR7
4dSB72dxGnZRKc9EwUt0YgAMeXMDWSXw/VJM3Y/5Xljjz22SvXJOmg3mA+ArtrvL
YoMESqJo02Me43QtFy+SJoGtVJiGr4WNVOwiJIsGc1znTsVhHn1WuHqxNB2rMwnO
ASWn+TLxVPWgGvhXr9vrSLyoAtltMiAQbnHAkvu0pqGntvcUZZkoyEoD4A6Zspdd
kPzKgU4LapP4PQomO3YEyCsglVJEXe6jhPEpzsCzU4j6rL7tBi4dCNy5S2a03XM7
cNPF0fjIaT4mH4hDY9diMPb62p+4RY9oEDnQHK64um68t+yt8n+4gLfmNKfEh2Et
jpJz+BjRCp5i7EcxocwTzhReeLlUBxV9cySY/U6ofkHNOPmmGPkMkjSsVFEY/gFz
cgXeM81ZocxUoiYuiuI+Ch7QUpWbY0O+L8PJqQfDvoRoM1a1bftwS0s1gSpyYp0j
tFqacnl4EnkfawT4eMEOgylK6L1jU8wVh3fIbCDwlsTNbXeoD7uEKdZrDUcBzBDo
XfIDR/8pI7O96G237a5U8Ow0E+DTRXIaaqJ5b+AStki6DjwOxmeSmYvHJ4fNhMFU
bPksjmhfscRGXZ8a/kVN2M2amhR0F/KV9VSFg6U/qWENOf2xcLq8DXU7HHHmCQtB
ZrKb1jUzaF6vNdfuxxP4jVICD4W1NCLHiwxp6t/cFTKb20jfr76rcniY9u9eQ+HF
jpnLn37bHX7z2CbecMTJCE38rT4r7ye8l1miEBYbKGng/t5qOCY/NS1U6Y7je1NC
Ff6N1gLBVI96J+XS+BT54z0QDmmLrrZaqUKALmNscuA3ni0RGyttTPXzNZ5NyYAV
X3I68IXxHE8XBLZZ/ukGS40EhSIaMLmMJqtNOm39YBM4JyDk/R7Fn7JUmb7117xa
YCiulViFmdc7f9BwpillcSYu8RPAz8gR3uwqea3jm8TYeUWguaKd3pHx24cQX26o
hiVcHH+OTnoIq0BU94KPSaw+69zns3ATxNkxXQmvdfjeek6RDEEkLs/gK1FfxJTw
/AFB1CDchtyH9XRXcTCelUwMg6Nrhjo62XSJczkTKpJB2ywLYUL+NHms6HkNAa+j
hH6nRWqaQZHuni8CvaglsoHSZKYlIhTrsrj3gf8YDTr3eSXwQxmfYMAA+ovrdwPy
6QejIodqO1u9g8TGKIyoyffIdzyyp4n4MYOBFYVjZ70UVkjTFnhkS4F8kdYfoR46
Bj9/vIjQib/LgMkTCG/dQfrkzrp/D9gor6V5tnW3Pm00He6Wcwkjvjgq3+tNYFzc
2Z+QiHE6YuLcKIboiBWJI713hqzdtd7gJrjMDWJMWd8henccJ6ZTClFOXovB1aAu
K6rhw1iQGleQcNt3nuCSXpMKKDy685Bb27J1PFeEKPum9m5CMs8dGj6XdgBC90tM
/M884Ipp9fLinmB7UaA2LLhD2Go64pK18sWLEbOivoOBmnD7ciAlvKSG9/FUt8FZ
UgLt7DpeKsLLSXLTBGVbK0rgfN1TSyvsnGi16qLzXOiHS34T5e7MK9ADUmbRpz63
iAZUve7zTw2KP9YJ6Hh5OS5Ve3X4KOPAlfh5xtOzEx0lnHCz5EAUOhUUqP8WP0bn
mM6w2cP41EFh5G7Ya7BLNBqV7EV4Kk3QYInRf47OiIUph5CNNnE32pbcIXvGWcZ9
goKctLkHG7I0FooSUeVUslh2pg3m74o8ZVBkH9stMCJ+FYbG2Fk5nENzWzs3phOU
Zi+VT6rdXFqID1YP9zGnFErLhPzbcBjCj4OnlgkVsuRtCu7oLkrWAgy4hWIM0DwF
+7dvPpRQTsLCb37LmtBMKR1WEFEN7232S8VqblJelCrhyBl0IEhkUgKlEvqMCH4z
rRZ6rk0PyE+Q/kQmXL6GOZXe/JKgq4TkV5wZVBEgFRTC50n/ckGsFibh6DDnYGbE
mXAnks82nuMGnWtZEPWS+12Pde+CRF4hZ636do3rss/6o1MbdF6FlocP+6mkbSKr
mftPmtJK2lbPAzpUCeJqP3M3cMy9oMC6WBs4nGZMcDmaqIMBHf5A3QXIv+q38GzY
BHAGh0gcUHkxyce5QFVL7NbQSDHxjYVgGTA/pXXM4Xdkk5p15BCDwSGWTN6AilIe
FSiIu0F1rO6WGr2h2h/GK56x4Xby965YajXNRqWWMEbq3Dne38aXp1vpcQq6V7Nv
nR+WTnA4F/J/5mFuxZanMHDj79tW2gHPHgBM2dthXOyQ7bRUK/UX+zFfarcxJ8YN
WADkdtcBlUea6BXr/asBdOx/CiOEb2Jc45UJZELjnDg7k4WgQjKa3vCPQT/K23h0
QEWTqGsrREsDNUVXMAGg4pFn+asUgUaeLqHHTgyjTbC6HGZUYU147qiKvXowiH72
NGk/HL3CiLvPrcnJ/0te4WqKtPo5QBjFCgkQg9fwGu9jObGaHo6m29wMONE+krgC
Z7LtEwDj0mVMZewcSlXGPhtb8abccX4LUxrG6u+dtpvOgDrGJdlEVSNpmSlcGB4B
u2zXrUW6nqcMcojFUwCoNHZMh3paNYWvYhP0vBQh9AUy6OvcOADxNtXChC3j49CR
rsC4R1an1B6kFisWn65stwyOvd8tAvw0hZLxkP5pPk3b8WIAiOl4rZ8MceYcYTMR
zW08efVJxBC66SvpPt/4MiWyegt/8Hhd5XOcrhjiVX5CbFBXXUFEHmjTJf1jgRQh
X0EZmT7dAX9eeTn0ZkmuhSQxVBnE7TUc6O4U3zc/nZOGRQBM2eJ5qwXsxrD9i0FZ
h86sHbEcAvAEAMjhHhaVVZQb0Mc1rLVEpReS2ZDCjovmj8YIKQ487AYVDl8kpYjI
sjsAc9hZK/dH/6OaM11S0tEodi2kWBqV2udBsiiXQXxoUypj3UF2dL0TNzPjQwUy
e3f7VQ+ZEzfVFoWfDnLHVQE6Ywp72wrkxElewHc5UJJ4czdm91I3O52bxnMS2zk5
5H2UsWjtZJrE+P3e7XLgcIh/C9su6L3RVDeXUyJiYalM46kBoDyvw/esKRe2WXXw
eED+BSE3twOMUI2+nc8HtpQMEvwyHhH1FDOdKXKq6rneZRrMyQ9p+WAeolrd6iRt
R+FktzIcJIqi8e+gsVFn5GQ2isrQhwzyOkJtm8iRr9zrX7tkAW3fa/V9dv3dgd60
gED1C/BcX8boMg5loW+ADCLj1oAs4X8cbjq8NOTxOG8SowS8lU14yfSlaXfkH5Gx
727J0elfjm2KnuZl2mgzsfNNX7HnxHq1o/n+AUpZM6keMlwtOrLjoFWgCsWv77jL
nSaQyl9wBvoyGLN+9kygX1NX2vrg/OcNlKfmUvY1OOdg+eO6wb303spDFtAbAGx4
JXJ0/y0IklN1ueHK/KJDbehRMbNVNzI8GAhG595f+Vq1i9eQ1Qr8sDCcFOcF2F5D
4mxhMLS44XyeWvj8rHaRHwgukfyUUCVpeToGUdUbMvD8atcjBZlsUQgzkuRhoFDQ
ZaEdqY7GIyOPggJaJVG5pwO5xV7uVC6k0O56z/PUF5ME0T9wMuj469Et0C7TLeYc
M+eDfHUCRKQBPcK78D+wSsk4niNh4f1oKxe69j5HjeRvH1/ssEBLwDg8boeVIoJ1
ZDBv9QqMPlbNVv2TsreBJhujRb4F+nmPq/D3j/DT7h8QohGi9FSKtPxsqvTjlawN
NV20HTnfHRV7dCNNKrtsBRjxWM6bkA/yIHru/3ZzDjnWT91xXbLMGEwVIMYJ+LCC
M/7XPiu5fnaSzrBwFQozFVHouC1qS7xYvt39AvE/wAeIJUI9m3tTPsHOxnDakeDq
JRySyPsikSMy0lz6NxIJT5iFXSDOnBsdJgBhJpCAXBOxsDPCJXV919SqHGLgRQgG
dTJ/W/FrfVewxdyEYkFXENxz6pBa5bOMd4FoYOP0QT1spBMiWgeIOMYSrFf2fO0W
crmvbaX+d1QXqdPugk5wz4QYqT5k3tRAbgxSXxbps3RiJVExlO2tCDB4mlNWR0GO
QNhB67UDbY6s9Qn6/1zUlfywQp0FlfdBrWVPGyVAE6Fn55XJjTVqO+KOSBIpBrSO
Ucmw93/pYZnqGQMJamaVbznPbLIYY2+V42MQSDZ6QvHieHRj8aIHx2AE7eY+zY9U
ms3LghPVqN9E2bD3W1hRf7OhnlEYB/We1x1xYGgMCuzu/vxfLfAvvlz3MPCZwSMu
rlaKgXN5AMgUzfLSLSVtWDV9S9bMapIlwB17oM/RlULxKZFaAd3wCmEjglv8jP5E
WELgyXyIrQg6VoSz9JtI0ci5Re4yntCiVaFC1UaQi46n8DOn4/GJbTmF0Kp/FVvm
u+iWVvlM5DekKCTzD6Sz3tA00I6Qjqn0q4/OVuosJEI8SITtE2ncSuxm67IPQPbl
KD0y3NnxPQo1E/6ZgQJpY9RsmJTjJQTsgT0B+uee7LEftku5hCEFQir1gJKVAeUw
1ciedojiRdAZVOXr3OB2AQXbOzOAQpWt57jBZfzHWVdnnNwZoXHrtgVM0o52jNVr
eNWfU1J16YgNGRt2o3A/PLJlvNeyB5a3r2Oyc+CD+uKHTpaOpa+XnVktetftMm7E
gGbFUxiTl436PUEfi7ixsK8wDm3Pv28oyKQkXoSERdDvPLnbESCeQmeI3quVIp/s
wP8LLlsS2K6dBTJI9fWCnwC6naE4B0KFUCk07ffIborf5XumAkza6xbA2BhtlLme
Iqpl5RsFoG9DjSjXTtNU+/k9MUC7lEXFD6ybKxHSWUKS/O0niTRSXB0xNDSm23Qy
TMYEV3Irovqu0nEn0FDw6hz/p0ZXN0QOH8+rBXq7Ufbff/YDjcspH6Tx8fBsybb7
swm9sErJnWaijRjeDpHRhmSF8KZxNllBsZv5jvOPMOyNCKG3Tc5ZYIpDZoprEi3e
MiIxmnhCPylMPWH/OiKDMP//UATdWhyE394G2R2dOX9nj71Go24nHWW40F3v33Mi
4C6i2NB4u8MnVXIwbRaITJRHrii3ipvSE01HdVtWlvZ5wnQifiypbFpeCLvXBt4Z
OzDthB+eH/G2g1JVr5V3+kHIu5m6ff9AcyTmT0ciFjqkF9jwMu3/yNowj5yQuiBh
zpptVoCKMwO1C37XrXGG4+MhPBQCflPtuq2yXc0b4RwPcjJMsyjCnFk4SQ0k7yMo
ThdcJKw3RaptrGj/OFhGjc75TTf87E2/z+fjguRzX8qhMwBdeBUyrYUdCuvCdqLf
qR2G2i12Ypleep5Dx2pmcccgkAvfr5e14wYu+YcI9CMnBqKYuD8HPzeIb98FHhnP
14dqhRngARVA9bRh9Z+sxbAEUlCC3Okp6LvwrKgGufSR4NTkn2FLoWzjYsXAsBuu
jJyYp1FxQzMmBUYP+18fFDmrP7iNdvC7zr5Uq06rL4PijqGlp5LkWPshE/hbTXOo
6GBdmhHHtH9XthzDPtKnILxFAf+rrPp9X8wVJvHnkTQOPd42g6WxAFZGMlLlASQl
kr4t/QVaJCo446ACetmHdYm/4T0I0HS/1yqWaHCB/FlgKCuR86UA7KLZzm1+YffO
f3aiQS2xXSRPVfStLEquhDNDM3gzhufaCFiFdKprVNK2c4IErYsCl2xa9J2hIQWP
o9KZkJAnYiu+9qtckWhGtxv+EtLZW1pNgCYS9bV0cD22YHP6OVilNsQJSj9BVFgs
4P3WfCtS8PuhBSLOoHrRGOcRrBgVyJGQDjJRsmEc5BFsSIKXlzB2mIxO//4Cg/xQ
ImlR+i5B9OKfhT6WjPRbuOHCSFyNyRSXGEQwXv+9KZ30rP0hB5QrPKA793Oj4ieF
AEPqyQ1sW7KwBgFW0gBddEaxJDU1AhPZMz1pvsTkMrw/hTWHnZDecSqaFW3SCDJk
RbET7TifKgQ8nwCB0AAM8YfCJ61xlsppfyIidQjUBureRzC8+vJUb2VHHs3FE7Q1
jvczrzjo6TnIKtjYHBw4sYpwMF4NaCX0OpxgTecH0qFX+7D24YJamSe+oszMHzH6
ZOyM2hmWwUcKLChzCkx3zbcMA9xLH6lv0/7yhgpt/NI5xZ7IPUoRWeSrQcTOXqcd
BCrNRLRARw0Q0WenQL3aHQAXHZIJN+LbITZ0p0J8QdmxD3CDnHEA4eAFgsaEpE+X
PGZTKTAUnWQAWaM1nZQjt/fNNrmdlfb7or4B2eH8fk1o/kzDWy3jZTZww9WAulCB
4Xs6s0tirUHk7aOOSQH+hymQq/x0u3DVWA6KOZ0PygUy2gAwZUSkSWWZE0ktevvG
rzQPXLIqxliQGYMyIWGsl98Tf5JsEs0UYVi6SugP191LpDQsLXXB83fs2u98pT+C
2xAO7IRGi/1SPk0fTBdRdNUDdi9vlp0M++htt9xNzwaZkRy9AewomgEd1NC7pTSd
t0lpmJFe/Ky8ry/iCluu56dZvbrZcx8fgw3eXhEsxR6mMX5SNl5fqU4oFhx63E8N
ofUXB8vu8EZggYoTe+MeZi08qX/znp1r5Jy2VlXQ+c0+s/upRZHs5al1JSqWhViA
YIxtJSKziVsmLePhBoKxBlaC8urp1aCSB2J0Ddbzc3+TpbFE30QmhSDG3sqUq8KE
hSK2UZftuFvbEVrql1yFxZ3XgE5vVnpREkQWDGnvTtr49Pb2ziSrVPzQy3mVdaKO
LyTrM/0LFBxWddPy+t6etBl2jxYsSK9ohUzbRCnmS19I1gQcPW8ciX/eXx7kypdj
DcGMTUVdU9DZk1Ga/Hn0Ru73r5ymjIcvjOZddVn1pspSNMt768yBcb9X4fiRzneD
e20+OMRLDVNJTBcay2PObv7rwu7zaT+D6VPejxqmEspSUugFXOkl+SEfJuhZnNHb
ldPTFoBs0dHM7+4LCtzqxsozWRxA5djxAx/iuHdSH4FRKCNTUV0cdhB/n3wVY+qB
KXVT9Jns7UGDGkrcOUrWr3F19NFUGqk/rEwbqRqAunb6YNT8KI0g5K5bUQIkoU2S
SKpXfqcnPDuf/ZlDrL3LfaRlziGk7WJoRknm16PFh9jcLExd2M8FUkeSZ+HeIAaj
o9YVsW9P3mObshucCXlVhHTq7rj/wwKFvvIKOCHTrzPZZGj5h+DTOOzxDz8/VkMV
b6g4a4cAzc3SuI8J9+NSAhyi+W/2E5m7cV255xezR6T/LxxoaoNESo9I0DoADVqc
sSMDWlE9HKiEiEviU9JTarVCHGUnVAysFQYkwFZ2zC0ZY2/CK7bUcBBuA+1I94+s
AlQvPcvzhHch72a8FcJtI3/RlzZ/e8BS2tY5tZOMvAhWq3s1dboZ/bAiZu2IKWGv
jkIrBxbdIqa49YSm39ggTuKrlFnADgnJBDIAzxJgzVc3W6rJov4wMa8Djzs6ph3n
VqRJrDz+rEbADO3L0gIG16/f7nE2mFZ80/t6eG9HH1UJDtES7gZM1ZdhzfI0unxL
rM3WAGrIrU8W2bBInwjPoZa1FIPAuQHjaNQOsIgsMR0kfNj8nydyibaTnw1CuVrA
0pbqj3AadGUxIA7BvBrs74Sizybz54F0NngYIfNQMUs9L05dAFrPmRs3qDzMadCz
ow7LJx/zdl9Zzl62y0GkWgP10MluKDOXdtFjpObb9jTLdO1+4e/IhyaXKXQ+5i9O
zkZlDY6gXn31zTDWDeeIyIdCuztL1i+Bjc7bGKfkMdZoG3yjpwD1VvyQcYwEhDCy
Zh0bVRv83w7+SWzHb883FsWCAn+IIeCej5REQ3xqTe2EAnBswUEJzfb34PgWz9xU
w0n9Jgjlh8SBpkxKI2IQxjn3sm36hdNa4vEvPX58Fi0nR84vto4fAuZMCF0maTlj
Og+9dKIszD+DtJYCU5A2nnJzFjO1CBjOZeGK9TK3fnSZY4szkHfN2acrACa7iiEn
t4KKpyHBRXn5Pd+9e0AADez7qJPv2slaRjg9/kgIQI4P5N0H3HSYVoFYj1xLWI+g
vvevP/r0hKZPVgYwvboCBI+dShWIgIsyR7eopSU6UoE9PLIA8m/HF2LnbkNxeCQ1
l/OGj8JhWsIySkP99Yo6IDesUB5xuGKqVtASIPsDVpoDp3gI9AdymmWRl1i9e8DJ
ZLpV6ucB9tTlLAyUyrSDL9RxUQHEp9HMRPPRgP5ULWMRD5RhgG/vfAqVUX3lk2j9
sGYDTWkhyCbwlLym/epie+oLEqDv8DZMIg9vgHKa1MflQbz+q/UWbOD8+dnZot/K
NBJOvIpS2R9qTvjH/3+dgT3JBISnd+ODx0kWFfoQbaVofhjln9Qs7+7QnZofdBIh
qgT2eTtnXxG4pWjAGChjjL1YGEtsRyXr28iPICTOx3ioyeP55To5iCau012csk6b
0EVL9QPIsrq7V2Y437awrb3KxYIwzJprF9OasPh2LU5AFzB6b+1K1eQq16HIFBn4
n15ifJ6VRJ7ztVnhWOuLa1tYyK6lcOdzOJep6oytNWvy1X0WEZdcaP7Xg19v2SZ8
p4D7Spw1HXVS0EaAyGWNCq/5Qc1/FR0hvKv2NNg9Xo83m0VS4L6ZEJQqesFDDXeV
fWR0FDT0QxhW+RcswaPflNK/co75mVWO7rGr/4sgjqu9aqDdn4Ov9mocU7/hyu2/
MA0lh75r9N+OoOewMucxYMYCnWlVmzCsXemI56jtSSigJuopR8kDVyaaoJEeKGug
Z97Oc0y+M1XUy5Qgw+BM5dR74M2o4BKGSC7Owb/ukilSEgwULI/Z27l5Tj2fbBG2
6+xqBWyMbtyzP21VZ9kAycKgKLcGGzner2AvyDcFayqC/CsSgpqRw/I4aeWJvl3C
0ahnwYCqTVFCaxgUzoJ2zNqKRJqzDHWXEBI8Z4Dmn7cdmTSUlbgDTpMqKSm+LDT7
3p2DBMPJ0DJTYbg+mTWiCPyJgqBLeIf6Jwkic8p2wSNsovoV5nyq8i+uQCji8tpZ
BMhzE7STXd71OXJTo/wp0KpURlwTt8cgtXoWl//gxSkvwlI0RkuVBGcS6jRtEUMt
qIuqcYsbyz/nwH4hKsJYmvOpuGo5J/EuYgDTyN1hbOrCyKvFwBklzzYbp0bOHYoX
aa/lCDuP4QuTm5H/hu9sQBr7mIC/+e0kRpZ3Q/cn/+yWAKg9zDJvLYjcomm3ohlc
OHdRgW60PGdskuHsmULepq7F4bh4fSw/qE2dThRW6T/2/eNt6UyKsj12YMvISbn1
SbgP0B4FH1Va3niiyfd4Ws90MCpi1fXwN6iXPhLoZXPdCG/8sB6OLUyihLlGy6J8
ePUvK89Yh86jfACKWJyhEFogwInPTNKZk2Pvb9zTqk9DajEe5RQDmPhZLDlmDEva
rywr6t9NK971STAzYZunafIgn6joo/w7sAF/4RMPAU2ojiupwPEml8aJD8bJOo0D
Wgwu5M/ZNhedqWncBRAC9QVg2B5iJsK/nlMAbLk0QsjonnxYfQw4p+gnacFfpyUc
fE+z7r37qsP3VZNRZyY1vSbf9ZY08FA0Fk6DGxEnzsGVRkEQvvNTsVAkadHt4EBb
0WaJ3NakFVLaYl8nmW1jBlODzRv9aq6MBgU7yAz9iJb9qXd1QsKBfrw6Us5ZZ4Kf
qzwKV515eS2nPRYFbTASHSRM7r0zZUbI8O0hhF3ZGcw2Rs2MpSIIVfX6FZpVp0rx
UAJ6Asq3zzEXhNmP8ckrT6WUpo8dZ6tJi43Pp1zoiHqKtp8fPJmz18jEQpUU+VQg
k5yeYAjO4zQATj3hJF8H6XQ7vGuBRkHiWZ3BH5VQomf3b4ghHwT/drcrMM6Zv4eZ
UTdi1wWMrQ14PHkgFqy1tXIadG00defDbUel8+wl2iNXFR4Ibkykz8qpUAtYbwA8
pcmuKiKbg61mUQTHtfrwPMKnV8LOutkPqiCtPaIEX8rtQfyS69TzRrFB3tR7alx3
SeR2ttZ5cW7EVFKr6Mf46MmjLHWKfh/LEnYJsvEMdTpALqB1dMGEa42oeiwKDitV
SQVyCsU48QjPaNhLKfXFp664nwG75gF4fzQDcopZXvDGMYvulgNXnoK07j1qWmUC
6ervWd+eIrqs42mrUSFB3jR19EpjnXdtV+gjfsD+RxmQsH6ffU7UeFW/SI5wsdkQ
BcOflK8S9p0uRi7uXYZTUgDflGKeotszPxQmwbb11OhJWSXbp7bR6ETNYOccRyFt
+l2hnwrGRnhvFBm0Laa9rDxidRzCUy1ypFbs1r6sF3quzPA4iRMEnOmJzGyRJIm6
4SHPDiNG+B5KgRubKc53oO0i4bv1cIsOXpv3/R/hfKdfW3V9kpLnqsaWEyF1XmA8
t3jaBOth74OcQmJQF65LohOhYAytZxPwnOpKLhdxl6iF9yCNoAEKvbecrxqfmLhl
8SLMsxKcovVV5qxuhIb9zpICFSpqeASJoqMl5DA2jNt3UvdiGQsbxerpeFNKFapm
RxmLd9Gbt3MSW1ADhK9Cn91hcvuiVEsnf3KJLATROASokXhTZwCsx+f7oOMTmI8V
jHM2tr+tCBpnx3eJYnRkGF7KBtSj+v21rKZ+g1ewQCygQBV+o27EkOeyUc7UKAmF
uMQ1HeamqcVj9GcXp2FTkvnHaIsYibzTW32Wr+Yqpc/Lm+tb5A0A5dsjTthupWbh
alfZwz4cGtFQ0yWjTDc1otMhWb3x388toQwDH+Wd9WeWpPQj8IxF4gEqYc4Mgmli
0G1NPOJhZfVdGgoNk0NRP2wRPLU8kSqg5zbgZQSfBnfOttfcyPtCSObo6mbIMkoO
QcbGrdUKDrZZrOB2FRIZyybns5jTI8B3D/6Os3qW6Uzj50KbsaBow7F5IZ7OKXKu
sm+jpcJI3BmBvZtzrXWnpvmBYw3lkHVwSp0ugu94qnndBgIRBt0gPtfJSrk/q5BS
qRAnqiDo+xS1d1rs1NsWGhSmgskBmq7fBYoJ9YTcOwDTOku2j4nqBRdH4d5IlBoy
w5kqbXijHkrSacs9zv9aFGeT2LwLRr8EJPn19lcuUUU0aZm7Y3FOXp/GQFnntyd0
ZXLwRf2XM4Y1a3Tm5AQo5qNWtcQYh8sGLfF4Q951JkvOXW2rokypGSkF8Z1OkoQm
OzEqPu90JuPr66g8KGaDjvf0VKWTzecSF75q3bBBp2HDPKW4qlFIW6MzPcw+YsY7
ay1IrWFDb7BD+78bBvDcgRuAIehVZLbZxayqCoQt4/M7n+M2hOaKTh/YAQaBktUp
NbjxG3+Jl03RRkky29UX1z3iNzu25Em6sdjU3yc6//lNDrPf70J7+gGiDFrRQI0U
mudgI9pxUniptsYNxrbGwtTmPBA6xkFagIdo82LNQtBYAYFXjRAVFg8IVAQln1F3
sZBV4Kh8xpBt0g08Ic3wBdFk0kxhp3Kw6pS6fUslg9zdIZQXasHSHAGVzt0WTZRf
zkIdiko/SSzHIkYJEVDKD0l74p7PYNgpfSXQK+P+IWnzLSfPziJUOsze3UbTjQ2I
smOZphHdsvN0X8Gft5HWKdoBfRIXk0e6EammWuspav9ril+hycppIW1/bQ2qjpLl
WhlRApmOtxVj8z3Wvqba0yuKyyC/4M2iXxxQQzkIAXqsl/ful/nmDggWnYvSdA8v
jqLha3ReXst5vZGlHF/V6opMml6LEAHt7QZwQYdLNqPj/XQn973x53e7sAlnA9WS
1uhsnlTNVPn0Of63/bUrYMs5sOvf4vKH5nusQTXq/zTSZawlFzFpzOUhI1UMUPCz
g2Z7qFpsWLpMvmcVXgVi4/WFs0hoBFFCxxrI/eCz46ONktNV5vacwjq2tzlSlkXJ
fB5dgKROa+12MnOPER/rWKpw2pNQqj/DVT3SkoOcpPCugur0Jo8HaRsCDZOkws5k
W87aCkGRjcmsTkrPTd9G+jQynZSCuTAM2xIBaYjmc5FtZpVWkUbjbG715liEkS3w
FXGZh9PB4NoGmaZCS7FeLPUttZJR9is+qyhJuM9bAmwxIDp7Jcp0WQ0mfXneLp1P
S/5hjuj1PFZG71axCxM4QIAwBRX5kuPrHC29s5llMovPxq3nxGXCRrkjUzEO79s5
jjr9bC/CYsasehTipqYaECHs7T8zWcKCkJNSC6DiX3SJicFhGn6nHbHg1EvljQge
Y1l0/D+kN1d+S7fojbwOEuWHQ04DZcpZ10YDpBwuIyd4/xmT1Z3iFfbzF09s0iGm
n99lfKiYNfWx4W5OyAsiooqYwnxAaICuGIW9eE4FPgXeKNOnRMEOReyf+Qo3Jic1
DSMRFHoJFdWD0HAK1IhoB9zrdeQbwsjUbMEojkDiFBan8lrxPOmelpJrwinohYkR
uVCFKnuLn99iFATEzX29WHSzUXPkcjVacUAXkbzCv3Cv00gbHRZeQcu5OsDWVjPZ
bJSWoYv6HNMSsTqExFgvo4QmqmybvEfLmbFva/icYg6i42KCu9PpO5cRs0jCegSV
cUDZocinRhtCwJuKq7jeAnJS3Mn9BBCUQxUzMtr7NCdF5Nxk2sBZH6cpgq7bhyK8
g1lKt6n6g8tUsDhA9HvgwTOTW5n5/n8oU3OYe7SL1BBNUfSL87kk9mdm9Mt/NK7/
s0q7PKlpbhEipmyVowzueq0BNXAJOoli/e9rj9IdtMAePA5JqjtH0jcXrAw0uxJR
BboH1T1KkhWIc7m4Kzc/hhxDLPWbRk+/H8TY9la86FGt//rDtsv74LnT7k/b3lU9
wtlm/8pBa2S2XiT4i7B9StC8aU8lpeCmY+feDnBHFSlR6SfxGbJYpw5VseAKZmHW
ZRq8ypT9qytGqGUtyx+rpYVwa1MMM1rZn4xB96AjSlLPiJRm5r/5G+mSc8n4/9rx
TfVKkCMx8Yvzg0kyZwEpVSQ0FdYZsmx9AQRBTO/fQbu3PsCqviO+1uDWm4Ge7Ziy
BXBzZziZ1o4opFY71MWm7Z3cdo/GP7jshs8g2ITVtyZq8rA3wlWAUanOoKtyjUH5
LN9ZZMdUCfTidUAu4mergPi6RJkQFpnv4iimgrFyEC8PMb4eRLZk5oZFb+gpKw80
OpphbTI1TpJYMzZ5/xmLLx+oTOa6dbLD4G9x8yip25yxC334ucataNNTRtHdZ9Xw
Ile+mho/Er1ckjb9LF+36zLnXfTzDEr0CAWpHH/FSDWBDZRQSpYwotD10MVEhPqd
NbfgCV4MQvdAAm3H97rGAs+41GzU40hc1rWPLIQcraP+4xRQfJ3Va4VxJz8VNWEM
ItwUS5UnSpsmumU6ikTcjrfhwcwsLjNcUitaJxIUwpVybn7zjIrHuH4mBEbXYBEE
B6s0oxTcGc2uMQueBpvqVJRGYO0UcZmGMkWSxdSDfn7ZMweUO7K/dI924ZdVfZp2
L2i/oAfrw3XX0+rX2th5yIyoAdMtXVR73HOZQgtYTsjMJy9o+cFoe9cOJfOdsfPY
I8zC0pp99sPWOxKgpejH6fI1BpqpcjjBxMRki6iVnmj3Oh80+wqvbVyaiU0VbxhK
XTaHnY2hkYQxPL0wAnHR00jzC2YhqL9CasQIvb4neZsv8VIsv3maYWR7zll1fpDX
OnCSk9VhCQto+58rJesXarZcxdlVsSK5KwEWGOOaq9wz+tkpwoIYm3pWSCDT0Gal
EUfxcAVuV6LtNWf/z64lc2I5yLkPKeP3WEAStI1vwojsmy2BF/HQsAJuNFEspzin
jMTmH2iETYzIlP9N+Ipcg+iPZ8NoyqHCvhjJv0HTcFgp9P57YEHoLaKAYsRL3eu4
FgBRMyDD9PSLkiopnpC31hJxHl4UOcNQmcWDaL9aUqXgGi4vSwKfSBbOnuQN+vEr
6aItpN3x9LQieaAtwLOkACSSrAlTRV7bm5F0WCleY5f5btR/PIv7z7TXPXnm75YV
LNHB7OR/7ad6uMTKn6WDau/yHBDWem9W/SuN+t8qMMC+BcUch07nDwJK3Pgee8sx
TEcDLWkMKjtGE6JHMV0WjQBaMU9G6bPnjlpLIGRAzKB/YlWvHIcDoPgooG38yRSO
RPDvhe0oSYU1vgJMh6+GJDSqjroFxnz9n5SyYCgQXN9x07WiohJzyRtk4w0MK0pe
NhAQlFC9FG1QurWDwW2iufpWqraZRIChQA3XcEbmSrB4BBav+GJNZ8QDSNZxzlrF
yXvsvQnAvpJyqPOpTJDQv49Z4O1dC8nxjyN9Kir+age/1mYgSH0QF5xfY68Zcfgy
kPss1rWGoTPQVg+V2t2wPi4mVvHJHFfVvdZZTqBj2R/uDnWcR2H5fCpvwbl3KU43
fm0FEhT4NAX3xq99DeFD1F184uFY4QPzrhmQcL8SoM74WJ6Pcej1HWmFHYlYbIYI
xxkz4+G1tH6cYOZMOlGixFZId/GtTUAE6CHxkJyJKbrJzf5y5tDOCdDIlVm1ghon
p/y/nilFaz11Y22F4/0DdCdK5VO+T+DyLJFZdp5kzCSR/Pp/B0vgpAu0mBbTqRcN
3YbVFGRr15CfU/RCndwbH5oELLOGaBWjjHAJnor0DEGEG8LfO0pdA30yRCN7VPIC
65gMiBBlrtgw5hWIFVoAtQ543wfy04f8eXNTlb8vywfQ4mGD/lgXooFu1QnwN6Je
ZL/i3g1gOp5M6NQ0yGE1ky7MXMJ/rZgV2Yn1UMmdQcFDLDcDtFZyXIy/77cu5hOW
DlcUmwnTGhpMthWxcbZI9qNIrqrZLCD+csddKgOiBE85XEY2m7oHiHsPPBcVoqLQ
DUS0b6OFOLq4Oa7MYiMXKnpfOuJ9TJh9f6O2Yua9DPhKQQkTLOfLFwwXwlDnTmRQ
vDqmCYG5c2vS/0CfK9FmLSimSgBPP2His9PV06L5qD1Rn8cM7yHXIr6452LOPO+q
v+GgRFUx+VxKM1nhoDmo1v5SIp64hLYLjrLEeu6j23kNvlLFPxKMBaNATuWfUReg
6JdN5I2kkxmnA1JqKiBuunnXexETno8LYZCSrv4Gj0QKuekzm/tNqOWGGWBHi6P2
U6VLy4kBhRm3pXNEEMDTnVDhqVOUXayUkKQ5v9NVuGqj2BmWKN9OqvsMURKz1j1t
4Yxz1GsBymyEJZgROwC2/3AnZqCLgx7pcW26LXfSJwpKkVK8DSZASGOeKcD3aVDn
XGOfX1lC/Q4pLMC9sHsZJTuK1kRL3PjFHJSx25qFdzQuA/Ag2TNPimi9Rh2eIGQf
DjhbPuSsdd60W8fGa67E9TXpdP9Vnl+TQv2H/PI86UDa5R4YioeMS+OSez8SFHwj
1UkZVyDRQOfW/LRBcyoskZ6vyMBuNpegWWABuJBYrcBDUmypzzlNAoFH8ceiGsvl
mM0lxcgL6v3sen934AH+hFMm+gBQCm8/vBP73PpwG2Q=
`protect end_protected