`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
ddtXksX2+yylW5zu6QL2Lhnb2d1sD00763mmSITNX595NcHTEkwn0zB1Dry37fOW
FufOhVzEJp80NC5qZ/+F0Vk7Ik02dIR0elf3clrjeJRK85K4e3Hoo4xn7YbFUIms
l/8VZSb14+JVGURjfswrIyCUotIzlzVYZ6gzoZwDXIi5gQIBf/gI+KxNXPaKV+PQ
Ufys/12rjO6aI/pPlqSm0hCvftmBcnezN2hk1UeXgOIuKZnogjOsf0iJVX2aOOWE
6pD/psybjbnsNB6kH5uFTA5frkzIzkzl5d9+YDm9OyC+k84E83I/7/j+rk4L2dah
QJOvksSIzN867/4Qt8qYTQ==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="MvBXkzurAa5VTw+1JJ70nePUfoQXBvZOku/SMmg4TwQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
oRtzZL4VJ4iwysPsC8SXYCzXS8Fw2gtZTOskLcDV+1B9Nzn1zTyNtlo6lNICRmmK
ZRVu2BmCc2G+fmzynYlNTnSa7C0Cuel6FYpxCBlOuk3OF2tzAmLAuDyOH3Z1Yjzk
a0aHuoCdIRKv7BrZCdALt03JeUmXKPdOmIlkVGFl8yw=
`protect rights_digest_method = "sha256"
`protect end_toolblock="Jn9CQpRhJt4rnzZPRk+dOpzAubz7omckX1MrFd4p81o="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 8608 )
`protect data_block
gD6l00tciPUa6pDNTk/+tzLxvdHE2s3DQL3/JqqujQBC/Ei+vcAB8wM3doqg5vTg
mdfn9XB1bLOis2CVSfu295W2DNwHfMSTc/8BhCDRnTlLIX0UCJs9Za0+LoM0rMrV
T7EjVWppbP+Em6PkVKCwlmIQ7JKaifJ+Y+kjw9HCGboYo5074hY+K/CBbfsBQY86
h7FrhVb0BFNFA4lVvsm6LxpiCshh6n6Rv8yNRHQIpv7vSLjgD+lc/anLpVphFdDW
oPaB/8mWxLx3M/bQTUDPACVHCWXHvtKTz7MQWBB0ARasV0zW54Jmqgq58P4kGAK2
iP0Fj3G/qzAv5gtwNTxb5GJRKSx7OODnLS62OqZ9mWOjhVkGStcqnDEyLD93unQa
zowvDOt5PP9JZtMYafxZKoAqlk/yl8iwuTpc3sSdxntcwmvJklnfsVPkKjWU7Jc0
YE+jxeLlKMVywzhXTw4z6W8E7hlCSPAHAlXhKFXAec/+3+Yk4MiY2oDBJ+DCr2+r
pOTViD5QEH4qWhPB9s22dBqSJrSd8y5hoSP7lvmS0oeExKKdmn94uvraZUd5Gz1b
aJvCKOE5+5o+lvOzYCK+c2WDnrkIVKw5B0uxucOce9i0bUtwB4JVqrruczP0LQ8t
Rzp8nkCQQxRvTRXYUQ1fZoIMvNoKpG3kh0+wsMeUaz+5Qo05+Smt/QAtVn3mJfsA
l520mnQlGJYqk9OU//SiLsvMafH3gKHWrG3rB0PB8Ev5W8ICy49eSjDD7/frVURh
keMMnV8WCeGqDMpYA3+1er0ZoqM38T5nZaRM+ODeOCVCTT7ZbPmHMVUYHjyV0bjD
KWn02LM1QqgKxOC33XyTyBIccvZRM1lC4zLL42dmxJzRhc7R1UHptwnbDw1pSJxc
8Kmq5tDMbs/6m+J/qPb6QnDZ5x3XFpJr35eFMXO3rldTMp2XPOtSCNR660AzJcxy
/YgX9T+jACyuEd9k3AxELug5TVKkW6GxNRKeoV/adM9EE0BvGzr3VGy1RG4HpZ8D
zlvK77OTuelHRCX3Jgh1jqtHs8r6YNdVsJRZvoIBYa3ey8xEq6xLje3ImGad0Cth
PtV4R73bJecsuGR5PNhnOcpFWgA8zMYBzfwVqmObr9YiZ/DZlrNKL42VLCuV72zS
eG875G5osxCR8TpdiPPgteJtMCIHKGoz5Allt2piB1+hW9oKow7nSBXZLiyQy3dK
7K3grBj/vnypLC3xc2a6YD+tbpgZahGHEZLpGDPnzj36VarEHeMe087VX3gw8IMT
+Eh8FgC1Oa6PLwMvw3NjYs6NBkQ5wHr1x/CBmivwUnfbBmFI8GWWY4Ca7d3roM+A
dAJVyuquyo3yW84L9KU6Z8iIWZnuv7gsztFqQ8xW/GUCNQKai4GvUnG3xFT9ZAe1
l8I0X5FgQ1+v6TdeP7uJEWox/S7GNUWgCAWwkPOLT8YD6mkRr1SexdndInujJWBB
tuq9ADT1+UTY26kPq/iagmNZi7Sv6Jz+c13Ny3zIxsi8ZYiw8WxZU3ysUAo8sX3h
vDp2o2VaYrNk+fBpZPHE7ckMTlF0/nOpU7B3iGdeTau612CcrJjL+j87zhFQebqM
6VSBCfMWvI6sswpvjP95DOjuxksaLMtYo5lQpYAagB++6+KEi9aGOv1l/CbwED8+
wQpVHUX0mwXitrPVEd9YHCPzfSpc/7aM1F71Fga2ikIKr8EqWBsZtpqp3Toct7lj
riQ4eYxl3qwi1iaqTfnsm7UXbZ5kNIGtsscFlSNhKRFUFCXcdBICglE2h2YgK6+T
iUwIFQ6mFw+t+kl3f6lnR7w2d5T8V1wRdCFkMo6PpvlU/c/0FYmKiH37XhcpjJns
aFDLykDvJhTmEuDuk3GVb37KlnA/1nIhTyMzZdKSBaHszstykZS+7I+/zlHC2GZZ
NyAq6zRdVrKvwS/84jaLbhqCww/iFg0NAxFtLP1kDxCTYGbhIABOAs5AM2iimj3O
ZYnyQRJayE8yfBJfBDV8J3AKWkiWcr5NIj+aoKb6qEAJSzXCur1oQk5CVtrZR63g
b0FteeEmK/++CzA18rngFj4okCswe2iDPWrBczxpGX+GsNTFU7Q71FXV5jBIIlKl
zfPgi5x8NtOUXyC0+az+RPYKpruMsF/rDHOdtjnxKrBI+maD96vb5pUXTFtSzqoi
AXw7VCetBAU8Ak//0dbvHWErTqD8YhLu+WYXSFUBxsYtTBxk+WuB1WzHZ+qVPxAV
sKuKgADCHs7Ek1HdbD1K8S6j+HjDldSZNfni2UQPboQq30GFDKMqRycR6vJjTYuJ
LMN3OuvjdGqFv5tTU00Swnl8eAVgfI0fz8d5JrrAPYqHsRtefj/ej0F1Fu2p2oKE
qPb9SpcI/JajvoDAPV0WQiJlCiWj3fnZqqk9xlioSkloq3vWqoY4tyA61Dewu1/t
5+29BV9Y6SNLb67AoVIXJbLiPeWM/F89jYXVd9AY1euJGEkP51QN24+TUdZNmasw
NaMCmVNJAIUjszsOqFH62md19l1xdBmFVQ7e3KXTs3nE0vCE1ELMKBKfaQgxJ0Eb
LxNWsVsLLfDO+UcP8bUZsgXEVZ4rO7rHrXneaB16JL/2gCn/Ywz++YhaxjQsSKOl
RYJvH84ak6/Ou0A2brJAu1aJaP7AKuFs+SikzT6FOL2PJ6LXifVioPaCvl2VK9bu
ghW7/prdeS51PWvRLRMETJpjcQYBVSKu1j9jYObA3iwsIQqiNSWXwdgjh7ligMEP
PKv3IGQcG9mIcCquuB3ghLZLY3OW9eAJY9pfJVEQ2kaK3ZE7ry20ZQ2EPAogahOp
4uPuV+ohBk1t+v/+VcVYBR8TyGCJ+yTGlluHJ9fK4LNQ06cQu3OQOU7+WvbFPu90
ptyQ1IgIwMBJox37DiynL3XJf1w9c5WyotjDH/heUaNK754W5l6jAHmr023ebIA2
LzmYDBtvN601cgqjOH8GG38LCUJXDKXJndA2IzKtKzEXgdyxzLNs2scY2/FalCh6
TJdszRIr3Go3Lanr8gwVMWKcDzqwW+NM4pw1EEC53XXRPJrCYIirI1MpDY36AhnA
4I49IEPLiW6D+qfzMqWcsacrIXkVjplIFsIsxC3YC7LVXg8UEQwWBWtQzeUbXp3U
WyaVoTVgTNKRZ3sfQGRz+8jH/DmdaTFSKe24NjQOT40v70gshecCFafamemSFtIe
hARUvVqNXA/6JNNdH+7LwOLzSoqJoj2vJwLLFImr8Ih/NUVEbEWNYiULPk6IQ3lM
ao7pxrM+dHREoV7KlV1pk2j2o6gW4AoDYqr8XyXI96xvCBFLiXa/Ufks4tPIFS46
dN2r9Hb15j74tgyZNOBT5wa8hPaJH2+FH+5OH5FkMRBJtqznPPaDYgHIUwQMyx/a
z4RaSNZqcqD6dNh5tNZjCrYJ7qpPFK/Do+x1fipLYKJY3Zg15YmeHkraMHew7vHE
QptgmYxbgzXaL0qt0DOPwEGVnm2AyLLAAHkdiqpy7cjOU9YBk8ee8LWiA9dZoE1M
oru4hevPavQs10WMFuVyiVwD+seklAGYbWlvgkrmbAeGAIXu/i8M+Vpqbk2E2Lbf
PH773Jd+BTh1Q5jpPx5xSPQPchTKS58UHSpk4ElRL3+8vEv6xLcWrtB6l1zFhaeH
JXzso2sZZ67IZHr3XmcDRDVuUt3Tw0UAI3+ciLP89XbBlYjsUdfGtL9wmbtz4gvH
Ld4lhxPGmjf0low/rdT369TtNJFurrMAAt1S/McT8bEwkS0a3ApPRN5TbStkedmk
tOugClH78qRX7zicHmB9Jzd7gUsnC765HWhexlgCoDVF5oYEl8DEyVViLdl78u5H
XKXTqQiGjZcqmiEkMBnL3bVhEGm0sn8eedH51JBlpCQz9cectAZuw9k5DNzPynu1
2Xnwr85kKRntle8cgTKJqfaaPpz9QK0m5yThT2uoMtuIqmWLG45QhFqi0KQuxWuO
vbD8SoBFS3y5hwUqUso8QtHicYrePi6+mPPeLq/BdtHYDMUf7yJQHOcnNJS/5fDe
r9Hv8OyCVub6DAX+6ILXmMRKcBdLGRKvkYQDZ2uu5KzIA+APs52lp4gbQzx9l33m
nkS5/5W8XZVASn4YNArPPmCy1oW9I9xH6CzhuVGvvrtcQ0/Yub5WV4J9jMZZ8MOe
p8ufO+orF3gHT/qD0UInpB8L5V+vpLWy47pcwAOgdn+9KxBCjlzKmSn1ZT+bTPe9
nv2lNMeSgAlmlNNSQL2ee63tFCIdtZHpZg6pl1ILz141kV1hQlQ5DNWzYH3W7Tpq
QvV47/h+npaLd9e8kJ9lysjCNcuBJ50+Js6oOJN4XyoUZ81ZbiAxv9vUfsAm6LqJ
zzIRndLwu3Ijxj9+Kn+aVo0czdsCMDE9y2UQWM48X6EZhF5wOAi4I+tzQKsn+HGQ
/QslGG8ezrDSZM2lCeIwjTt5RG0Np8gIoG3ZCQ2kXVCRpLPZ1biHz3hQ4pSwJCcT
weZ7n7wwBEJ2hL7LM0c6rNdt7R8CkiCLIyFDaF0bMxEn1OAwfDu6Oqt6BiHZbjW0
o6RcBIeUcbdUgxd4vVVWXS68USosED8q86VS1VM1FBPi3J8YjHlexlV8hYnBoUZ0
uDFUj3zhpA2+hXN/n0yfyz96P8pYLO8I4UrDkO0V9ORdJOSyc6AZddx8pRC51I8f
8BP9uR/4ytED0biNNusqUKoLcAbjfRqCvTu8G/YuisMMvVw/8juLfMcgIg+4cAgQ
QHxyd1M4aRkvawjChh7WtDFO984hmtCPZ1baZhS7IG8LNEtpowK+pb3E1QXGI4WA
2d1Uu87FAgw1NuwzXvuOYnvR/3ayg2Nu/EX2nHI6TZF696tqqvJLtSZRdLIOHP8S
D5U56N+zWGCxOfiyUuMlUTlxVtRPShnTFFr40QmGMs4rh0mAZ7CfhU+x8aCkCPe8
ESx+Bqlgcqqq6QBapGZEOET4mJlZPzxi00tYEQKQVMXxpE3R4SHUP12ip2c00c0s
lNYH9LXE5yXxBe23mekW6DFJydM1DqE0hdKi/R5N7i6nbaFm0j+EeI8HMYzRDTW7
AOVKP1FW/sAwBr8/veXXdnZUfZhUyNLg0S8h/eBt8z7kMfCId760OD1g98NYWb1A
HFnhMQT5XkjCjeSDK6WxcbESAOeN45SXDZRjhR37rsouBmgW4ukIx7DyYEI1UAmg
iU5fnOqPnfa9nut6vB0FKncsQgoKl+o5R6sRshnYiBwj2HGEfixcbgIR+B8haMrN
qS4Eq8n3IikWGof/6swM2Gshnsp1ElJdKWd9GHmDCXdFCJoKKK2n4H6y3Ex84Ur5
KD0InOyYUMCwmer8yrP2IZk+cY9vb+QKa87zV8JSXmDEWG5WJ1OMfC/tjC729vur
e4T8Eib0x7DmYdrQ0aeU/aR5uKSqaeUfwCynWYPoTTuW7pCZhHkxpuOYV4YbwpLu
8gj2OeysQWVNvbeeyC686ze9/UyRPbMEHTTmd4ipqOu+lZhfp4/bX7QDPAwDX92v
toz8VC1h70W0VCODWjDsHORmVftudFOfmg3HlJqzuR3slzLEoGQ8oaHfpjnG+ivt
PW4P48wK58zsF40DNTJnyxE9rDQOH9Lb4E+93+5hkSnL5a7HiwY5qNs3GnqL+PYT
RbysvN73vpxTDGY1AbYVCULFhTnOm8JDQsPvVYoBkkkUUDVz5Oc65Q8hcAduC3hp
yIdW6q9RAdJc1JRzuzkBYqwWuXAEhLqdU4RY273mKeQ2NsFWNVIJZixdQMIXChuM
S1zRuAQ/JKmkDFsj11EIrQFz2iK8BHFrVWpD8CsMVn7QuC5TVXsjvJsbI6cgeho+
X6BB/cpHCxsrBTDeeqoVegfO6TbgCkqi4Det7aMNklXqaJXkWOi0PpoUxlVDu+mV
7+rXUubsEA7fjd4iRFS3d5jrAkWuENopS17rBt05K0ta3CkzPPRqBMEG1KheZ8R2
VbbNgUT3YpB9fuDVGZi1hP647BYsr71/jTXo1xG/ChrNRdznhjpd6RsEJCmzOcHP
c+ELVy0dU21pIpJoOKQgcuJN/dNRMrn27vvu//dxIXn79z0O8ST2ma62bvijqZtS
7pysE2w9GCoDjE/LQO77kFVOF+zV4llmDpza3bJf587Qc7tJbDZNIaRchJHy6pmq
IehjnqtzDacueB4ZMQ8wgk8QXEIeXuBRZybNXFKCIQz19ZjGDrgJ64EN70XRB0Rx
Ktvf2vZKMv6losjNVm/5F9mJ2Jb4yZNkgCzmtmIDAXG9CVcyWAgrNlNmpOBrMl5b
tr0Uj9SBG+yZCwK0C93sjGEpZjhaeTp8hRVbglmtRBtaw3NrSe8vp4kHnUHNs8gv
wCfbjsOOol36tAYlqPdzUwz4Xd0VGMPxX3QwkyxS0XPwrjWo38BkbEiVQtwNl4nw
9QqyzM2kJdRVHsQhMW4xUwrY6iozJArmJGml6ru46Qu6MLQoSUDKk8E36A9YoU1m
BrHYDy3R0xQHzbZIT2+4gsMdEO12OMysVAhJnMg+U2Kp27mZ5Zlr9xie1X42LB80
K3No3U4Tz3YIPIUEfV3Fwf7PLM7Zt30mL+tXWqSLlcUICD8TYpAwaKFR82vkDeR1
v5RfmaOc2UeMEQKlGamUJm68ufKFXuCRgY4MCZY74IGQLyn4FfEN0946xopyf0SQ
0dmuAf8hy9JQ5rd/1Qqnr/1996BLRvQsmSjSXPPrSxnoxpUC08/ICXo45f7c8EMe
C1htHUNYBFMupml8PB+BnqFI1wZ38/IpoBJ77aO0b3RLKWa/DWW3fkkepzoGqS6W
YOXYX6pgBEcx6PNxXr0GxTydhKr9ZrpjOvBTqXcN69gSBM2W+daqznTwB3ua+pl1
WFjr2Hh1qqI6zJX2+RoxnuZtRCfevKsvgYK0I1OU/P6ZvBAzVxl++fSaNKE63tmV
neIxcA1dhLTKOZuu3Fd6smmeInXl/pP7l1TSR/nbAXoaUnH8HDJzmopSDq/DNI+t
8ZRtrKBmeLfURctHN8lIgZlnX23b41smKWZf52WX68rTI3X+u3uA+gBbidqRI00t
n0wHa6iPe0xdUO86dLaGL6+ZJx58V/BoKK3XoU873zb23JQTzUf01cYREnjB6S3n
uydYwxXXLnDCc0DIqR9uC2N01PDyZz8/rCdrIx/3p0jhHWJCezX3xk0vNZ9Gv0LN
LXJTaMfvIepw+wuapcLetrAthZ/CygVbX9WZKbzL82iWgasgnixJrDzfkrtDGcB5
QSq1uz1p7n14hPHJWh0VcmGn1S6wDv/kW8Ihn5mFC3I/jGxwAaHHpV2Oi3IuXb7T
a4z0n75uH78sku+kKoMHutSAmm+/5phuApOhFg7BVnO5XD1N95HhFOgW9xOpTXc5
EKfx0ZhhBnlXc3gPSi3wsxtnO0heVIl1OYYaMvARUTJxM2XjTsOXo/gUy+Y624PD
2QjNXqbySji0rP1jjDoWzmi31p3cf0PPBneydLyD1ABX9cbyYk0YTafK31PYSHqJ
u7XSzfcU2kfsth8dU24YSRgkvDuAsmvfE8ODedK68U+pWkLB7Md2NGWLtjbHyZmA
LR2IPyiUsLB1BKKHd08rjwFFmHHVT2jD8JbwXKuOWNwG9wOfygzpMz+MURAVHNQK
tLVvROKaDfEY9NxaW27qglMfDI33j1hNtrZIFLBunDQPsLgxnTf8xdEmnIvHLUrq
YVzD7AacIET3L0eTqa5/ZkDK6VcpR5V4Ge6pCVw/YVWc490I8ogpq0Q0+lCEVvgU
pQ8usZ/BO3QaNTXIvKxbGvQAk2/zMMeZB9A+Km42UcMrP8ZKnSNc4KTCyFWwJ2KG
FOqTNjFyxbQSa9EXn54KjHW7XJUDxCttWkSv5dlwB90NTYulzY31cQC3n/YU15B0
rRXiQnSbi2qgEDyfU/P3gDqrqv6eTpJFS8wh8v6PW09vHkuDa2sM7+oc7L2dPHeG
B0gQU+t30rTLE4N83E5K/WsmCKya8oaUvpsuE2nlvlPLVQ9igsAdnPm6bIpcQhZN
GO8C6cQtyYVjFS859cth0kA0G8oHX9lasW/odiS6e6LzOEje5XB8JqEpt6Pni2gQ
mEvyAHIGzeByGOh5onvwEyiLcEHHuB8/uztrNzHbEX+G8ryyX5Go7ptQmRF3cVwl
XG4yo5OpoR7Kx34EAFwni5x6vIxeSmL9zuaYEs4RdVrw8eP8tPTNZXUxAsJLEKqQ
PakQmercQd7E/4caUtfxZ+20O5iGN7W3GYW08I3soWEJYalV/+ayP+WKA8j5J5k6
R0p76tgzbpjhzNGhY+ctPAqm9tX/hnGGVnvc4pOn1qeWflQNSmbgV2vhRHQv2J3s
GnHBmx2u7p+WDo1s8/NC/wYEkgYLgqFeHCq4ZXeuzFhsbcdGhyHoK5m2AvR1PPEf
uWjEABrb68yd2ErNyRQmTO9Rz3hTylgIS9DgHwWxRn9x9kM57VxtAWdeiHbOCtej
yw1qpK66C0imKF4mvJ7Y8GdaLpy5biDqdqVCuTPXXaBF527msnjyjk2G2I99dyPP
X4VUhcLJ9TxhC2O8OclVS2LDmtTOtXf3eHqphCRL/zoGj+UaJa12QFQDbDKIo/Nf
tom+5oCo/JdBDbmgDnlTs+jJW4lYB86/MPq6sGcFqBjA5q4dQiE/PIszcCZgwpDe
/FfD1/qo/r8kwM/qhkViHkKgA5YAf/ob5YnvHkKvJ0LnO55BoVVAeoK+8hxv51L1
LMOqlnN/nH+5LTcso4qScDNO5wbIf29e5YKyt9CSo8K0z4x8ooYPbZSO468BKEQa
bUU3S6SqmVu3+OqU0V4E6b7UCAt1UvB24BvOj/iGJibWB4422CxmLt1wImN5HIgZ
Xl5N13KvT77cLWKT8f9A8XOxDD/xCQBSAkg5+ozw0t2QYAVtr+cRAeS0wYje4SoD
xHSSjjJr7X7JR4zW4m1nGTibvRxUP5MF6M/e3X8kyq/h5a0jnWWSn76BdPmoRpbL
qj+veAaQV+1OcTE49WI9ZmqwkNg02VFuIind1PD44rRqLvneQQIzn+HM4fpCjKU/
VDYjMoWQbtn2Se3KBBhn3ebYtqFo47EXS5Gc8AvxtcQo35K2RB8V1sdmL+o8/GLW
N2Jftyhl9JyftLuFnZhLj4cYVrBgVJdbE0eqcojIPUrOAuYq867ykT3U1GXrKp0a
Eyrk8n8V+eqiboaOnlwR+ZVdsjARflLULs+HrgZeBiyuWH3jjpQYFctlGd6VeU3T
C9JRBj2T66g6kZoPbnxHpzEmbyoWt6rFQJ6e/nfTHrLVqxCs6Jw5Oy1cV8+blAMG
Ea7H5IwQzBxSUHQgftKbKDjUeGRp1QV86VSPrUYYT13Nt8/r5IneT7Q8Q7UAVGQx
gHv/67q3+8gqOsdA6W1KOUpI5ve0HaaBPNpP3dSa/TsCJ6dhfMeSukgu8lmk0y7q
QDrClWOdsGi3eHgTeimFeWdZCltW0OTnk9yUMM6oHoXJiXPsL84edMP+qRitBaBJ
hNA5NZ/4XsMl0RvUAWnxBIBTrUBdU5Oab2Rj7TNoScfOgQQEJSF5D5ZWB4k0JNkd
keYBX/9LMGXqitxPJrzXjeo+2I7ohxhQ6vLPWWJc59c9Ka4pB7f0Z8J1a3iluHo1
k13ZrQTbBmhBWpyesg3NwASqXUhb3F1wBzhLf2Cr31Ctkup9zjPXPzPaj7AGOLU0
hA+OI5qNWqCkEHJDV0rlMp5/bz6h1Got9/2mI8D+6T47EFR30YlFTVOthkIqzGKY
Lh5ETL92xTd4J8YiCn0xmoGA7fqdfMNIx4677/JGgr61XKKfdeMja5dWkGPCE+ys
WWp78qKs3pIym5APtiq/gT03FGHtKwY378Kp6ddb6w3gYPH99+0Yu0tjP+nDHyzp
GbFFoR3uE9wqOpNqrX8DO91rk/iVpdGz1rmJvkxfZTLRGH4CF+A6OT2nzMfnan1i
8gSE9R5AoYNktgYDrybpSRgUG+dFPtjbp9U0tu1iaB3af/3znOfowRmeuGc0olp+
0uB4ge7Eq3SgIwuQuhDYixnK1rniPBmgLoChoKGzKgHaIEvfsnvBRnSzeheY/BHm
q6hlpULvGiEl22ebJzVZeG/+qA/LAA2o11/r37VnWDorQU72cKjKVtk2pXV3Lpfb
f7q23nxuMc6YR9oKgjBFO71Rfj31kEojGz8BnsCSQTicbbt9D/xWY5lzkXqm3A8C
VDuAwVn8DmitGY12BcOjD81rXB08SwCLX0Z5x/AT1O4LdHMxMDK/qhHOWiVK8rd7
liHwVzUtFp/EN3/137+n7lFiRv7T0FDsNjLadKlWhzEk+hSR3rFHzqvngMR8xpnh
aB3ko0bNUDLhv/oWPX54F7EewIvx+TOCAk6vdC4IiqOxIbs3YFpX9Ox3l4ZT8fWL
tEHFuxKk3v8UqqYvCbClMTnZsEI0HcawCstlUX47ZsBxFsazLCXoR1jecijgrIca
8KKTmGwx8AUIFcNMqlqTJWzpeLsskFVZZa2PjC8eFgwmvcH7IRkZZrhCjhHSLXw+
kNWNQFKdalkNEDI0gg8olaVTX5ECz/8rc7dWxkCEbYYXJ2uRMFFp8BLRdTcuyCi7
XPFUotAOvdazhAlPwB8RisSulUGfm/3PSJBSro7Xacd1dlHIZLkOsHqw+s8h2hnL
R3DoPM+efQiMeafizsqHRbzgWqfAqwnRPoZzIBZTM1gTNGncBBTTFUOOgL+zH2SB
nat+r4qwDTrm1jhU9MSWcl59skfeqprOig9VEV3IyRz7AlFTnJHOMGlmDOPxdIoa
8savOUnLV5/C5CEv5/XH/Zyoy/ABgHgcPh0IqLzpkLpyVkWCVn820LPd3KubjhBT
xCbonOqxg1vSiV8gXUTEpGjF78d8pGatnu2Z/wdVD6QocNS8BT16Hv9Sal48650Z
F70IStx29goT0bNyID3NqNsVdvlaCSpZstfDsB6lktuGlTNdIWuxsCAApp5HeJNg
Q4mvyG2nKFg4obVGbqDifC3nMaxKrB17/faApbjCjcrNJjvre2oP7fmpQgr3hn8c
NalV6AjU5pzX0vxmMrsNLGpO+jQDVDBanb2XIqggvQCODBOhaIHdkGydp1sNzBLV
0PToWt70F8V92hmLszTTgyMtOziDPjMZ2xULRVI8/w0eeuyOF3YF6hlFDzN/Cgad
1Tty+zKuLYlr2Q6OJfUwC5a4O7+CW5HViU6FI54yUye9hCYczoUv08PIls/qYl3O
HivRIvJJLQTpVnD5SDHaqZZcHFH7c4+SQ+BeRnuLrd+Y0C1jGhENDfZjvZdenNzZ
1XCUOU2LTRnzxBLjwS2HUiNsb9RGm+FbBSpbRCZ79ETEXNPXxEMEiCzNZDDXPodI
zV/ttwB7ub5hGRqYYATN+vF4tyTfusN8pMQ73Yzx5BsBGAujQMNYF4In+VkOAw0a
SE77PgSyHPuWd1a/M/3Oi6XSNT0Ohip2rZzQUVQI9cTdAL4WMq5t3qfpGp4ZPVy9
50hEF44DweoRS4NocXoBlQ==
`protect end_protected