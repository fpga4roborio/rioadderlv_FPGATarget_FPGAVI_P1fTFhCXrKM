`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
ddtXksX2+yylW5zu6QL2Lhnb2d1sD00763mmSITNX595NcHTEkwn0zB1Dry37fOW
FufOhVzEJp80NC5qZ/+F0Vk7Ik02dIR0elf3clrjeJRK85K4e3Hoo4xn7YbFUIms
l/8VZSb14+JVGURjfswrIyCUotIzlzVYZ6gzoZwDXIi5gQIBf/gI+KxNXPaKV+PQ
Ufys/12rjO6aI/pPlqSm0hCvftmBcnezN2hk1UeXgOIuKZnogjOsf0iJVX2aOOWE
6pD/psybjbnsNB6kH5uFTA5frkzIzkzl5d9+YDm9OyC+k84E83I/7/j+rk4L2dah
QJOvksSIzN867/4Qt8qYTQ==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="MvBXkzurAa5VTw+1JJ70nePUfoQXBvZOku/SMmg4TwQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
oRtzZL4VJ4iwysPsC8SXYCzXS8Fw2gtZTOskLcDV+1B9Nzn1zTyNtlo6lNICRmmK
ZRVu2BmCc2G+fmzynYlNTnSa7C0Cuel6FYpxCBlOuk3OF2tzAmLAuDyOH3Z1Yjzk
a0aHuoCdIRKv7BrZCdALt03JeUmXKPdOmIlkVGFl8yw=
`protect rights_digest_method = "sha256"
`protect end_toolblock="Jn9CQpRhJt4rnzZPRk+dOpzAubz7omckX1MrFd4p81o="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 35984 )
`protect data_block
gD6l00tciPUa6pDNTk/+t1gcgy1iCdpjTkA/bOvU9JA+cpFEv5u/7dp25hHk7lLT
6tYtR8HgwcLXTcx68BnPlzdPHkVIv0lwXo6yhFVkYlDWBcqD9ubowgKij0UjlXmV
p4anbpVt/gKvAYRDYe8Q5F2CQ8AIsxOuOcJ2vhCPchS4QF3n7+oG0MKU5ZyzxTu6
XCtaTx4goSIs7c8jbVtrPTEum/nVIOZ/FHiODYzHs8/XxC4TKl4baAfD/5hIEBxJ
W+Gzu9msjc1W0cH/P21CV98ROmrtq2B6+KDvLW4YkW9qFn4dlWsTINucCRnwJmp3
nRaYAKAcdrRP0pxyfGHDD3qucfOTT+ixbRANc8pYaqbJwX8nf8k/Nj2GVAk+RsxU
xJuBmh4i8YFGnHZcl4QXTL3JQ/3qnc4SgItQN4eS9KMIw76pezD/4uIk8gUsV8sm
0eu62Zuix0oLjGLNY3aibvQ5dElJsMhKQqdnQQTzUs4dPHy1QeZ7rzPPtsYjquYB
j59d+NSJ8GeY8bRq6I7kvUadCE1lln1U+SH/+mX34m6aumnYOLW0TtjRTPQNWigT
m1VUWegAFbkfWHEtxY4Yn/MMrzGiRUnvxTnj7nG/PWTwv2JtUWiOL3lwTTbI+lGb
jKIa/Hjum40oWQfpHFW/ur5+S369HoxkScMmbGyg8QefEoFuJDYxax90jwPJhHS3
2wH8lELw/aA4qZ0QJHhlNdxxiUW3ArwVZc0mi3Y44e5/h0zgVh3nyHrPLR0PNEVU
olLPHgQUibgcPSJOapbOMZcwJblAQsb0A2+Tp5tYP3Ojmo+UXugA0AFEozgm6Htk
z5woFfgo5toAtMirmVdI9TQFRF5y8fKn6NbULHuWGYuyKN3zH7wJsptjd0s8V+HU
Rh2obgHfIoiNtTeLeiAh+9AQVEjQcBxN2dWBVKyvcVulMFv+w4RttkQcGz6PRi1F
vll6ue5Gj0Z0+6qoiSWyubqVjnskwMAujbI2nqx4K8DQY9Id/IPpzNE4JdmAxltd
8844VvW5dfsKfeUfqpx9W12igUFLf7DhuqXUBsm79KsEVKxm1ZDyObBCgnP5v/gH
q7zUU7jyMwMLMYXcd81XHBQ+jo5IJQXLVyI0c3ZDOSJPFx5YNLnqUd6ohJNOJhDH
34IVNmGEbZxFNxz8nV6HAJ84P91ti55tIOuhI1biRoey788eNB5c8xYfTk1eMIsk
9AkCiKvSVIC0v3izDV6x+zVBVIZi3HOYb6g44DDqtC/doaYgnZCF+p6Qm8pPzd4o
QF9IRpLhhXRWpCwdmHWnO/LWPB1iWa3QoegDLiWDqVn0Gvm5PjsTINtt6EPrkuw/
oV6zA4qNr80yLaYxWWOb8IXTu1pugP9pgsZ4RIIWY/17o1EwvXFjpO1uIAGfRPos
Z1Q2n9LghoISQ/gOUquNYJXEIW31aQGfAOFvoAb5aRJx7kaOWdM78GITmCPlFrHG
/37DYJJktqPqZJmwH7fGeviFV1zGPkqs2vuVBlToNJbfA9cfcDS6uj5hLKGlkpL+
gzetDYS0i3F5kJleIA9M85c2dD+cGnxGr8qqGC7H9vw14CoDsNk1AF8GQiPi9z9b
cy2bCyaedHour31VC/iVOUHYAwdTfK9E5KBlZ5wlES3PIVeGYj+mloHY6idpXtwT
xx2Z5nstiXPyS1eSNdYINNqdRgCHJFiW1hFPy9p3DuE0ZODup3WF32XZjxdWkOxK
pLV898/Zg7R9iHDF/q73ooZhECVN0KAjZbKseTmGsNy6vhAyrmpefWeV3pv99V3n
dxV7Q3Dh9vXBix427UkECAR6qObbaB2gpD87S7Q303cDiUsebG8xwKVXgb0TkS6X
IHZw6Fwk/xkpkKBSRYhsPz3fKbvn+B2dPCDOByhmBSosa7rJJHyv8qWQfX9mu1vo
AM24+u8XPuUvm3FuTOspo345it0ZBwfSO7hyXCkwgZwyvFPqLJE+mKdb/9ND3LmD
gROzfDMRKv7fB2wF5wG2VdQPIQ/uker9J/PO6Uy/7mOlevuFtPdgZ+seln+D/UbK
ofjMzn7hngn9T29Eqgp1oU4tPiYIQfjPwQoyOgVDYMiKNgvOJCgnRmvISqqKq8MS
IdTYlTtpwKeFtvEyTWcyF2NqFKhNVyI47RjoE5K2bgAoDOGtD3FzMHD6JmJ3DfxF
y8O5Pttfl9KYIeprVKfMv8UX2ryX8mR04yiyAMTf7QqCNB+6RKGRYnOEm6Kpi+H9
jQzrNb6IGH36cf6jb/wbfeJ/wG9gUTd4Z1JzJPK5gCnsJCo+sXHFajRA2FEyX1SY
QbhVTvwxLaixnyfBSw9mqgGfp/kjcs/7z9YpmuphV90Xs/gnmp7iW5Y4KJHGHvqu
1XuEF1xrOAcCWXXt0jPer2rYds1ehb2j+ziiCK4cLr1l6f2KJEIzssGg/6LzbtQa
66122jtoRrUzLhU7f23eMCPk8DFz6WJ5bD1RmRHKLWpl/alSwaC0yvWUggQACwzw
RGW0A6Zvk2fyo9QKYKtDJtRIvdihsos+xv2vITq4YzWAJ8S8rh7KrKApVJ704XbE
rtUK+wQyduzyBHWv9eShsam0PWy70hvJi5XwSERTr4cCB29NAqBOSuryVQTsErMG
QxFKan25l5Ps6YhQV76PV724qXfMSvnvu5FFHg6Z4qSXer1Ho1VIRnoJe4+BDCUI
Nq7t8Nc99uQDBtRzgKVZEg+M7xGn+ZzcD1d48GhXsM/uABeGrk2gciTZxzs7PZjR
GvUnenakCeqtk9LyG2oBHA2Fc6ZU14Xvp7uFu6MY2d6TrX3Iev/09PwfXM6J0HQs
OpViBX24pCKXQRqopQHYw4FlsktJFsHuhXyOL/b2RpHoZcgJfG1OKA9c6F2XUt7h
tHzaGoa83sAHd9OYS8UpmxpKQ8aet+kPG0P61AzdJnUoCvYBK+F7LOqv6VsDjUw6
2OBtq7PfX6AvYdgvU1A78JIw68nNuvAxqWH/Yp/3mCtR1+qGlNjq3fx7ZVp5wt0U
tnkPsVlTh+MgFRdIv9Kl5rxrsqzpnOIUWnOTKp0roGY00Gl7JFC3nkXzolM2QyOm
7ybn31GGRdUG8zq72obg3gBFz6yORZuQtGLhb0ODrLtUavf1Yt+9r41khy/MihD7
HAYaByUVS5C3XUGRilr+hid5we0wPsTWtIC28ap9bpqKM9CHC1rbNQpNMNa1C7uH
WoiTbQlZ+02BnsI9lmE0Fp3zwOd0IQSv35mpagwN+nt/6y2h0yVMrfLKXlcBEi1V
N4RgNlTYni9R8LI9ltfYhsKP6uM11iMxAEPYl18kj/+sKha7I0xhWrXckVQL3nCa
0KyPU2paU3CpHf1mYyb6An17Jh9SO/AMfQnY+TyVVKFCowtm2txtuG+0gM+HBjuA
UGXINFIlS9GMdRq42cAZm6AYJKUKrQ78jBjPGAn4CQiQlspxS5M8hdfOSmLywK7i
iKasRaGJA58Jl6id7LmL6TmmqVk2Gtcx8yiza+xkImC1RLla+szXd7jgoPt8xNMy
E+RY8ARjcBnCBBYXKNvIbTXo5aHfm1xpD23AmN+VIEydi6cnRpTBckZqxq6Br1LS
fru282VenIXQpsKL8YII49M9dTvawh72OLK5f1WmR1yxcRSBVLIVTcOjomE0zyGM
xcIIHTqWy7cAZ5aF1p/igGs4UtMBNKjvuc/Pk0aegSdJGS5tXDOiXGCKSg5sY+37
dLQ/3V/HSkP03I/AOeSWwsr8t7LVJnQNKPKLQnxgZ5ETZXF285ajjzliTRuK9Gqz
9l+PW2CKKd7uFml8HsyeukiJOBKo2dUMzOD6eEnRhCmxCa/LkmGRP2uD9dgXvQCq
lPNT5ROW1LXiD7uoHn7+bsWCQWr/cwOL7RWstz2SxCA6J9K3XK7LbWmGw34CdBVR
uA1YgWIMf5XNkUNXZ03SP+xUTgx7HW6RZIoutqZ4TxKvJLqHXdtDDPdBhQE9DcJH
pIMKw7jkHWLwElnDo95X5uUbCNQqXkxcO8mOgBkF7j2JxRdPAY4h4jmzLiOZycgO
dSBhJtmHPXZFMNF/oihleAaASBqpPYdM8PnY7ji0okI7T82iLBOhCvxBw6KEsrK6
bs7ddPY19GTaLIKWBeQMMcvNBtuGAu7LPpCbDvlnikoI/NMbHomB02DWdVBBQjU2
tInpntiA9eNntSdtkcpZ/+T6uH8bPD560G4fOUMnEWlNBFQhgXexjJs6h9tOpuxp
/+uWXqBdNOkg0tkDBK1K0TE+AWH9xn0sD3XZu9PnKbTfJamESlL2IcCA553pGiIP
GaWGWjLSD5ntdEs6j9ksVUXh61BfPOgHJzLpe6kv/LIiQ2KzniFoFTisiZvfc7z0
JvNF5gAY8ORfRhJGJkCdrO05SXEHCLQvJaINh9RKanylXMmlrR7BnKeEFK6FWAh5
+meer5lfTzUaXGyVaCiePFb3wsSVxj7Dj7e/LDTO7cR5YOwAWV7MKEv1/sLIdUBE
lKnQNh15GkrRXqTuhxyB8qgMfE1IK86IeknDGbPJw55WYXe1ieJLH2U/zCyxOa2T
ccIhj+5+t4PEHGCzsff79pFLuUIF/3zza9fGTNkvnjIvKCbXm4h1LrVvRiZ7qWof
kpBRe4ww5GQNa2/lsZ7aBUl+m804sHXfM93uCPX8k6cbVEZs/7SEyrK/h4/Eqm5v
pgzfmD9gDLAh6qrO+n/NyCItk8kacMoqoS68uuNRUhITZGenoWb8dofRPBe6ZU+F
2G06Q7d6vUi+Q7NxHKljgFN1yOL8WCREm6DhEMWkzx6o5byW5e/8S7j8HdG+m8Go
vWZIjeNBl8UY61Lmb26TTWsPWlXzNJjqIZSPC42+uL2Z3+1Fazda7nUnE3vcd68s
+V2yLWUK7qFanRgpTQ/Pf090cMRBmIw6igdxwwQtFCIRnI9+JFfsKK6E2bRQdHIc
jW3ZRWq5cIbAVIz2g9RV0Rl/7uSSwusXWg6VJRtn4lcWO0duK6Uilx5CV6xOeUAt
wm+y8vCzV7jBLYITKGDKNubjYxF4BQEO3NGDhct8PXQDMAJA6muF1nBqbs7OR1/+
qUkKkmQX8SmUvUTkmPR4k2Jew5sIdN62c0snoSr/ejcXZjnLomOMgqjQNaDISPUZ
k58GtvneYz5p6dyIrqv30QyjOwrV46AKySXkIJzWsEzekaCMkW+yfSnD/BD7bZLx
EJ8p50frsEB/5iw0l6hiFmGNHzsxQUOpLs+kvanu3TE+KorFcA6ktVe6SGf59uPb
enxPFlfsoCVWsIe53hGYv2MDidZnEjub6m4ZYetl7mtKYVoT1ASXWjkLt8NcOTNm
OYeSqCMB8l9HwegQTKTA751fZD15MFsX/zSxB462ch9mwZ/LilqXEb8TqTORSDS9
m/Aq5dykIGEIJ70SwMmXR9d3nFWvAdyqoRoMKG7EO2hB/oRS1LESDZYb+XNFkqUs
EqWhrXOjTLTDYBUeJ2qRSu9toX0tLRu7vrLHVwTEu03g8Wuaxr0iKu3Ni2fjmdTc
Pfju4DS4DJI/duWYOHZ5szxygOX7G32u0J7g5S1kUcICK2oDjQFRzXCgBkdnfLpW
Rhs0sAyqIoQoKDWLfVrv0NrZTTUQ9e0uxGzciLpf7ca4ZUxRVa/2g5l6GauqhubY
Dir4QG5e+314/1gcvDorCVHQuI6LiE6DSneIzqInzNgCKNvv9I/tMKwoVsiGEX2P
/wc96Az/3ycxLEvBIATouTeF4y+SpvEJBl2XokG4wTCy6olvC2niAOSAtBidrjs+
zENn625R6QzxL6sK0zBKypC4Ayo28KVikSg9Ik3llzJ105/duPFo37Rnv/6VRQcU
CnYv8p1rxFzpq2wdkzcHsIKp284b5rDcTscGwOhOLPbDqyxyJ4fCoW77otD5+wTf
sESdkgUYr5cNAmQa8ANX3VlaD9PIUvuGDKTRHX4JSuCpr1xiRAXFYUZZ25Y2F841
5DAwWQRsUg2/Ni3gf3lsQ2jVGfsI0ME58+GlGi2yAUlJaKcfl9B4jLAszroADMZw
YFPoYs9u4v3T4yo7Ml2QR0xJHCUXk/YRHg2QYWZoDjKQZEPG3hLgTaT0BkPB3EL5
3I8+ov9IZ+Yb70+UnFqLLSc90e7zrWEncS6iDxnTHeOXrmiCWKiqegDyHZUt8+CK
Wb7bxXgh/a5bLAlYsvYK6qZ45dGjhGBb+c/xoyPRsNGJ93Xj+W6FankSex4M/E9v
bWLu+rZiKRMd2mdF4AhrX+AP9NCDpbXvYa3JR0MoTdJNlgHdnXcx52lC6Vxtjrtp
o7a4NcB9mwnItnOvE5huvTcRHy0SMvxBREXMEEUbYMXKPnku8Q6TGqem/RpwC4G6
BZ2G8E3JnLgVED+TMgqocoXEqG7zy28oz+fRrtUhmh+2YI1oVZE24RJxLvR2LN6k
ajQkv5oN/yAbEI6Pris9AXl3e7s+nO56IwY9VicdJiBhY6sWbK0P2WMtyCi/tWiX
y6XLH88gUKcXtzQp6mbKfwQVolhLeJAsmc3TSG+ZNf5MswKNFgy2PeKxCc9/IO/d
FNTWgloYslhOKxFwAPBAtD1Y/2HXWZs6pbLlUBacG1+qFzW6PMZG/cfZjwGqieIl
1rUbF0B7LP6xUvKY59BLnEWxZnkPO4eyIrq5PveK+98ZXOv6RTdDQqGJRKR8DhXo
vruugp1MaXe82z5sM5mVVmM3oLdSeK32wyD+kWwnFRv/1+I75qegT/Q9f1bJo93u
4qB/S3xuSD9m+8shpMDs9Ex6RvkDC3QA3I8yWVxcQvDjwjHlxQ7bCK0CYDhl0/7i
kaq20zGywhBNpwmUyMEd7ascPWsXS01LF8tAeo2HktOHlpuX8RfjaJC5Irr+Gi6q
Jt75UVKdZF3iCNnUCZyii7f9LhDVE6pyjnYyb/Mp5kKqZtxzcBCQHmTpKYCE9YpQ
vhVZj32iwE6XXnO5YmChYEgqQdTWtouul10GVcRhuQB6+6Pg4SYecj+KniOTciJT
IdPPhS8kKL/d1tWD7qg0vjXcGsqE9c2Qrt46bTs6jpllejBoV9blXuA55Kute18N
i1iZtN8p0VQB2XaJPBNCkKzLEkLl50A7UL/E/k5pPRsqKKGngIQ0T5hlgcDl9fiU
DmqNcoif1P2XOMPg/tW+rc7tyt+foigzu/sWkTVqujHijeBjX9S+yCH8ozk3b2tH
hbSZIY7h988/59Jb2J5OkLMZ3x46acXDu5I9GutTSUxeqlUel8YDmeGvmbX7SpHn
L2qloMVfI1DDeWcW30ls36feTitq/EGTMN+QF+fFOOwkbpvjSzpxTbYrU0dZj+Gv
SMIRfQ/KZVXd82CxmWI9tL0DTPEijKP+fUs6pbSv4eo3bHlSsvL8HB+mrZr1SKtH
Ks3XkrkFLBsBphIMfTZ3SSEXGk31/UKad4yg/X0a/yuP3Uz76McKJiDGrVnYaCcP
hOv1nu65YHVl267/ktlcMNaFICUzthOf12/Ig2LfjxjEGL3UCmCHBIaMH+JHzotO
gXZWIRLy1TpffDJiZODA8G3Ladz3mai3wQSAuTRHRlYcY9N409UbFJC3MdS8Cs/F
MJl5bdrHFMc+J+JVCxvVHktcK9x07xzX1M0liWiqxQD1p+I2skphg4p+Y/TQqM37
aFH3X4OanuhRFBaESgdDJH/9gna08KUnE9Elk70qru5UC4U5k2JD/vYbq6p1yHt6
tm3VL4NP8pC7JY33/mGAs0HkGeRqzR8q2S6PT3EvcelE/sUR/jA/XMRgzk0knbh9
YK8mVUS56ZK7ib8s+CihZp+BVuPh0ygnKa3nAr3nbA0OZpMcKtPPamGzhT1D0kYR
qbAsTMsTrqFlK3i1LzXO3JCoaV/ecbMfuoaQ0Ymh6ZuecLLCweXuF4qcM9oMtYlc
d6uMeYMCzjru87yntLsTnYEE0dRwPGOcufM6XbbslaiD8Vh8f6KG2/Zipl6XMwjn
RaTajVZxWFEcQDkEnLWjJxAWEtlluhwS4VqxuCZac9haLSeY68ltp0rhrnnUL1or
heVHn6j62esHFnbK2oZzA5Y7PD4XJbgXIbIxWj9JS+1/xJVoUuxrYzkIWzMlIOmt
HKPF1VP2MtlbIygvIaNRb9U3O5Q1ty05E/Ijw5S//WAmlRvywn5W9w5uFo6WUjwu
fg1Kj2SckfK11G4iWBrDEsLjV7HCX1geU2YByIlSwAH552uyiBHyO7geYHO71NfY
sRU/d+ZofhZjukJacnoU1wqMZIpFqiRA7YNCReJfrGgne1BNYuV/tRs2EXcpS5Nd
7hnDzMFhl8CxMjJIxiWdD0Jgc9kNaCz6HPwHfDCmtPOneBSnSySGguUFuVeihU2a
gwGChotf8J6F9INogdxXX1Nc41A99y7kNadf9jeMoQaA1kdOOC7X5Cz8nsHZed46
GsMUddUHXY1h6JrS9VQh3P+tz/Z54RtLFVywtObzhdsYRhtIgFec6WF4wnyvLnd5
J8LgF3f2wHB245uKEadHgfcy6wLOEYCDZAFkudem2W41uimb/UIPam5ZJWRhTQbq
Rb1dtyisfCIm020msOUGoIuAjOh+S2fYqo4BGimIVM+2x7wJ2TvIeAyijvK89rvG
pyV8DtglSlfnSmewXwsTZFPUBaMs86j46cz1ZshSoEv3ofdvCC5JXMUvMpEJyau+
2UaxV09FEbiqhbwRE8rc1V0oypwNbAEjGM3FTfQf4v0e3cjZ37PR5dVN+h7VsVkU
E8U16caiy3Y3kWbmPqnMggXeKtvqb+UxpNVfrbFaTcNb7DXljJr4ZqB22jMELBtm
y2NzC5IFs4opFlsQPhkJnw9n0o3sofmFWOfnGL18Guqq/RDYBw9V2vqGl1PgqEKy
w9QMC9FsgXKApmXCI6B9jeASoL5ofOAAhXDlsLerIyzxImwcWODC0qp+ldYEXo2k
HCY8Fp5IFcPlg4S9H+WFs1gFb8RJAiilb3wONTiz6Q0Ho15R8yYKjIp6//PNgVfv
BX8ScUetk/Uum3Ce5umx+Re+XUYUboxqoN9kXncAz5DZp6liZfX4QhoF5GNDeYZ+
2zwL5cWWGTG84/jp3IuXkFf5fK/5jE7P2u2dxFArefR0U7HLnM+MDIVpuF7i9SFL
7L7YEJKZZlcaUl5WCT+RKd/0B5s9scVotz/KmySj1b5IWbyKTljRs0JKjTRI5aaI
6ugse8JO8QFi3cPcKZx/8g+4k/HiUrKem5cKXB7TyGvAaahenVd7Y0grD6zJYVza
G/CZbSC9cQhxqSnNM5Uygg34HRMyiHaE4keVG5c7tcckUIIEpdxUWHMU2dCEixWk
+lTSHKHSEjQE5+Nb9fimG84ioyYPnllhiB6kmkhrADdI9gAbVjjUKG/LBUdwiw1s
XoZ137u9n3Woici/dwf2ej4d5W8UIp6/bqQxfBQyhzadVdk7GISYk2YptSAosPFt
1tMyW2uaiu43D9FsLODuTfGxWE6jXM0lPWde6oWraSlWWqQpBkVcbPOvax174J/6
2CUd6CmIKvRrXIlKJtTGMIkc/DnOUC48Ttd8LFWDgsPe4xujSMQwl5tIDIt8ewMV
9uJX2KDC5/8l1ez9UVTnkMjI7oYm0KexhHi+L1oH+o5DEebisctlhVcWIRHmaa2l
oPr8oYMqWXsyHARQBuqCahgANO+vJnrhMO6VyitgEsbFjFgeMhVOMeqyoCKHsr3S
n/yuPlDGQUBmIoZdbOy9XnCUE/dEwh1zQMVQAqx7XhVT4T2YQbLcShUBc71XPAw4
Fy40GwB0/9q1LfrWyFND5tHySn7xeehIlz43aRtW2fXpJBsPLcWGZ6LmASuDOjLd
HtKsKNbBzhvoEggwAGd4yGuw0xTqrT+9vXWQn4aEf+pNOitR0r+gouaAV5Jkh5S2
vEublnESMtTL2PPlrPn+7+9s6GqV7v5+nckJy8Rq0yzAQZANVwSwKLsWSXkPmPRD
Un/88Jt02YHqgm2UvD8fuRKQsZkj9MXBHZJsYCXMpUV1URaJvFW7eE4jxFD6vPX8
itYOpJr1iMrg6zKwJCKTjHc99p58fpicwR5SdB70jSR4n9DdqTmFQn2qTa39Yj3s
FNpcOWDNmiXBSzY1Wp8occa7q+fcb8YNc471ac+c3EVqffC6Zw6GgUIoiBtkI5mn
vTMUVZ4HjNtkIx7i5tsuYCV2r+t65vMmRWiLZxpsOCS6JodP8Qt5T0xiFXIkbZDE
Twlw3t3GMQnFIQGjmKctAYzFt7WN5SD0FssoJIYAMG76QoeQu/RDgCGqMx1ZNv8H
ATNHqalBxczRyqWwoLE2f+clq18TgjODLZ5vzIUmFIpYu2R2hba0Q3OH30oxZvpH
QwV9+7L1gTdfb+ALe26tKzAP01Mzsl4NpMvDo/g2ZiY3/q3vQBa7F7o8cLmUJMqV
twAmx1idl20DGdEm6RJ3dVIXEHaOowRJ44awjB84wTTuJnEfObZTSLUhdRlB0YfW
Hqsk5TPg257fmqIPlyDw+HTdMGx1f0xHG3yi2Zveh/UJuKogbIg8/kV0ucwkhvEj
5CYRMJ16jDiwOPbsE615kNUqA/GKAQeoCegOtWwRayjQckhixZjPEr08RopSLljO
aGYt2Hn+mHZMqGZJ2AbOCtz/cbDS53aWRU6AP+9/6M8zcjFolgtRVpSldca2XDzp
Z/DXiELYY0B/WKuxxVP7f8/B4HjIiNQfWC75ZhwB8siPBC8qytFsS/mfTdMFlprL
ps7HkSqRTnNfz4wTXJsiXNLNaflwSYqvDSx58jOio0a6iZGQ5+1LUQ3OJTzFzn5e
JdH4jygH/XPqJrJy0xsbGNoM8m3SpfvjBLlTNSjKnhCnHwPArpcx3DDyuKVoeYEn
dB7coOaOq5AGAdLLFmiw1ovybHHyX84ts90MFiDl6EtXe4ESP2+QsWFJTG3rMt+c
CTjRejDzm5OaKByf7H5NsYVXZTSdGTHeVn+2rALTj89RaoC6jObzqbX5ZSFpyYSB
2S9dWu7bQdOZm78IWZ6dIvRn37sg1wwe/QR7Mw/9oq+7Ud901PADszuuXeOS9nuI
8OR5o1CSg0jCiSAZQhurxDwoPcNLKT6nZ8qV/dUESpC9l2GrxQ/4DLk1PhVIVwTd
hZqV+OM2XI870q/eFE8gx/P3njJQVO/cPefcVhd92gqMbtlo2F9RlaQL5KfiB+ot
YOPLoyXQHUicFwLh6erRffaxIGwKuF6rydzLf5Pqp92qx6gBWhlRg4NAHotV+Day
mQe/IkHLKtyI+SG8qebdBFzxSzD0geV30AY7YSQkECEAPP77wdg/xTpz4vRHbD3b
6uhfhJfFUwasfW0RBnJyMh8U/DkNgxOr/PvvLbz6RTHyukrnA8FRUuc7r7l6aRgW
m1Vx6GZYDkJ6RpT8OiTpTasoY+cLYwygxPGeA9YHCdlYRnXC1g9KHl6fd0M3PJ4F
cS6kFAgK928rQDhtJQStfdyFAbb3iH14tL4ZqKCTg1IentREwFZas4rQxJuOLxHJ
APVTqgqZlmOfUiCsOXOlNBBEAnFou7ftJKpfQxjip9n0QGuLb5yjgyfJqUl/A+oc
XqYjtKWyvVg8qhb5mBDgG1sghVZ8v4XUdPnbgo8fzt3IvlrKWjfGqoX051llN1/Z
ULIV+Czgyu8m515WJs1aRNpKnkmJhx2cwjL8D5vgj7MxhaKQMmg+8YlsCA5qVBrx
vtSc34UyOtRDjdhIi+/tsjwSEbFj5OgWKjCbi+17GPbfVfV6RQRlMQ/AuuM9u7Qi
cPDyynS4edB8GlNkW4VZYSpCS3oFDZ1/WkwslsICz5ij/VcSKq3uvimWqD2oNBMU
tZAoEmenAl7G/KXOVcn/2lFzeqOCEXAEKr+IpdtyPPUrvK0oNU+sZnlQVCfcZ1JH
s0vbqfamPu4/RKuj9V7Huz/o5Ei+qK1PEppRHnnjvMjbS7WoXd3RyFaAAmT2MbP4
S81kCwM66tLHwBqjWtgg0Hz44lTef6z0CEwnGoKWOfmMn7lZZxDxHHuuQv8t1FF/
ydm2rbtzrH+hBP4Lt2HdO0vf53jmbe9uydNsEBLpuhR5D0hnbqCGHsoVafFA5k0S
ZnT9K9zoriydiD8SuuycCgxlbus3lbYFgJ2q+TzHw3HHMj24nmFhhrG9nz7KK777
t3ThN81hnNrRrdVz4nSVx1WNQAKIh2eXb1yFJISO8IfLZ1mniBkiJqC2HFysoCJf
5vTjUvCObf8tI6mzcceniNCriCrkfKc0GyUSTlKPBbxQt/DHFIGdHiqtwh8sDbDk
bHMBCJSYp9O7bJcwVhMuL2KRTP5ma9f87tdaGbyeQFCxHs1YrQHZDDJDeVJbar+3
iAlu9kWEqJGWzmPBJ8iGfHCtNReTKn3GXQWn4aBfntNSU2VX2mwldqkio8UgiL1H
eLOVMzOP+dPdXpujy8BrEV6hhXYMMFmC3+4feq9hGVAr9C/OdrZjAovJGCE40x+w
0khD4u+pZKObe9j6+n4Tv1APx7NK/O0XD+8LFK4dZtz2tR57FFucE0tJNNznvmn4
Bagp2hYWgHTAq6r2wA/XMrFN+jHwWUrKWvor8untG2TzPZjHyZhDepqhNHGSe9C3
eU0x1sxwKq58z1hUZs2FV15Gb4isu8puntMIjSGJpwlFDRxX3pgOzsnPbhG9ST3r
IP/sRvjq34NGqfAnK//SFqcndtJ6ioRtfYtWT2CzAwkUttY0/iK4AGOArzzQkHfk
qlgQMZabkAvBinI62c77m0vPpKaFsLsJmqkB8fiLaQkxR+Q/mR4EjidCUA6CKp9Y
jGImeOnAOykmh+DW4cdCg8D1c6/lmVFJAPTXfVZ27rEWU6n0kQTF0IYPncK/PaYr
g/5PsIpjUXIuul6r1dcewQ766849cG6xbxBt8TimrWfCEXU5IwrG2WqHXhlxtnCh
1sgJ+WYVg84xnyD1RaLI+DtFITbKkpvGxNk793Mvk25fsE0Ye+d7r1ScNHvcgIJu
00mrYFqccyYW/eH90xXUz3k3CVJD0J0j75TeCbCx9eeSzLmg0qXWHbU0Z6qcbG4t
uTH/T1jKOG1qIiEoH4GGizfJuOSbMMifR6ab/dRfhxnG41W1B4yCFkYJ2XxzkNaE
wxm3vbaIoRtg6DKqa4mW7lHQ8HdpK6S97ujIUWwn6zv9orfnzgCVf+d/1IarcBlX
KkN8e8tHGrXo8XBRFCgs631DLakT1Wp3q9xDb94cEEwwhKHUU3Qlzc4hrxW/LpOC
CdxNQOGBW2OyoaSewE7FL65YHl4w0YMxmPrEf/0Cu/4rnf1Fu+DP5dVQ4Qz+brsJ
IcyE2Nj1JtKkLcd0F4Ztbbk/Eb2ZG+MV4uvZn83+93ka+b4n70aZpDfYRIhHjYRA
GIoJ8eXxniHxEhao4N7rGcraLA8a0X8TFsoaTgQqzzH9MdajD8/mEh2Y7DzSqop9
n7ugXkebCe5Bhl7IfK2ro+YEvZT/X41wZ7eZJ7Eo0GNY1yN7KeGwrLSw1zGx8Imb
WS+/1Pu0lu7vdxVGVavJfgr/ykQqzBG0SSfc02ntOm5K030SaUTRfHmCxMc6i1C3
hXLPEZ3yaMUOhU2YekXUa2CoZ5Rhd2W/ZQSnslGpI/ku1p3pYW9Zgsh9GzKfvfun
KS6Q5RrqwckbBVxh0vP1sCK/s8JWlcopuWyGxXMiJOgcdijLQTKgyQIjXef5Ysbp
19dXr98lHU0pPqzutqkHsQbO7Cr+ubXx1XUdufvwcXWKY4mixs4zE2x7mObv7k+e
9zzO5ik2XqlTZEiFqpp0O3WyABOKDZsh9mfZd//DgDLrfwaW/+Ts+yYuIDRhtCPR
VzNjIgUl1IcNO7z9l2s8quOH6NDmabJ3DYXClIWBz1rpeY65ThaX+45KFSO6hZr1
Stfdmg6LL40RM0qQXNPtDkWoe6wFgDPTa7qXZZDHJyXQqHuEX4EuURWVDFXkWbsB
eK4aV3iGdYtbomwPycg2Cidip0p+1SY0YgXQFnMcKhJ6aTdEbEzwn3jR/niPgo4M
alhJfWyLDOS4Yx8Gqewf/febNo00+jYemFRW81QRS1llAvtvbkrrYZ4QOQivGhmZ
eITMkUltfCG5vNjmKzTes6CtrdUPQ2iVrhaa4+307M3zqgEBIAivkxz/z8qhAFhP
pkElBY5TZo+EqcAV0wuTlyrri1mBZHUHTEwrSl9/5YydLHNhOoT/EMjSu2Y00aqp
Tir2hcWcrAV3q1puAK+c+dyydq6SJWqPvGq/TscV4tlp3aVim2H6LWB2LOVtKP6k
w5GvNlvdjmu2xrcKobK/9V+dHbKiuXkUQ27Hf6z9ldNgxjgvJUE/yGdCXXmWPnYi
l3cu5q7Oq3+0vNIzhgv7sSi6nNXUv9qKvh/5fNtBKYvmP3c0BTNALiFtpCvW3c5K
xITRMyQ0Pimfs9AgQvEYTo1QLCotyCyaIBKy2++MiM4Ju93CLwnwc3YX+D4NlGeg
TCfDDliJCBmZqS9kTPmIwtnINQov6ZIKHX7gW/EjIaxBe/rLdk+eWRo27VsP/EKM
rT1phXYB7ihkZREm6SH/NR+ykdInSRgJQWXsAX9zF9TmJXTmXG9BrGfmiDxpuho6
m322drLfUkQon57t1d0GWueKmEe928C+gJ8lcBaQTIc548H/kCh52ZlHDgyStlnC
F7NB2lsC664Bjrugp5VxkL0qg2Po+7HSadC3REPjvvvWoNtnkbB2GAycSts8ma2n
tw5y43lnbazq/VWJxDznK441/hW3M/OdZYht7mrqEvKD4FfhDpE9KhY3XT+HquGp
9T7ODvFa8CBjmEwQ2g9ZHSvWTmT3LsOVlWtnOM5biS/3sOAENEJ8EKi5pl93YFXP
o9aJHhPEIe0VwckQMv3Po5s2VcxIjeJy4fd7kWLlfev0UigSEPHLNa1bTgcKzYPg
C2TeGD88lZHajtcxlIlvSSFl5UcIjNOtNESPHsBbjx2m4sJct5vXfpZ+ki64z6sc
2KL13zFxHSMitm2ywnCTDGc0kQbCLHohZm6CssMvpfFx5qsJ897WG8MFdofIhT0x
r8WkTChinmjP8J0NuuP/CSWzsIA+Hzipr3lp5W2y10Bg4nuJBgn9b4wyS+dzIRwA
x0Lqtsyv7RJKQyJOlqFjatmlNKZX7WPjS1UQrp5thxF9PNQiOww5uxHqA9g35D/E
R4j8QD8cIxY7LvHXucotnEHK1L55FnABaOOI6bMp+Gewy8d8viVJ14xMMLehUrxq
KeL8eBPh0KaAlyenrn/Tad2MSCeIIOTrx2MBcYsXFA689cBqNf2ROHeCqwEvItrO
B0E/NmfbYowM91SAvxpV/C9NQSpu3Int7vodD3Jje0ESOCFhUuxlJHeKCIHtUCym
B3K5HuXfOSgsfQR6KEtfIYv8PQX1mbMKp0DEHrDr4ip0uRTs39gdKF9YSLy/coHV
XIV00Qad+tvleFdN3qC3H6OYo8qoyIrXzahZlbkY/J0DP+0ZhCSN/4uWDHA+6ZoL
gjAxMypM6JeP0O/N6EaViwY3sAeuacaJdsYxnknHlI5C3jipKwjWUlp1yn6rBpfO
M7CGEnogvwN/mg46wOCl87ce0yabqd9sT9GEQJVrNcXc+b9ZT7s3GkVGGZSkdATT
Goz5uldheG+yTNKKWh1IzQD2XxoL3lXlaGC6EaNHec2syQm9+aqwFSI/uui3Zofp
xX4qjo7COs/Bds3iWRa7uvr+miWiER81ffOnQqgyW0PTs3i5a/n4meJkB8pMx9a1
3uYYxet+i7ok2dQBPhZvemhDXYmLQT1nSfv+QaGRfkv/Z1loMjmf/1Wa8CA/ZvIo
L95dibJV2bfeal5l75pV70vcCeto8lTwb5x1DzXA81AZtEmyLK713+TlPQmu8rnv
e6z3QzEz9sCRB3rVmRqcVUxwaq3Un36r3a9UV8XmamWf8dwWEKJ0e9D5ksh2f+zd
oDhLd/RQ7wdl7rud7u3HjhYnclB4V8zDkN/ug10nsxaERma+M7myLgBneIM2vd02
cOQTxTlSCLw6IaYEqfmUt3P+sDDE0BEjdtWCcEdPHI4KOaZN0igkXsuBm7+1kl6T
eaDZHIJbzo971B3TInBqoPA8e7RzVdPU7ehy0W1qP9YkYGIxs7+r5+ZCJXVD8kob
gZak7bLYTr0zQCf4D8VIm/0NNf6vXH+yJ+bYXFXdqngUz+8Pj39T4LTNCil9W9B8
us/SUCAvaGZfbSF2pdw9GesBmNIWYOA0xJNMTD9+mPl3Gcorm/OVCEs7n81VywSH
9PKD6QdgvCIyW277J7an7H/6G8LnWsnJ/7atfNV7QMaaRr/fZLEijY9B7bUfNEoL
WoHw+HL/1yUlZqIFO+EhItclCnAPotCvGyOD/2cTCnyHa867mRg13EmuRZSOHTe2
hU6turPhPvkr1fbXbJxLUsNGg8MyHmqhqWuXQy8Y9FUa3XNJzleI7up1EoHMbeCo
Xhd8bB5rqPDcJdNfqHazww45OlTivk41l+md4dF6G4WKU/3H2gpqODTEsvOqwB5l
NMwpZVuOLotn+u/amdTis3BqsnBn1vK8b8NHalnRc71Rjoi0mRnE2MS8abYjMTfo
RH9U4w6D1H10hJyFwFE5kiO2/vGKX3gtO+kzmugDqq+GxiRAJUtx06PU73LKPMSt
/CXz3/Th74mbQf4E/0lBy0TKIAGEPE9nO3ZCuRGQS3kkE7m4Fyy5r2GEa3gFUXYV
6bmV+uTeodwCdkQNUAAqbv2EcIKLIH43UkuvgKocJl/5SL1gr7SeD9qElgMFDbd4
Q6ifk0fdVePVSkdKG7aWQ+jEcdQKC7QcHOYCKua1E22pdQIKSU8v/Ovh49YRb9vl
rAxeZcLP39C9gjeJDI0MJuk4G2leHZr1rfmN92WNNMQxwTqtxs3kg+L4pKnWvVkf
VPdzWKTreVr6MS5U0YUvOEhFbNAXzc4dBa2y3K0m0atDs/Etn7D8wKstAYoTzMTD
CaPQjEfA3lfzQ/n3iVA4WqD9gOkEDUPdQHZd1otRayzZPp+SeQRxShCAclwJlKgQ
jlEud2eE4gg2/bNm+kAmoFkwXTcmRfd1xcrXJZwxjQiodO2kOZlJxB2uz3gW3TRZ
31XVvaCjtsgPWSgMF/CSR1SOVQdrYGY2UWxhDm5Oj2kCHCky/TBai/0JKhwDSNTv
yokahValGb3dE0QGWo4l2QAJNf/Aw0e3h22HQaq3ucl0Z6QI7ocsu9/BUMMNlnNq
xNXYMN9/6Rdul1ROvhI2T3bcBdV36eQO73ftk8x6eNKZgbm31Hod6gpQx4KTVJsl
q46iLmLRgtM3EtH+wjj0cQC56X83FKKvXA/fyF8jnUoCbHrawhbhotjrMGttMDbo
ZnUU9ARLxHelX2TCV7jXKvx3EmmQVnWVT9AZKmgVBo3J/OPemtJZXAcWIhSyrmlU
rNqnej5YltFWeBQNu2fUFbwNgaskXjeTGeTKPrGY8ZYUjiAigMOOZFADsuw7aQ9P
a5gIG2TquflxUvTr92Iq4J2EuNRVqoLnhsAKmkxKPcpmMNpT+hjKk8T2Dq9/wfdG
8drykI8z5Cw/1fDl1AjKuxCDLRPRlaST3scGXHOaS6oKShltETPKl8KKl2y4FT/c
6OSaI2PaQITcFahnE+zg3gOqntdJYseZUgEmgjNCF0GOetE9M9FxreW6rWcAuXOI
/pgiySPgzDH8BfECHKAIUMYTQN5wlF2bRTPXZQxBtrkTDzV3+679hZ7LA52rPdiC
yTaqErM9dte4X7C3hzVd/KPOmT/K3hFcaSG4gd4HogylQoHxHjMkUCIE1uiizQEL
zU7006opOizpE0K2zrOMYGGoq0ryVicgNb/wHSCKco6IunR4u6J/ysuKx6aZ/68w
1BhiPAR7oSXpDVm4aOCum5qy1nCiY/z15BXncobvzRXcKdKWduB8s6QSq/HNt1LL
Am1IZ9a9ExvkOr+CO7YwhLCDBk6of882hJB2u5D+qcknkjV+kYJs83X3NCH6Agy3
yHGFMea1Rl2bdvmzFbcFmL0R24lqv+bLR7krn2PCIM8R08rhQRbEf4vjd0GZhFB+
Fd44chmI6Uo1Y7zfWyBsFcH0uTzz+rjkWA1r23KkeNZDsuUj0TCjH3zsDLIVBBP9
k6JEmeRel0cVR4WiBJASU0DKgO1ffJeM86ZbaTucos8QskU8W10DibvcakQXhCSZ
0R/v0YctF1W9q77HnYQNA/nS7UmGa1qqfz7oauqbEL7qojL4Zv1FX3RsM7Xzxpef
AyhvQww5XkJlgF5C1Zr4VZDYf7IEj6VAhp4enQgmqj13J1sPn6CKJakpZ3y4vhXo
6uQmGqr5DeSMRukqLt7tONqL/xCsb4AAvtgmftNv8h8DvesoIoaiUEXVzk0HpbpH
u9u8D0OhYU42SPc1m0fRxmQLdXBJT+r/fbMfK4724zX4UbHvo2zqXLhX2IfSijSp
MdwEiZiXsfTQJ2b6ONH3d8+Wb2MDDilyr3Ymq4kwmOu2GDmen4cYIbT6NvSDRfTR
t5B5nr9Swtokx2gtp8XmJ1roDAzwp55PyHp15J+Pejy90ZuN2255MyBKc8HESAlm
SCTNnKRdxiB1nSUl9Zf/HzdlweK4G+QJOLmDY5WMxpX+0MYZO7jwVmgvkEbmUQFT
9gbT/Oa8IX10bp0hPXluayptgEz0Q4288sgiLxioumcC8C6DRdS+x4c77QYm7Avz
ocFBgX2dbFDyoREH4UM5/mzJsX5gqILWGVa2SZTCQd16MlcBPFv6whazQDGx1ED9
ywM5U229pe5bJAMkt6wIP0/ZFaO+cG0lSrX+hV12w2/EmQZ5bRqfXGQ7hdVKGxG9
bRfRigEwjM+xZ0l6SA2yUMwMH0ahBqTaKMjH9wSMynjmRrATgW6L1lU7mtqqRX5T
f8ycSc1j3iQBfV/QxQ6O2azPtbWbTB6RiFM3u47hIdI/WKTrk+pa7NQD0GBF3Q99
paWTOubCO1Sd/ZiArKslG4BLFtIisp/PELAdzCJe+T0JFaTOvjVEfDU/269PgkEC
wcyBUnAiOI4uB1N0BLOcZ6a/uszOcFYRKim3EOwa3h5+LYhZ+bgSI6CDYHwFoMJY
v+lAlyx4NImxjmwJ82xKKwf1JpKOkG8qXkkrgwql+Tr2uV2f/++LZwrz6fhyHfsn
aVOg9lsd0TgDFa1UEdGJ/Ckc1XXFaFH0rwyVEgmG/drU8KfHOQ/1HIH/z5G6gOYi
ZepE9RpzJ0EGDeLgvx7ok5ijijvXuOjUeJskrSF8Kz52jllWZtrmSQnBeWRt8gu/
NhPOJlIi8O4eJRdgYdsIKnqdNof3cOMcoJxEjxHVX1h6dvXFZ1N73bhdFVW2aKAy
T/5BaJAMOeaApaCN4BpIZR1159tHGJkLVlRGUG11IT9kCDZGAP15mI/ASqInEKVD
rpLcincIbhn4ZZCR9oKV1T3kooY++McFMx+CI5U0D7gHgNHX7i57Un1yhTHIjwD7
kPli9akIyZPWD2GUlVjWK9/hiwKaAQcAkSaXUHYzz29MfLckUe9WiXFPJvls7CXG
ORu3LyZdKJbVCeTB5LJRqkBb+q652ASLLY87l9oNauEQMiBTGeEZWAt6zknz88s/
To25VNWuPs51WzuP2UgVDSFGylc+ltv9ZQdRwSx0DDYqHcjw5I5yIlLf+ln6H8//
9lGcTKjwNpc+Z5L5TI2r/gvrC8Se2nMk7ThKHB0sys/bFDVnxdWd2ysk9Hr7KDLC
RDRfmk+CQQQOJJy04O1pEGrMaGBu/PnOkHPH1GdUBJDhflXkkHziwAE0DILvcjOW
1d9AJJQKOY56d9vAh/oKLqBCLVAwXJ/jitjLUq8XawArbeApffj6zhcfYrjK3pJz
YB7IKWBEaVZdimWJnnfnC3jaF4xTxFQINBXRXXzCylFT+4T9u+BpUs3O+B30VxS6
ol2het4R1vgH9RJKuWdrpbZrBtjCYX+jpZ/mVHLhLijuz49RU2rXFxyAbvWubscR
/2KwSPM0kyS+AnXI6ekUE0UTv/xwhYWKXg0BkP+2QpIffCoTQUw0f6yOKypwpyEV
UbFy2b7NqzsHz0hZaeEsDqPG+/to6gWuHXNp54a+8yIneNLWRn6PQNzGjyge/SkA
6xyxa6JVpjOQJcs37JkBFYg4HEnN4hdqQ5V3kBcczVxa3VXdkwi1IK9h6qwUa/8g
LxWI496+N/hKlLjbP2bsvfsnPUIVwQdgDQR6/rYM3oFYUaLCPShoeuHX25ryUlgU
wd2xH4CBIPAWIQr/sBsq5ysilmaS9H9SBG3T1Eqgy2bgC2bLcMYCBMufFi2XHfat
8EpLECYEycmsB79FWTaxUavhTPb/CB1xjkPmrcCFviNILPt1EMpFia9HyklgVlkH
4JRotQGU2j9H9nfCYRIC6fPiDrHNvSPi03HrNU3AIXACPhHvO/Vt2Tgl7C8FQjQ3
dkAtRnRVqIQs5TXkpRPU+dlVdCuqJDYaTHxzCgcxjTjUPFwATnzW8IAZ82BoxPNg
X3I4hElo9C2J1jDSScv/WE7FROQ+fE5r0p9FDSoHqOre8jRDse97VLexjDyU44hi
fXi5V2Fh5QL72Q75sl9/TrR1VKbdtiL59gWiIxHFg5eimmOwAu0sbuY2+mZFkuev
i9asmbsr4Hn9R4GAMGzX3VUepDf+7U10zyL7kw8Yqpi5h7GLQYoVIkMy9DLrqULI
ONqR5XHwFg6eWP0Fcg9W83C1zN0JjPV1yIBSbVThZp6SHJd5CSNHgVX3poPYBwkC
L0ipI0q5aboEhF5qJK6ge/L53bmjV7rjQ1wxDHEzVwrZgam6Fw5OQI50u6EzD1J/
4kXbNDD6XLpSMZVtC89O4vsv6yoViv60hr0fYv0gFbk+YoIsYdqCQo5b65Cxd/xt
FTn3a9IIJbZJzHjcNB16MEsENiJeq+Ea5jGKKgVGhaDfN7XtvdoGnrsbCzRNqn6D
aRDjFWXKk7qUwy8hxw7gx87a/LUHIQ3oYTOMQTKGpLarIcITg7NNssDb5px5S8OX
sdLIDQtQbaxsXLAxdJPDuMutf6Y9oQfiJwBDba6EQG9FyJPYM0NSqgbqdLVVfX9z
NGK97Q1kkNMLRnbVJzpUu6HhG+J4KKy0ywHA+ThshF/KP8ihL2XyzD2YZNCf3XVg
uIx5Q1kbTv5IembOVWtAwzBekqUUd6tmav1XuppN5bGJCx97IypIEaAjETL0mabh
lDweEJbMf5O1Zvg30/FDamJ+qg8rdXMaRDsXrximVAvUMV4NoYmPJydT/f4V6upf
Rr6hGJljg3B7h7dbCqE/A6jbpgc6nnp2OZvRq2eodSt9FP96ZGtuNZaLlMBWrRSc
knOy2RtVZCKazyMO/1fvlKMOOCHFICNvoNPEoIiDHPf+HUJ3WtYrhCiqdyZfQyJ7
n6PvctfTtAtmuzL9iKq+maF+vmDMh+xESeAY/k62YL+ChnxvXc0OwXhMP2diuC0Z
T3xlocU9fMOHDf7oz/JJJME7/uRYUxGC3+8+ggznOYH+ukqDN4IYsNOxjWf6Q/hZ
uoQoSOTYu7W6K9YKGq1sWSstf2gKZArN3K6IjhLb9YJuDvdIr1cF8S1286lbgm03
J4ZFH1ONuANnWay0aq6KAwhUaEYhvVsohVFGmiAJrt1YEJ/1QbmHnb2fn+bJEoZ3
shFPp49sDierLqKWRVhFjX9rmQhEP5aO1JHpmdvTOAe42jNu9fq0MpVRLTgmxgGU
ZvXZa/UmPChWckcFPKDvgBfgJgD5T/5YynKKq+KFRozGmOQEMiybUfZnLbB0x444
VxGjgoC0gCXYqs4fHMN8yC2RmuRe4q5yFoZd1HwhV5eqEjk/tfLeGsIJexxGX8wN
Ftb9pACJSroiKoLMZx8tVXgJ+rMIfvVc0/hcOZjgvnc72x01N/zDhgTBl49y0Dux
IusvslxL+KOXm/VpE/65QH33z2gcCJd9Z4j0LbpNS/e6MVNIL+QSV9MApJDz/LOI
rSGnXH/b1XbvFuoFOwrN3Y+cCsoSnozkyC5gfvvNB7eOMqILCNvXSMZ6ShBNvOtR
7AxEBA46t6H5Yh+KjJSKOc9aCMw+Qh2UmiftfV5+OGxkrT+lWBtKcfNdQkXU5VOb
XsnUKt38YNFmampp9u+c+Et+37FbtwZDt5enKg7Lyr7brGYtELODUa1HQpfRQLOn
ZX8KtG9U8MohT6HE0XuB43ymz0Abkxi+8soWRqmxgpAbCIt6+EvXAVo61Y9W8MdF
Dk4d7YjW79JxVUBUcveZ0TW5pIU87XucXsMWcfh2VUYuoGLAKh8mNJtBs9LIqqbu
uY1Xixjj5AWWk23WV9ZmwXh8R8SUQqN73oW8oAMFhitnyp9zdI/9uCO/bnUmlyQi
qJzrxmSzvuBoyINoj7lWIn72yxfGuFHwurOz08YPr649LDQksowsDAIN+ycN8g+E
oqz9VvYHTZGL+prAT8B5gKo9xLiGnqLAv9fuOrhW9IEtEARYmBpcOdIiBy6hdyiI
sWCIPixkwnJOhwheF4STmeCVCJfLkONdN5oaqoJEFNxE74aRN9XSy5AQkxzpLDIt
PVFYEearo7YftkXuRVTbZEtTys9r3VViR5eYg1732bhsWNNr/z7gvJazRLXwaFTU
ryTLW6Q3EQB11TenyKT/juwH+psbNj0NcREnhCcJ2clJPYmRVUeNMPBWyJDdQd8m
hHEv8cdYbr9kW+rvN5NbRZ93M8qAFlU13yIh3nbl2VIYJJouFOWIo7tkRpTgWz3K
bSHVJJ93aK9GjpZziWKifxvh9fUFdvwQp9nirIF8JLJqDajOlgXil+Xzq7f9Bgg7
u+P46oYrtKa42FsPKVmwjrM32gpGj4fZpBhQMw+SQ2y7cCt6USsUYISPUkGe/xmO
368g1vgn78k9pLaXTCuSXVhRwhHFHa5TC0gJCMPpKNQqIYGamFUBZ/4+iVPJNKF7
8YxWkq5FryfsX4U3H+KzqMEni4gCYRdnSAQ8vyE3/uyKSnNSX5moldIxqOeJ69CS
BwLg/vmYdiUvmYUKhbrDt6XvqRUdse1q1Hre20QKrK1mcNzIBDusyKrjemVYaxrP
D0+WD7V5k2giqAll8qBXJru55xZsdSf5hhsAj/2Muh+Tkk/rudixzUNAdmanwueZ
A6JVCOBstIp2FEmz1mrqMVGUjb2wu9pxTHftZPLi03cj+DNYMo/+8YvklTKDElP1
/BK4zsPGmxcYhvd+nwA8rhnZ2I/cUZqmbHy9898qB1pOtHhINpAqjhKAo3z7GNLF
/JHIV/88qjCK7yCPsC9HWg5ztHg6lDL5C/sfCmtv/oZ8StuCi8Ncl9bhL7JNo+yq
q7vUHhiMGbIAW/r+ALqeyFjcOJWkQiz6yQquPSTIckSufHnVZiWNOeKP+Unn+2cN
h3/kbVVrtTpuJHpPkqTAfBSlLuHKqKewh0N03H3Lhbqgb4HBHBQ4yk7JB9VO8Cyr
oWLtAYwKqae4yefV5kJXkIO54coVK4lMPbF69ygMHheGsR2EZsdS8ibMBWIMMBCJ
so1M+hPJIvKEI8kaxIrCiiBmagxkFosXxT13TNHsHy52myJ8Q9+VKvdZaIT10KM2
TlizC3U2U81lkTq6soVIQ6G/zMrO3DxWcZFQAVst5jpoSL7LqyOgzW1R8zBtMTFI
kYQ2ijrXvF0QheWk1W8mKocPPQyeDe3Aby7xv8388QuRjAlgramhyjta4WMEg8VN
Gx3aigtoeUMoFcHRiqZQe/q4nR1RoGSUQZdN6Y7TIKkImZTSiC0grAaBhP/9K6MP
W6qgJ1CPJQ/VFw7kMhEaFkwHFIqA3ABr6ta4E/CWA2eZXIvC5YWsN17KI2ZvLzzY
CZ9DOdypfSqgdSrPiNaxMZJcn/2HHfnPREUyMUlxdQCc78qig+C6so5tr8UeIrsa
oGiOcqxt0eVfzmUbGPEi/di7n3Lg2kf2vnDTzKYlt2GkZEpPvhmOwzca/LlcYL7U
cZ21X9lLPVs9a5QoMExCGXtXZ4bHpS7n7PgN/gZCu49mhESdFM6wguuQVL3MFTUR
JSzA8jpq/7G3tiQDiwoCN/Cp7qQd8rpHtB4jfFnps0EOn+2wg4m2mJCDwGXano0s
UbUMgnEB9H7RTRw1Tx9Dl1h11gHMpa56V4DwzTGzyGLwuBbaK7rJOulautd1cUiA
V4o7lMQpMO/pGkhTObJRonnc7XkbboRPob+qiAYdiJLNoCigsos3aaOqGTzpVR+4
mGX64+yx/9+6KDMakFeveg9m3v2MipvshRufTG0EYJq7jS3rFscOWKZX57wmArQX
fMG1hrnyxsG0X04bQcvviXggGvFGSqg6mGxQYzJP+mMGBp2cy0INNHfltpj9JxeO
tqB0QA+lt/2cNDq6sIgxxbiuAGlfY0LPBtyR6FC6mlS4Ai7ORc9JscNKHC0DoC3l
iZfArowiFhq/SjddcdP6k9XAWDW/qZmr3VdlOiwRYISRaO8TE4xZNo1r1+uJT91+
Bma7SaXvUjWZLXiRZl4fRFfJVbPw3ps6NydFZY9nHQSB7V3xyh/oYzqBplwE2Gv4
mVbLEgj3kcCRb+Dr4C126cP/pbA2nZMCDSlBvaKO0TPUVhFMraW3R6+fxB1CLMJ8
15HirWVn34xRJqyCF5gm5yMc2BAO1LLBztVJvDTc+I2UlKGpdjtcWBrh1r3ec9SH
vTCkHz5MSqxeeGsbvVKLyyheHqAbloHxJnhaY/j/Fg47ggZ6GJCqP5e4AWrS1LRE
xl1Tu9TpnsvdkPYDC2lI5rPdjQnCSxWhMoA6Wpb6nTcXDidlIk3HjBTiWXAy273Z
a7Uh+RcjSMm45EPNL+/yH727i52mKcl4QOp5743L16BaCYkAcWp8NIQzM2/WLiu0
opHf3qzLJ/Gf40ha7o9rZLOVzhiOL2GHDmIgefokj943dGDSGcCpIc/3y4Ok5GNU
JTzq1CuTaIIHcl7su/RVDx+kJXwZJyDh+rtIEcywEuGJ2705Vkq9lmcHtKr+KPZy
vKxF1F4Axzs9p1ioi5rSHul/8Du0m7guRm2A9axSpI4upvkAMOUPF5w88l8t2IJI
88TUcRX7pfBwroQDuf+U3wuQloZbr5WXwp25HU3eyG4bod84coMoRFYvP8o5zcuo
0un+KkaNS11oT+CobnSHOCsXuZfDTHHBL+F8E2WEzoGK9Sc6l2FGwvaA425sbQrF
fT0dXWxZnwPlSf+SSNoNfN7+GYLPTD38WnrBVJ62igl8btknzb4oE9NEDJxuW6ly
fPUqIe9ddb8Xl3RfIzcn6s75OSwmJgIauyyaukH6Rd1+NCH14HPNDdMJMK8VnHWG
/uEUNothJBBBD4sJiPQR56pBEbXkzkX48BEbI2K0SCT8l3BGu6n7AyUu/XducgQG
Yna+pxc+3Tfv4RphgPWG96V91LGHRgNIg4jwOUkdA3NNiEMLeqJ5a6rXqRmBzciw
WVp/ET+6yVcCRjBRLiBj6dIJclUNAvrpgHmcGy2AQlrGvVHrtqsnMxqeBfpITvUH
goojjLA4YKE8qKzCKvIME64qkhFL1FHhhvYvUHX/mCpVAHJQnBuxFJpmWzQ+O9Pg
+0AYyDdDNwJ0Ezu+NmFLAFi2F82515JBe4q0H1lpjDZKzxbRA7KQkI55U+35IUyQ
zMGIKwxG0w9W1wwxz3eCMSIMbOpsKejEY0uDUt6GKUAm4dobqnMea4PHZrQcUvcn
2uI+6SzXz5DT9L0oIvFiJZJYuNL+WoH3VjMtGHFS54fHzy1oghdfC9SfLhrM+3n6
1JgUZ+SanOJK0kl3dA7MbAgBWUoGwzUPjFnpJUSJjlYjnPmxIcnfsA+ix2WjN8Wq
RkjTC3d/0Hc8bXiR9JLZw70EHLWzsICEdOZkr3LrF++ecOtlg5PgiU9CE/skwA46
oRovcUJ6XL8LosTvJM94EZTeLbcr3mXrQUjEI+64n9IWmNEI9Lp2JhXa7AJP+V6E
acjopusQmfvXsMUCvBlWYtXF+pvm3C62JQguiIs6SWKZ9fXkA1oG5wt1YRCcAl16
MgG6iiUrL6R3Zp9KfOi9WE6VURTEToDyusBmqC4b5UWUsm30zDOWJG4pUIXbxSnB
D9Q1ZeH1n9/nVfJ4uWlt+F6/54Ml5heg7Fve/onD6COEf+JJc7tOoGNFTNj/UGwA
2MQSU9vL2TPml8eJfY0PGM1zGJ095/04CMcJ28mdNCUUB1oIvG46P+ANxByviwTQ
63KffBAoZ5NeM4NnAK6SdfYERu1YhRoYsky+1OyIcmCNL5uBwNS1ifac4dD8fv3u
8fT5jMqRPc0zoJapibH++U/fjwxAkV+A/Ny9RM3PVE+W3nu1mSdkegjwNQmQX0nT
Zbln2xSzk+A5qGSP8Zs26Cq2zksZDgj25vVKCd/jD5hEUcdk85qreec/4Q49aS4n
bq+VW2e55DYji8Iura2rUJbmfX6PiU1HdxAIkbs95xJNW0tzSFffOpKONtleHSfP
sFndOsOBOYI7V46rQimoJitXt/Xdg8MQwhimLWYc8dE0DWAhKtaaITyH89BIQRP8
4EiJJnVAt1Oz3TVp0S/o5PuQDhyI01VPNreLAxCcsnrnTsyOR2iXJFLkT5AgpaOD
eXR3Hau6vBGtR4uzBnc/TRjKgF01OgWTiGPHAwi4I68H0VrApjaWiUPJzH6s7wH5
kjeJtwuQK27lzTTI83JJnPIsYGIBasbk0txtppF4/mQboLEqOxft+qoiHxuAIOx7
XFQfBuu6MkJjeuDaUpvo3uHDdJNQ9GeMlGaYd7TC+72cqBdG9Jqy8/kRu36hiS+q
KjzjO0qOLO7whLLJcdipmGSq6/Ng/XRE5uJd92bbWvT/TEtk9hkbRleXsSjTIzbK
gvJgXiASemGo6lCQso7trfRfZUdM1hAh0ATX5wrZXG9ZVQNyUu/8JZX+vPBssdbV
9qb4xEiX1nBoff/xFA/++/uBJmBrkFk2z1JGfLR6srnROphE7TQTEdX85+pr+8jU
w2liFIk2cG6+enJnBnYRbsZpi4E1unl+2D1tTTw8kHJ5VFumCcbBvxciTwasqw9K
48mpMptEyaiNbPYmJCW+TMCQprgWoERmQD9D8OSYdy/i3Ns/3nXSG70zeDsQX+BR
TDKXU2RtKMwyK/naKw7JDNlMhEmEKfAQevAev2OEts9lFNonULtEjcMWq9w9pJp6
753o2OYMa7t8ym/nTlAe1ijFjmxCzAkDf2HnS/vFSBRSEcmjgie7P2K22QuTmAhp
VjuLoEdhFYM+5k9canfwNJkBvcS7Ys3ROkij1nWMsjaBY2iU+ZDKKk4D3wSFaRB9
1qfRHr7WMWkHBIuFWuH/QJoAdLDlkImJppt6Q/hpzXoMS94ZYEdLYDwZTQMGDJAc
SDPO31F9dBf1r5C9lKKfg1isl6KfHkY1JzFNiMWvtK0Au/F5T7KfzvSFDgZWcq7l
0vd4n0CC36H4kB+Bx0rJ7O5u2AvUxGT/bJ1+QylnFATpo6ihsaS10HfyZkfTIsdk
gyjSmRECOw0aEQuyO22BcN+Y2M1rXbeghOO340WD4A4MNoFdRL+nLeCGwHRFo6R6
/etFXdrwvVQZwljHaJhKECOHTis2HFy6IS2vy+9MjHxeK53JCOBAypv8eJyVl1Ir
Wzfcmz6kZ2hX1q0lSZM9pp0M7JYZ2GVpaPPnJGsLy1JoVmD1Ys80CZKFwTxDnwSg
sr1g0qsR0P6oqdwKpajrBVoo57w5vY/8UnqdFy0PZ7deHHz4ZK+q83HdQpz5gQRG
SiqsE+Nwy4qqaTQxB2HUpYYPYD+PknIKsnf8QglDHbyZV4t1AtxS8jnU557uh+fj
by1CKPfBwopzrG47oaXZg2hPLdjBks5KBe1JQFACJdJx7xWnjf4JACd0Ri3VmfmF
COr7whFgMdFKeLA21BXl2M2WXvLvg2rybT2fm9a0DVOso8vr8fCev7Nugd1uJ0/Y
KhQQKjiJFHnCwEbuvvftWvlGh8H+22kbUitw+PPQ95gJee8VJyBEig1x/MWNlOFk
ktHnW/WukvB1AUdt03vfZeCgPLAiTPI1nk9BNqaBFqczMtKQcXWf9IY4REhWB8GD
KXGjdyUpgVIVZiFAebe7MAQJa1jCMMdACaXnYYX+cOQUB8ODHLhNFQZnJtkx0+5C
wx90ruDEO2erpOLUMzHPLIHmnTvJXOVZpKaACaQgTrXEwlGcp9EtPeag0hHQmsBz
jYbOR2lUJrU++FZdymp3aDIA6MBAuSZSmxdokxI1gdvacAaYiNk4Vs02wKOTiCW/
tql1VNBJKa1CMjxjrolfmyBob7XparNLSCzaCMSRpsz9PhB7/aD68BkqiVV4yiEU
fsU/C6c4g+oYUetmP5qPrpr8x2jpodHgBXbalHi7vYywrglPsWtAxUIbY15z1LXO
hvmaDWOrVlDM4hwv7xHjrKQBcl+Xg1/zNcfD+DIhBf4wbsJZGTo9/uJiKrtF+X/e
iE3WYTW4JSV2/J0/qmWWsnFHi3Joky2TNNa6LLtyTeLV5ajkAjKx9YE9P1u8z52G
RYMGT6OlERIbEQTi/0ujUt8PxBDPdsZFKO0nqLZG/+zLNoZHXBq2zhD9GLdBSiNJ
ro6eEQ61WbO2IeeRlcADXEuNj26Bw29R4bDoB3I24uVrgxzFsZGXlNi8si3U3KdN
hKAku5L1Zg/JKKTOox3HzdiKiZWzuZcwtKjIQNHteOOLdlNTUVguv6nAvlsho8mf
mEKWTwBvcPNvFGuUwJixs7KVHlcZLo9Uu3XZQL7oCdNqepv9B/I50aOGODsjHVt8
ZLxJahfBZubvzt9gUeaeIWn9xUALzGr+CslAFcKcIi7+iF0c237eD+SJjFC11hJ6
ZwnnwTpMaIT5m9N/vhqF6P8vjOLA2BjSB9YbMbq4Q4TtKIZpoSEB+JPZzomrG7Jv
KuiD5Ccrg+EsU1sMkgqdee/E/mkRGHzLPeAq/Cw7jQjZPVpkhS1A+gmHkg5FYvoX
Bli2x+4rqXF53YRCpNENU4pmgblO0yaBYaWYszPte/gt1bGV2P/9PK3NIT4YSUob
TFflmHgB4d/ETyWqgdPc1+ayL+1TCFNtuns9haGN8enjuk3PHCxEwDACxmu/Phz2
RApYHOBswfj9rzXG3CRcdcsYDhtuI2gg3rFF5fspdBpGvNI+HlqkpKNXMiN2IVFk
u414nhIYEsSa6Qm8TtZuyta/zgHczFa+OPXvxbUkJqSEYJQBZEYgCqjZdAC3pL+e
4Mk/N9QYwvxB5UkhIm7miYQY/GShstXKKNcJCA8Qrvl1fkwRo3Preda34A8mXDm/
UpgjlVH9tv9og7d3Xq0Qe/67P925bVX8vZx8oxp+cjAscEBEpcp8xKlnbH/SPgeo
U2ZufS+cLK+p0Cx+8JFIuOl6+KedX/d2KfgnHhm5mxsuJz5+1OcJNCcGwFFT7+Bd
WTTE47xl+nvrRoNijY7QZfPIa/6eixVqan7iawStEigFYIHo1G+yoqAwgqD+x2PC
TQaNJyC1qubEjM5I21x2AKoHtrIVfCTkfiFVVCvTDvZaTcO1U1IyUsZd8o2e3LfY
z+SUefDvG3M83i9kk3QmLptRE3MVSVbqIOcMKCHdjWka9R+R0ev0Wxwl4ZiI4VjF
14Eu+UQxH4ddkOs686alAbOb0GJWHCM8ZD9b0dwQWoIMEqRnsdICFztCYDa1Vvvc
lepBbj1LgnHEz+eBZX2FR40GAxBIgrwhFLYujp04vniVYwFzzWIV2LwR8HE/UAqq
BDe9hPlSLm48PiJnRZpHK5M4pEGLPYIbwACK3maupEE57Xuo2iGAVDj6srM1DG56
EHWBHD/3PKN5/l5Vpi/kNXlkfP4THqWBDgclc3dDSvfmEwi9+B2waL0azL+yyI6G
P/BkXfOzofr1w2Qr4uovYVqeV7IjBfppVPQX/ge+bFziGS0JwXeG5II/LIo5fFCT
lgwoJpCYjBp5iuB3zE3mdc9CHsrirkBvQ1htatOzoXTlXNmWRBcLKA3FT/z1Wyeg
fWwwEBkzI7vzEnu2IOy+Rr3MgvCYsHNXxIXf/Ualeg4lOptB7+9Xhoa0GE6F/M+6
dQdXPeFxHcUtvlJ/UPksj6Kr+8Etczch9xTGeER/+hjPcYecalp6fd1QEbtMP+/C
6fsV1vQGSGIHpgcbbAGCt83iQk519bZ5GESEaYljssx69dloJlOC7LA9BS0EisKh
KugSAsGStNuFViyy6WF6pO1xsh35qFBrIcKXK69V80epUGIT6GcPqNHlKfcHrpQe
h12m7tK5UlLwK56olmmTvwH3JEsxb3dg27Lfn50NxxwAMUAlXSZ6hcykbYz8j7t2
1uM1wsOuLNhuOj+2S4bn68qMiGMahY48p4YiDn0CqXFvQ2uAacZmQaJ2NeFGXqEo
8SnGP1Sw1k/Ap20pVRLhsXhObupJvVGjW4k4zyk/gPPWuOiD6EFynB++GzknAs+/
MrQgOuxczTVwpaA6Gtd4xXQVpaclvy+l01L9pXhDcthwYUta3Cd/RqMJXgZvjH41
FSasMa60PDQJRa5gYd+yukgZlfsV6ExIzzHtm+Eposng3M5FMbbN5L48W4cZoP8r
MehQ8hL/YMzfOGO3wtyUW8t4smJCp5pkuqhtfwF/4Yr9h2g3ZDGOQvYlWbIQDWpo
J7wB1tjBGePqQktzcpTunyv8X2Q7RxgqVViDQKYLtNOgJGCzHjrG2XzdZNkXR8Ny
OzbvMsgtjzoLpIOQu7Zgiu4QB1x07v6FJxmbeDavrOXB153tk37Z2yfP8Dnpta8i
y7rin3ZxT5fYK9uWFv+30B3dpsKtCs84tdcqcf2ZOg0ebPKZ7Ql40nuupOTpXrsu
2e71hk+ZgUfUnkhohjVCdTo2v/BHZdyWjkF0zWgYNw4GKntpZMbK+PRdf4O6lb1m
jOaEW6gG1GqBTB2tLJARcyjY7mz/IlmNGdySsBa88b8/LEQHQSqsVkXl0IczhlOY
mr4+TZBghf6rAdbpar92dMnqreIXyXlzUboZDcREVSNHgoksjGG2xTadiHrMOgDS
aM8jLUW6Ayoxtxil5w0bnEngOTQXc8MbQiZ8NNee7h8RB+5Gptvz/azHMdu1nm3M
3AxN5NKWCOPdLa5u7vivUfjmuHH/tnkeBDCXQbB4Q8XWjaf0Nnupfea6ab9Obpzh
AidV+Dg1e7pnBSZIH7NyNEzo4P3CO1/obxxrR3TD9NxhFceBRnsT/v3uaX/3PoMa
nTQICxwMCAeq27eOdXc24aYCmWPmiuXnRZDv6JncLITP09z8NHDcK7IO3A3K+c29
7c1XNqm9nQ8oYvD7xbcdb2L+6Irdnri/aM2F4/YwRjvGIIxUF3DVFAWLGrG1Hbqe
rjkv4zXh5X7Ox5LcLxx5MSC+e5o6VT5Dc41zjEXl/jLt7G+vucVYDPAklhRhpITd
7+dzfgkTsGX/q5Jy61Ygfi1KzUujgscg0BPqXxfdRmfZri+7PzSnbJMXjVXc0cng
GrGcZs4Hy+t8PRu1yuSGQhPEFuW2qNSV2ZNy7KayHh1lySbwY1xsXVnshq5AG/jG
AyaBhqMgJ/gtZZ3JwK9sHgXHSXz3geOfrMmzhr+NwjAeYACmm9BSRSyAARAcotjU
mUeQiVRBIZBJH4/0MyySdv7kNJ7WMWTyr/oTBu+v334R49H5aAzqyhDdhSlT/cyD
JlwuqP8vr/Pc7eRwedMIpWp8r867H5aDLKLhzqmnjialMvDnkzTySyDAPuEduqHd
FBNQnBai66Bijh+QVI+OWz4CeOOroBIXLcfw1yP0M5cRCYAF/thmvjLq+ZCFiQwB
I/o6lDEd3hMdpvbaDTCUxxqaxdRz2MqAuy5/KmA19gogpjPHNtQCw0fsn1zq92JS
R3opWA6YDSWLSnvy0LYLuJ4Vs9tr/uXRXggwHKlw0q0L9XQpsmftTPTbTqNgdz7f
EJ4WVRMToVknrmjorCOSbbV0pn2A2P/sHuPT7zi1CEN0noh5CQMDGqdrZDDCXE4T
qocYMPrS88073Rzh+sV29rylhsIS2pnab10tihgxNZol6S0ARt5ywRpXVgyeSKyp
bxWQ5O2sLmNZ0kEZ2zeJaXwsbJgtewNvRz2KH8neEWDIb+ny37dbamsE6OU3YfVZ
JK3uwRzrR10L2QCmtjCcFTAYxhLvB7h0lyMnDCPss1sMDAzN3guT5msCpQlQsyyk
w17mcTBFV3DrNW9RhSodPmo74gS+ULfD0ByhSDuUSXH/GjnYKAgucDnhbREN1uMo
Y+avAEwFRH3fMMrShk65jYa+MeMWiwAvxXxdvcQlcY9tqAmgUTYYAAzty7IXES4L
WemsxrmOolcddcMmFR4ZxtWLauaqIp6Fh7akROhglKF6Jc7cFzCxVwhx4i7dMn91
ndERfG9GJoodKVDFrYYFiPCSvmA/REOotLvQlB+6wKWpE+y4lbDX9gBlUoq2hTWB
aCXwtpXOpCVnHeOu8ZedjfeuGVm23fE9/Y0EzwzbqomTV7C3xgxt9SmCjNZjhijo
M+vL/BUQNAzfW5hmR8a7DhILENcr1VmYNumtw6UeVAK2/hQR1uec4cQqpHMNXUBJ
F1523/1uBpy+DnkWZlQdFqy1KWSsnkEM0qxqf+rkZAJXjvno9a998aBulFMonB0B
JkmjCofjQt3nlxPZLzJLd3dKNS/CpVul4b2vWY0EknoFSAbwIDdzxzFf7tqSogBl
5JXGyZfKeLTsTQ0Zha388UP3g4sWQI3RiP3wgWYEfknNM8LmewxgnFRKlZK9OLfE
MTWhsYfGawuNW/Mu+1f8mAd1XFO8fteri22sEwNIF7c2wlqlBF3oall9OS3LsZra
uzSnvs+BQCTquygbzi3tCgpjAW5zCVS+mWXju+xDbKHcDJpqU2sKC+PC81cXEPFG
d7CpEXTW5193IxaMSueWwGegxniKvCw4V7arQfTBhMwbODxg7p2Epf6RIlrhHFVx
5TlN5r7N/4MEjMQWEZ35tCOopMrlZxPNU9Q41ihHuUQBhiYN0lixiD/9xb1kaMYn
LE5Tazs4lJoFsEXBrOWhrGwdUbptnNWu4SkQYgJGAz9I1nAMyOwCZxL+K8x/hFQ/
Dntczkh+AfwChSwzU24ytmDVRTckJocxPcCKDccONzaAWJooN7Hq12tqKqQkn/S1
rsHFDxLfZHb1eMfGoU3VIQvqu9DsUJjjaXpC7dboHYuMhbZEMSn/RWbm9j6DQp8h
O4xzhc2ac2IEVutQp6PHrbqLcNTG85V9xQ7KJsmlsAkcVno43gDjAv7tJNA0AHOf
12lpfe3DEpC0Ft3O+tp7Pb7Gy5IPs0SmQE/qFC8MW7WMw2MdPcAlt9D/GyNcrw/G
ynJwBRlwAq8ek6+Ofg+wQHDdZM/oauszfl8R97rshe/XjD4Uu8QQCOUMH9IpyKFW
OIKbZHhcStyee1QV1zcuneo+7qxDRhBMxUVluRm5gN+seLj/HH6xyB4munNDfuJ/
oeKmd8VfUcuEDMaNKpGGFOHJQNXUyMG/o4FwambYGP8Iq1bjju7W8AKI5G0bo4Wr
INhzvbrrPlza4FNSBOmGk2AI7UMIFu6yxGIiuVhUI4XeOyYc1vV1RU19/USjbsvU
Ttl8me1LlDc5QMPvj7qQrbSiVH7W1Sdot3kea0BjdfWcWekIDa6F0B5n7BJA/d3T
c50EHd+W3gqrhDTMVz5tYPHEHpwXzrHlmZ/wI/BT9eRWPS/VFXIVisxK4B92nbTw
htoLTldsl8rkMsYdXq67JtdwD8DGrDy+Mb7Lsy4YYWIR5ZnrEKlP9d3JOKvJc9Wf
InQSeaTvnsuCt7nVWDRasGZB9KSTDJ5zB20J4qN+S0f2/RMECkjCHVNme9H2H4bF
i58q2h5ehDqx/EuVLNC/g7n2pZDHlF+kZkAMlOh2G4S6Ys73qvu2XGhYb5pgiohm
XINFVDj32hrKIm12wiNFY/VhBr1ObCWRPh+ywYEISjHOuW33OT7SiYEWhpWY0Y5Q
9vNPA4UCNhTPvoFEj1JtTSBbZiA84RUIu4VNYTNGcrlMO5tFFZqWsye3N1Ok0AS5
AjnXETOf5aTdTQqOVigoSoODE0OkwJaAJInBWHHlmduIioJNlsQUAoFUGFPsVzcB
6QTFuJpfw/Zr270Oyz99UiiwngWzG/BQjjW9D3H4RJG6DJufuGje32GW06/OkJem
bdrSFvCHvVJ2sboYy/ML1pcAP7mEunV9KPwURz+aR4Z/XujQm264UfNSvVsaKmgM
M/dNU1TzOXP0Ft2KFRpTHkphOfJ9RTF5YGcDgyETi1rSdNt9rVH9M2+kp+TVxC09
UDCQC6HhSD04BUw/+t5fV2bcVRtkh6NaQONPG/JRXmcxgRFB8wZ1q3dwngvdeGxb
PShSrOnSgdr+5Q/kfLtPiYADwuyFZB59cPuQ1W4Ypw9V+M1RDd8oIQ6GgyjWW65H
7hzbrQboqjmvTcZHyxsz7Pg4Yzk04I+LmIRDaZKDlDkErW9Xy14o02Q676QgkOR9
SSzrtIHW5/QMxj/eyN50B+TYvXOarjuYB8b9R4GAlBGRBograO9rlOEkqbV4HnBg
LVBqk1F8vmzmbHn3u5oDNwMEZUxhoIeEm5jOn5zov87SAwjcn7QPxM3iBkIVC7rh
s4tuarqjyWmlYSnMduS2a+b101d/E2WyzPoNs6FR/n1Xb7YiZojAZyFzLtG+tMXs
OsT5QMYDtkMLkoUa1XiFrKchyHhWilwpqNeUb4oEvGbSErcUsQdwF2oB6wPp/sRE
w+yhUgV7n22lOSeotjTsDK3LukvNIRMgMEA1McV+ysrLru6vDMgYVVEHDKo4ju70
8h/a185MZOA0SKWB64C482+8LPPtTOzDdtk5m4JTv6QEWHoNhfAQQID8RIa5okR+
vCHRFGgZdlkjokh82oG3fugcs7d4cg/p8ghjRuqaRdHKby7CtRCDOv/CPrvKO0x9
kvEKMnpQJwgxZrWXdxx/0xsz1lhaXTuK2QjGxyv7X2pUoMILCQXUy/H4J6aDg6h9
Ni8qTbFy7C+FOtxSdueCI2yimLbpke9bHQyXQ54vhM+yuj2DRppv81f2OH8NwJZj
DkvFqO8mCLqLPjBrNM0eEfXwX21Wwr/Pxfb//rZxSLdMnkF83hVv9saTjNf83aoU
T0DbiJPo2FixbCnp/TIWsZikxJQEha/ebwVLPqaVzYVSNhxbVV+C5KvcuEYQXR2+
b9v1TnRNsyPuhudehAr65G3mPMeuBJ6g0gkzHNAiIQ0gZM0KPNa9lefRRBENIrlR
vKvqv0h3PMXYFHDrTaeg4kw8fG3zK2nOHACeigXdIs46Mi+EmAyFryM2SyDPZ2GL
Qivu2U59nwo178iYCHkX+WapEzw97//Pg7n1LPZhV9gSZeKDQCbPNYCojNQs/pMk
gU3xeD5W0VWP8679N7hzwubZ5yX0Ugj3b6fmiFGjUMkdUZdkSLcj8evj9hKkWycn
OzYlRKduMPqjMU3ovwfqkCbs1QzaD/gaARbO6OkTndQ3cIKuBAIXfUBYrjQt3MYW
Yj97t3Ple0/42UtegkV7C15qbFVB49gb2RByKagCO8AbHegrlPewURlhbzR20n6N
Nr+qFQF2JOnohwaQZdWMLJChhcnlRPmBw5vjPbJO2vJOF4UgarHjMyWgYYyuiSTl
mSgNZWjZfSss4BN4KFR6yUJGa2aWppKrlv1+f8ZTxikBRBKqHAkPPLy1c5zJSRvG
sTvNm9JDbVlYTmbgfI4+TVqo8fUp3eD4OeV9m9WN/hTxenRSDlXwC+BLRRvxixdC
ykyLnYszD1TiGlBnMJS4J60GGsEkBvCBqRJhLLCHtx2KB9otS79uRXDzSQWN7c3s
TvOroupmSmuUsyuCn3jUCatcGid/a5FVYBowzWTuGfFDIU5GA0IpkEnfe7v74AZK
+SzznNDKvpRIv+U+vYpQPzOL+beHqCMTbG4gAvPR5pgAHSzeDoE8J0rf/myar8Fm
1VpMyB90+bajbJ5XwehRl+KLmaqRMFlIgbM48NLU+eRlLTFNc+PYMfuwGtrWvQ/x
ll+j2OZlFmQdfzppBx0RRWmNZhOKVl6z6S1PRQW1XJf3+e62B+wWcC1dMso28RFV
oGoEx12SDUJv7129TOLQEDarvPT4odZo18CO+RP9T+dhxKBVVWHHIIEjdVkC0mJ7
Z+4Ss54eDRsKORnzA8Ia6S/zWHTSqcg23rYp+RdqemJ9CisKdH7dAF9CBgcT8zH5
d5zyAQBDegHkwl+CeQlUQcHsL75dXfs4ov12vk8xZv3nxkBUEk8F2zJU2dvHuWt3
k8sNUERdPmn0dpjD+ilnvZ4NT1AgLFuWfgHH5Bs+io1P6dw1rJPK7v7Uylzr7P5c
FnoMuocsx/Sd/7ze49TJy7al2YKLMpvlYpUS7OWqL3OXlxuzcKcNzHp6GSOLy6OZ
nAabru7FQI2FhCwsMMNCm/nTpqV0q7IYBaj8xunY3xVAN6rRHC+bhMH6b9KxRL1h
m9toJF9QpYq93TyWg7WkbZaK43edlsjA3WN6V5HNHf7DNceDCh5aj9XLn+HQafip
hR4PjjXSRZx6qVwpMfKumBNwvtZGswqorD+cY8Ay+HVZnbvDOy7T+p0IOKJrZ1OG
hUU1JYAeGHPn3pHubh4V8i1iTYQR7cjiWddo6QCVhtOPnA1DO8ia49oDvpR7kLCn
ffAFSEqtP3fPOkudZ3w9CCbiKDTO1vQRz2c12QpHhwfmdalyFC6GK8TXvZdcTuVX
JkgnBVviB7bkvB9UK0V5dBQqycIKA92z3KGCar/SkCzZ9AOKds/oa0/N1VGZ+QEO
pQ4KCp7ApooQvDUvvE1rYdcRdxOveq4voRaYwJ40wfvqKvViQbcnzMZY/e8ehEe6
xmtspuRqyHf4R9b734Nl26UqExdTeog7KHSGEo+/niANxCAORurJYKytsrZ12rz+
T4EptwdWqh4tM5Pej2HGsOch+0Mj3bZMUQGEiwZ0oANMbMeQZNNteD208JZm72RP
gQQVlWShYJQccTHIpi0FGaKa9fgyzantbmxHvzt18WGn7hSJ9QaOfe3swOCgRTDU
AuQTGlje7IMnl+bGvzpRxa4TIjTh/kyoYpHJvHxmY/Vb6wsIdSHejrCIPjCae9z5
oCSGsPP0OmSxk6lCiWKa+LZW9PXHKyqPoXUSuRRbfL8FfT9cpvXB3UbtFqPrXMuC
yogLDwvXy0f1TCr7TxiM8OFJSIkm5deujvcoLUhePOwpEXgeAocYGcmBuolDxuvZ
gydYty9w9hNZPIXx9CErDTc/Pn3v5OTY+khJU/l6FtzYAhxNXkCPWYiyE0mHRLFe
X6eLhUilgIJaDUMKZC/3ac0IIYejYA/5sIcDtvdTmZ8xmSZF4sFwEbZOoUbgojl7
blts+b3HY94Kc53WSYVLlavEaMjCefcX75/n/TkjqHimvOC3UBbKiEhwBst5k+iS
KBf5H4CYIO5Qwz/itFYlWizcZ7GG37UuJbMx6Wa3C61PpbeGPwIyNhGucbY3waG0
HwYfodDylOww3yZI+dsGk+oI3r54IYfou83FHBLvtjWwy3vGxYVzhy/SRs8zMjSf
+q3XGVfisXdODRZkTgbtpiO0dz+LXMjf7r1F3eUR+g1RHDZXRwqLXl0TyJ+5FjSc
PG5fxwxeZDm/m1rUr/Y9tR0lxWPb39nljCLDQen25tPulEI/Aqm3pHRROgxGsF1u
3HDc2p8UVJRt1rSdv6Cp634j6C1i9xCGsx2koK3lGA7znSdaIrGwuxga2eSRM5rh
+dkkj4q8jEUdqJjLN8wwZY8LSmMFag9IT0qrkhHXeYiHlevNpAGPnNrkoi5QcnS0
WfWp/Kb+dYZ0xb5bCDgJZ2G47p2fq6bitZhROkfqu83WUiY5Xm21pO+lqQXYqZMG
x36lg9ZIUaGiRq06uTFVMKzoUNlxeVuFMpiMtrNolrVvVGtQkRn3An1n2mLFfPv7
yelV8fULYiMSM0E7R+RmPYBkxaRQsERq48nFRAYJJxF/slXlyNZEnDgVuJpvkhWE
h1rzL1zUogs8FpdJX5GDe0dauKFBVHo/Nz1+zVjPTqcgJ4V7/DfLMpl+45tGXxaW
KvgpFWyHhWTVr6ZAsTXqhzivxlqxcNcq7tsrM9b9/qOZp8I8V2a5KgahqzQYVS82
CrNKw5zwsJiaQSpAAjrLlXQICSJngmajzuM4cXuxq4CKm120T2Rq1GpbBafJZI5N
jPTZ/AuYiPBgW3x1IPsL+vQaeQvatUm8e/JEnTYSsQiX09TDNfi0Hw+rUQGy1qkh
FwGrowPgIxMRPLEZMPlsHIeYCb3F7eQ/nqj4eg9X4K3wNaALFu0MP6+Wn5xyZ7Wb
RABwDEHZza3Cb8g6EeFZ4ZHdflQMXnDZevX648DXxhZz4H50U2KuNDcQ0Z2Z4GCS
W7RAZqAmRxD8sosxpk1qLntuYxpo6tg+NZVRboDQtp1okyRFvgla0jRnv/XJUcRT
BzkUP5vrT7sn2lDcPNBe3CMtmEqSfAtm00F7IAVsJ6l9IpHcKZbAY9d4gh6BlvGo
pnKPx05ASzdBydCmuC3mDmxWQxhu+4YvkFRCZMt8JL8wBhIVYTh+VDqzwE+mSDR8
xYgjVsE1d1zdLHisQ6/e575xQHWN0aVQeuXrreQpNMuHX+Jp+QOHBiZrBI09NQAs
xaNjYV65ycxaLZKolknARfgN1W63HUeBB1B8xOGh5RQsCRqnF4GmXV+fJHoicT9T
Tt2/hboWLjp2AqLznPqtQYHVZnbvPg5kgDQgwaOT8GATJpil4/gq1w1VAX0R6hcE
ju2MMwsvjrVxcdqx+w/vWCDYOThYj+I5S8G5c6gjYlSUDayL0M2lw6I9WgybY21m
yhUz0vdNpQqpY+aDfWYofIltrx8JpDy45k5DNcRuKtZCT0RWx1txSJPReaC11W+8
eSbhswTuANeVuHVAl6fzIhWT+d++zP2czugzumUcllmlq6z5jP/jxNNdgTujMTHk
M+XyK6+ZDCCwuCrmzMhUlfH2DH277ZVz7e1FS7qq2u0Qik3tQpzKcF7ITXZUKzoc
HdF29thQhmwTdaiA4bpntpRInwKrmneYYeDjJlswOlQ+Oj1WMJ/coMYPkIv9Z2xM
8lbjqstDOwjFY4KXqyVGUCJTphgbpD0wZZQmopMOLNX03KtuC6eaOWE+FGu6UxXR
jf1ICOlTAHE3roZ1FHwS2I3KCriFBetyXWmx/YidHGjPb1hq9PaCbWgTKzY5S2S5
e5Ec9cMV0U4WwrSEu5GtjSAN6EZqoidW+G7lx5g6FB2rizCKImMYYCSePuanZpYs
7EGyHRG0DNbX4QEavrseeFryE12mGpfoQKzXffp7+2zzRaQAzhjXXMHSBF12cqt9
hKQ79gCWU04R81mKaqwEEiZIotn4JljCLAHN9efzz01WEEeUz7hOUfdiXQrFIRHp
mXvzLv/NhCCTcuBZrNDFVaCUxObB1ossCF17mm4FUeJEE+R5Fj1kTXaeduQ3xJ+E
gUAGZkkvexEhwZDkh8SP3Rky7STpuAW34uC04Ie5XHWFuHaOKvuoRFDGUcMKkthk
YhfyqJtbjEulQep3uhMIT9xqY86mke+bHpj+q6ez+YFfpk912X8maWj8P4S2k5o9
DQNpYN+O4dfajBfPJzoZL/gY2YKueAIinU2pNRuClpPGxMTZhlslZDGvPpiJadZl
L/ZRPkNlfeAyyma7m0fLauSxWnaW2xKOVRBZuDmlL3HbDtfPDXHFUx4/WnwB6E3y
JXlchZ0HDTZ2VsaH3rn2X0COcwqYJC85n9RdAjkyAf+yDxeNjz+MfQ5lZpewSFTs
94fDshjqyQVEKsTc3FwyaTXqrKLrrX2yKYDr4MzOROzEWe/KdHaRtfTkrNRZNdTT
T/OwhOYrRcdUKUnlyOxONa6JxTOcmji5MyHN8jUrF/VbG/oFFoMF0iat1QXx743Q
dydpXbFp42VfNSgLgtTCLekumib15384yZ7oernEyL6hlemMqq8uZvRpbfR5Wf7A
MB99vPtGkU4Z0LUTcIXyjsxbAMPgc/GwEFa2MKl4pn6UbWrGfnK+PIQb+KVtSrR3
G3QF1bn5Kx9/BPQPC6ZSz+oRI/EQ/yDmTfcnQQf5ZMbPVrbsc+QjB5SenWTbmWFC
2FHmeckkGckZWMaz9dWYqFRG2KZNvZHArMMi8FoB2IgwhPwNGTtlNPhGabcFLxye
gf/3qvZKg/RhLb/6QfvynsIm16A6bTDEVqlVGBHPnR0jiB3og6dKjYz1ZRUiwh1H
XtUNy1x/QTjRh0vpW0B26ASm6wx/c9J9kn6340dUuA5C9WheGbmDv+qhDAd4DE4W
mBW3LIbD+XIHqrtrSjD/lg2bMzDaEJxnGd54R/hnK4ZbTneMx5RKXHwyuj5ZGH/k
0jyMKGanJlOwwo0ij2ehArefGboS2zObNY27ZenxHgN3+UaPCIP/kWlooZq14+9W
XZJUB4vUmwoD6LAf5cpODIJRQUC1ZOBEmwz5IMCzBvpaz832PjhT+26sJF2z3781
lxqS+PtoXtrqxS1GqD65o8V1u/D0cAPA7a6+x57d+UYQQDM035gxw5p9mNEeGOwk
kjdwBanejDRAF49y0RqC+qtCLzQz2APFQ3IAdeG3d5AsshgsuoN7OTkr8e0j0iGZ
gggulFR8zcKL9znVAQl4Z93ydeewG9RI/vsVVESkXZyM9t7VPjqEOU0s0V9K0XFj
7M4VmqkEtK4Hccx+/YqMytyhpW6L/uEe/59bgoVjW2pDKq+GdnwS3/3aPyTgHMt2
mkXi0i8Pnd/FbVRaGMLClWWqfTzkw+uhlvEMLXrza+pCDEL4+SN2or2FIfJD8R1N
30M3flD4eIq+LYYBOgGDi5fVFRojeA8u1lNksKT5SniXxj5DLyYEHagiUJAdj4ZC
e0fmeg38iOlZ9h15sOXGyvYKprwjc+S8WSWtkerrzro45kLGDKXXevrj0oxrMP7S
qgEIbnkmTO9Yrm1skkN+ZqGQT+Ayo4lKNSm/zNM9MUWUVqVfmWwLwdmHTEIlkVFS
0JQsZCiweN7ADVNEOGXvApsto2Lm4Qq2UB+GeYoIzilb5tLYhCwggtO19bG5zI0R
1kRwQ7aH2c8HKHPSbbmWnxMgzNQSJKX2OsyML26NTs+oFh0QVKLAEb4H+qeoe+Dn
aQa0GeneEN1wwp4CAI0IOYjiJl58khFA0gvvw9fQcpNxkgmdFcMz/uL0vqy0nDl9
iBh1x1qJTwJxhFOzwSitGlew+8egWfy4i6vqhLe4MM/M8uL/vt9449rk5eDQf80J
d5sb7XY3t8GgNkDIaP2DO1wzUGez0VrRqg5P2NIdiGo+rzt7W/GY08JneHO1pGSv
lTJGRK6EZtBHj36JHDcmhA0n8N3pzy1DtoL70rkFdBsUg46LlgpyAy+Achchig0k
n2q06GY6OVMsxDj2NupFdVnSLALpPY74bQ9eUCQBdvin0rygNL3rCZev65NP7v2K
b1JEw61J2ldmO6QicZlFHjvwiSOgIFnWwi5IVFK/qKOTfkBS1tfIeiBqRndFO1KB
PQ3N33vD5RVfQX7RY8D4sG43o21Pso/mOKAcUmFXOyLIgMOU3TOvmN7jGBiJEDDy
pb4l3RXLLm9v+JO+ss/zwt5LV6WjPTvWkgaJuE8PiEECLL+3z+qjgFJWQ/NJOI9o
HPqiSep3iq7JdHGQtBoUTeVIPsIFCkHdreqI+SJshfKJ+ykz9HrlRbgYOtjnSsNQ
LcO2n/uISVdCjxyszaqZuoL4hfOIIU5sbJ++mzHqiMkSqM+n6Vi4qvh6KMBR08s6
Oa6ZfoYa3TURsuuWlkxQvhQ8W8Pd+qObwVaXqZG1WHS4c+gS/G+XV1YJARWNvv2J
70Nl67OvY5bO8iaJBBqNSolp7FlTcr+bs/BSu74U5JeqJiZNcTqwH03qJffVCYhv
n6xXcSpxTpE6GiudbmEX3UlX5GSngh73XKcvgniK8YIFaRMMJAO1FB0A+qexUbdB
m2jDNdpyN386wlYngUl7V0j0Ql4/znzxVNhdvfoqRi3EEakuKqkMhJ0CkhNRheRY
7xbae21gMI8AAJNKwW9F/e0ZYQ+3lPjq6d9T1h7ymmb7swptYGQD3CzgHsh19Ofs
bS1jy4+0DqfjKJN2vCK1S4LqUTt+sqE9Y0Y92KNy8q7sqWzq03nVzg8WEHe7HalG
IaO1u5lPWj5CpF9jqK9SfjVqRak3UMIaMovue49x+84jFml7a+pMllmFOR/av1V5
1ZwQd0bH9xCkwQV4vQZnP+XvXRjXiVqP5I0+Zrt4gIMaaO+eFCJDCnY8ELkl9k+d
8gC7+Qhvx1oi6r73Jzdo14fRZtHOm2xmYXqxQgWbzt6CbYijgvdn4S9x8VDlQWtE
CzYIZdtHbzgtqbygnHnuHJ9nRWxFBKwUseYO2iUf9nkgrdThGV3kNq6KEQ9mRGQD
pB+oLiY1EbT3SvgDv+b3Ra+89z5zAHMHuKXtftuaNAY4+2AgsxMTv++NN74m1ZQh
Pbq0SZdU41QaI0KwEydH6uuQFFOIpw5UMAZnNg+L1LV1laNVqV4xFl/jKmm60dVY
s7Peq0zeIkLrwNQrr8icbP/dntZ+oa/oWz37vvoO14dhtatJ2iSi7BFJHDMnLvRq
FCVhJKV1nefEx7xQLlhVoILnD6OJy9tSLfWGT1wEvlSnYoyIldC3eUy2W9RnBbWU
Yx5mQJHfNF7a5L23v7WjlMv5FHHtWB0i2U6D5SPgQwfUJAQc4B5tN4NwEBIB9BF8
yORx0OTiTFIctThaNEQqGamuGGNUYm3UmH90kOu4Mt+V5LHsu+NBQWOzoelrzZlw
Bb8RyKdJNJUqLs/G7KZnKULz6A8SwsldAVtU6Xrndwh8kNCxI79qe+6UvWa+BGfX
shfz2G7WyaDASaRGTIgiLnPmXDqbCK4maE17OuEhfxuEZAkFTjA7kbvmtsMwz9KY
B19K4AieMbMAEHH2W50bSdj7UGOFXP7yE3kQpdMmepz8hHd9Gt4qtpdOppUosjRa
SlIxxn9ROTVIPWG86WG0DbcZ1mYuDeZ8jmz+Wz/em8K1XwL+yo2S1a10Vh6McXAz
agLYeNlSIo1Y+V0cGlWgLNWIS+zg1etiOtE1nsONR4uAX8EkmPZcgpi3xZWLoAqU
j07fmBkxcSlkqTUKjFgEEkTYOvBn/JqfCczWfXikLx8tsZIjxtX88PGk3fwXyr55
537VrS78uC8e8q77l/k+LjzpOTkLit8Wq6uUT1KofgkkT7itfp1qZrz1EvE2tZkd
F7dRm4OsIv1V9xdeLgocZk7t+8YxC5DW4RDYhrGc5cAWqKyrsKFbTp35UDhmd8HD
TnyGLiFcNy9397I+KYVLm5b0rmQWPvhToAxF+0xCs52F6DlUe62etpQBRdo+v5cP
BnI9Trx0mXrxSbeb/9ggJGXpmUR2MD7gIgQaIR9mGmEtBVR8z6leEAHd+dBhLXL7
MwKB8ty1bHHkWpcKBMaLhl1QXuzyzMd+auLLQYfZO/xCTMDNkI+vfvnum6o4Aacs
wL3tAx7O+nV5o7VHhQxZE/TaKHbRrkXybZPlcGjQeVcVU8s9169/Yf9XK2wktnlE
dovQo/wBl9iyImgh3capdCf4Gd32D0fZDhFrB4A6Pj8+OhI9wXwDG0gjoOl1xVCN
K9U7325D422RQRuiIVnEn1shZ1W4EhwVysNY7MJF7+b7+IlgyF+gvjo8uH0kdXHe
knigongt8eLFvgZ+ZsZfc5ydV37ikh7/neNMZmsHTrUlpwFeAuAcoXSKnzMYT+MS
Lj1wx0WEWaH6XxheFRhFd9pRsfQNt1h7Ej+gLhq8I5OhrnraYTHvFdVxScSE70ms
l9qz206i64moCF+DLSVy60Q5VzLU+MUYWRyqsCJF4OlPKWQQD6vXz8G9a2L5B6RJ
r+s9Zdrjp0kLVNVoq4Szu8sK+pIuqFpIB8Ghx7/2PgqcgjFiXJl0vLrkoaXCgowP
8tLFQajZDcbgzj7eWDVKcyILtsIzzNPQI0XOfT8LbDLacoX1I0GfW82XDQ4lTyGd
vGI1w0mtinl56hdJo+04Jf0d7LmmB1doStbWnw/jCkMxT38ZxtE3iNfN6f2EvGjQ
zXiht8OC1TVA0jku6bejgVU9tYcu+8juFOLeGGWzXMI8d3YciCh1wtUceSSdwi7R
0jMuzw5PbkTrOhzndUpVPmJT5e342rDU8ZV+2xZ9OFAJTggbhNcsFbO5VhpkK0pT
y7H45TkMWUKvlAKrnSUyVCfGzGZoxQIlBUlYqj3rl1XcyIZvMjHl9cxd8/URwI3d
lNnBX8BHRhKCRIbHqi039lNyXkrjQIStvWDdpfVyDK2a5OKq9qccsq+oI82rnYcz
TaSiYsTKKwPBcbYXgPGlFEWy489TUu7GqXjY0x43tHKAW1OadxZzEOzYvj1ffvf2
tQDWwuZ4x/WGqe9iLe1czO646wdHSTAqIEtf0pdAJdr6cxhHSmML+e+q9mUgT/F8
Z9tSxjg2HEqpL3UKTPRI+r/EaugJH31Nmz+OtnKRiolpR/D98pLkRcFmeXreKbIN
cvUmfdVy01Q7wIhseV9KNcySwfXN7L/K8pl607PinTZeb0XHnRehtHIYmZ50N5qE
C7zHuvAJ2Nys2AvEzyctr3w00oPVfNQN1/3ygJzCmvuSDx0oglQ8ujCMoUDZHRqD
aqm3zB1P+pUrFzybiI112ffaTixx8FZ8fNicJ3cGG4PV1uRgjkXOzVWgwQ0EzNDD
GJ8KxVdjjJdyJ5JE2przQP4sNmMY6dDHuDLk0ifQ8WruXyhQlZbYqaH/25ju15Pp
5hMAJjoc2Dn3biy0VePjZVzbfCogwdPFVZEsHiCbWBjgV+qAVOKukw6+I9O99724
mxPEDlNdtTMz+BSthBynKd3vRC1VUIwnNd3FTOh1x4gP/qWTgflMCJWnHo4kivtR
7zgPBp0G7jexKkJ5UmNVtpxn1Q5hIyhEPZfsH5XHpnP49mexaE7VQpSDcZKvrftc
r0LmiizrFeIcQ2rantbGWD1pSaWEgUEFmE5bu4G/V5Xeg/2xsG0g+HQk3yttHQbF
UcmG2LFOtZM9euJFMdh8wpz9SikWg3w1cUNqDdx5O3wBBiIwA7RHyCpY2PsJAK3x
Zh7UREq1RUSiPMl1de/ksaVTnfpSxrIkz+yHW4G03JgCybHEXHPHkWAaxHFVdKI1
UYJdCBZlOfvJCXk/oB2qrdq7YEP1QCIQH44vFeYViUziRsDcIvcdRrLEYwwrrdS6
hnhgX6VJ2GY/p+PqdHUIWOaKvdLxU97isEo5IGEyLqA7bCaKZf3VI0A2mZQiVNfC
W3fEdtNj3PLtxmy5R83b4bQDD52NoD8IjvI6luGOgg5i0PaDKIUel25Pkys5F11u
94AQOpZGSVNuUwf/07r/ZUlJ/PYQKwkdOMe75LnZSCC6coIBqNExGjjJI/9UUGCc
Z2gLA8TIlzadNGxxgAfOGXGDhCozbSm7To3+Ifl+jH8Vulwv2c9CtytnAWapN2hd
OS8j1NET+c0qQB7YVZ76w4l0/733jQCC50iw+2F2Yeba0tZlaZHv/obj3UiJVY5J
N+p0XRblzLRggFl5D0Zc+5LHIwAsimD/Kek6tcNza7tD0tMufEhphx2Q8tD9ZLDr
6obknA87PnoDPusuMnhM32QJI/6dWIPZlvMxHEyAudq3dSK2NGiLhs42Ajpo2KCE
3a2yOzR07H2OVJBYjFq/Q242/xT83uEg5Ex2+nywBfoDyq9ezNRvldPJCx/wHCJ/
XlPpHOzmBag7i5/8vbhm/C/+RsldH4fVQwCBFoW+Z3cdAVDYnm3Pw8YJqrNt6trq
pQuhI1Rybh6URPTT66weP7c/OD/HEtPHm6rbpuiJITQkhLnBcuyeNHvDavnELULi
G+LrU1+kuBwinYqoiNoxJwZMzQxoz/oUhTJGifFvQdZAEJsHDqtBvGv3D000g7tk
enQk+vxo1voPm71up6aV+wkXI+5re28egPEjWb9dwTNi6aaPdzYEakIn1tiorvlg
5OI7iCnDnUX8xZRJuX+J7YHr/IHl9Y+LsIilkEe2jtVDPFJQV8ioLGHUILboqjNI
LwlJb8FVIMoRswEHoogSu0JjNODkC7/2Mk8ean/Jb1aTiVq5e7oZh3d1CLcYmA5V
SUfJlPKSJLDsjsG2syskkUnXuKoBbrefqFD4wW4zM16PMlsn/BhGq3y008FewQoT
DVqW+kmK7u6e+VaaBRZG96xC5Jk40ojrR18EuOdo/ZAiva+L4CElADOBrfU+wDNx
HbxGzSN/4c/VYF9SSkAMMCDp14J5O6e6S9zGwPfkxUvKAi9nplVUjY+p16zzO1zG
/fyDTwcSiStoebCvMDj+vewSA++Con+IawfTy8B/jb7iRf8Eeou3psi6cusV5sFK
Rp36X69GiiioXimI9iViTtG/KThAeuTegfJIF2aDoLf6dLM9PqNJrqB97iKPP/tv
679dwW5yVs5D7fN5JwCZip+MfVRTMqLsb1/TsRqStM+MSagUFB/uUpR1087mEXf6
d+zCXsI8NhNaeFKJxImPRe8tEKSaaN40CwyQblERz5cfyY4On5Vh0tmczhivisAW
gRJX8ZttNy98Y8OxNe6NCk6jFtDWUoIpZbFuh+39maElJjp1xyYFWBzknBQMNRCg
x5u0TFrOySvC4ggMz1XzKIWWvn8uAUpqUcTS0Pcl3Cn5OICxiH+SWKBWdNrzjTAr
H4/KD8xG/vYA1jgHWQFHLanBzf479xo4UwJolIQ6xmbRdByglv1B89I5IeokXm46
nAmaQE8oONvjTyZQPGF2J31O7V6eRcD3KQAWQwGE+8OBHkujvmVtws+lyxPxCI7k
UsR5YJPbY3kEdTzCqQdtnlgwaFXJxfpvNIy/gwePxJRU+vkcToMXRKcI/O3jsjhb
oGTHkyMrmJdQrOZwV0Rm4rbgdS/z4iRU/v41Vi+OcmlCjZZgkgkhqzDim2od+10a
m620Y18HyTfQkESykIunX+kHj+qilkhVziGkOFzhqG0r7kqrX9X8l9KPSdJfc71+
+MRwfDtYCDW+O4qM+7BDG74+Rqqpg41S3NmsQ4+eqxLLa8RbzSziqwsVsLnQxc43
8DA4yMEsIzy0Tiki/mVI6DPBuWEJrpY7tESQXWrzWjqhk6h7+fgCw28Nbb1MQ5Yw
wxrCOLuFLu5muq7s+gqLa/MoMbPlEbJyFZNv4VxSlBy3Lj2mKJ6ToKOLOnhm8n5w
Ybhumgc5gAm2rJcX+SSaAsNQzdExWqR2MT3bJdJFCBDGbUwyDHVzSWRbjgkNiFHJ
9BehTHWenJjNTL6LKROd23745c1z/tFUyNsEL/2RHjYFLLDj+axVJvyvGPhREDPp
amE03y38kp5wg7iJQ/m7y6gpTO1vwwAJTB1E02EFl8J/vGRIoNn28SNbKsHRs7ZJ
j69TG9HOUD0zKCTNHXgepmFKVLIoB7kR8RlI7u3HN0YlKAqRClXXh7FV4dFhbXP4
AUG8eBxpJFeRu7JzoJu8Wg5gXl9saQxUxkJwt14sTyQEnvA1QbZa08us/8SXQvjh
nMiw4wlpcF/JoZYqi2NnlymRc3cjejM06zZXKyBNWdVYv5izU+eUG/lyxvg7yJCx
MJpKlth5ohBFcbJDDMaFnMwpLXExpthTDBur6n+Bh83bfnrDZB2L16KcqA7Ib6+l
Awd3C1zP1vLFWbhu94boHrhgwAsna0//fOgkguhj349/hsXvPI1EBX+WrxIWV5UX
bIpB8zNm9GdZg1WM7WmnSMeaR5T2c2y37a2GWccjs8mJtJ2GuGR6Dh+zF0mOet3K
JHeFeW8tT8OUSxvoaEKaSFpRBUvru2+glg7UFOKluAy7+TVs70e8PJEX+Owi41yh
tbfWOVhyGwQB+c32ajBQXJQNI807ycQK/HkKnscvInGjlukp6XBHdObB8NkzmuqW
PZPpzgyfXCqh6wW4mZDgAUDr4FNMTmpNpR2U8OZOlWcah8sQA3ceYQW0wzPsanma
MyBr6sFkzXLzgpRj1Ffkwb240UGRv3Bqsdlr544NT9DXoa0yzKe2YXmoDgreD9P3
Vp/fj/+q9cR+6TQrx/tt+Pfjuqf/S/fa6Zj2fN21yFs=
`protect end_protected