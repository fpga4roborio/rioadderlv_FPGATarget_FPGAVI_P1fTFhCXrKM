`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
ddtXksX2+yylW5zu6QL2Lhnb2d1sD00763mmSITNX595NcHTEkwn0zB1Dry37fOW
FufOhVzEJp80NC5qZ/+F0Vk7Ik02dIR0elf3clrjeJRK85K4e3Hoo4xn7YbFUIms
l/8VZSb14+JVGURjfswrIyCUotIzlzVYZ6gzoZwDXIi5gQIBf/gI+KxNXPaKV+PQ
Ufys/12rjO6aI/pPlqSm0hCvftmBcnezN2hk1UeXgOIuKZnogjOsf0iJVX2aOOWE
6pD/psybjbnsNB6kH5uFTA5frkzIzkzl5d9+YDm9OyC+k84E83I/7/j+rk4L2dah
QJOvksSIzN867/4Qt8qYTQ==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="MvBXkzurAa5VTw+1JJ70nePUfoQXBvZOku/SMmg4TwQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
oRtzZL4VJ4iwysPsC8SXYCzXS8Fw2gtZTOskLcDV+1B9Nzn1zTyNtlo6lNICRmmK
ZRVu2BmCc2G+fmzynYlNTnSa7C0Cuel6FYpxCBlOuk3OF2tzAmLAuDyOH3Z1Yjzk
a0aHuoCdIRKv7BrZCdALt03JeUmXKPdOmIlkVGFl8yw=
`protect rights_digest_method = "sha256"
`protect end_toolblock="Jn9CQpRhJt4rnzZPRk+dOpzAubz7omckX1MrFd4p81o="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 28224 )
`protect data_block
gD6l00tciPUa6pDNTk/+t0OO0nC/UTtBwLB41d4inuAUA3i/ALrNyoJVcBnAmEQW
ptbcNp5fxEUJjnOxnedyZEuEBxWRieZFQnkRdF269oNh+Algn4316Ap1bNz207R1
HiiY2pWmGauqo6QNQswgL2lJrRPz9W4Eb27l28+5hPxlZTPEBsaQkbY5oy6TWuIm
VFYzKyR9u7gYyzTF0C+Uh97KqLj0Afhs6plGVBSmB/40j0MO0Fii2jr9czKcspXG
i0O7a//qyhm3KVUdL9jAdp0wsR6PPeO26kykp7IunhGRt4q2jAHwi8dnR7rQnkc8
oRoagKnVtLbzOj/zUWcsVyTkEYuVI41QYOHRvj69IBnzOCOHjEvJWaiSJHDTwgF1
VixnH/SkqsjKrJkvTYiPHVI0vK8k2yKfQnxVf6JGdRBTB1dGZFIVqFOwQ3snAELD
1q917fXr/Uk9BBJC2N2oh8+p4OySUapXw0IlQa/NNUIc+OZNW42bEVx4pPRUmv3p
xnzFues7wOSb0e/UrawLPUbVE4v6pCVTYEGzZv0X1XxYz7mqPn1bDsWe8HQtsGD2
42GmzFo4IcgBr9Gx6RNrEiellBBLSJXvvx26U60p26bKMA3MRAuI2Ui9egvoc6Le
KUGCt4boPtJJmZdijL+U4qxac2w1o4K3KXfw+n6ZCrBJ+w1TfZ0i+WHEQdzXFR5H
oRM4ys+3HRxGTlvE3/L8AVtDZPiFi788h6gQ7WHpJ/gxajlgqmdmpJuzMUCTG6qf
/fMRPTF2FTvzPRZq20VvUZSJxab6rfwiM+ZEArE1DEZqc8zFdRzwVeWZ/rsF/XM1
xu+/XtIITpnne1xir3UAMqZvDqJnG02hrTBkkGHkYEXnbv7+Ghy8FR3BfNlt10uG
bxLGK1rizI9YqLJMwKong1sBU+bkXgiiuvWyNO9XHA6rdeohawpq8hT6AMjlev7I
OqHIPuky2QhmU9VpepfnG1KKBBbaNR1kfN+W/svIACevdMtHGqv43sa7DhHiVasd
/W62ZNK+tckmMhtCHUk0iZorMhK/7Fg4smYxnZEXG2AG+WDH2Jovb7sXq4asDdyz
tWmNbRko0pppw9Zl0yLUmmzhWB/iML3MT/f3AHZYnqYeAspPBJ09wHmyntmkrYQX
iB+mhq758y714J2Errtp69LhlLv6KzOH0L58piYsJnl41GSYPNHNyqLbg77iEQG6
Y0uky3dfuYuoGs64+ja8JoIbDIFWxC7DbtSDcvLLs0XCASefDZem02yLyEPW/UJb
T5YmIQs1laY+CMs7KfXlKFHERtg0prfjzsFunMNSSYmx2CMtvxI6jljVvp3SrrCM
4MFMAVTQ9mxCyEo368Cx/zZO9EIoPddUemyKFc8OJMwHDoJ9/FqvU5qWiker4H/q
w7zgjgkzqdWbBxvhmIZdAdj/Vuu8ZrHeoddOtEwhv1VK1vUMAcjGhN641V5068KA
T3VVBE6Zam9awFhWYJH0jgC+icVWwFiSNlk5XctXFW4I+X/hTBCCU8jEQYkzkPs1
pLHeL90XnYZBLrAxRAMV53kPESgWsZXXAhjwAwtFWNlFfosrt0PR5IuRQDeUNqia
CBDQmu0QU8VrKm1o1wwaw5rgT7zQdGSGl1CX41jyq3wl8MT8bjdFYfhx3yPs3r+5
wl+cwM7RMZl0Ca5oUo20J79ZyxR0vevqZLa+CW4+CN/RmTMIbP/ZKCEKGXwLby4t
7Hx+Rlq2EdgpQpVXn7p7hhjglyWqbb578K4dhLGPe4CQL9lrb1tPs2auQQogJPpv
aISbBwUR8yT6RFDTI6bQlLuPOiFXZevj9LDyIdsTVehWYTT9fs9GbCCZ0erXok4V
5LWm3nYJr6vfaKh1q1+H51njPj40txZAjeTgfCfkHc+XRyRxEh65xf473QoJXWGE
3aBucuYBWIzu8uuESO/inKVFSsX/D/7FJmpAO8dC/C6PPJSWGBUqv804hT3g2GDs
LZo7aDkhUER4tAFBGcjwSWidcf+E9CqKaBULkQFmOeYAZO8rq7d91L9woaZ5Rqrg
XrpIxsN6Ysh95OXQZ12cQXMgpVjy/MLtxfACoA4fFg0h1Gkmtalt6yQwJvdBnSai
1hJzZBjdLY5jqNDDJaDVo9ESsu40I6hsfRlVNLnSG7NAo1CGQIJvCH09+ro28wuc
4jyNFFcJSD+u2jupldUJstrKJw2Tnc9b8piV8NdIR6h/qIse4gaTFblJI5QDKYnB
GfwaGTB1RjrwCpqlR+lxaOgyiYfS2lf0x3nHdv30J1ggv3pp41Qeq0dEK9KUfT1g
i41PeSa85RHrWMDCmsEVMCUa8X2lUYV0VlJ5h92Sjd9G5mWp8TzMdZnlcl+1QQCX
9p32daWD8zdja760FE7wpurxKhlmlZtDCY9ku+PBv8IVtLvjL3Cw0SyhtDplOcWC
8RTWWAkNh7zTWJue21aGbo8AHc1lhD5QttU37WLCAUvFm5x7Cp+DIgbTZvhd/N+8
DqWpUVrqb9LAgsQaiFC3nxM52lA+1QoPMFztHsYntQHu5ujxEHQNmQM+/uuZKG9j
rO8753WURTbXruhVtPyjEaFf0yiARHvIeHnimQZBTuyC4SBpzHdkgtcezyOUJbI8
WZZ2MetbbWvZLLkTK8ColH6iCm5YJqv5gGp7obh6rZt6G72ubC2Feg02OeGJzFs2
FqNsT1S/m+oee+9p6xH+krq4NXgVgB5JZV91JM7D8vj6ENL+1GO/p1nGeQcU0c18
tW9auk9kUM5A4+uVn3RsxpuLvmrOGnwg+l65X8VzaKL+d4YH/ivBqDEtdn6Knwnr
0+EDom3VH9J91t0hN/kLXHzVrCPk7AoK85vLTwretfKQERYhrtuwkVlV9NASSm5Y
zVqg2Gxkd2cdCDmqKggjMLDZUpj+1sloGd2uI9yPH++qoHhSWAOAets7iFvd22Pp
L1+bpFiJXFJk8t9Lni87U6K/tQouRhgnA30a9FrOuuE3AJeu6IlAkhfRKZELlxtb
N82x4qIMjwCt54tQWTmEaoWZ+lcTOKN72nVdorOwghjCasN1ud2KDaN9F1Sm/6h5
POsqR9ePfnoN/MCgm9Mwft0Llv5+5IRNtUELZsFWkztKketGUvnBMmzhTFhGIEO4
y0Ms9fPmshlDJZjnqVRkon4ZVUOPjGIUxTUzIL09AGqc9gNbF621/8w+nwxZm7p6
TbVj8UDytu72XwzGjM+oMjotPGcIUilvEFjMkAc+nzCIcAwmYQsYnEalJFfBY2qo
aVywBsqiJfeYl+z1TfAOdZZgnVIEvp0QVO9VAVTkGFdu8sgoV4VV75PnR/erGQ9A
dEqENEZsFld3YxzJZd1FOZ+oQHv3YCWW2ImDJ9WDfLIUFPGCmBWBL4IIekyAV7WJ
oLyQ7TF/suzepL6hEf1DAaLdh4b3VHK9BtFVgkZJY80gp+Aktbk//sjBJBcpBu4z
DLBZHKC1JsKtYFdVr8oE9GCL6tGu+XJNlQHLNFrSxzMWc6E1FxVruzhMt1K0r9iL
rx+/3fCj7d5Ck54G1+eGKeTKSrg92AdOfcWgWKjSXXX0TAgdw886u2y5GClJirRZ
g6/xWm4s6U+x6TkxasatD00oFQ9jUiU079nN69qzo18Fur7sOyAxbze0EZwMfg8p
rpSK89yR1+LCc831bbEpMOvSHIxeWy4dI0YXs3dQmRqyu7FbvtDdFOXJobadlnqv
r7wUyzIQdvD9GtpzOimwgTvlUUIlwqe43n1yH4pwcVolp6GIujNay8h+lLgHDc/f
o6FTnVv6IiyZZYUM51xAvHFxz92LZrd1liZD9LQg+QBQWe4eXx5kQywpBYX24olv
PC49YMSGo8u1ZGZJHruCOpdT7E+//0wcw+a77WN8kHHQDUJr+VVVLO6lWCJRp3Am
qbJkbl6iW6u55lFc2cJT45wYoEHaEKhDbELGxsgk+Vj6j+/0uBa0/pPO4opjPufw
1hk4pzDk4qtgXXbLdOpO4y2RE9MH5gcoRGjh171hV/iPJgco50gAVWOMkUj4MGpc
KuvItgzGshQLRT8bXJyAEAVJWilXjSKMv1GwOnN7lu1vOtVugTcPokVrELia/q96
rUQIeBA+xYTqC9ktdNFFjsdD7dUvh+9kq6VLXXfgI/dP+15n/4qID9UvhJykx+4h
WrviNdpEhpvqOX2xkPC7yZsGTgaI2XFgpFKeVjNHHklLTXGQVZ4o1E8fFxIzLuiX
bd7q2WxlClMgAbeZCvj+kwyGxrdav3G2LTR7r9mnli7HTE1KcnJsGDDnR+ih9Gvu
5tPtHzMq/i6L5bNzl3zye4UENRT4ITxPyI7GR4aMqh5xqu7VJ37tX8Eh2wLYlVEA
MhklDy7rQHfA690pPDyCRw2hEptNmrdqNd4rIAa06P1B7J77FS8CiPe+pdE+7lCq
Ude/n9dBDzuIM/SlWmpOZAEVvrpFq6+fBOxFo99/2nRPLMwyS0T7Qs2cb4LINlLS
347cvkA1oXpWU+XYqluAEuBmrLiK1wbZEQKrwgMqRIiz6P3RT3SLWPFK/K9R1Mp1
8WudDALt9Shhz9J6qn2y1a1rfeBZsRGewTwvr5bqS3c25DXae++TU6qZ9ZuDBhb4
mr915q+asgZQchpks2p091nJMSNUfRJ3Ah/HPCcx+c9Kmtguj0OIDkgLePCB8+F6
KnN2y5vA+J2wFmqrhtjba5OpDi6NEQbIXrV7g2mHyjh5bkvI9r5ZHqLrl++m5McL
Fxre2fq2c2rRZagt3cfwC8Qdef+CIhCo/iKbu/i/TEs+P2VVUa2hAMFrVhtCRKsK
D2zK5jeKt/xPIvbWVtdxEMqCa99Po7ZrPY0s0u8UJ5R9GSeYqjUa0W0nRmpruN9M
2zZmBneV4M8c89bm7GrWiseJB6x9rTMupE5SHBwMsmHwN1BlLNBkSzzq+NgtJrhH
k/T8aZt9jWTZUAoCBP0wXvnFtxDxxrSOr+fgQcBnpqHpEvtqMweud7NB8FrpvW+u
UdewjrCCuwV8Pl4qwt7s34gudSWHsFsG1ckGj5OZBGovV95o49i+Rb9j0XClKRbv
dSOb+Tkm9N4aUEKLbgMUDInJin/tTl2eYUxCRuoF0xeSM0sBt74P40lxjfOw6haj
GuAdFxUfI0nG4Y7TtgXDW6pYXImFK4eLK1W+PiAYooZ3pNoib636NqpoFh4/8GQn
d7by6gLIuNRIqurKyW61D6zaBdDcKfVl1Nf/9mN2bL1lLWuk04aq4XriFduOLM4x
4QvzT72AK8WuLZ2l6vE2KfnWW5qWghQ03v/l4B4+S3ptwltUhyHBDC9Q7WF+JUfT
dDZPFBxWgfvEpi4VoISpNrBwPywgvWow9nhH6tiIEn5+F8z47HOPSRLywdpZ7FM5
adGSC+jmgLAP9oXJFlBXcSvYbcT0ZVakOjqlIgjZpocZkk0wyOgOUZK+27g1EXSl
zUM+knu4+LdkuKlX/OIPbqHBpzA9MPimz9GwoX/yFoThy2Ob66Wn/IxwayCQMrWX
Ah2Z6wIRiHEikJFJEVdUyl2SFGVqh28yVmugUh1lMfbPm6lIyuiUvE6l7BJAOf73
2o64wgj1zFL8Yh6ozFOgFxx1hSbgG6AQoVaELcXX30SiEv/+3htOdJWpluQOIh0d
dJz1SS1xGKHrOle52Fdtys+UwdabYh65CnVegwwIoxO/WuGo/aziCSi234vrbpKB
gB0vEK6Lm0S6rcUd8vOV0XDpjKDxY2nr3s3COF0uJclL6SKwBPpiIFyUqhsVP3RV
RItLERcvHIqr8MWeaTABujYvbsYWCJ7t05STAq4063CUq80BE4TbuEeK+cdjjIZU
C+rl3C14ZlFFqOBkPFkjDNoMy3dnGc85Blu90VGE8p1o9u+zJoUcNnpOfodXJCxw
Vgu6ip+dqOsrtMmE97MrQ/qbZt7V1GwU/2i76rJjjOUaZsurpfSonrZ8KUODRMaP
+oGgWMXslFi/O5gfhATW80QBt1KkBUMCyYK7y2pGywXMpJBz5BiPNjz6Ng3z7m5D
6pREXBtQdBF3VjgXXMO+uM2q1uQHPpj463jz0nYFxLswh2S5xOxjoMZ/lTm3UFB/
miFbXpI9dF4fZa9ba0MfifEq2dJyZ9VVf7Kiyhaj98x6/v7+GD3cvNE5zQI0o4NR
X/XznSFwkVETRnGxcvXn7necsUcb7eKEExZalvcxbg3dC/QqX5AWYOWv/FCgmeub
Q4171UMw94LtMjJwirj+JquE8DU36EQgux1oM59BFNbNyxRR8KZ13eiRuEU1WrFM
BdOZCtOaP72EAOu8yyLGAjOBZfoEphLKe289AN4h9e1jMCgOlPXNHRf/FYrxypjs
Mqz8maL5sRvoULqNTrhsxIix1ts803DFOA18mzcfkJz40klkc43VcdgdM8HeLtZI
En00YtKQGtkFIW94cXcLhmJqniS5Ee9HdAJOEC0V3mqGwuK0Oh1ZA/75f9irdnKm
YMjBBnlhBAFH0o0w0xEYyRzpCtnekdxyXInJz8G4O++/2NwlCn+MAqZAIpgGX3uB
yVolFCTS/D20q2QmU/jMcntC+8j+ZtC5ta6twh9cCtDJeFOYoPtK2NP8sFr9wJKQ
3n4V1LU5uK77sqFXy1l81Zs+qovj3I32hlrc2ZuuKRUV4slpEBXE6J54DiZlG6sT
V9Qx751vLa5UeSwyGeqqBhQoV4q+ir/3yP1dNW8bChRmFe4qqssXPhmsIuMu3ero
jmvzraMpkozdSm6bM0LhQ1m1D5vS4K6JBHwtzCOwJUtzXOPzxSBfXurjQuckz1kZ
7BrqtvRZZZp/qzX8x5g9oHfSTFxABMyNTLHvm0468xk+LIWW6SLvi6tS3UtSdttU
fMYgYb+oBqc7BY/h6NWDtICqjWziZxWOI4kltJPZB37Q0oII6evtvd9zg5tNp127
MggLDVU6wkJuqOrRzSawyFgDoSda/th/AJeQpDYgb7vlSOAHESyMPGRv3VqVNhFD
USKymByzfOhH4CmyZ7sYuCY9pFnJsIW1ZYWWooVfpa4cKemotmqbtS67/NrgP0S7
uATbYLARB8RmX/p/a8NyFIZ/gLHcAinJvCm4mOiKfqQLznpX3DzTtp6RaBHo7pFv
MtctxZu5lBFcMpUv8IJX6d/J23at9In6nYbgtg7Ov2nLhUKlNKumD8TeZT07BWgU
iV/W4PzYfnswmtxRMtKeGukHu5nl/xZ/yGUB5PY1P48ceYmweurw9cPxu+FTa5R3
hqmnEG3lIPfJ9bUm0m/khCURtG5ZBFSxYVAGGMgxTZtkpQYFyYaqNhwnjy1mQpKc
XWBNBxWlxpUE6QNsP9jHyEZ+8MZqitMGDmewF5zbfQrBEDDEtFPguOry8mfClpdf
WNC8W/AQPwBli5hKXNV+QJjANHXejz99U9QGDBOn6BG0l+YKZy0QX7fbetOqYHrE
g+fQo641M2kTEaBUbgHHJj+C9zdMRl5huz+/BAVQ98P3vKWdz0mFAv/vUmQCncno
yw4Xti0hr8zl66VtSWrBpqMZgkaL7t5zmPzMQwaWxqfqnGUSHLMZUL19zqC8SU5+
KCRWADl+h+ZfRUXeOJ+Pf5jcJcF7gofdVns2UaM/texXKWV1bRP0l56IEjPpCton
2T6Kmly+wb5lAGL2cncZjz1qmPf8eX3HsW42LB9V2h2N/VsJDS3zI4qedtp9ErR6
D1YYpKeHkD6MB+RHUDfUob5NBKJanWPzCyQ078U55+0PAQRl9UGQBuGh1TnG9Hbk
MWcBIwIC1yzhgbeKEJhJPgVF+t1StSmk74C17Mf3Kij3iQkFOmeLeL8iVa0Zrcx9
WUXyENbdYybUIUa61zfyBvEVUBTV/ny44Qnav/5wxRHeULZF9o5bTWblelKBju9+
WQjAOHlHCKMFxuBoTsE+1Jyz1bfahhN/4mROz/TwdHxHWucWeNm7Sf7dDrxU+8Q4
x47nMdHIs3vNGsp3lPA4XQXipNrLJOPpWcZKXgcHeI/ccpuxjnlp0Xk74hOwS2tf
ebInkIHsSm5XaXEFqpeW1Nop98nUQc77EkRAuNDZsv71i+UgUJWzZf88VFEg7Mx1
fduXlXFeAjo5l1r4hzT8A8GSRQ4CkjPN65nBobK8k+Hv7RKwZ9IXD0ZO+7l56j6g
tu0L7n3Ln+k/CgYMEHYlz70j4tu7Jm5gfLzJhWvVSbPaRz5AXbEFVeN3MY9jP4xH
p1PU778UDigmQs4yrswDE/DYsfspnEvV0DK1zBVP1b/AV5a45zsL+86+toIU3+Aa
pabkVQeAwwUyjLSJpA+dY133rHfHTJTkJUPVZGsSp3QCNGCzTkai0Uo9rMR37iSJ
BYYQhi59z5X1Zkobyn7yNDffNvYqiNdfbL8S0sII4xjlzOLInyB2nVaaR9RpuCbU
1ul4gVjMScK3DEDQ3I1Ks6yeBf0BW8CmKQcy/eDHtoYXRb43V+se/ObWcXzhth8k
bmp1zrRT/tPO1I0kQT2VPGwg9KVH4t20V5eHQz1GZaIcBe3n5lZPNk0xnJV8CK70
fYdO5xLqX3AeZrXlOApeaQsPKTDCVvrH7R6QAJVeQQF8H6Xl5YXeWSHLhrgt2UMx
cnKHeAH+l5q8+MpX+1ar9nYALkn8jgeNB54G4gDh2IfwMG72vSffqQ/i8iC2Yur5
oNBYfHE8pd3brEl6xN0sPp0ZhLzNR2XAa4+IlBUilPuyds9UjsozTDo7ZxbkYVOY
TIwwiw7IAPVcJ4MfI6200L+1a2YF9IjnwBQNiOQhHhlqbXLDycN2lEuAeWCb8xlR
FYQXr9sefoyD0n0Mtc5VT8krouJ6jqQiKDwHweXiQdqQlNk68z6iACH1ElioPKzW
HEMkV/Ay9xsFRYoD3ULytxh8D88OU+aJoH8jW60Elst5h8WmKcfcbtE1+wXU+Hk0
wLpv7EbAMlfG6KZigJE6GPyICSAr8SoDg1sCQqv8pT/ddsz/AOfjCrKHpk36s+nV
8XgLBDqTLDfQ5EX2ZmEPQMg47cuRQfGAm02FPyBKsRODKfXShYNod3BCDpxZQ1sh
MAZWuKLkhAtR0RCbvTlyZY0i8/HCcIKYXx6swmJwRhsBAUUxMSRumX4iFdLutVPz
0LF25iYJzFch3SxWS9I42oJxh9+bWwd4JHoK7MYhXF4qQd8IF63+UZf2oXLSo+q6
aRUW19YxNInXkH8L7467DkFyHC3HrojvD3i2iokehvzjkTkcgmranJ3Q4YmsSqEK
nfF45cPh5z2g0mzKnfBDteP4vvzAYhHAoVgnb4NOSjzSTPCKi78oqj6+yhmMoAFV
okS/myepbHorK7rZ9gjZzMkW2x5v73HDXi8hmv9T0j0aNWRceRXr5oygsu5fD4Wj
hbsbUNvdMmtVOjKInfctIYmQ0+y7SriaL9tEXxCyeR5zaHRQ1YapNowcIcUuThr0
RsdsJynmhUmOOFdhT39UTcDH3VKj14PgnD1FrX+9unVOdukJqrNUD1xWTADkFy5x
NiAiwPhxALo0IDAgBAmOo29NGceeoYw4c8GRUfsA5SKGuMypnYkjp7gvAPdziZBg
wpVjrD0ItNOGZh/HlFMsKdS8nqmHaFgeRWt+tnuo3vI9KpgPsmTUolYcgLFJh3k+
ea6B8G9PyQQIz8yT7VATmhhg6UZxn7Thwbsu4gz38+vGI+cfgQWI8FkIJLyjtM9J
VL8l7RzrGjARsDyWhRHniB90E1yByJOFCt7LCH+EDe15n/ZWUPm46XxetQ6NGav4
GxDu5kWmXklt4wUFriZBgGXjj6cOTGwlyiaWcsCwsdT8Ihm7Au1BYk5C8AhrwqDm
4tHrgAo0sFpJOr17b4kKFFvU4BDhOS6ZlcRAoYZUyb+67elixQfmyTqDk/JZm0xW
AYlRreDf+JrBmkCl+MPOAc1VZGUZG8zAK6/aJTVgepN86boLyGjUDAodCmi784qA
461VWkSPH2hMBIPjPgGIZaXevLcTp1e6lprql6AgskUGiEzOZPNuvWLXkN7xx0nE
XdXQb3thgR1TrhHOGLZUWndefqiQxI62D2GuaHIBWgmb0dl6E7hS0IHih9iTsNhB
YPOEUZyvDx0hAnPvzAOVzedTmZpkIkR87+qpJhCT8ah6v9D4/koHW765gN4aYk2M
9gZIaRamA+ZbVRdARKKgiUpVdJuzoGllnXA98RPLMnECxhhEHstssMk02QTwEowY
gwHae1DlB7BzJAVtqTj905K4Cue+2g9mWrEFos9UUdnG3q3+dWrevjrfpzd5QSet
aCYmUBeGNyIIeZKpkJAugzt5t1Vm1q2E3bBcF+oKR/T2sw2LLfmen9FZswERaUcd
Ws9Lkh0phXkbd4vZl3vJIjKoIZCMjYl4B/9k56SpCog6dxWp06QsPihkvEjoxkC+
wZy6G/9GVvR5YKAhed8pSvTs+cEi16XQUqBcxbChkg718zMGDflMLg+GsxwJXyAZ
fW8wcl3TXdHntEcySzQ4SqZbYU7tYbAt4oSZkLYb3m/QwFNHoe8v4MM9a0/D+jji
yRvyAV5pG3OV/NT3jDi+zi37BMJKkUSaSTKAWENi4seWRKgYFb1sI0omvJv1fSyn
uuwsuFAqdy+B/j+LRaAsPOss5V8V1T3Mu8oZ3fm5kDIdLtJMsx52g3spsirKeNvX
4TQIAx/DteyVWs2Iv68e37Luh8skqKNA+U3NlYcfKezQRNPSapDyoxl1mfALqaj+
nEO0P01gMU4mYaAlFEBxw8+b+rh3bnc2K85YTKKUT2W9y9hQPPR5u9Ij4VHCx9E9
b1iHuwHvKIs3o41dV9ge2sl2VoLYB+NzIWhnqg98GCpMdY3mz7CWiMJe8KrYMVbo
R7fcn+YOci3BbPAdNxiFXqK/OaDG2PgsOkN08PdfJ/dd+7z4qNoMycSqJcO3ZZgJ
xuLWYbaQCl/vY9kVIjqmH7OPgBr3VA4A/HMzBi0cqTT1KlseKaZbAtOWKir8TgTh
N9GEVcl9gSzmBdh3QILqkrhi965twu7c4x2jfI3I8c806F4SGFoM757bToX1e7ad
awJGkQ7LO1MM4e6TqpheS58qwt8ISOe7jgfCW+Vgpyr9eTlwXFsj4ke5hPd4G+e/
bjc2r3OjJqwJvPJoJJgk9JbPs85OhHqsNqRxDtGuejPG+y7TyvbdHvDRKf5xXEhl
YpXoZGM5DQ4iR5Hk6De1WttVmTPL2Jfj0mspWs5QMGxPXizzX1XXny6spobIDgy1
6ukCZvEev0DBtqNWBd8fATMYkQdyUrkCKy4T0cUIe4GIoZRNRbD2ueIVdNMmBWZe
H9t3JCFCFW/fzc8XUBak3tI8xYhubP4V2i2z31qBWafx3ocHX3a1sR9n5Bs8S71X
RPPsWJMgU0gXEsBkhDt6jo9+7uFR2aZH5mgWKYHad4E89q1ol61nq3kU8mx9E4PC
buNI2TJtxVO65fJLhgVNyn7TSEp2YT/6S2pwt3HXSt1KS2+bPpcOpi7G0ShYUDnc
q1wyxBosqvNK/mSNHhUFc+Bd9ksw1e98XzjeqzlRq4w4ElD+rS39OzSpTcs3/PoD
zPIEPboJ5MoU2THdZMpycSsaVY2EXqyqlKJQny9lIVGC8aIz4c59ZkUn5EunL3kx
lDCGbBJmPTR2+YailxYFe/Pk/PHbXvSPo4W3ZbqIG7JfYUk9YFwmzyOZxYk05cJY
eSQu5O/Qwb0LrEABlw7VkzsouVCVzedYZ04kIqf5bMZZGIxkaOBcKN62ao7xCru0
L74LOZaOJ9YsPkj6CwcqmEVf0Egd0BVToFdZhTXNmS30dO63fg6b3e7JZHJ7vHvL
8UpfgJX974Fqm2KvgcMiXJqWk2sp8+fneJOqc12gQqzpczJSEU1zZSqta+AvmSr8
MsOZQwPShAYXYriq8LsmWiwPMO4cEgng7MrC9rTPt0A8hQ8JeTkneF3cakcU2OU7
9KqwMULKBnLYtYBiE+TzE1WNtIkllu72QUd4yTK9Yhv2zPZZxy/E24pW7E88SQzC
quEUtmfU2Gp4flQmGumrn6iCnnB9fJ/YdfFRu8xsuzJgHKP82Bls5Kql3nHKQMIi
KzWCpR99V1DMmtq07qFva+pKQr0GEKFtQa0Qz30qnUAFVD09ablP/MZFrYiHZ65l
6ehIRjbFzuDSPJqzxMhOWOX7eOPrrBAJZVXpQGQiVLIo+2YyW25d53v+ClOurD7f
RYUO1j55qXyIndZ3dqc1UI+i1DQwmjSgHMMlc88oZbD6AJGLfzXAjVwAFYgoVJPu
pUwv6xCoYtzk58e6Z+CqIjDFD34xRQM4PAS23OcQ42RalRQK51wFisUtQNEWbrvf
GJFitXWFg6myBwbz3Dly094JwaiVcMXbWzemoyOD1SeyIkRplmhFCBszaffEW7xB
U5po+2MtnlDjwXyNuPt0abp9azZJQMzTcbiobd8QiFseSLqLa3TUWNjNTgB4V8DI
ZqRmY8nojDjT4e6cX6BcIsZMJFA7DNuMJHtD5DEPTjquQqeiILjeunqJJyAcbROL
AXdxxMUMrIRx7P701sLOLkVXQ9+TGvBWMV2Z2shKSRT78QHdcKB45OvlQp4cglo6
1Na0piL4dYeUltvrbKA8kUfNgUxt7GCS+hB5nFKPA4DjvAF9Z9FxOxrkRSSkISfZ
GvlsbeZMWYkImQVt1LzudS+pS6d9RP1/LRhQFU3SITgJztAoxxy0IVdRNoCbDVgq
LQJMDAzL2euxaCmSmwHMltuDzY1eHJ5+YNQAelw9r4wfc0eRQThYvuz/LcjvPpnA
UNBqgdyS3RxDTiDXGSuN8Mwu4+lqXVqZTuQkTM7prMzQ2moLVmRMhVrVdlDji9cQ
w4Dcl1RFuooP9GCrNE4l1w53TQFS2JOuTM5MeTg2cIG+yIqVmX5YRK7xVVy2ZcUU
HKhU5DNQsLD+uNu3741KEnM6V2cL8Ps92MMXzFiyo8XsLwVJeaDNglWXlPc44XOm
mJ86GOix7KhgGqr0YyXpoP2vy993S62Pwpuvlpq/sZHnAp+RjqtB1XIhJAWUJ+/7
HH2FpSWq+e2MTtXFMxm/LhJdukkQKAfBXa+KOOEZv24EKMtRS0rR9y9jcGb5QnrB
EBBC2PeY8Q2DJKEAz0hbAoSJWTs6NrYly/fbhvttsghILal8kop7wOtjjWKhdDPz
gTsr+UuJJPjn22DapD3Qyxus5mEaXTBkyiS1LtUQ7YpCrN3HmBRTDO7IIWToJq3Z
bkK6rsDMTiRXAJdqR5uM36XZkj7d5ONYwyPLXmvEWEUpsrhs4OmWuG/e/mtJY20h
J3pGrDCHgIRZQ21vxdXTrX0HK6XAslUXyUoMSlMQJXu5dKFREIL4TH8FLthTpogS
uvws5w2a4djsFgC2LPf1yoBETpgH27RGeax4yWRc2hzTh8Ye9zqGbdsX2YPp4Ud2
mpb40WpZq0BLVOaoVPTEdB4XqaJ1Qxqea61cHJ+gfBQcAgPRvc4ItUgFNCRxLSI5
iCJwbcmah8C5ZiRjiL88pBgA97KVdyf+RcQy4/p+JSKyYXNWnh9JKXPUoZYiBkTp
U3w11wMsjdGvkTiT0kJaPXSDaIvIKpu8BHJPe+HMiFTP/uSuCih7WKfoOEEiQ1Tq
4d6bVO2rZgkS8lIp27wZiOaCvuF/GSF2oN499eB4c9bIwjDbaHt5o3a5caBQ8HV1
3y3wSYvQKUQN0giAEXPEudEhhJwAGo6ES1IIee+lrF0jGkJLeRKDxCDAORWEJrMJ
Dsj7RdzhMqy/BPJFjd7eVO+LpTcRvlYF8M75XJTVjRpmXMbDTkcZp5BZZbX86+zQ
hXnOTP7X4uUI4d1264eXg6eNHVpl/D/MDM5/87bVIwVR3uBdzpsZHAMB1iS3K7rV
3DCX1RQX/U5XvnUzyfBAIkS8AQUI/YzEFUOGsqQooeXvowK4fqeK4f8PbkzjkRUZ
Fa6YvGFOVMLp0S4hvY7LJS65BaQx2tOqKWV8wlYjRvjPWc7Bph8zOAEdLYLRaK7e
Vdx+gnwWdkbFImzX1WKLFli3vph4B39pq5Xttfdo43HNn4GHEPYiQxfAmD4jBMLu
Ooip2WWJSUJqEVUaT9gREMf2zBjlVdXQU6ML7cUJfhz8n3lzlG9QHAUVs1ZYRhsR
B9D6UqzSpi48QonL+YGw4FxvS985h8/OnG2I1dRoBl8FGUlJj2Qg7yBY05iB9xW+
dhtTkY41r59JUC2hZdDDXzukvlfEmvIrYM0mNCqhsUurONWxGGt2so3yV/Hg7Xq3
BAkOHHkm24fHsE8yUcOZIec43zDu3uHcU/zx+EmeLLd9GEcyWUlh3w+LgA5q8lB3
c0mMmWftLYMTrEFtXT8gLBEoUfFpbCwzCr9UBFANosy2YcRKejV74xmtikenoa+O
s7KAa0jIkx44RzooXLLMf0D4k0W6gsELIndVNmJlRbU6azjrp3F7CoIClgh62GC/
b/oPX1lZbnMVdT2OY7pZQdSK/3DixhP5O7kWNEIsdIxkCFhTrCZGsLXitYt1a9Ga
ICOA3t8P/LLikpu3Hk6Hyx35/zVVyXvm/2sbVDvfBRuYtdtbtZJaRUWBh+fXej62
kEHr0oly/I9SwpNjTTrUSZA/EjJrWKkvW/YzCCKH/kRrlMGD9+CKgPkyFF3ZJv6M
nb9SdJdXH5vN4igNtuaSQhVmphMh3WLkTNaPOyyHvIsU7sYuGBdgL5O8+v2mIaJP
ZlYOguNtA/hV4QUEetUgRZXXhgbhPT1/Z6egP5mFFNrZXrk8xNP4QWpmlGzgo/fB
D/1PEBanlx8wDrAjxzcQQZ62omkILOcBqL2PxQ+OpoE76SCgEY2TsXDtreYPTv/e
6pm66WcRSk2p5H0tcvOr1s539YJUcU+0KZnA9SDY70zz+A0m7u51u8qWmPgEpTwH
gTdwfX0IJ61mrGNmNDEt0X+/y3I+7VVXZeBhRwG74Jh5ehBZJLeQKKrQHn//9BPv
Y1Zqqey3o1HL+7Cy9bG0LkdPaHRcyRs/CYv8LvqoxaCDVdq9lsYXBkhhXet1xdlC
nAGW0M0P14J72RXn6ZFqo7kuY4jE6qTZcHFjSxG6K321BTbZcNii/0krWF3jbg8q
vil2EbgK1oZI7bnmiPJT5NsjFhT8f/mKWodLmTChajmfQyZoqXhf/eK55LKi9h60
8axOViBzVQzMcVNFSvlmt4Tb2GXpE21YVaXWqDrcGtq6lJioezs6TzTLle9gvp6q
dwh0txlYUqwEbnaIejjMafXNan0ENMjt41eCFU0y2w+Nkg2VO9isvQNpzgvlii3N
x4khxzh/RmLl0js1H7vpVuh7YqKubqCIAqmFmVLKXGeW2E84/3o+qKqchsgdzNYL
QGAU8kPOdLfFCcZODGu9Ik14YCPdvXth9ubD9ogPxY78GbY9Qhfj5xjTds6p8QB4
2EWCRObZgaVXwDHJM64EH/6kCKrNNn4RA33YJe33KAKW8khI5mpPR6eRGjWWa593
Ra4JYUjyY6bcOXu+XK2dCpL+lqyluFXeEsmOw6sYDJz3KnsqN+FnW1yY/DlvJ2az
aKmKCRWNZOTTbRg4h/Byvjzpq+oJfxCa6Bl6ID0yvmN4+vfwWec+uZmGqjXkYPwS
Dwt9+y1QOTdT5VZHpRcCv6JHXNlOfwkDBb0/dOiL7lhlEITGywCVa/ysn4eFN8gX
nhw8cQLJ/WqialdjzmRg4CEuHFAZsBU7P5HB2rLR2hswiWlxV+A06wLIdbkbuzh/
BWSK2rcu4blja7DYZFTuX5KLbo6SycWXdWyCD6zYO3qyUGL77DiwyyCYaQaILJR9
mRkAxmLgnfX9Soxe5RpQLykbrsOcWta8fLrQfklYQe7SXeAppBsjUG1GlzFMV60l
20tn7Yhs4NqmU1EPo0Uo+YUoTOVGRJG5ttZBv0491VFNHf7yQ2NbzK3Cqz+OZNuv
yzw0wS3aQ6agAOs/HwZQ5vI73Rj/xgNCbBCHMtEQsb1lxy9p1jEL9p3XumHy8te3
th1juBQotgbP5eqLarJGZSyOFmf1q0Xe2LsZi1QlKu7Dvci43UAyeFM7a+pnaU4N
5lktead3nTOX2Zs1NDM83fnArAQHZYB3Lv0zMnBlDl7DsQaLm50GuW9+6eK8LpiV
mAHbObCnHJagcZzb5hGWqFMQAfEW1U0N2oiQuGPnMF0hBnMyURNd8263TtN5yY8S
LZ8oKEPA2Gj2MpP4rw24weKAcVbGOOuLob/ttRIk5f2gGFu6ZKTbuo1D/JROIW6W
wJxVB43/UznjxgMJx7haCqhSJmZk58CTOq494JXHYXkzOcrmb62J2gw7b1SRyvCR
wqnCqDN21SpzDPzjlApcAXxm3Jm8VcKsKH9eWmCbz/gd7NGqwd50L7FDt3uGp6Yz
SBxswM4NBcljMxjusgUvUzkrd2JPV+zmkiV7tx19h3pNG5BclvtqBzY/F8EsENB3
UjAOyfnEYXpqHt7gc6N4nUHy9ilU5hEmpw4yoRMkVWNG68jy/vh5yCXs4SlnJ/yO
FZGPn8yroRLplnf/328mtVGbRjJdWtm7DEkYSVyLGPe1QNrZo9cCamPgVTSOQBQ4
oqe/i08laVnhSA3lWs/3sk3xItL/ix5TsyJZyM2Iw/Sy5AoYQuqkWqlB/GSHQ4zb
ru1ZqkZQZmvm2qrcwlkUQfbWOQhUrpQeAuMlc3++Ilp70ry4nRkuaJGWlApQfRp0
iHpjQ15F8ksEYurTPdlAYvMOvJSWZnZPD1l6/DMf4l2WUsUQ+UCDNXLECXaVaQVg
NQpX6RloQ0N/zK9A0u2LxkT6NMwyyjTLLtfaJmOZcQMjOnX7EPBTCG8jben38Kgn
uH+cyys0NH3oAj68mDJPvACzVbgHQFrs15BFrNf9SXWFjdiuxnPDWUV1g6zm9fm6
t9K/meyQBzGA17k9qrEfeCBWc9zalJZCQFC8acqhoQwguiZbvJxloVcYrxJgaOgv
3vT16sG8rke4YfVyzlUIou427TUbIk+y+hQfA/NhXoPjoNV0rc73aY4Ule0G4++3
P5Xu+lRCRcYKd7HSch2yRBIJZrycD38S3xc0aajYQUg8MKjsWLCBtOqZ4u2UI9Ta
2brVOz1+UlntEKwJCs7PrXa9pYPxRBUiPe/KEu8lr/lRajz/gGPFmTTxGEBj5VXL
OOrWeQK7oZwAejtzAm+0DcYxOl70umUrWrwqVOgGNC2bOv/bsZlELcHNOuD3Zavx
pGjO4hHB6maa1dk4RXdyyWcPbW/Xap2dpxQ6a1Jkq90IBJwmX/qUy3f854RVIu2R
q8nHFpOG78TKVeooApfold4yTtrUa+6u0VIC7RLZRGwJv4iy/0/JBxmUrIUjVid4
rCS7aRt7zou/mtCZN6gErbLSlv4qajut55wpgRoozSa6cffNfRt0i0FgRdOv+d6I
F5pdSPL5gAe0FIsgmdVQqnkgxDK6t4zATLaREOSLz13sC3KoApkRUdVd93aheXZI
18V6c5WLbnOBP9fpkw5evSTlhdCBstXVgxpD16rq/74C1v/l2X0FSORCN6wf0zcW
3YYzE8pN5U7rsyJ0O5N2Pr05kwPbWrVT3XlEBykUGfM7jIVbWwKkspETWbs8FVhb
d7hzWMldWmVK/AVIBM0FgsROtG1nd7tUEwN9uUju6WKzsDbYb8ZXSIrpcm9kogxk
sbOa7euyVJuwCHDSMJsNAtPstp0UhMnvP50j4fqF7WDqU/T5lYqiRsTU5aso+yAn
Jk3nUMeumrOSy/SCQ47U2MJQ7Co98yZNvDDJTnRqFxSQhR0JJmq7u3L2/erFunTe
8JidLhdAWGHve7XqmGwzAWJQSPTWx9QlE8cIwY+kzF4pwu3F26nDrioEbDhnsz5g
3mpIqAfZ6krq5Nv5KgyU5undKxvBfvh0VnCjRmTQ5nETxmN3NbbEmpefhuTJuZyd
60+UGoiVfMTc/gBg+ggQnjGJ1k3x4Au6Y+XwMRCSccmj4e9HwAzcelbAYje9qhtw
ZZxcPgWt5Hu/Li/UzMEMBnBKJ5J0ZPvS8iZam0ZnszlcgtTOjMIX1jeJSdCOSOhQ
4wAq76LGspUhycci8w17rPxqtGp8QEfKXOGJbqSm6t3DwmHQPrPhFY4RmTKU8q9H
eLqCKc36CQ5MLCPYXhRiLcW0xtTmTjNKGlF+o9K/058HLAs1CHR8EUHrrqkp96NF
mC/lRfiNyEZNigaa7BfdJuvh1bxiRC6/9eqiMyguo2BnfwebSIAxuHp+3DYGDr+b
8fRWirK9uQVHDXkOHQuKlvcXWDKUuNAlz0SHkYu6JMiPcLfiAFhT/yzIGHaKPBl+
OZxM86YLXL1JpL0CP5gBh3We31hL6vpnpWM2PrIDmukqHpoZNDqhO4paQCTfvTzO
AmYVOPXs8XktICLYRQ8TXQKxHerFUcuo8kC8+IuDyoMV+p0UcAcrs8X0pOwrPk/F
P4Tv9j13ftKZK4P1MUrmODj2RYT2QFzVT86MoS84ZPY3R1zfDwJ2adR9Tvtquxyg
FMF7XMbEfA4xNjShu73X2dYDK6lJa1OrMFsnRf9P5UESOIq8up8w7rrx9H7bhyZq
jMF2Il/jY5r8vdAd8Uia/H7uUbItV2Mz1ZYRO2c2SfQ8NZ5vBx+SjOaX/aQKgDgp
CN3qLuKgC8xlWzuvRrphC3FYaasJT5UNGN3kWTrGIcBW3WF1uLcuV6G/ayWQKaEd
FD9DKS2uY7Ns8nWQvrrpEF+6gd7p7z/9DOe6ULwYz9REQFX5rnwVB+m+WT8o1BUM
/X31xg8ag6deZEsB7hcWj90FHLKFHQ8+uNy98ZZ/LPHwY/mFSVLo/69pk95TlPP2
5MLEctrg6DLfIfMoPAra/hg+6qyHjoy4GGN5B6iCFNB2mtJijfiCJbobhp14pwU9
qSXwaXzfhYw/gUfpVwBgdbWiXZN0eewkszjtjTC1PrD/iDgmXLFBnrtiK8cu8GIu
d4Kv6lbbjs0c+xZg1wne/J8dft0Bydukq9qM5cErS4ZU+xSzGsA4I2uncfb6fpiT
qDVxUztNWXW+dUjVPd38AL49xbkqrNUNYVlU4N3eAA9dhKcHLaSVwQKEJIllp0sI
ZLnDRGEJU2QqhSTjaPopEMzjZq5r1sanHU8keoVOrP808K1bx4OJLDHMlADoEFdg
v7NqkQ0SftqIs8AYpZdkw8UcfK942q/QALJhKfE4FcUIqCE9BGc3RsDy98q32KYj
SAqVIsLYe0mpNv06dbrbCZ5IHzLd/0GSQUTIl+f2kHgGfFehEy73DlgbfAs+CVV2
ThumhK3ujlUrCIT8bMXMczO80lbPSvxXtv1ZRCbeS7/OnZodOqFX3whCMia0zCTb
Yiyz0bZ6uqZOImtBfumOhOG/UgwfFRTaR2HP9Azxkcsqah8TIW5A/2MLIlI35Bij
T2Quez6FornMq76Z6GXDOYHwpu+hzWadaddTb/DSddmXlhgXodjjALwGjeYVL4JX
g93CpTFVh5K/NPyyTiSi3nKsu3hD+fe07ImK1DicUqDmljhxIR9FqQ+kwwPu0+4g
cAh03nVVhsBSN/VHo+Sh7iE2ZGbXFo+I3JFgMKacg3tFeIGbJdnURK/EmIbm4z9K
9vIRjfclJHQMubfDxOdU/2tPNSA2pGqdJoi8Ozt82VZRR1N8A70RQQpXyQrIeY0C
HlpjfItobXf/23Cgc03HTTEcuKWYRAD0A1fHTJx06TJbFIQ881CiASqyZwP0JNIt
0CSM46deoOaC/L1uINntOZmWP2YjzWAzU6JiR8uzQIHqY/DZAlrDF/yCqWO3jn4A
UPYO+G0WCssuu/7CbfIp2TmHkBJGjIujMA3jc3MhBPdCHySdPeWR+w4OUqIWOft8
rLDTUKRiBdwkaq4DiT4yHf5d+/Au1Ompem5LT8Okc8K1JtSxdOgFJVsU/RYZuSS+
ryVemD59okl+zO3HQynHag6eE1YS/vHQzsEFVKR28Y7rJY8oNtsh0bXqxDXaaR7f
iUCexLWIQMgg6QfKYSiolDnxUPIKoqMbKIxRH2/wfhRFtHNPKRoUVA6ZJkLVNLXW
ZD6A6wAp5mIiVwBzvmagutdKgshxHIDeYi1+yT2rezA6fr4Yokv8FI4skn+7atdY
Hp2lcMNXYvRseGRY+WJZex1qNdbNd8vVth6YSA3lvbGgJi13sOBlEFgrmKDdoL8g
jI1Pc5zwqtBOddIi98Fz/23uLMY5FVbWH+5e/qS8F4Yz2VoOzRlaervXjPImr8zu
RusYeLFtSt1T2wflxmYdIegrgxo5vJq2UXLffJqH4WiwfB8oVGOUgjQLXDGNTk3Q
r4H2XpajOPe0iil510TQ5pFcAtq6FHrg1i2hSQCpcPJl+ne1HYDp9wIWuHyFydNe
WdDnKqNE5H5jfMV9l2dEv8NbQYbwAYTDKrDz/Qb1GNvgOKL6bltx+pwfoqgIpMlQ
Q+X9xdE2smg6TYKtqtyxM/tszg8jSxoi6kPLW3z9/PlBf1AEmP1Y6Sl87k8dSPdE
4AdgNDKsmzUM/GsKWeMuz3dYYkQxXOXZhanRTIwKXseatX69TXi4AksSXLmuEaNn
gURqyZo7z3Rx2JXRveLz/Pb8RZz+JXF4plF9YhqX0ZIbJ20SxC6J2b9r8mAS/zJ3
bn1mEgpE5wX/LDb/RZKuMyaAmdezGQF2IxRa77pZpJHdr1JGvTy4v1PnnnGLtt1J
mqxo2xbp3wjd5QZltl7zsmq85FBps9CnMq5cGMbjnb52Sms2cF3eXQvRCRNZ/1o8
9ICX/cdzc5PXqDSGRCoT7lSXGCXBgO3IjLPTTeJAkN/mhq0wG/AFIjSjxQzCakpK
bxyTZttw1zm8YOhlEmdvnTH3PB+eOIisKy0Ph+JPbbWoEDr6agQPfOkTr2CaGtQV
Wc9iMBBuyIBZzGHh71sVqwUWE0odmlmZn679e14e8hiVYttNC3Dxj92Kqyfp9Cpo
bQ40PLMoIzz7G5fjjPdpbHZYVF7rKZEvpz2/6VK2zR1ht+HosotnK2X1QFc/m94L
jZzvhRPgwV+TEk/Q1zN1+OkOn9OjaJK+dQnUdOrL61PjUhnlgPNt0FT6eb/BkCwH
pPxhkkuh7UppMdkphI/tEQ43Bl820C10FVqAKjIu1dFcDyGDc/mxUYqqRvngw/VU
K6qs7++S3t024GDD8rBFpUO/3rdFDm2+xNjJvjfcA+jAjduwmj7Gj0L6K//4GveB
2MejP1JHB6cktfi8INV1vrdjTvyoU9vHoRSkx8H+OoD1IQUy8GUGnfoWtZuioeNl
D07vMdLUBlq+JoL0qJJAR7Bb/Z2K4318pwa2Ox9wqs1s7G5blxeoIkhj7o7XG19Q
WNzF2FCvMOQgI8zeOjUw6GgqxAYdpdUsGtsd0rWhMi0aths0H5MmOYI+B+bMguVG
c75EZGKqVpKK0gp+hwCIoj9trrhta4xoSX3zskjjv7ucAAvAqgNdfD04i2LV7J98
Ual7b2xL84MTYFI4T8ne99dapcK0JHyFsIbdeDTvLWGnJaiPL3bYE5YqAIObz+TC
bEofJclzDSpWHFL7w4VKjT6817pJ4BKrpzPeWfemm704FbHhRhJJBRcVB5neFDWu
mK7D56o9bLikQoH6KRNwpYNCFx1D5FlUWt78QkzgGIH2nWkUz5s23wjQpoAhqSgb
ygwJhVMWAZnR4RqBKY3izoDuP0IqKK/MVvICkwmmYZ3HOpDlTe8GNXJ4PIjWI2cs
fqDzgXztRmTE2iFO1GHXbgyIDz9U3Pl3uLp7RfsnTDZZUdhW5ZGOKGx28ni/GpKv
xm4POLSX265ZC9/M4bLL+ylpw7hWMVtRM1ptAIUSFE50RI66Hv9gogKbOToU1Xpc
+/a5PakHA26K7WKWNdbb7Dd/GwOgwaUPwouXQfOpDn1yvDtUDzLPs+JcQRBODqnu
lYcvz4NXqnlquT6WT5E5kz3ThGPUW6hnRgD0lWy4IAZgeZ4ygpW9PoWP6LV5KOiX
fi8YB2wuBByHNcPkG0wsBTO4w9ri8LwBC3ANrQeL0537D1KPJRwpyb1NIGZvQEJD
tCo9Ro7AG/DotmkyxTc7znJ6DHQ8KOnxg54eXAbBqz24znB2epuBphgixC16x7Bi
oPUgYovkfkns5OaAQXPxrnTBg72imwGkwgtYQGhkzEuKknGGithNNIP/pm8tIRMK
VW84g12godU3NcDL810P0Fzc/xMI4ikZYgSzHkmt6CwWL1QYDXvL6ItwhJVKcTks
GZwECRu9CrgGJE+3Sem6ZAlbMI/HidsDuzlOQMMI6NaUOKfc5oBGNRoQzlyojytf
3KQHgdGeQ4jZX7EQXcygZPphDSe/CZxBbZj9NoVO4+1/t6njr6nYh6EwX2sLfEwE
Gkni9BTc6P76BkxOejVV6pprJ3PheLaoRucpai1oQI6vFGwNwqzFmF308MlE245K
sorDrUduPaGmiutvA1WY33U+7mGF4SG/RXlhcvDG1zRuHFq4weLRY2l2p9k38J9Z
V8Eg33TL/rLgIdv60tlwYYr/Sq3Av4XOi9umuvJR87GuXdedLn8cbDbKWjzRHNM5
Iy3pdchVxrvO0BykCvwkOe+BblzDhoOW14syiWOMTPVKdrb9ryejZB/TFlSy3hzQ
9apwsUEeopcFwsoyAXOcJCpzx0CNRBrswNN/u22nmFx9zmH33VzgrJ8cUOwWfoEt
2XesnEm2stxVh67pv96QZ0hlZvoTVreZh75pCMzcaXfv+0MNYVSFNbnwLpM+9R2F
4myHshdiydaD2rx7gqTOAmbAucwSeSmImGZKY76obP5cMAEW3ruC/OEK+7ri4rgg
ohA4h4CjSUWPfNs3O6Qzvcb4lpgf6h/5udVKlX+u9Rp+cTM6ZK3q0eG8hQB+JhEn
TmXo2/bf5rCQH3UbekdsamziMfbas+E2Kc/MKKxDcQa8ytnr6cxsRbq996uOPh4e
/oYIsM0HrLK7Yq6gx1GY95i5mkYRMiVwkiuKRceag8AvtfdWLdH7J8yFIBaxMz6u
/0p+hgAe/z6i8R09+d6UT4lNHlJxabgSV0iDGWc+gC5mgcediCNe5PgPjKi4Lm3x
STn8/oou10HuiG/oTSSTRyt/jmrK+Ig8QDoglx+qBsujVBZGQ+8XH1rx+pVz8w61
suuhxNSg6nBnghbGM2GOrCNy4vUwnARg6qS1/Trfiv/vqfPaTmbHgbpFPnP80mBl
cuhHw2JnnPA4BeGiB76VoVYPcBU5IKzYYVRvp0xkEsNQD5rXcpR5IoKOsoXW1bk3
xqWX2VROY+jdaicpzVEBG0zq1EwPwg2kNaTGSU534FMf5q0dALRio5hRyEw/ea+n
IS/wqoYLG3c0ixN3ftJ7CS3G93tROJ4QmVHzj6wWfCrGDnTjlpM2l5L1xV0doAKx
J0h+MO2eiADCrP0N6seOnsntejIhWDtQs1/uoT3/Vp1zFuCg1GIZfyC/7qGSYxac
wsjXr3M70iindvtrutuyNljrG8Nj1uvTozJH9lMNhgFYAz+gzy7jY+ObO0rra+ge
lIIsf0zeRqq9rEpEOrnE5Dp4w6ZbVwLEQ9IKihnLrYeMw4FXwRxtWV56R8iSQvs8
kyjW9Wg2xtmqD3skLK6v7N5KNhAjBOSDUlWHBngJyDLx07khT6Hz32QucbtuXFY3
S0L3LsqTqJtYm2/oSfVRKmMIOCFh61RYXKA2kVSM+96Djfpp6PF4+nxQnmFSTmKP
EwZS+bMFmdFF3TtYEhpVNNRPN2NbcGMalTHb+VEjKxCPviV/YG4UZZpGObe9yam4
9QtRdxU+bp0hJ3+BCieC951PypiE9DftFSW0z1xKAUJ+5IqAKKILDhuzsofoUfvE
c7fR4qGbPdRxXeNBcS4PI2tEjH25aVQnx0Hq15ycZ8COx+tEwWnY7kmmMohC4nFC
taNLy/zXQJvP+VOHiVxAODf8xF0x45hyOaNmPqQDpQtj+fkyTAcLoJ1QLd1KeLo7
H+bw6TPXxuVA13aZhvM0baBy125q8KtyuowpL7qH5CjY3oGumEOiqcw7tXtnO3I5
AMAn2zN3ifotcK0zmNF5H1DyA4VLV7MCoOUPK6w9oAXi1QdOPZVJFYqLAXji8fY3
f1/iTV0lpvfNRfVFpmDhVdhVBY0nXrAZPjMcaMaQHbtOndNI41Li4GWrPFaztTs3
7BSpdIDc/+KuCCed4AlA72b+DLkz24Lh5uAX61llCdqqq4eEUWSl58KMjihdnNVJ
ipYWjkdMxcqhBe5l4LbZLywC8+fa/7O+W8HVgcM82+utkExZe8WkQNBLQpmKhhMM
9mk/UdpJeqn1KrBP2kgHArfN8JviG/PgUfO1UECcRbxqT5E0OEDxVBuXKAVxHVDP
d7QsucAuxZ444P8O+vMnuhL1Ctoz5csKopSY8oqM1IphRrvXQkzgMzl4tUglEIHw
WoPcVvU4jpvF9eH0N9t04y8Xhc+rJP36+GaCXWvBMO5lkCRfleRrSZwCivfB2PK0
AKKfOOfN3wCiYW2y1IqrX29QMXTaKgduItI+psrtC/w9qugKJUhmbW5m923b24/F
uYHBhfJDuzTHXwSFvW1ICwfK948q4l/R15u0xiKtZJE0P+FXNbcB0Jyw46pRkd3s
tAIJSQcKaZdfZ6NFrjYgCsSNYhXmHbS/VHTl9w3HFwtOJnuHRBbYTtC+K5Ko6a1K
kYRyQ24dKrJmf5vI1VNZMnj96R1GekP61Faa+4nNP+7KtRo5iUjhQ+jT9gWJHMvs
82pJT3831JxTw03Ysw+4RklVsvaC4cHpVdJswqchcgkK5p+e70t+Py2dLoHyt6+6
Y6+OvgjoGKaYievm2mDtbi0+EMKVM5AF2QuYs0yjw6Tx+cImy4Tll/J/LEczPmJ1
Yl9SPOrpDuVivr/Mpq5QGsySHY5rmM+wcZtlMLgO2ISLF3oEsfCyMSPHmofPD1Yh
4nZNRAGKEuEha/DjgE/OD/Cy5vebYDLlQ5uwRhdSMRqLP5/960wbFupHwhRLdjWT
hKqaYxGhxHOGwixF0dajL+SRZajBelf0a96YkHkAXhYV/Gnq30hWwlRg4IBYWbw5
+6ovFuFvu1gWx3WYceiMmOQzn+oay2fBzHjfDyn+usqu4129rbf8g1jaEmLAgeI0
izrrZfVpsq90bs7d2RVc1KRTg69y0YEfsyaa6BquxWDI9ZuBQVAD9bVGQqtmuVmG
0V95KK8T5uUHLf4IA/X1QOL0oRr/C9QWH8gdFAaEDlbJEIizoLoMH7xjIbZUt4/J
SJUJB6l8U+5FUlNvXRa6S3T6zZRnGEBWWYNg6F16/i2sSH9p/j8Eu8gF0PLmNYUS
P2pRbGUMpkcyGDM+DZvtGzcR/LF7D/Ld/CVGn7jmRcYl/iHm6U8wwi9gk/hv2F3H
9n8p3frR3FJ2FjGMkleAftr0qLMrjqNeaAbP+aYcB4dk23Ti3vdVKL76mE47+QVM
wwJGR9YVTHgudjTgUwpKvxr7OKwLCfnalZ6UHl/h9FeLcTyuV8BGQ+vIp7pO2Phi
794sbe6EevTLGo2eg0prCQnUCYPE8rVGAJ+TrzheoeibLlQYi7T+r/pEsumLlF5G
Dvy8nuY6QDbU6HWhXK+9jhrLdMVnXkZZzEY6fZpdKLah+mo9oD7SMp5F5aKmofFL
sMmiemaFR+pGG/ZE5Io3XT8gp33fhd9/uqgcBpM0Vu4087NECHq5PwHPwe6V8lXT
oLuyjcO2AFcyJdNLT3j4ExQZsBA0J67r6kUw2zUkKcHWKu1mk76YSW6laiXdtiVq
ZM8d80WuUG4riuvExTfmyyOs7H0gVW4kEGBkU/yDSpP8RMog4M3/Z8oI5dWJF1Ds
Bi9dkboo2BhAZRKmQNgqGOTvqdROCqps6zqrhNZ6RIdXQ6yOOMhF888Q+94ogRRG
KJS/EZ4d83PGpoqhT7aSaYSMSmmKAxP/5jYbG/REsiyc9vWZFPJIfwicrpcwWBoc
vtVA2J9qCHbxJtQwSg3dq0cCX8Pig2PGTQ3b0xixdyuJ3iUXC6DazGCcOGRUjRHA
w+eyFwWpx0P4ILmeQ2e9EIOw6ExArufLFjV1IixQ9MgWtiF+4kmPX7v84C0RvFlm
VhN3XDL6hM641E4APvkCf3Qv6QjMt6fDL2uAYZHWsl2ZdtiNg3LCPeQO7LoadH+T
NZ5q1RWMcSmCPwJ+9WrRf+439nDRP88UvzYFa1zg+OIvdgH9XvHiNIqlbM2kabyS
k953x+8LLrqRW1tqfH9+4s9ffKkPg1TSG2cI8BUFTfPQp9vpA7V7V42poaYMTrJF
V+9YfBZxcFqeHTP7C8wcfcZBvfYNIREBem4V6odPQNL2fzJjvIWXAkmNr8bFdW7D
e1nIgDxskbZYWu7bfoVKkhIKDA8ZGx1Ha/BicGaigVVRpVp9U8BMJJJFn5RV35RT
ZLAGELi3pGh+yFXqt0/yL4FHhTT5BZDBctjsvo+rGbtg3oBPrpgxii8fSoOufl1n
2z6MLrxx6SKwnK2R3kQLHY2sdjF3Nlv4L6GRMoPXUXrX518QafEMgNYxhj/YQeae
+JEKOjfuoEWcUrKKJ/ynIvPTv816iku/utjv3JumMA3CQ1ogXho1w5KIh3Ez01Gx
KNSsMuz+rtw/YzrzRZJhfOp9iI8kmcCUGZypYGzEoVFAByUajQSJJvME04COGDDQ
5q7D7fh7n+whuOANzCO0OAes4wDUwptiyNUt6Cm33vGYerVd9yfVwem16+KAfujf
0D0av3ph/BCAGKYs3R0n/NIvxzIYw9tDgxeVCRpbmOfpVMvQyClqvA1lp4KoHC14
izCscCN4xDrQml+8zjZvrRVP/SeWeirL8QARPktpy6GfNTB5ecP9iBz/ywAspDF/
O1BASiaJlJpmY8ZzrsekbdqLtvHkB213mzQC2JuyYV1DVtHQuT0fBWaiOpruazui
PA+gxcVXfGDSnojg0h2SNpOxNCVI+n1WcgNUUj5vLbgV0MFn7ynC1S/h6GKYvhS4
OVEOncAVmAr8kZ+rjGDanPcK810T9Zorg8xE1IfIM8+1AOGXWrXG34NQ7MrhNhJW
TCxutkjeGbpMiJQP32zqRbPEQvuLOSMycMVOVPfvYrDpXjB+qP6JO5SxEOX1UPfh
BUtctDq8TCHwgh1bNKC1sRn5kPC4jleTEztGesjyoBzCcyMeayjcuWixodv1V5pd
tYWUI8AIvHUJyr6ifGX5jnf3a2wMsTfVCISpZ6/ltzYxw2Q6+hAUXxWKSjBCA51I
Gqq7RSWesPle+urTuK7hQNAz3yaLyNKk5MOdZiOI0PCXeXAII/Gq24eIpoyHMUgW
+SFC0KV5VnOZUyYp+kVXE/SS9oP3FM6iyjwXIWFAoae2t0BV8UUFW+4M4QR64vCf
CmNy11vTdGVXngjpuXHydftxp2f4IdmnUXLKF2BeW4ziGPjuJyvl4+8ZFTeoSM+Q
t7cp7MHECvKx+jLjXjTo/pHEtTIufTAzOZ4hE8VqHwyudBJ3EwGFx1JNtwd0dPaH
mDJdBquZrOiLQPH5kJusXYnCMdiELYISSj2wu9mBweTB3Sn9GaxJKKwtQH4jv6Te
74o3gt3D5ssnCLgKL5igN+mQxA+g5Cru8+8kIm4hFPAjewU9G5KQ5cq/gPg3uBRa
2KKFeJjSNBLnXDYCddbRJOEqip9o9n06xXM9MQYHH7y5cG4OdPHtu68ok0P3pB7P
leeHGD6TN1Bvu8CW0PnmPK6XXH+x15dtrSVke1yru4eVNOegCFigaEcJFgQ1jw7t
DLsnlfibbNEk5nRDm4k7KrtLgC97a27YZUBSu8GjK0sgWm2+aD8FArES7X07UOLT
LuqvzZdveGE48QbLksL15Fuvv8z+mAJ/NJy8/4EMtZ5IXFeKpcaGlDK+29qi0r+m
MTD9/U4MnvLTEmhIXdQLcX6PRVXeTKxc7qzn03/dQjOt+0lIMVPdRHG+pNKFHESS
bg9/SLxeQY1r8CP0zA4JEgtjsIHKg1Qp7vG+hjGx/LGjH4JUhg3McxJHmyduUjqI
+NnAjdstFtju3eH1v3TtKdbPnX+LnoT62XRK+01KZlf1H02by/WJd5F2J8VMvARO
fZO9bZJy9YmErHBvwfR2EvvSUrW0mEy+hjDm1cBS74YnOkjX8J9pHwv0RbgeUgLy
9NRtrkgtqtNC+tYCLM4e0xzcT0wsrlXRm9i9QQZ0wyXzacLr/ZNYspNoAsdr3Xwp
4a63clfjJKjlE9GQF7owLJCwA+nwBKQqKDS5A4XAgPUXA0bZq0dL0LcGVuimqgJ+
djAjxiQdPb0X8YYo8QOi3SKOUdWb6cU7LV/B3RJvSNeVhbcLuSj2KpeoVceuDkxk
5Jf4rk+g7e9hMjE2i9FgQGjUgxsw3OzilGGcQBnsW2yxn2PkO5BpI/THq5eDBnqo
W+YSSQWCuyHhLsQ2FRHvS8xvfD0YKvYkvsEfVbgRhf/NFurBSGuV2UFM2t02Cqr2
bigEP9lhk0NJDD+A1x1H+kVRQOzpur6Oj6l1GY4w1JXpNOrgNk7SVi5eCy07Rxvx
vzTaGjUbUggJKO4miHTBRHcK3AtuHzwYw+FWRT50MVm2QcH8VQ1tEHTX9vkmNWSY
kuHkeJK9YZh8NvWljecCD1HQt78Y8bJTdQX99Rur2v93Ft6c7Z09loJTBqPaX+JK
5RL3QyILt2aoVr2o3YkP9e4r9FIVbr0k/YsiouIJbspiJJ9yLJ4z+rgWjfxLmhgc
+rv4pf1wq7FA9xzgGVWnt4qN+qBb/UDvP6Rcqv1BA7UaJfQCrbvJ5sF2inXlYKoh
VycHvbxRLIW6F3k5VHbcsiXejSr2QZ9k9Xmeulno9vElij8hWVkxRoLHMrhe2/q/
fU7VVcBiJPqeLpwSF9jsvpUDt4QXhxGuSFsB4a7WAOOgoqrTUmZNGlLthxFxEVuE
iSCF+OFAUM1IsSN8k58ERLaG8DExahbKaLBDgU2IjabYSrSTJpIDla6AfKPbJRb9
nCXkwEU2VkD2AKodtnnTvrrjrl2mtQ+cTLRGQdk5YEFUGI2jijHFLUvworRCnNNx
Wcw9cOk3CErCrLqopWfVm5sAadLUDET1gpSzhkiL5SFhYkRDP/OU8D0IVDz/nxV5
I4VIPNvPDKnPIttHikI2ZUv+G5yC9O4cn1PaynlSQZgQKjBqmt1IyXbmSYzzqA5W
EUL+8wjXzXDmLl6pzvvQn7FUFNGraCckFkj7vMZEaZI3XwkOQHQofBtXecl/HMNF
Ufcozw5EN0uN4n63yiz0kqBljdOmptRpk5gzYTWk/epgInZ+XHrXRS+zR+PUZahG
3af+rVl56QeIn3jKbs27H+31pEKaJGQNKXh51xDSpz+BmIsUuMeEwE5pVUmtZ0M1
r+wc3s42VTVEh5T63PzXSsnZGId9zecrKcF0RMldA4o+qWyMKgrLdeOhjcg5QPr4
BmhftTfxAahM8CO0T39/FvvOGROQTlcTolM0+w8GaSo2AIHnsCEkn7oeCrELRa4Y
e3gcEo1AeZn5HmmdmgK9JEOld716r7jcV0od2nICadgtukdufw+4Em6YCiE75YQv
cS8iER9ld2/pLpJrxz1AzDRPArZLjUeJigx4kJDu81RpFJQ6BTRNG8TQ8XC97dmu
qv1W/d0JSsQDuf8vg8LbSYSDoWHSqjkJIvKiBYUqM1IQ8yXpDHdcSvvTSGSF8wEC
Eau+sYotg8ppTkSLYdmhnkB1gqYjHQdBFs+/EQsij5NdysijB2iklshynU1YayKg
okhSi5Phlo2y5t2tjNon+90fGago4vTU2ULk3Y76u90gaYYp9cOmG6bM4KidJ0fE
uvOQAJjRxxR2j0Hkna3mwol8ATOCkbWSKIbL2nJBEWY8i2r8d1zNYHpXJ5kDtmPo
Nm1EJruBXjdI4Gwxg4Y1CVQGwsW8im3GOB4RQ+xUmEcFHRgUU6WE0/VAss2ADYU/
pg7aIBI/0EKO2TcSFtgD8CuxYUF+MvM+Cb8CJwyy88RFihz/aauhq65pv97dF9AC
fy6c+4sHE+cxZhDW8rZKHnInY7py7/el5IjukZvRXOyiYuSkTlSS70uMexOEAuHe
ZeNE9Mrjv9gQSTUrzYtMZLLdPFnJ1fZnk6dWJ1WE3yC2k4ytMnUsh2eH6RDcrRO+
Ucy5u44awY4O8VLEEH/o8fzikySxB+Q8ReuvSP8YajiM0BA/LNblQT6D0hc1NkDT
P+pzep5jZSHGZcnZM7sFdioEmtgXOk8b5yQTwvHZRWxbDmuLnWFHJptUXbEeUpCy
xONS4KYKxoSceH+ns+gYxH8lDZ4bCPFxiHdhlIbIVJGmU61+ZAtlxvMVu5NyXKZE
Mr8Ig8Ely/iplqmVwN33kl9AjzJhfdS1Z90EEISxe4FhYxt9MYmRFxm0Cb/P7ANd
6Ox2YkzysUQhPWKp/V8A5x6AxCUYTmpa4+rmF5/Z7GTXSD1UVd7JUivafLrPF4lD
97nWVbWx4ze7utMAFK2FFV5CNHGU2Bk0DR7Bj9sLDEBaLRdM8IYobckOLL6BrqjL
ESyXZ0AwkTm85XnDCliktrnlfbxzNrip6BMFxY17/74zKC0upykvSlOABOK3BtYW
CQfYHalvbT+ynOlt/UpF6GufgToyQk4TepFx6oJVMubIF0eNy0sddajUR7Asb3Iv
wc7Dvr7JPSR1Nuur6gz6xB1EFCX0dMzXPZShKVX9Aj50LMW/fb0mm/1m9uxzDjxk
UfcMWrMa0T+TElzy/GxkyL3r74iYP4W1XfXwX3uLkg5uWflYAFGewrUPIl77VBif
iaMIcfOWfICarsRE/5C/6LnCUstktTOysGnbN5H+SeftRO5ZdpZ1dH+sTbVldUv6
8+ZBC0g+GPvr31yCmSI13zY7PfuAGlA3RX2A+KIjHIvHaZSYug63qoU21J4JkGAx
ITfe3Kc08MkHMIP8L/oQ8F2su9h52eAIGIqrRtmSZB6vse1Kf8AFwQ93mVauovwC
0oRCVrUaWKHxuoW2oTcmtvPn8MuPPD2qniavljYWL0H4WP6GzliInLaMUFmo1yWT
YGI4JTZv5V0MePqCn2Ff26HDRZGvtVQr6cSn22z5bhrW6/Ji4+W/obN+bYT8+rgs
/R2fbmt4vkVgOD/apUrvsaMYStQiJjAdtIYgrqqB+cGb6oILouOUxvggaJ0sd2Je
JFwbCXJaQjsY9xUGU9CJ02mjxjZ3kEh7qDFD1tw46YMurf2xk5H3f/jXfbHjv4Bi
BcpQ6zVueCFhV9IamvdtZmObuZpow0IemW24llK57EbTDK+TIo93BY8JtF6l89u8
A7Qej6qd7s4/+alZ7t5dYPXzjYFLwRXCEc+50KgrrcWOjf85MzxgN2DQYujMaZSQ
OPSDZX3mQvvoAF2lt39SoKxk3SveYXOswkX5oNkskPlftWDovPr3jQNrUFFYvyeS
Cn5+Wkpzbaz5nm+EfEnh2iME6Z+ZmWGDWtbqSpkulwN25IaF5TcJKWx3FL4UkLoG
b6nhBkyHc2ICDbx1WxCcAByD9egfcXVjUwcxo3InL5/hF7hmsq7KWXFyhKFfkr6A
yM6s420bDaGg6FyTAqJtFG+1i/LZZdJUplt2Y+6K+dbg3RONg8k3RP6ly/ROiRrd
z+Zn53CfVXtom/QKdpVOn26AL2bZHGiiW1pzgSVRsGS0OpueNI53jzLX0MF9FO4B
FAmu97gWpAcchE1gvKS6phrdZtgW4hpLZhlS+iFOl2t/WL8nlxd+xESqoYETN47K
Wuo5Yu3UTVmDr2uQQ2Ke3MQ0adzLKgFBbFZ9tkvDd1zcKCIj6NwMrxo+nMpYNslP
HH8+RWyxDdwQScI7jj1A2b1wrHy/4drh+MdZ7FQE04i34ekwdU5MlPu0R1s+zlf8
zD+m3sn+3PmxZIn8e2gVpXbjoOgTFnkO9ynr2tbiVdbdrmaQLj0hW65J6zA14/aQ
0+aAUBbGfVL+LBMuh9Nl+M+XVw4O6Gk9ntkhk1NjjdpECTlmeSebmBSrvpLcYj6y
RJcz3FFW2QdWXhGUPeD3C9WGkF2wE2b+MEBqF3zvEZ8kbQfRx7Wcel3RBcDWgxnA
gz29JWtecaZqsHY8PmgUydftepATJkskkrVNNMHOI6iBecSwh5mv7EHPjUkLCODm
mshyrUUvhZEueB64xS9RIWfZC92bwKffBR0jPfQpwxAcRZ9qEUj6ZhtYIfqKiCjr
gLqf6ObsNnu9WNUZjZRc9G1NHrO5cBZ1Dm84Ujwpi9zQyUjUOtDX+Z1tzA1b3/Vh
GrbuPl8vLMOnPyrFyv/wvW5QPcAQNY254DByEZ760fAReD2PjW6MSUxi3epVTwJL
c1cjqkGw4GN9o7FgO/yh6XcCbHIaLGMH0G9D6i493TdCDVh9McXtCzLhFEtTiLTe
UuhojrBasn/nm+dGtVxWSQgPCNIwjiCy9dXmSPi57j6KaroSslAte2sAohQNTNx4
Jpds5tq6/xfdM43mRnX3DPjkp5EGABAPeoWyxmhYUzt8fnYo6G8thH3xmsoCu82K
0SGSJtayHPfspYk9Qet9/nSBRn3OHWevmmOEDp/Kga71z+e7kMI21O+u6oK2Zy4+
Na+SA4zFkHPoWJ/xHlW7FzWAM+hkN0rbSVLHJwrYI33+CAguaaFpO4u4Srk5o/TP
HqKNHhuodQcnubfBEotob8m7sheiU+iOi6J28jYQHRXXedWVSvAhL2mME6NB/ffk
CaiUtWzjlY1R7RSLzLDu915AJsNlc3msxs8bbyZQ2vuZ5dOUGps9WboYXonu6pU+
xxXs/n/xVefYX306h1GqfArzeKGhFD2FeoL7TlInllwABkLLzzfrJzi1whOS8jQx
JqZwMO8aOHDjyefCHzljRQ8szy77EdoyNyvPVmuBYNWYTQYIxxnVwpTksCyGjW78
uDQ+COx8GqOtcIIlFAOdWa+9ekIH0a19ABVbUbsl5SqK9hDve3eiOL6vbDIeVIFd
Lpiipz1Vlxok3B8KF/RMm0oml3c/DBWTlxSo2j+qCGh8u2zDSD2KnoYc3c0MmY9e
G5QX0UUTswCyAWyQcjzo1dkGC2q8Iy2Vk/wehnUF50vbDaGMBkAT+Sbr8/EG3S+S
3c66yGtnwsOoR49NC02q32jFyTNH++/riO6hPtCukBOgCATkk2dYar/uj+39IhdD
34lIQH9W18EZ1AyieCLdSdVYhbxj7GNZG/CpuYWhYwzHfzi46n/cDiqu6Q9n1Byz
C1bdEpvE9LY+aVzAMbnrSAoDMIrSQPpb6s7pbnDg0n6ehV+OYPPklCi0USUJBt1E
K/dwYwwBnO8HuxZDJhsnet+OwZqHkMTBUbpBPj4p0Dvgsq5h+WwyOvkprigTsRPB
t3TAtoXHnZq5J5vPMROUHQdtrjxNV+VOfHMIWVUAL2Eey7/gapPEhrEgkpu8ruV9
+NkTGnzIbFo34/p8ibIEK8cTp/Zn22RWsQbB+umCb6hbMoFjNj3ZvzKBwFLR89/H
u6wDptAPvvE/UPc2BqaQ3/Rsy/j7nSxdIk/2myjGMIVZ7aPT2S0GUdXD9qS6YB6c
6wCtMKoLsERPytuCyBReDrzVwLeJc0KJHpL9FzG7W3v/vf1dg2gnmWv5WWxRvqS9
ay1I4f1cd3lOKIBcE/vjgmmcvfXIe7s0pRtqpljEZ3hbc0zkfgmiAxy3HIgO9al6
mVvSgprcEvYaZwB3V2VmLbj7+lyiRti3yYuC3FI1g91VpiydLQHmLKL+HG4jpOQ8
Au+vve6LxZWQ0YgGB56ul/htmywCAQ7C9TVpw7/NkIK3orN24WLc3OP6VsgSLXav
WyWFLEkt06K+qJUP+ne9pqbpVAEoTDmICrCJLsldHpxBRs5QS4B1Wrm9cpl1Jxp6
Y7ZBWCqL6GoNTB92DG+ejsy0dfP0HeDTKEnQyvyb0yhSC6RC6KngPY3IKNVm0Je2
OGUgwTh1cun3ZS9JpMyCXPXLEaLs4ZV9EywyEJo8D/OB5ANkhptJv7zarxmVjibT
NCrJCT1eqUr0Fs6/AXAPzR6rz1RosGw0bTSz1BRyBFLEhZu3jh9m1CwyXtLQYefP
w+XXxdEZSyBJDsOfsFMknHoDSbv2rAhYzWXt1pI4i91wm4XotWaSNN75eJXQ0l1c
eXjRjmk9k4mdQUJIEFgwoq2aAnyw3hteE1kPVvPh5J1oPwSrAswj9LGZ1O7p2X2D
1LQ26u5ggL/K9VF+9u0ZxR3+T12RuT039poQvZlYC3JjFDHZKM39LTo3dv1m5aI2
7G6NLBwdktt2KuKjV1i1ovZ7TiIC7qP0rIOLDvxp4+SYGyD1KDrOMpBj1G8roBQC
t19x42ww8up65C7ZhTZv8uhT6dL19W8BE8ca1Jb1xLe73kMhbYXyEBt3QEecOJkx
KBIUFlZCzyMpy16jG2GxCXRPgNxmXre5k06aE8dI5tfpiHbAa7uDR4nzPR3wwSjh
msbLJyqpfcPBXVJjX2WEr8HLHuzLSEWvbBo8xoUtGlva5ubIYbdyb3xguThZHIbY
oPZ7RJzvjnL+l6SLE+YSoSjDdvw+9w2U7EGIr0d8j8zJpiOFWU7wwGWbxt9TrsE/
tLULc94Eoei2GjLF5QScS1vVG40KrAc3dQ+npeu2wvn3yPBurrBD/nWfIB/EDbQU
HuPS9GyXLleNyzeNVDzcBV3BIBvX+2ao3E24C24Iwiesk55pybkLJnP9LsCmFmaW
yP+IDmQ/3F7FKSoFvXusZM1Gse5IlN7aKurBH8o1+kMMrAKH3LNqCvnC/oYvKX9H
e90fDJmar7TBNvuWMPmNxRyFELkrguPb/n4rSzDq0nDVePbBoqhsCJIroOFPgmdc
Tgsz/G0s0PX8H87OR1PyF3Mx274jWAl0Qezi4zlYt0g+7i3c1Tyg2UTh0y/4KrfV
zMBRE8+rh8foKjbEoB1TN7+Bbqz9XgfJJdXPqQaaixfLhlZ1aFJfuIGUrjjVoO+q
5lovEuWC2ARX9GWDFoq5G2V/2v92n1eMNzoqjFfOlgiosXZNbY+r2gnT4/c0xYhb
AKF0t/xptxovjsuG7DNgovC+vrzYeNyW69uhB2Cozs4fv6aTS3mYgHHz+Y1UbXOC
jtw4n5ZEYYOuK+s72g+W8S3mQj3xUlYW8/EbSfzHLjfpETrx1QmUiONIMlKmRmth
1cdM74hS6sVGjM433uPbCb1UmKPp4sCIATuVFHobdrUZus1G4eOqpldEyzBH26TF
rahu3D8exaQYTvraIFED7rBHPMFDeZTB2cCF0taHIuXW3ILE3k+DQk96m6yy+FZ8
uEJuX2/ye2mH760l3Jgfz9EYH3F7Dj8849+cpfzF5bcH/3ZwS7+QIx++gMI+65RZ
l8E2/q5PuG5wVvY0e5Kur9mB58OS9BnPyWY5+w/u+hCOL6Fz060aqjYw040YlVCF
0DIbKh/IUx9VTJxjXIZy2fivsjKrCQCU74rbSRpYe5zENwEAVLuW96f5ZJnHhoyo
95GepSbmuCAv2/+9zBWR2PoEDMv5BkxAwfHJCo0wrpolOMzDZaFoefFWJyH3+N8P
uMj3NK8qfIyGOIGopCPyvN4qMqACucYu+kZkIsRsKtlz3JIoXGTm65TzWDw/GqGb
3GXUCX/Lfv2CkUEWqQkD+w48rv4PQcxyWAVjuRGuUCe94BNP93fDLDMQ+zf6GOr3
AtTDvmr6NS+YMSiMEp9Fr2z7ULr+VR0OBDKzj8opy/KCqX3v+g2ZZW5KkdrcidXJ
AHN+k1vvuKNkXeGe/PhaypVN4dah87k+Xi5lyOr4/Es5fx93eqSqV0sy2640LX+H
jyf0nZqisG5jgc5lB9wxQfLLySpyYRvkbKgVcW3UOOvVo+RqU/rEeOzG4ogB9G0u
Tm2Wnws49NQayvsJIscnN2y24gql+EZNZPRrd4QxBOal9y6J7ki1sqvTLwBWNtKy
s6rt6jb2pk4BphlCqzyu6kMgYcjUq9zlTsbEzZLTeABpDTM987aq+CAopgFxxaHt
PVL2C60InPVAcKmWJAwMzBQrfoQJ2hubzsxGwBbXbL1UJjY2KLDoeARBtFj/jpEK
zN2s6btu7p9h8zRgo5K75HJ5kl38RDjZKBWzo0UkaamxdQ9pLxASht8C9hv8zyIQ
NUQIHT0QZ85CFOkAnUOsjbr7SK00q3uEIkwjZHClrkVJ7bXr1jm1EFIqxN3p4TkA
oBQUdWYaeX3EWJRpsTB4aHrehDryHpk/SpPzVSq7+aeYCb9NalKskOAVqTv7wEvq
gZqQBnDHCqQ8Y4vVpBa3auL7VtTv+p7/FkavrZr8I/EOFYskNJmKS+wXxcOwMV72
iklL/5IoL/FVrELAsYipTEo87xNqJ9jgwUk+eeSgB8RoLGJ2TIghA1ydmmfkrKfz
sgA5R+4SYj68J3aGgyaPJlfc88wy8ha+s5RNd1BAMEjlJxxA9pkHSdMxi7M5RsKS
OQ+ILYCrcJZ8e5sveNbqj8q3TLDv2TDVb2lbpiKTtrNQlg4YcSHlPqYah78LG079
H5n0hms8EOyEKOycHgnjAUE7Qqutl1iOMVeEjPjfdCtM92sunVNH7Nmd9znUG4jr
TSTN6yJgSC9nWWMLqRXKzrNBB78QIr5D5RARbc2Q0AddRC0uBDMale494ZLnCb3v
wsgnX20+2qtAY2AEbnZ1KBUQOJ+Ac/8KnADAgXRz0PaLgDpcXe3a3fF5fMEpmhhf
CFuYlMxSnE5QlI6PSwlmgIm59K4jUkAjcwN2gi9R7nQaD4EXqXLHPhfpFn9PxLUE
Zst33m4fkdTCzcfW98yWXf5NjOCuenn/F6xEifGV61qcFJCXCTbCM6Xycs3cjL7l
Q63pn1bmoAgeCdCF3Xh6Szpv091XTrwumiPjhkxQ6MfpUc38Fwt/f66Od8NOO9OK
670xjseZl6R1/IFBJZ9yR5Z2vU93rHN3+wbmheYvU45H50EF3dhE+kvWYyLgeT1t
wbQDEBMm1Q+ODASY7jDHlwIS0QQMXvpdKwedgsePtpePwx8bkxIjFX2q7aiRKA1g
2fVzXxLYMUZGFUjJR7LxYefh3feXgqeM1w4MExAnXytlW7gUaLGid35nHH61QTqO
g1FQuNmT/DkE0jcIqFny+riLZuyL9vFQiYNFWlKl91tZZfWrxBiHbTOHYHagBOd5
0rSPgfXvndM3fTTjI6MfBXB4d+QwavKdBZyJsuFOJXommQ/ondPnwl5v/+DOBzcg
J7RYsL8s+zXFzXgzeFcE1TvuFXO2UOiBCMCnsXNGkMUa1a7H3QDNFPPixfk7obQi
MYjMhtNnVU/KQsf3rKg9Tivp4yc5OgoVIAcIS7Ny5IZl5eyxyaqoWMf9RySokYdO
q2tg0U9LHVpLX6oS1WLUTWEQ+Pb1SG8r4P6zNAt4hxLmXB45FTGn5SwyWtVHYfrJ
0AbNcWUgw8pYUEhJtvsSneEaImfsPN9ERwbLrpIf9EPLbD0TuO+OknM2b/rbo1U9
LUYBoXSqHuQmTvHTlFfYcz74/Y2sd3qZJYO21VlZL+GKfupppHtERHXDRHnGDjrP
STkrvmo/JAiWV3ImqDcsoWLsg1ZdmlNsDkDDxYiq4QYH7U25RePHRSiic8Yc6ssg
uSSTyIHy1vdlWfnva1El8/04YKX5TPxFpVe54n03Pl+F9LWFv8DmfZYNasaFC+Vu
oxuagJSgpLPTm1p43MErITyCALU+rz9RJmpmngaGTyzOkOPNgSW+iioRtWeGGq2P
cFsFRL4Dk8wbTlv8l52weh2FabwWO1GLCQ0GL+MjyNr92m4gjel1YUChxPcvZLAo
`protect end_protected