`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
ddtXksX2+yylW5zu6QL2Lhnb2d1sD00763mmSITNX595NcHTEkwn0zB1Dry37fOW
FufOhVzEJp80NC5qZ/+F0Vk7Ik02dIR0elf3clrjeJRK85K4e3Hoo4xn7YbFUIms
l/8VZSb14+JVGURjfswrIyCUotIzlzVYZ6gzoZwDXIi5gQIBf/gI+KxNXPaKV+PQ
Ufys/12rjO6aI/pPlqSm0hCvftmBcnezN2hk1UeXgOIuKZnogjOsf0iJVX2aOOWE
6pD/psybjbnsNB6kH5uFTA5frkzIzkzl5d9+YDm9OyC+k84E83I/7/j+rk4L2dah
QJOvksSIzN867/4Qt8qYTQ==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="MvBXkzurAa5VTw+1JJ70nePUfoQXBvZOku/SMmg4TwQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
oRtzZL4VJ4iwysPsC8SXYCzXS8Fw2gtZTOskLcDV+1B9Nzn1zTyNtlo6lNICRmmK
ZRVu2BmCc2G+fmzynYlNTnSa7C0Cuel6FYpxCBlOuk3OF2tzAmLAuDyOH3Z1Yjzk
a0aHuoCdIRKv7BrZCdALt03JeUmXKPdOmIlkVGFl8yw=
`protect rights_digest_method = "sha256"
`protect end_toolblock="Jn9CQpRhJt4rnzZPRk+dOpzAubz7omckX1MrFd4p81o="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 11040 )
`protect data_block
gD6l00tciPUa6pDNTk/+t0OO0nC/UTtBwLB41d4inuAUA3i/ALrNyoJVcBnAmEQW
ptbcNp5fxEUJjnOxnedyZEuEBxWRieZFQnkRdF269oPW3WNW3i1UjaF8geBNg44x
LYP63kHxhcehWQC0muUN1iHrXrHgBnC7jDJEQOKST1zYv6EZXcfNgzEdaUEdL0+L
C9FMd8dQ5WbEv7YYZPcqmBitTRatIX7mG/0ZQavkv9R3/tAEmFQd7zkWITfB74dJ
Zlcnch918VwPtfbRCGERZwjSsHAEh0PPYk0kL18ckki1NURziVgGMi7rK+sga6mv
dt9qttNWCGbOtJB5AANsvAVGHKBQlocpdJI8WQXGShWbBwhajXCfq4pxJ9diUfS7
sEosJ3K3Gx9HxWtew/QR1tIq0+8ZMnTBgJHgcTNFxtSg55AN6q238CJ/+r/1h1VS
q6G7hgXJkvE85qlCWvrTaLuWTPEZZU7psrKBmnu/3wdOaYZxWZSGa9ZhTDOJvwJj
sJJcPEikSJOTA4sLrbeCJnWq6wv3eK/lzKWgrUIbkrxbp9KPJWxJHUfPId4RZjvi
6egUuwT1UzLn2f0itdPj0LlE5Z4Su6Qx097IsEx/z0IH7aozXFcaQPHGWWiKyWgG
7xBHaj3Vlhf//ytz05DHGiZAiDhosENQwo5fT5MAuVKzXVFwdi7QHaGOtoIncOGy
xGmiAk8AvWKuyKRwJ1Za22w+VqT6yLp/AEPkHocdCnUGiI3oQkzWayy60mDuB6lU
pMVPRssrEjlYG+cBtT6ZFf3Q/KLLsaUvkdC0a02Zr5V//G7iquLtHg1mcju3M0aJ
m2DcK7FvHv37Dw0o05NKliQwvt9mBOH3zPNvuPn5tSz8vBaQcP3GMKUS4wTbz8ck
lYlW32KA2tSRocrjYiPUtoAbR4Wuddk1dTCDsyuUuFtsrdjqgIs36qLj4T+uD9a+
35yY39x7Yhza6k0uMKtMrb3Qe06W51+bbKLtGPMlOxNDNav6IwxWIRnXIPrzU65a
p0WJwjkuYs34Xx24SYnp7G3KuEQBdJXmbGS8N6V50rYubnHZ5aoEX0MqxlXxqu3+
1TQ9zwdYYmsBsl/72n1Rgb2JEY2HAQaLRf016Z94eSRd+EnCK9zFyuU6RkjFQlTK
3E8cjo/aji2wbcNGu2XTTWpgsfmAhkeOlkA7QtQjE8ISeP3WabQPPa6rrAEkafGF
3TgNOxVtC5+W0MWOQOgJ58yA5SBQ7fdyhJEqzNEQIpxklTgChIgNnmjdamPp7zar
8T7taW0bRosDHhFfNaqDr7CsQuAmiUv9bSkqF2gq8xvxRSTotzZx3XWsZuXWhtQ+
qw+VUpDB9N5IptvL6O0EmCu5aWEp2au6QDHBmnjgz6zj072pUrdBxd89kcF1cFq4
j40/lLfQ5AVlYC1bB9U6t1oK0ApUYVRQTa+I9EbAWe2Tb/xTu387mP6mmCEFQA0+
kqVK2aVjyXX17w/1b9it/F48s1PnxawYtgn9ksWW6YP+j2bY497qVrY1gB4ffP8E
NTJPbvaKF8Ux5/5SsI4BYKuEox+cDLUOJuzxW8YNzLgyyKR82+Rf96s3r0FkF7J+
RgTlxi3yuCH53ICJyuegceXg5g0tb2h46/lNVU1/5b5IvU5/q3QDwRw8ZPBul1VR
PR+tbMxJMSq9TyUU2viqxyk011H60FVstsbQ0BDtU3o+sbVj+r89+tvhN5RO9SMQ
ba15pU8QkCwJfSHGCMZ6G1V+u10O7fp+PxDNrNxyg8ik+CJfPIKjqJeB/97MFIhE
QdrcZUeVj72h13TYjdaywqUxUghyPhCeSUTsEFN7sFY11kcpo6I8YmpZfL2WfVwA
AO1ilD8/m3kby97oUP5dSZOUjZkOxncjmMLwT0b+96RWqOx/ojiZEJUoFbbtxx1/
8R1kGDaDnU5xLA7exbI7mGiXhbHQhUzD65RB/27cVoPq6Efra1ALtGWg8FaJwBKx
nIZa8iMn+lixkOtD5XTU63mOkf85rH/Q4syReHnlFQNyuakLpJYY+JSOjHCl1chu
dA3sjSBHnszkKznBKrrKCmodb5LoZFHRRkReExRuAduzi0H1BEsUKNYOJfczQyz6
kru/Z594hCIMBM5eYx8Io3Mq3LHhuBB43R0ZuLOT22CUjwSgfPVydAeQsJ4axWfU
Ckj/vwjTcLT4sGvit4uVA74wcjxqXXV7lEJJv8DpPy57sCq8rlZtVT9c/Nt57ZIO
NbfbZt5jVx/0NnKpB688cPXDdFRgDXQKHhIBJXzu1OoFwvY0zofPnhpuWgkgQECq
H4usmPgkuRk5gl6TA1aO1fqH7BK0p1oupqC2XFhTrMTHQuWpujvYf2uCCVg/yK3y
bmWegwGOliWT493VffF/ZkEkjdzv2yTeBohf51zSt9dk7/heVDyKjYpDAUqdDB7f
41prXt5dR8eF+GPWQFgBm0XQoGFf+sgJo5gHVdeqerG0JR7e9C54I1D4QkpL1gHI
32dw9K1BwdRqDCHTbW3qjNf07q4uTLVqYZfucPgyWNEO1zYc6qAfQniKbKOD07hM
ckt+JIRTVFNyuX57sMo3gLOL3QTDOmNVh5xEmafFGAXDjGrvUfIMDX+54T/Y42XD
vNn51QakL1VrbYTlJ4ItZcl3m3SP2z/GKIwFoEkEsYFJpF8cBA8JRWsU7L9cUUVt
SVdESYJHr4UgW5Qa9LXr5FuEmpW3g6oI+dKakFZel1d37jdRVaqF8eqOXV2gd8XH
Cr/YhQygCR5nUNybfjwzAvf2gBsybj5CilnEr+o7/48Z2RRF4U4NVcEqdlcZmEMU
4ocaPvLWTScpbMuDArdLGbjjDcCeT6oLKAjvAWCGMhYKMsKnhGWH6puf9ghOkXIt
8oFE7ipRyf36Mt9Z8Qnete9yxl1rI4NL525hT8BFF7FJFpZ7/U0WKwLmkq0YEpun
J2YAWRj+s2GL7ia5aX4yTo/j+dv8VbCj9uBpUG1oC44CqUh7qduJ7UG0Afgyf2tz
O2MBIyIXJjqyl9rYwm10n4yQA2bYW8nvM6Do9RBSzrmLAYbeJ+wsoNFUpi1AZPJp
mGD5pNyoSy3+lMifXJsEopZnXQo67FFoUn8r14zOkajaqkI7il0akiMj+HhzwvKT
mwLEdeRVNDnr3IYjDclQVEcfoeu9YSUzgoEF71nhCubDEaQqNmzOisMiYc1tJDUt
h8PnSK/tl/blRsLVfBe1UYlQTEzjgkFlPuTBhxR55q5YvefKD5CQ4zhrd4iJEsO7
oQCwka3SKadyOPGe/tlN/wf81oytNKJZiXM9hyIOq0WDjczNa7Ft7Foz+znHtpsm
ofSUThrAqKfUezHK8F1bu5MnVTkm9Oi5Yp6or29zNGTO+6+68eqckLXtVgrcCudb
+PrTsy7rcF9pBypHcDHDyfc+g57qZQ2u4LYz9FmVrHuQTaPVREEEt3AK4BdU53Ld
Vik/LztDJOdZhnMjeaLmBU7uBXw1XuEvIQV69gM77K1ixz8bF0FZpmsXKlyqZuo0
MHrG5RiwxqhB/x5dcUlryOtftjs/ifR02RmbkQiODSfpuU/gbcfPbdEsOxeSSIsE
afvW8a2BC1AS/hzfCTNfVbvX0QNclxg2rBwE3XsSWqZWuUv3ehHatImTdABjuRHN
9HiteLYFTm0CiL01cbN+mwmwOshs8lRw19AkwrTM7l0fIgf5ATCGaQVSWJQAMHAa
eAd2iVHigR1rP42zRexwM2x91W4OkPl3IAV24v6wcDfq5DbFETezP7rbPRI2tJH+
oolTd88QC4PGkPtT5kqsZhFxQeIMPZcBodf2o5Sho3ZSwNXX1hr4sFwbhGk4bFan
ah6lWIfbLv0Gtw+zCv7LXFmJczY0zfivaOVfKWR18MNKSF5kzzyr60XzSJSx7fXK
b/tscNqu6ORCIpzcAKkyD7FmSyE9eZvAlcXWsBJMqByRRQ1Io9lnaKjcPskVbcrZ
tWvuURDqkh9V9Xt8YqKEvoNBXfDiTDJZO8DFxWT24WcoeLw0AnvieOL5Y+kgEC2F
NQLfnwMT+OrCsj0nEqDFdunua+khcVEIZYy2DPR/AJ29mk2l4arLt7r6LIG61yJc
Q8a6vasuQZHum3S9AXCN1Bnd3xJmPgyszXI8qaiJUtnhKPoIqSn/nekBAygxePGA
mAYdH2K9GDogR/D69FFxq0lQpMxbzcTcN9lsWNX0lLbK9TQ9/XYoJaN1Y42z8tCq
7CuOCUxHSTYPtpBQfTWwiTukaEwnHnFjWGwhLzNZakj+jUERHG0HhQgkw+di4L4m
Tl+rj5Yzxb8nV+giull7EJy41fH9ErxyHKBrzdR42UJtigv7CrCjJs1769kgJO8Q
3fg9SWinNqGDkEzOxQIX1KhCxKgBpHigP9NuC+vg+NgRydUiTT4qJ/AlU9Y+5Cp8
sClOirBiteT7PsrWootQ0Mz13Lxo1+tikM8JfboGzVEwvuufuLtUDJPMQDuwhSMl
T1lTj57Gw3MY+9aa+Pzx6C6rdTi20ih72BZvem/eF0dSRHbKhffYSCylxyscOueM
te1eAyoVnOZMfS9ofKTZxSq4HaqkoILQqKJNcKqAc3q93EojG3qDin6hru+vjUcV
fFl9f5nVJLcoMWFbJBCci/2eWyAVdLskW96L4xa1vYJRlhnr6FCdaX1qZGm+C5Y0
arMqt7MTiZn/l0UIbApRbh7iT06o61xXRSKYnG5/c8eLvrIomo8IsFw4pDU++frY
hKGOMcVPja+JG5Fz4FiZbDjspe6WJpn9ETzPQhzddLk3ltFX6Q7/XsL6/0ESrDsK
OS4TPYNE4lcnJ70vsLdTZm4ktpcd4auRJ0LANxDHqoShiNedooe9x/fkYY1m5RP5
m4mI5BxiGD2hDsFbcTA1jbrQG1RusOIslDukLECew+RrpBXXNWj7FIhllFQJ05F9
vmDEYPohRasYxYDHt9TxiDnOK9pUlrwXV23grZO7iGPXPE6z51QTiM1CalvnMHxC
IoyVHDH9koHxxfDJWbzPutgp0wsQl8m18lM2ynOVbeE+jULB9RvYFsh5voG11yur
1ehAbuQP/LkxzC85+ahrRN21IhZpJu/gZ9zL6e6Y10lAIiibn3sK7hPDyg5nCa9X
UhXGZpmViRhwQfqSoMd7Ogs7JyAZcdULpBVKVnqvylawpRE2Q3xM9+3LpBwNc5dh
lNfQNrO4uFBGy8JcQVFNhki/0Q/ScZ9HbtBWtuGIdmcT5uOi+cRGxeD3GTzlDRKI
9dAKuM1wsN8A7bSUIiYZTAKk+e86tq+MadsYkIs00XT4E77HePhLN0HZ2fb2Guya
Xcx7vznH9/GIY07pXaFzR8uB0bGgTFHlmsQzBKDJqibt29h597XS8eItmKQs6by0
t8pOSkbsfk3weTQBm9XOXBMA6YW7+VlkBXSYCiimPG+lF7gPnMXef94oxFxtQOhe
peLjLiRqZr0IDqv2IXcvPy1L13ax40d8rZlN+NWBRTdKtAIq9JvONUbLkYtlLf9Z
7Fe4cOP9n514ti62vxdWr2q3lzYfwg5z1kc+H5Xkke/IwsRaW/wQnYQ2s8WRdYD2
Vd3nOu5o2KyBdW7ZheUNH6JI3PmR/FfEC1UkUChGgaRbQXM+6Jgt1no+mrkXFW9W
P49UXmh1ZjDy0fSKoKiOsI28CWbxvoFL4zPgmwEUQQ4sM+DdlbP9jWGkhaaibwVC
b1P2CscshN0oXoKxCOo754hnTQhgCE3uYyR254tM8bluyeelD3ifs7Wcj9mteDL2
Y3qumVQhQXZmj8j8fVYgsTNcVMv+oiNvxQ3ssUbEa6jJAIhoKamCtK4exTQQb9tT
VXc5boqITnbxg1pzSugFiT5afUwUujBaf1Yqs0JUUxyAKHfHzZCK8n56cId8p/cq
PYtMQgcU7IVumxUF6qaNg4d+KkHCFGAWn+/B8MqOajVKFtYARgfjoe605GRCOpPO
jNNxKc5VaDX2yJBz0h8uUufzazlpnxUGsOacHJP2lKJcdxL77TzaNZMMEElRyWbJ
ya3LBhhkZymFYk8M4gtWE2rEFlrf5SPFhnmTvqF44iRgp8CDadTLc/LWSNrFLxXj
EnQkODRZ7vzrMAXhhaNil0ZLEdpMYiOpDejMZqtMKsQkNTTm0gsf6DAMx/rlhLiS
GuWM5varrM3jH3VlaAviZWPQJbfDtlnmfDHYkMQTHuPPjrAShQrDfbpfVPurjyld
MtkJrdcaAOjBUxjNhI0M01P/U78qeZ/wIMPOhT6T95lieJNIMHWNBycspARQtGZm
tdPGcTOxSl+JjcpeRBOnnxcTt6Q/gO5io58rwR9HdmUrU1WknzLRnGeEOdwLe9cZ
tMZ2ttiODkIAYzWTPqz8asO3GMbqLmPV5/bJPlTJuUXqbzRrlt7M0vSXQ5eh7OhX
lWO17S46gD1OXR/8iT0v8BDzOKfZTllRTt+nbfPHHqfKo6IzR6dCJH9y1AH7zk4v
CoaL9EFNrDMxdNbhw3XEkd/FXn7nIXbkbs4rBPLh+nRNMCeElqAqNA0PmGZ6s9k/
J2waz952A3pVZKbIk56+2iMhqk0jEUUCFD1fND4VzZ41/IEwdG+FoJeXxIcWA+lr
9dNWLScYwSgHMVzm811qnxOwLD0mIroPDG3AwPjK5L2QUO2NL0eCN3BGz6d+PJnm
S/baMyHCWVa1lwGvvlK0XPDxvHakZ0/g4F5hwmpF+iPx+nFb+MA/G7qlk/tKKIpd
zH8XCsazcnm6S91Bjd23ZzdT6fz5mXObo/CeKnQ6kVeOuuQg6Ba2VjU4q/P1W96H
o9jiEPIUqXXqZmfaO3+bwhNIvE51FyZ0/Kl/ir50zsv0kIAH2oVCQtitTnSZXM6s
RJUEwGXNSu1B/Kt7LI6DrtlvsOXwC1IWXw9bUyFrAx2ZXB04MVuDqTaSoq4rLjEm
g0/psusZJajU/qAhcll3Ryqi3EqGF5irTxu9zNyeTCxJCf5Q9JsggLtRvNqvqZuT
Xfh+VoGo6EX/3gx93U4L6MPs74dFsKPJSd8CHZTSpwex+fuSwF8jqCiHTFvcuyzJ
lZWzZlEWkKUH5eWKFRSI9pclHxMAhekcvTJm6B+7kDHRTC26eJSDjHmZs+MumH0V
agiMHZ5eB0VxPoRsOD1kjXQrbUaWad38fEpq6YLCnqFHbpjSwVA4tVNMtAiwbWhA
U06oNECcQ1+1EmEVl10GgCKIaCEjtHjoqznCdqF/+zdcq0w5gRJvaABY7wHcc9WC
aOHwt0DKtrxX5qfVHXh7y+ogDsvQ7WYVw+5uOcr8F4b+GbbMPQVcCmGNjpKAvHbQ
2s1qagcf5+vMtbCzRJXdJeVz2EjYhAoLPE6aCF9ymeuJsZ0NQxqyEYOkVF1n33sr
cABIsQxQF6LEN9+y0lS9qfZnAC0hFG3somHshoe9qOjajzrJBPVWFgSJ416Ybe+w
2poTRhz9wtliJslauHHkYZHP3lfJ+DwQVR8wSx/OT0ngfQduSGXxL7LxIj11AGJC
1cQZGk+9My8YcyDHu6Q1IDwVEI1lf4GH73Qne4hznydH4dSfC6l1dcVldk7kGw9z
j/QhveSzSI8EsjjjF4ZFcz65A3bQqOu/cosQQmgpE0ZBbzwCT1HYMlIxZC5ApBCU
kF4bHksBKOsdRH3fTxKq//Q0iUtWdQLww4euJxwR19XaAP2gbs8lMX9TOd3cdUWA
3r0Be6suGfIR7ddL1Mk5JPF6NAjMzebWGCKM9/VK6BedpVDmPU1uJITLq41RRiXm
ukfEqI7TFOlNulZj3XPrehqg4oiFWkmC/uA6XkOVFbWQzofHWquU5wNbJZuy3JYJ
wXpaSWnDiMF8pWSqhywgk1rnTtSyITzQ9XYsN+s4gZNLagCQOhWD82osf7R5b/tA
Cz/oRClPhv/qPYJYfxL9Mxt0KZzs/3VEQEuB4BAcmQWimspFnsRyCYncsv1a1Ntn
1fQl5InZAILZ+B9nsTCEDWywzyFebRhyW9+eopY0I+uDVSOqF79pCM1tEjyE4QlZ
of6BXCVz62/ziOnR1o7PFeR5CrpPSn6lY+lliyJzwEXTAYT3fhYuaaJFGqiJgEla
RE1PMuYFQxf73G0DhZPhc+qnXcKEoe/QInwQwmjhv2ZtgR35um2dFtEbxzGVhDqS
8kghzAfQa0isEOKthq+4Yo64yqyPiUMxw3++r01nfh8Iqz4Y7wWdhfQJBik6P5FC
bXI4rWB2GnFDIUbGhd7j9exFhv7cfPChA4goATFyBQ57l7buWvI+hJ7RAfCuSjih
FzfkOcTNK0+1QPUDpJe9lnsY29Ml5kWKbr5bAMRbk0bb9AxmJcKftOYqYyxAHciQ
Dw0lGl4ihEMfZcg1mE7uYsJysGQQFgsCCoxPWE+RLmDsTF3aM3FtNwAI6Ewu1tBF
YwLYQ1Xyr+Zr/BQ4Klq5bbqRF0fUnxdjS+UdXtwk9DOv6QoCv4yh2c2vQYyZJWy6
dVpziP8GsNeKz23xvDqJBIiQQeNRDCsnA8hXZGCCY61A+t4faQOX3+oxJYxQ2gkJ
jeRzgqCkrhc4C07eVcC/Oo0LNBV5QFCqqHESDN0MqRj7uiVBExTeDI5mi4BbNEKB
DxODaA9TOX0fajjdGk6LGNozSNS12iiHcKdsJJ7D6iNYOqyFn3RoL83c0tcahKf4
S1o2q3DOtphQmGw8kmj+XHd5k+cpEpzYitI2t/pcS6Xx/8I/AJjuEtr80na17xGk
K/B5LgJ6XtVsWS9ZzIbGJ0KduhlMIeS5VJoLoLDnFPmL4BBFt79A3L6K9NSXg6Tw
sUjMoxzTGd6dtPysVPQfNFzUYTxMXgaUAhqzgTeTElsEjD+0ZdzmrjzI05KcpnGI
jSn5g2AMGCkPEm7ItctJzxmrCSMTPFNboCAm1IH/ZgiQMJwu+ZxryIc5c/sGo6MP
LAvc6PPB+GhkI/QLnakvIFDh9VXSzIvQ1jdJjC8IpIYAvx7HWSieS9neNQG8JW5L
5iMeQwl2LH3D2UHkWGTOXSD8MEvj7FCqqmnes04Bg8vEqGiXe7H8UuO2H37srMWG
c8ZAti03HJSejsZlRIVXDBy/3PI9f7AHsqS8ighqpw14cgTHkAtyoUitGEgPawpf
+EDu023SYYJ8rNIGoQrgcuD1xikOjSTdEMbWhxdAKHW0BgS293Xyi/xIpsenyyjS
xi65konqfXdL9VPifhV2YNw5XKhvlqKWq+Nk+A/Am2lbP277Vc3QNxiociKLw7A2
B2V2MtRJwAUnr0Am2ekS50CAYp6bZy2+b/qheWnuTSA+eleh5Blkp6PYxoAhj6Az
t3ApijzTtr39KWL9EplQhWoa/2CWonQgOe3ECool/GFDvdbYAzpoioqkVjYM34En
jiZu76DN3QUoxdGQN8ev60eajibctmcoQSGn4D3Ib7Lc78oUXdawdgr6yvYUIetQ
WYhponp8N/HEFUMTkvp2WMVuIGHH2GuzvO5zlUFf0uGfEbC83OcqabvYLwk/JrKj
2NhloKt0oRIt8DeITYrEIOftBXns2OXuyyXsbm6wEtJtwdLP7Is7sGo93av3K0/d
gr+eeOAF2NX3vEtKHQW7uZDe5aimqGxliM1ico7C/0KBjxZn3zYBtGm/lSb4mOwh
FyVD2wGPw/GvyI6ng8y7aG7nFZ18H6Y6Qlc9Qpa7Vl3iQE9LFzqFNc/qdoR9fSer
iBpXK4iZuiLDvgCfR3OBSXiQInjgwB2JKe4drN/wwRLP7xoSqH9C8TzvaH/RdIGc
4Yv1oeGb3qr/h5LxioWg5139lGioWVo9NpK73afjXDP30JYxvwJaQJBans+yw/BW
D7Jzw5178ikaGIRILjWqaQeIHreqwBUfnMYOTkIm88lJM/9M2P7G4cC3bVZdaZMp
ytX+H/YHShQMhyOIQIOAY5rkNuMXPNb2PZPczVOEbDh0fm0HRlAfErCEGvK1379C
RzOF+vJLjRZLgQzZKWEjsgm41hyrTgynuhe+NxdXAlzmFEntMw/Mrwmev1D5l5Js
/eYSTWo2Ps/blV7Zf70fcO0VicjjUbqqIAbf9GTQ93vN7DPLfNtRFc0h/oq+uNo7
VC1mClUcSHtzoXFW3KKTne08n7BvIC63WNziNocqiFHy5R00d3Ra/vBdqQOJFkFp
Vtg4m0uIPb+zLY/hkObuPzdFqaHkzbmNcgfjecl9quW7iwVIDzXYoSyLdmU0bHe0
1eb0kL5sFa4V6dlVotCzmTtewzIA/vbwmnWGvWlqlqxufl4sjbwyZ1nPvSO6xMG6
mqHonMRFD4LisdyEKM59//IG0/McvdnKsVcsZhoUdvyTMMY7uP1n7sTZAhNnRLJA
vOHcZRSu20RD1rH+/+Db4m8y/GcCGhn4qAeZzIvyNHtlRrKMjenFXWae1F1AitIb
oUsb54w2MQBfDT0txuE3vx0dRkuy8H6ess0s/8LTDnT5rchrLvgdNnxuN6Qp34n7
e8QSO+qgMjdFK8NYAYzlzYjaFA65FV28bj/hHqIO1dpg1WKvfvHWdG1JQ9HtCjtL
HP3dhXnOAz/ylyOQyey+7oalvT0/s8Z1J56icq940bVjkxW5PsVn0ixFo7+O/OZL
oYh7I3rpaVIOalvgDxWX0F09/fQdXsrlZ1QZ9UlRPHADJ6CYJxqC7jgSxrQqyD/P
RqtnBa0Ak47m2g9TgEx3eJV7TveqjEKEk7r5ZK292xC7+FTDqxLGZYQ6UUS7uwTT
jwSEJHg4iLWA0pNcaIoX3wZ82IlM1bWl/DFhSZaeEzBGPWkfSnXpB8+8BRFNKVFG
DLSXtNVx3ZJ6A4z9oi8bvPE3Lik1H+a+myclMrF9R36GJPQ0tkSm/OIkBOSEQnXr
XST8wtO4cZ/ppDE+AcFkrx1S5feVntxUyYF9zI6Nf1ztKFfT2tICqOP8Q1EtZSRA
e5og+eORf5dwXFxSmP1pKf4ybdzeE6feNF6PCX3QuHkKBFyRigMgudFXZXppdu9n
o/LBfAKGcwAKhxuotifB1XoQ1jQRxx8T9IRZ8bu8pLitf/bCx4u0axPXQeAiTlDO
ROn3e6gbI+C6D9Qo0tRlc9vHdTmWSrf6zUicc2YDyXxk8pzKYqPby6xYoOJyLR3a
ssiuCBbF8w43jOc2i8ryVlsN6q8AeqzspMia1mwh3hJlOscOscAkhk8ujL5QdEeG
MMMxDumAY13LwSbsIPLAXD/FNkNqphrjRpLngNuHWdSyCd+rmCKgH4DMx2v1aZMc
R1HWAE5D3a1hrjsh66RjljGYvqufxMdhKSiamwm48xcGTDj+3LnyZzzaIC6uO4Lb
3FVoV28hGuVHpBmOYdChWRlyNA63VMIGm0rTBH4J2do+TdGPg509NF0CRoxkeeIv
6GZoolYTSSP9kO3dzByTWOwzD3gM5n74734s8Fi3vIOe5q0bmrGMEeyEuFNaibgw
RE1RKFOIJWOKRIyIiiF6w0yMiK0rsIR9WFLzrn3fjqqh18gqZcoK3AkG7dYXM9uF
+z9TqC+cOfXFNnGE1hZhbz7xWwU4K3dzDrQ4IOsup0rwXv3dw1PJvymMOxBZ3W2c
a439VPyg1JSHsdl5RQYY02dvvjPSdUueH1bv7Mycqv0EVMjEUzBEkHgrtuhXyL8a
9h7tvryPgKVtXa2M4ZUEId1GzvZshc/GbB8/q1e4e4N/MA3K9Z/DuSNImug9HG7h
bfxAzKAOlR+qj6ldV+E3tNBE5hUo7o9FpcM6UqCNz/cBdS7CZvmF5QLB7YYdgd8y
HtaY54w0ZpFr0Y3rD5zY3IgkV0nNMVdq7zJVc3Y8w4YAOMkM/VSvenkCttmzdAHY
D+Vc0RxB1nNH8rv9ETU9Sy9Mj+qZB6ttdqO4cdaOf26+d3w2w3cZY1Sgx7anaaWW
DHLxNPt+REqY/AGGl/VpUIoA1eh9sIgI+bvayYSLYVrsPZP1j0kEfIsl4rR5THLw
Sjog/Kn6wLY9J+0t/WhQzUbg4Mbx6b4//+XDVS24dxXRa4vFS5pnEVhgqltMTiMT
fSHj/AW3pjPFjb0XGyRwQLnSAJ3ReKaFE36Tl4yPtAHu/6604yEb/bVDJwi/ieKc
i4mUoo6Bb/taFghBHzXAW5uAoNIKaCNR0j/jB1ociXZXaSsG4NHcDhBWM+7cgA9M
vw0NZkNBhJgKmMa8kjZW8kCnLWy6XThlCmHhYTVelizj36EZ7ZSEZqFracVsCLK1
oue0x6/Hy5QHenM0OepioxGYVQUoPGx2hpkY1hMq2/3rm+tS43ZielEFI+k9Moes
wG9/ukSFttOMkzCaGaR/KpwZmAojpy76iMZNrRBXvsIrdEsrMouxwz0o+x9b0Ggz
nbgD+5775GMyE8BKg8VlVtkePE0C7n5+m+HTS6XWb91JphYlY0loHCck8owtqQT6
ZgRVZm4SI9ey4NCk8k8H9TTlTLiyAnA2zCdQbuXMERuald9Kuz3G6ZcJbYkqpfGc
h4HvVdTO4QlbLldRK7+kwrT88yabD4GAhHr3QfFY4e3GR/TJxHzM8vXAWTLRLHgy
fKa8Q/JylHP1WMLwJWn2jMe05sZMLnUdei09uhAh9w8CoBv5qhOFH/jO5FUYY8B6
LMTsgPyckWaVDMRi+UVbW6XW1rb0LGWMoqsN5ufZsaUK5aZT+rhXgySNVF2r4/2J
pzSO0T+R4Zn/4DNNvVfUDOKkAegKZHmhOSW98aU7xFC7ZDa6BYHNaLGfYwKFL+tg
gK5N8d+BTHGk3UvzTgsT4ndofCVM0sNgaYb7KFygA7tk2i1ZOsAPgyRmZZgrTEzG
PGQrYZR/by0/P2i7MU61Yy5Cqqk32VsWwvgMi1J0YZPKKfK/FIsRwo5vDyYMfx9j
K/QwT8yRTtCnodATM1KiKKFNR9OYUduN1oypDhNjviz7+nFnmJeQ+7jBATjwl0BH
RY0BLyajxKXhngClI3H8gRhvmaPXWf8XHDIRo1NRjxckdwyJGc2MbPWBz7NcSePX
2ZvNgfoGZIDoQr3Jw6OhIZQqiPD9GUxjo8rymeyAfEiX3NiMfAcwbIsTuQ4u7vKy
yf+LuFnGIdZnxeOxnBuEgLFZQZFnLZBrfCDE6MhvwSZVVlBgBIvQJOAxW2C/XOX5
buK62it2+8lvNUVxuK0q8BNYFrdTU2jJKiFcg4powZZcb/SmobpurHfxySQ5Kd+r
jmtRr5KZ8pJ3uVli7NG2rZC+MJVzGfjs1jRG6j90/5WMQCMqlmgZyy/nwxyexWT0
lpE8CNY9jXpXG/1mMd64Fgy19rCUDxRURCM1Ys3B9Uk40cW3qXLj75Pxr0smlMfI
WY06ltRVmSzMTO69YPb+j5wdvFKB0Yi2We9gwNlfqkw4VNasqnp6VNNJ16SrG9Kd
gGZ7wZ1OzPx9+S0I4uFA+P0PKcIX18arS6SrtDBCloQ3zEexKQ19ZrOc2uNnSX9d
AKmvJTWcYt6zx5nWhZsonUQpYmTI+Y8X+KHim0S/nR8sslDBDp+nv48BfselNtqM
9c6qmDN5fnKbU/LAMU8/wHWh0TiWsRmINJUmUyXKHn2KQpro3VWv+OXBlXkwfrrP
549YFJdJZM2LNsRlGaIN/h1ur2ASZJZ2e93/zJVX6LXGVungDOYmJJxCMBUIAt0v
tRD6tGPR1nSTAizZiW0xN9mPoZcvrmXmjiySwkOta1zq3YiQM8/U6oFJjhAars5W
5DXonJACkWOikufME4oE6IxsDcI5DO7y/VoH9BAa1MgnKCSTdcV7bP7xXIpoOuYZ
vCHFINg4z9Wfwdf1wvCM9hDfLf831lf+pzBlbO740JSSpWxP+FOYnCL0ggOJt/6D
rpiSKeRsodP8zziN7hvdY8Of+2kVWMgL6mepkcEWBDM4ijA1PeS3gBHhoGFmbAGA
uw/49pTGmZ00vzRpcljlb3BUHpo0sePONOl1lO+5oOasrq9gq19tiVCtAAfh2oQh
MwImyVx8I8lhKbEdW3a7pBQW679vkqVyjs8bsh/yt03UclFXa1NAPVpqy0Tgfhxj
3HMh8OeBaVEZvx/AA8RlqfbYupFsmq3TEAIZwuW2ae+GEtGywyRu1Twt/cYSU63R
xufHYT0W0/BG1PDAOtsVY6H7sgg5rE+ldp8jfy9YHOlBzWDLo2VT6pKP66FUExPK
QA78AhxyR3qFHjeFj7iFYj94Z7Artodqk0OI1sHHmRmSYa1QRrIH/pGGeVAfFe09
UO6RfRouWMoTkMgNi7tlD4ep3VB6VvP5WyVSB8skAD7fvGGkrZavsz91/Sp6DCSH
Ytg8DgupnsPYx49VQECjAeKSIA3X1XdvcP7r2NKTC0dAoKlKi2K3Mt7yaQkGSe68
ZFWoTfrPVdIj2+3alt9Dyr1ex4xOS4ENYQ+8jNrYEFP6IveRMczG33HVQnPXUJI8
dj2LwiqSkNWbJ8SNUa0M+lrFrhZH7F26+RAO+Kc7qx1FIQxrJs2tzq32Cm7NMSvi
4J/QSu1QNgrZ07cY2kllZFnyyT3yAMy7gSf1ijAz5l8uzrZBRoakWe7vHfyHXH22
/c+URwH4DfoRX3lLDmdVcDP35upPfjjSM5xRH7KpoVFv1z6I59W5jZCxi1VyfJ5y
I+fUCDyx28wt6srL3xtyCLHKZ7hgP0ysaUPwnTXWC3BvFzvimPOeUtQ/v0C79scq
EdRkExvPabQiXnxCa7BL1mJBxFoCV4yqsBWW3bCwxwMljZ3j+iIf3verPi086cAT
hFkxwoAN6YCjfRp256mjgwoi1QOlBgYEh4YC2H+FDHUE6K2h+Nt+boOSCVBmnZ/I
`protect end_protected