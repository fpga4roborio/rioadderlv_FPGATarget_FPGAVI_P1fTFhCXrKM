`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
ddtXksX2+yylW5zu6QL2Lhnb2d1sD00763mmSITNX595NcHTEkwn0zB1Dry37fOW
FufOhVzEJp80NC5qZ/+F0Vk7Ik02dIR0elf3clrjeJRK85K4e3Hoo4xn7YbFUIms
l/8VZSb14+JVGURjfswrIyCUotIzlzVYZ6gzoZwDXIi5gQIBf/gI+KxNXPaKV+PQ
Ufys/12rjO6aI/pPlqSm0hCvftmBcnezN2hk1UeXgOIuKZnogjOsf0iJVX2aOOWE
6pD/psybjbnsNB6kH5uFTA5frkzIzkzl5d9+YDm9OyC+k84E83I/7/j+rk4L2dah
QJOvksSIzN867/4Qt8qYTQ==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="MvBXkzurAa5VTw+1JJ70nePUfoQXBvZOku/SMmg4TwQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
oRtzZL4VJ4iwysPsC8SXYCzXS8Fw2gtZTOskLcDV+1B9Nzn1zTyNtlo6lNICRmmK
ZRVu2BmCc2G+fmzynYlNTnSa7C0Cuel6FYpxCBlOuk3OF2tzAmLAuDyOH3Z1Yjzk
a0aHuoCdIRKv7BrZCdALt03JeUmXKPdOmIlkVGFl8yw=
`protect rights_digest_method = "sha256"
`protect end_toolblock="Jn9CQpRhJt4rnzZPRk+dOpzAubz7omckX1MrFd4p81o="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 3984 )
`protect data_block
gD6l00tciPUa6pDNTk/+t0OO0nC/UTtBwLB41d4inuAUA3i/ALrNyoJVcBnAmEQW
ptbcNp5fxEUJjnOxnedyZEuEBxWRieZFQnkRdF269oMZnYMEDmaj9qnzq7uePXyd
bGArXafU0vO+1xqksgUtokMkAxhL4flAaAtVDVNuCHnIEzqZycsQVfAZleWrKXfl
wUVZEeZ5N9tbEXN8TaTyaaX5HuCUvc4UV/UbqXRsmcrokxxW76sBry1xKg3tkHhs
+dt6Z6u614+OgXxi9enX/NVGHxZ/fco7qkQFrV77HSr4MwC3dUl3BFIkh8p6FDw7
qmaHblwNfRKZJCmhJyIijE8e2xP+M3a4hiSUcpefO3vl41wLxpawDKcwA8L1MgEG
LTQMn+y0BkyzTreAdAfRjkeZoGdMO1zWsNRJejAWA24A4YwoCK1IkRZOZpasfUa8
eRvhksmZZ87D8JFIdGe8X5JJfQsT7dMrhsfBmJxyO42VBAmH6hndLLTp0NVKxAKH
1xjsB4cp5Dyk0o/NRvBac20dDOGnth+q86kHYcbPKtyeKZMkuaMOUtYg8x/o+wTk
9njtn54akOrBiurO1MKT7HBpa1ZW6ly3ti1R8NoA2s4Og5hnlvreSjVMcLJsiyNy
CVuffHch5z6jhHugLLlwiaA6M4bW3nR8Z7xFeyJ0FnzF5sfjZux8g1fksQ2W0fXe
igZStBlV7tIsSP4ZJjLS1/IakN1T4QNptCLVPTcnGTEmbOsL2VXeC9gNu2nJTf65
iAUVVU1oNWgyhD+q1P9UshOHvMIoMB1XlRBF7ir10RJSkwtmtgaRWvK6/GZMmwnu
EU7CJM1i/WwFZ9sdYVPg9QIjOGxqBRLHXtBeo3uRFpViZNGaI+1qFKi/FPUjCT0z
WazuTsDpheY79NEIJAqc0g2iuhrkwU0AVFFdx82NIGkAdePd/OpZTESO8IvCSk3Y
KEGwYQMbO9aEBGSPjm4+A/d5cr0vDWd73BPvZDTxRIQnTeXQXL4qcR7jbnqb1mFj
bOwLBjFlGHqL19e0+s04Op0YNvCYXquAgnRKgXVGMo4UuldAr8JqeQWKvEUXF8mD
pFbq127vU+FRiFIbd89+S6V9PF0EhhC/BHp40l0DEpDbw6R8opgZ/uaK39yogaAK
K3FPC6N2j7+8u+cL+h6dJ2ChzlIZqWzRf/buvCkEvDKpRIczQkmnwe7eZO7QmpTa
dkFyB9FHc3bnb4U4QwZ0TXKghzwgXRN1WM4LnQySZFTg9nqZujwzZ9ELA7pm0YjJ
Oh1LD+FG9Kn9FAfSQNhrgOY3CkI5CQCbGZDbYzPoLS/WaGm784IwDTdBSygo9Ql9
DOU3DmDOqKDQv2AIM9hc5yRcg5kzhjpQEaX7aBqe3nak7YiqoVYEZcj7wyD8RToy
aUcQQ58fm7JFu3xAkCKBgS7ZfG984RajPjaXMLwdckEcEIsLB6fI+amUGrO6thnh
MEEohyz+JwF+RG/J/f2fE1cmRs3fjW6k2CmeR8W+fg0my2yHOUPxVTS1Vhy8S3FR
JAPF/UYISIT6jWGMv+iiJ0cZjADr5zvMCmjDMHO62OS9D/3EwmxZMbbJbGz7WmDq
EPjZ0DYx2mSkIItvfG7V6x0enh89HpWjhdBm6dN+lOy0f+IqJuaSSLUnhPvTW26S
Y2kDyWtfN8cDcapQe6zweJ7v381X5Gn/4xdGAkkMOu1CyRVwLa885dTw+QwlJLzp
86UXmrGHdlVBmp2zdcUfVGjnYV+E8VLYtzr7VDP/rICeWFoYSXxhoocbTT3SMdYu
hA63r6xRn9O89M1OjtIbcm8BTCP2lDbb1xLD3fTVVT0KWpmFcVNfKaEzjorziVat
syimsdEJzZpwG4pAV5jQDX/V3GJ5MeAPGGeSJMQh2z3YmMR2qNyg9NnTJDsdj0pD
t1LkPoBEforfFcRqtN8UA+0y06W7Bj1pmcG2tyyu7vdoj1RqghKbR3ijlWFgedoh
6AKCT5ueKcOZ4GA6xL6aS8pYB6wNXgQjkrFM5siZ14y9EArMUhvnZFjpteDJAyNY
W4kOMWaXEED+OziE+4yzncMHhXiMmae38WJ/v77Gnmi2nEMOvWI7js19EWp1p8gI
zs12vCgkvTb7gd4D2Kc7naDeGDDf4dxj2AX4fLifU2j8KWYte37vR1gWD1m9J4lw
Y9CcAppOoOyAeZkxVx9jGGZPMg43ELBga0lATX3ruYSnPpl7gfJ2LqAqcG9eAcvw
4BQKLqtoN0h2XdmyWKamhkVsyetPQV9ZMCFHL4+5UNMtL+Jd+ccOCWr+UTOVVQsJ
z5eO0IbD36lbAGZgCMMeJhdUu+fOyMyhaNDUGfxRhvBTAL3R7WZ0wCVR//kjgu/p
bxGHR+l7vyJuuD7UO5WYcQvMKfVVs1HEiGtWjX9eKmj7ZMtjs8lOlXViFMeFsl3I
6XxufKHDII6eLSmZ5kov+9VdbH1Wp8+FZWfflj01XwTM9vRLxfeuZOddi+QYf+Tp
OZy/JOuSms0rkXRFetnNF7n1sC3VFxYBRsuXbG8KDICze8Z1R3G7DQ/fRpIduiV0
Ng6w0hL2u5vkYDpef4MAPxaaXwRE6IlEQxl/X5B+odtCvjUreJGBvqxOicceguqQ
2cMJ0SZQKiF35ynDRcZAKmiDpwgqBeqS9BlvFbokWFiuHcjPuztXdp9guJaUvLXy
T+NlQbMyZQs+etT7fEfesIpSNohi2i4XniRq7UdQ2OjIEB64H80PoaNiMMdlq5zI
jK3MWjV7IEkblzk5NrFXxV9GOf217iVJTYKQjjMyssbw3bvDBLVwUD+ZByDO2PhQ
9pgf70xnse69tR7/tLQH11nvQD6BWJ+5lLMqXQZBnNkv3EwI+zubqSy5fte6LECk
+1d/gcPUgxdHA+CkxuuVpxIZ3YzlntkrsHHk/3kmzqByVeUupt34jt8H/6w5gPtb
Y3IENityfV+fuSVSHW0MrZSFzNQu/wt+24i+G0we//JikJq4x853ymo2GYZ4370n
FGPj8t1UZ8Snu+TkbPDodh3Hz4K3Y3Ul4XfIAhg0VuXMRpJtqni6SUQZFNgwemOD
8qhFAXarq+Y9hkZoNU5RWm/6BWzUAdTbn64mTGXars9xNQe9fz8vrTZNshjbBb5m
4A9hW9soXnjXijm2KlGD7nv8XtapuXWyxjZ4/kWYV5Mi8BepjL6med86D58U2Ze9
OyCfPJ4cNeD+7VKDDcaH8vA5phUXz3ed4mhRq+whHD+0PPdutBTu1SZ0j7O182HA
VyoLupSELrbWUR+CpIM9tPtp7bnP7fDbXeaKheEuxhVbIRiXUwVeqHjagNNY18vZ
HIFD31k9aAHC67BSJqdIOpO4+cCoHVdVsv0HYALQKSWPfNAdX7kQUzHnfQIU5cs+
LP2ui8yoL/7MaEXYwGYSN1IBnWJciWhPK7jlLdHMYN6LC0fv87tYOcYyd4jsNRmM
MX3N63VntPchVTw1pgsYTy95Ab2HOpav2ljbRUKwkjZDsT/xemPOMwBR+PqrwSeQ
CNz+UGEEFy1whl6503Vp4S3GTePAl/5g78P1xTBN26uiuDA/qySfKrUulXhmFh8f
ZkKgeXTSWz2KH/RR3keEGLxpOQ/LRBKOupNH+QMLpygD2T8CnEDUN1iQln0oa1wO
6c6S8eqxveTbqE8CdiFi/t7RNE7UBhiHmMQaSN7m/7UWYT3S2AzZVVaqK+U2JleN
LGic4kfdzPEApfcpjEE6fpjzyRpP09I1EAfptfDHjCckTTOUfO+McVMScPnK4aAl
ejRjXffy11uzh2SsuxP/1JKecHJnNHE5n1Lum7JB3acwgMcjE/gM6+Tyuqf8yCg/
qVnUvJlj7EwY5nShL9jjPPqx7TWs0fNTL0W/760ye6VQBnog5L12GC4k77tgKxz5
hQ2kfd6SMZQOqRvRmNZOgbitn+MRN8Y0sGiLVpytkHCWYY1X0vbazzxO2/mypjiN
nx8bWNHdEv081RXzFhVts0rl1Eo7YsJx1a6QKlvbpBwLtWidTfA4qIXwJyW+Kjg2
f52YBWSBv6UVlZRIQOVp2UVC47Vfmy6t17Z+8C/oUuP/fBpmXwuuNkXOvA8o9ofQ
rRh6Kc8b7+lNIkSy015w5d6i9C1ntwG4b90kWp9eq5UT+/XMV6H2P3gQztso5ZHt
Kze/NpyQCBOjmUNj3P+RCU8pdpxarjC9U+LVTDQ7WLFdgmoVXfUMfQHdH7W1fyz+
B8cZfjNadaEnuXRuEJlpHwnYbqeJj2Zy3jUIhALQxkUxJVVSza4+ff0mwdemqvrw
5cvIiiX9EvC7x9oKKHEpa1ZlrP/v41ROjjJnb3d9/sVA1bkAMw25BGLKYmYvEvsc
tjO5uLu+tqscPMLGwHtokwVHRHJr3p1nn5nj+eU9WQBpPgpIFzzCueg3r8ARNdlf
FQ84SAnXTEvaj6El3mjt2P0A6eHE6Hj1B9yXg+K6CSbbub5Zp9EsXDlEB+9FAEH+
Uw/878XJefarhVBXjRXp4BphBoiv4h6KUw+JgkXZ80Poec2Jw4L2ka67Wd2MQwRu
OvKWAN7mn56KUA+UQvqSwYjvuo+al4LJgcx8x39wU8V9PGKhbybzExNwOWy8EAH8
XKM66lXWbve1azP/kW3zEk9YRiyU7d0LLvG1f3KAxAVX6cCA3/+ITPLUuaBDMC9K
k4mYuVz+DdLh4J5ahhLc4ElrNhH0G7rOJZrxnJ0YHqS/rd2kJH4BGadMY5F+0BUd
soRb6WoCCwMls+8o1pC93T0W1wDshkXLCFV/x+RCQU26vwk6laVJH03mObevFh7A
91qIkQpumrjjoN2IQCXBhI46CXjWx+FfJm0KdKCCIuL8rsfmj98qSlU+GSqSFtOx
ib89WTGit+KKTFyIiix35zu8O1cWoZmppDU4aWq54pGoz99hoBEdsyCwdU3OeA7/
5wW6CnU8RnHe9UBHOYEIITFPZfNDFActYKEhz0USe6vw5zvUDPL6lRux6PsvTaFC
93Z73YgkSf0i5JCUcCn0VNzZE96q5d2vuNuUw3M/dNKob4zgmaiuoTxcr6hTlxsn
MJmKHeGljWY9JIO1Y5NMt2ud2xl5R9Vme+MYMtk2tsHYefiZHq1PkPkVZr/q1FJ4
C/Cn7/+ZCFFlHd2oZwzh6G1WNDbCTIEhBRdMvDjxsLCh5g+oHw1O+Lu4Kn87pd+z
s1QwnoPDkHPXjdEsy9hftoTE+9uJ7JXqaDllpUlmNHR0yjEUTmaITEEt6tjqFbvS
mkqbaGiOcx+xbgoI5An3mR8CX9pObApaA9fjMUxnQt86EIrQrOkA5tnMFM7Bj+sI
`protect end_protected