`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
ddtXksX2+yylW5zu6QL2Lhnb2d1sD00763mmSITNX595NcHTEkwn0zB1Dry37fOW
FufOhVzEJp80NC5qZ/+F0Vk7Ik02dIR0elf3clrjeJRK85K4e3Hoo4xn7YbFUIms
l/8VZSb14+JVGURjfswrIyCUotIzlzVYZ6gzoZwDXIi5gQIBf/gI+KxNXPaKV+PQ
Ufys/12rjO6aI/pPlqSm0hCvftmBcnezN2hk1UeXgOIuKZnogjOsf0iJVX2aOOWE
6pD/psybjbnsNB6kH5uFTA5frkzIzkzl5d9+YDm9OyC+k84E83I/7/j+rk4L2dah
QJOvksSIzN867/4Qt8qYTQ==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="MvBXkzurAa5VTw+1JJ70nePUfoQXBvZOku/SMmg4TwQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
oRtzZL4VJ4iwysPsC8SXYCzXS8Fw2gtZTOskLcDV+1B9Nzn1zTyNtlo6lNICRmmK
ZRVu2BmCc2G+fmzynYlNTnSa7C0Cuel6FYpxCBlOuk3OF2tzAmLAuDyOH3Z1Yjzk
a0aHuoCdIRKv7BrZCdALt03JeUmXKPdOmIlkVGFl8yw=
`protect rights_digest_method = "sha256"
`protect end_toolblock="Jn9CQpRhJt4rnzZPRk+dOpzAubz7omckX1MrFd4p81o="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 12864 )
`protect data_block
gD6l00tciPUa6pDNTk/+t0OO0nC/UTtBwLB41d4inuAUA3i/ALrNyoJVcBnAmEQW
ptbcNp5fxEUJjnOxnedyZEuEBxWRieZFQnkRdF269oN86nmdlAKAigPob0M0M+q1
qDaSQsxI3aTT++joW9bMmOzro/nii9s2iTyLGocI+jKiMzSTIzSZG4EstV6CrqVK
ej0lfapJ7A2LAAXiF5NtYUCbiYmrk4O1AlXGEw97xa4J1xOJ1N5gizcXCDW8y6I3
STp7gkHmi8bocpch8vGerUOkF0FeylQf4HXHmo8+g354T2SrJkzAOOToQlBdvseD
DGmkNB5J/of5RKTKRb50JYrOGVX3Mvguuics5mKdICnTi52q8v4P18vFsP80F3tL
JlBrcoMKD2ri7mfLU5kpxMblPobsgBi+15zYAceeyZXmt+5U86ysbKeZAYmEPgnG
lnBTUGXgKIF2Joq6ZOfutbe6fHhwJ97xTKXSf2FJr+RJbExg0jfYy90SBkhsdgWr
9DwW3jnaHpBU6va9SGPIc2iqYrWSKpMxfG2at5AnHnwpCMfoUvkRt37+sDOLdrTt
pPNdZPKdssgjKk7x69x3hMCDOXe2mWTE0A/z3NDK0FVqvEfpwtOQdJIPnuaVPnAO
TBYuGvKG5Rhv30HuX7uOW8PH/6t4F6WY3Vdg1I2wMvD0l/WYnIeam4bWoNC8TK1N
i1iZCnX2MxTzf1JbA+HUhlArqfHw/Y4DaMlKR4NojIT0QYORtigLDblkEGeAylYB
yR4PoX5X4s34WW93jap3wkWqsIS7qK3gk47uPIhCITHjWZFajHuntm03b7vi1+bQ
TkUS6R7d3j+IUCfT+vrWYvCDIeYcg74j3LMHVGx0+4g/3EYtTMqPDwhzclUORfwY
fV0wUl2PQbPQgRV77+hKWu81TpjZ1uuXsz3dM7kU12Qhz3zb/nj8AiJ2sRD9kbdT
Alg0Tc60SEGAJkNeezwVh2+xyl9u3QeqvhWWUFK6PWUxhYLcjH7XLf7yFfWCXb4w
IJEbFFMcuMFrQSJDUAqVJgD5Pxujaf2lX1/ZCpvdThPVC4t33JqDsr0O9iX310NU
FBim1rN/J1ZC7NfG2aGt+dC5Yn2QCg1ppTSzasxcakPLRrEnqGdutRkmgu/4AdrV
7/8Ctjtw3q+W6dLQzgbkRNXti+f1OP50hmlkx/9eAVzxDq+Oq1WKaUgEdWU/SlDb
pXlvJSkmCOB9PYfQSgFjB/0XzWYIp97mNzUDhX94mngTV7J3GJA2dHpdTxt8PrxL
HIfogQ6hD7F8Xph+89yTMSoFDE1g48PlongTtcEGZdy95S0LEqH8N4+WNCDjVAjC
3UsscXARWjUXGCpY6Te2sk8UUmDkbYU9s6+ACzWFy5nB2NdXub0T4aSG8ZI6i4+Z
2vNmdWIw/zpvp2rSv7/2BEt2ysffFZ8C1oBkYEdfRkKxU5YBF6BuV8+rmBoeK8DO
wGMx1JlzTOqRv9t2akXg6ZMSsE1ds9DD56WOZ7zTqJM64iRTQqLpbZQE/MoRw2tV
d4CMH9fyDFzdCrW92/x5jZ1hbOlshAZiQRJZh+Wvsk/QZ3SJi1G4HHI8v2m7PaMv
/91R7f6ndzzJstnwBElCUydHrN37Q/Lv3LbQoNC0Fk0dkp7Ziy3ND4S0mzk4zLdX
Rknz5O6oa1YqpO5bXND5hA5JQNwfZHuDnNc7kDaBVVyTnLAqGhgX0TAarrn+qeuS
fCgyFS3fkgkD09LB8w+uJwpFsbXShucqPudqhxkDUiOnrIYTqlHU2D46X4yczsoD
Xbpb7d+YQOvMj3HRwAIhUJe7dDal3h78Cgj544+8cgciMVezzky1exzYWDXNkEhP
Y2+WHJhQQCtFV8MBbPqj9Erq26wTYl+y54xOuoAvqOnMaDFIOaSlOaNLTjPIPzMF
TXl7z0PNwNQ+R6BvODrsooFwY7+i+zi4GkGXyQM++A8sDImLk4vUy5veI1Qb+Mwk
ilTh2ziiuxor6ykd5D7VhGo7BAQvG5kxFzNhZtSCJ40msrwVX50n5uNyi3f3hAMW
S9QqUxPeqrVAwNCIoU23uybZ8jJkoS+SjnTn1DB3rm/3SEnAP5CYsGZ1CWT9SawV
QHSvl3G9RHHbKlzDPypxMJt1GtjF24NNCC973qUDS6HtlYTK6l37kdrDrqXjOCFM
6mKYb0Xrz0TPvL5NDWmx8lh8v1tKsfq10Yr4+uqA2DRlmFybuDakXVtvRAqFnMme
aPHoIn9z9XiVihlvZzJL8LOfbWzLEmN0hnrt9JbgJLC+dW1V6/PEBFlBwgMEtUZQ
7lfXms7oU3sTkaWsJU2REAzWGi0iKMh4Sjiqwchda3O444F/GTTQEejesZQbrPRF
mvq1Supz3M742bTtXpQ/kHHeMsDtzc+U2Uccc+kafnd/vAzlBEDLBCfXoLtXl2Zw
lUe12748oVdSdrVEOpt43VUBy1ums+5L1NEBP/3lsaHK+eueHIWPbbSsXhUxra9A
omXFsYbP+DK8iCEST87dRbaKTcNhDdB7gv+Z/ZBj0HUDP6DY5oeec39CKI5a272B
m9L0gHFuJjfT7JlaswDHEfZXaHb58eT89ygTxxJ5HvMYkgvbTuj0Ho0l57rBdJFI
nw6mGCFa+BP+Zo3OClfok6TCiilNOwt2T+dysRLTcA1YBM2qr88q9rH1MaOoQuyv
ug1ryc/UR7dCzIzn+3GjEBQoTLu6yQOO7oMoYVtb451/o7L7nSVRHkxf1zZdVFdm
YSBFt2fXYOBVtCMbeGpx9O1luLuaz46IKaSpTilVI/mS+Ih6ymuiziKkWEjVoxk0
aScPZcNgro0xnqeOWGOIEMnq3dS/+/O/LAU7W4Lsis/9XNhZaAR9Sy/1fMy3JvaY
pjZMfSdpS2lLvhX/yUd1JGpMk16k/KiPbXoTo9KOs5L44ESWZeb8KrSItkf/E0Hv
pyisEUm7qYze60K25cIfQ824VMe85+8gHuvCcv1BPWNSnU55xxO4reX6x3on/Cxk
FHqkovdjtRrrb2TmoBM82rBKrrcBrkpoM5PPzuWdGlWYhp3m81d5IOpBj0eI6IPg
pH5WODuWCw61zeZeDFxbDxMqHm1rzbzB/7XSf/OVT0wuvmpWST6sZoAoBCvHluof
TeczaBvKKbobf9xYbQAYhfy/RiR/WrC4kcC4awPecvqTgAYfJzrC0op6boW2wa56
0cNsJ/1jFo5eJgpTK7tEb0mUDo3D27tZxs77lbewYTPpGSSSjM4DBGuGlnmqfV0f
1MPlV602oR30X08CsSX3+42DYAdM+vy+fBjbman7ibfC5FK6CNUQWZnzV5PpuwzG
NWxqj3UOEHWd5rIzaIj491SlmPNTQwKLmrGrovQtJAk2CnUCv1uzCbrrRiuyyIon
tmRC3vY7wgeah89XMV8ou4FvWh+9tVuyXZv0jbVSiFriICdmf+eWTqz9jR+L7GPB
kUum8NLhxo+MrIbQhju1hJzjSLLWZNjKsBVxuipz5yynymTEsdwdDZkBxHeNpdB1
6KvRbecl0gnXC8YgE6jwgi1NdJFP5juhEduTFGVRlD+EDyyqbh7pJI3G1uLnnwDp
nWb/1LS8Fw70nJwjq8BYgIUmn5SWJKm+ajXW1jfb4S0EySZYuP5hrzUgnKm/maa1
mkARtpBvGNX5YWDc0koSWhQKA7Xk1DW5Djz6BGaSsrhQmMlnzULoboYHB05wdc0E
YDgYW+tityQOH4aLpRosG2XINUjUB0rUIMr836TSfU4wx2iuH6dlkE+Rt8iqlW6D
H+rbBLE+ZMtCYPV7GZmW7l5xshuAK3C3+gX3I7iYXHtGCiWI7dprp6sP+5WXQM+Y
5stWlFWTzOARngvTyXXkNT4Xrde6XJvTDa+mxBUZfzXZpEdZczunvBxO8DasjtpH
m6o3J08AfMNVzBZT7JcpBsPsqe+DQrscQRs9UQlcuGORXwuJDLLpitHBbaDEbgO3
ASo43ZozTQAxW6JbgQMghrP26k8jXpOkjbo5DMv6/83qQs4BP5I/YTWLr9d0KyEW
+F19JhYMKotePrksWCpMWKGtINM6PteGfbnsCDl0uDldwoS2rTvjiHeIxkOcsGwy
oTR+BLH8wu5y6Pg5RHquTf50XssQmSge5ZlTXC/KBstY30POlsHMFdNZBDuA2tl1
8AgZGD8KQJIJtdW954ba0OIMpDlWgc44RS7efcXlTmMp1akJFUmivzMT97VrahbL
EXdxug+D6GFBCXyhSHLcTbFjiGojWsRM7Vfd4ZXn11CntAgQQKgsihZciFdLhn3P
nr8734z3fxSzwHhmdmhD4IfGDktNV6W/si4Hr3hVAwX3awsg2QSYSzMoDnoHW3MX
ZNNuxGx4qgMTDiOVy/GmVGUmK7OeoveYp5v3t486pEuyvyyg/LuIjkfih/OTSZrW
q8tlOSg4dS/C110Vbvs6lq++vCg7szCAnwihKdeHLmv/1uUtiEEeY4IIkg9stz3+
Q0dL9JVb4XHhT0xAGr4etrwWlO93h+ndd6CMdmY4xAcWzww4/TdiptJUKYM1h4SS
s0o5xW4idzi9JGr2l4bmYetIyVpAJEPdJkICA+d5LQqGLQ6DOJo6DU7Fcs7aLYEy
XwFwS0fLTU5NQaySZHXfK5iu9F6B8uQVpX6aOhtSOImTgoYddwXWShM+T00kV/m7
SjdelytMDPPCcyEIMFgkmK19nZapSpny8/WX7OIYrDJZLGkbac+eHNTSjM33boaQ
mIa32/hkRdoB9D6r4h3X+sLJ2rhTStpobGeXq06A6KK2TC3kAtpyadbb5pLd5Xtn
DD+D5P8sBqr/0UXET8dVoKebgxytBb1ZFX6022oEgIj5yhLkPMm+oYdwwZZ2vF8A
3VXVjjbl5Oq2uIqKWCJuCG8BjcBfBkC6Gy2UWdXby8janCqYsWxeTrv+wFehBCXA
wIZ1ah26LWs/x2Fli+1flnEq3dFXwetyu8vjB82bKa8chPeu6j5YSS6PtrLuRMb/
Wh2bYg+Etk1r2zu0YzRtljHj7iCm0RQTQDMSPPtbeGzXi9QozUKM28x/H1Gf9ajD
3HLuScahV77mL54EXKDD06Ron6cpxZF8HlYYhPJWVHwupaDdTsc6wDQ02bRcq8fu
2sq4molfkA9JO9SYx4Zgt9k+VOEWuoAria4iOubt1WMpdYHP8MQidosOGj59NiDw
B+YkLXS/gqg/RRHWkGMOnPvc/TNDqypap9KzmyKHmEaBm2p9O+hsd/gBlcvAMIsO
5DcAgJVCuKWzWhpgMgFpFXC9uoqNtR/ELZrI4/314aemASMrnoD73241LoLwTv7i
GmVQK0d84tcZg36Mn4R+6nHlwF5c1hW7UM3mZ7V3vN+13HCCV3iTeZ/vVF8b/xYx
p3sRJdFHufasInsRJhnMEDsdS9PBqr1T3f7Lf0hGQjJN0v7OqnVyTvClWMQzYlKl
goV8Xf13+lgNjci1yUqfctiNQo0Z8jqc83NzVyevmK857apkkINJp4acXGeeZOgl
1+pGpVT9cyvEBtzc80Cb7Y+BiPyKOJMc4Gf4XxlZeVBO5n6BVVTthX9SkXThC07u
eL3FFoqvtQ3yTIom4+qCHwsIc8lgWy4cobNTbQ8S9gvxH2HmWlPV2mdumAAtgl8P
PPSOoXRukfrUpxPygvlXRGWi3sZTwZ3226AUr5RXHEJsk2wcXhrvI46FFWD00YNK
guTtMj8TTAKRRzarQxo9DsfoRItk7JFNbuzjYOU3QUEqnOJ9zwrLF8/VdqmxxFoR
9PQCbk/s3yQ2nQz4vqdmVSO2cqKGiT8QV0G1RQwI1/ImnL7E8bLQvsEwbvGVSQ3/
kSdsUtf12uZcyYR08FKx94R+ApPo/dBnNoZx1EeyJAMqxz2e+6FpvWHwXdjjWvbG
AZ+MbGfr7erlY2dhI3agfDzPevyn1so9RPlnpDwn5p9u2uDAP7YCVp8/4wcnp9Ah
rWWPXxhba5ZD+GLYphu4AWYhGtInZRkoPmWLYN96FQn7xzdyJYeuJ/ySpvkBvdUJ
5edhxKzuuhJAr3Oq1m4m+c/MOXawgzxJ5qHPjFf7UWe+lzWqssCz+ZPLYaRjBsWu
47IQU7h68HFd2tyXwewjbBhrCBTj0npCFYEFa3ZJQuf9uv3lrr7w7/diXUeDVIPo
eRR6hnwSS2upws/MO+Zh0Ww32LhmBbyQIky5C6m7ew+iRbvSu3BkT+/MWsUK7O8X
HGn9hrUqnka8m0yvvINDPj3PkJ0Bk9xo/qd0mjz7tI0Rfj0d6ysalEfQwY7nAdEi
VLnGmNlUNYysAx3CaKr0w9O+7obaC00/2XFjN1SEtSRgB8hhwXgh6YiGhC1tCnhP
bKKf0scT9N/smivIojhh2lSARSWmAL3lxZNBTYVa3DfPig4V5XGSkHWjTnpSB+rB
aTceBE9dLnlFqvmEH/fQYB3G1JhQTgFaMEOl++j4z4+kf5fks0nx4lKfch9K9kJo
o6007Pa0sb7UjKgbON/WCL8mfqWS39jvhgo6RPBYVMwqOjzfeW6ah6OMM1lgN9yE
FCv7Ma+Nxn1eGDvZOxZNwRunpiuR2QTwt/d3GI60tKCm+kIcq36UTCjiL749uLFu
1NO0++lj4IOYZbWmXEDHCuyxuIl3sgzE2rEQq/EIurLdZUMlbZ8SHGAIGskoAPpn
yA/pB4nL4EIO8Aui6aSRuUUMdOUbYYq46Kntx0Ivj2s+mWtVXsgSDps8OK1+Qlhe
auhPIJHewg6z0J4LpwVDIIpHhmTjtcHm5SPABqzoEck1f7AM+FGdujeBHiEMBkQF
ypmB2zt6m61YKX9hZeakP3DFOfz8OF/lzNaHHXu6fqjhCTdCI4T/AlfzKXlU6HbG
sq0QibOq+d4JTRlxeTFIt2PNF/U1OmmkpIx/3dCAre4ay/iVWjJYgYci7EDqNxyz
ondM8QQWRJkSly5zuzjqns9GDnl1eKLVMicdO21FHv+JSokwrQwOmcteClNOu70E
bXXgBLmc4E69hI9dZQ6oDojhgvO92QNYP/r33KDuzf4XGdu9FZcpP9muQKNDyl/I
tQYUOA4F+bO4eOUQ/+oxPvdrF7jrZcLCd/lmzo4Wspx8rrR3/PSApyoSzc5CD08X
NQYWWJUf8TqxjXxZnHYZZAJCDiYGdZ1b0UbqRqJ8fH88FisYxcRD9iJZe2fxN2Qi
bwxoGooLm0ZEsK8kgUddepQDeQ7Gqan78PAmXPQv82pl/6/Fus3j0oqS5b8dVpwS
oOpK/5eEbSNPAXJZA/l5vrYGYo1xNdi171eoxwSfFee2k6EC5yy+KYJkzVdvtsEp
Dv3BcIXLKbwd2WGIPdssaphVUjdt9WWVaKAqQ+uJS9zxgr+k0SM5IyVXI5Xuoppp
ULWIlKMJ53uMa10igTrSgW7lyXoSGSbTNmcpMl2+tZ6W/4Nim2fTvYmP/IjDlO3I
q/eI9Z/zKYhc6drsH141vlrsdz7EKXKdi4ppl9K4uj2BCVhG/CNGDtmUwhOv8C//
rrAWaguBzoiHYKWIL4TTw7FW9lIa3RCaOZ1rdAsIXeA3Cx/71JK0kiBBFMk8xsVr
B1N+gfjcRD2235aoT88Ue95fQDBdeychqoPu2oTrp0pOrZdi5zA21ASoz2D1fcp3
Y7WDMyExM+86jOLBSAZRLylrIRs3WvXufSbgoI4wJ+oLfpEdisZMxZ7/ZQNTywmT
4IYuCfhRvodnJQr4K4AaQs0bTzHlgxYrUVn33dzWLDLFS1dyEuDxze+AKIayMUPU
oyNrfCF4RaXytxu5RYkikfZjGrjCEyOQ6/pQXTwswiBMNMMrilLNKaFxt0tZ/85D
2Xvs9245fbMmg+KZJfCnYT3Dztc58KTZk/qY9lgA3fcMC4pt00jxLmkpu4V0w8r0
4/UEcU/mOTu0sxjwL5kUg1dtcB/G3bxoI9qNaHyZ4wYcejLS1XcCwXisJYCUOS1o
bQSEneZyD+bqzT1paHoz9cytFi3aBkann3rgQcKf/BBYbpfvOg1TTjKzKTnVf5Cx
+ENLr7N49GCTElYrwOEIx2WtU0UoURbRrB63QDPqdjGbYVhH5A4LNN7QpCKBaUjG
v9lnqPhFM0r4w9KaPHwJiNz11Z9Ik3GLjfPGUllQoYooQpLRtPUznWoawivlonzD
/CUqxCUo6Mt4dnuA8n1f5BmbP9PnKcK83xuYiq28qtg7exauFcvvKm5d2iP3ljXL
SV6jL8P/d2Al8L/qF2QGg2mcNwgpcSFEUBS9ina1AAjdgnGxebeK/uXk/0Uf/YzN
6WUobQuINJItj2DlJrcSuS5fV8FjY+nlENBpXzwBlJozhZrhmf6S1DDm11jPQi7l
Daas5oDamm/VE3+GRAIGdRE649RhqLHxmMtMU3Yt7jArNCkMY4MRNx+JbD6PWjTL
mYPj2lMl6lIrk1aAXX6/wS0KBJWjZEXrXJGY1mYn7r9kM3XloYYJdeomoM04KJ/k
am2SNrZWe0zfPHov4sbi9JIMqRQ04lmOADkrGOJPP7baTJAJUMcsipP5iIime0AR
IbpNi/JpXey9JJ71GfKYnPffe7C0b49VASRbIZHEIJgSoDVe5ClcTnUCGEFhVE9I
l60oMoaSZKRf3DjzQWYin6CTAjxR9EX2qyXPhTl1xMGsnvohmyRxLsNdCZ2rxGGD
krS816FUE7eRETlRUAIqBu94s1hRSeE9EyqKCeJL+OmqpcnlUtnxjJf24E4Rl+71
INwz+KTHYDAEeDXpX751sWaKyihC8BYflD/Mxdgse7s/CuazUZMRBp04tYJXaX04
9hmfW6UlHc7ZGlS9qqFnFqVt6ZHRm7f6E87UOf7/s7VvGUgjbJRow9Pm9MZq84Fr
+2VHtg61DdrbVaE3ptRJFU15iRpSVhiF7ioTTlEhwwRvlkHtBw+A1zkcNCsS/k1x
ShjOZm3tu/si5UMtJX1YH6YhVm4NYpeFuo4I3PoyP0zwtRijk/QUIONwzKbn5kBf
FEcWL5maIbmxnb3p54F0qprb1SW+BrbcT9Uo6A6Pky2jcOnZPx7op5c/Bawa8aZi
VmsXWVi8dEk9bpEjBb5h7AsrCVcVRw25jgifpzJDbOHiQJsAhvG9ochst1nLDD2G
SY+xWuB3uiLH8r8pB7Xrhtq1y4jIg8aCMeJPojwK/EIMJx+L7YH0sCVZ/F9gOqT1
+j9mUY0dtpKBuJ40m/QV4LNgkzUiJftmQtGn2W9jBftKMFRyqij8nUnxGEltoeG3
HifgGDvKzbfkIqOvzUlRgR3yvWSsSlDn6uaSnkmBTTjqgEa11P0aw0PAVZ/zg0WM
mUfdYXfAJGE2Hx/BJKcOR1JWpKhexIq27TCoCqIgtGXOzNI0IUE6jST9nqACY0mW
oEhstt6wuRm5BMSl1TLwvie/mNdtY4qJdlPwHLL2PqeRaUBjHlprxrkRC2kk6MPq
EEixYfHA3+b4mM83pDCiP9G39nWwOQwrFs9NkcAKrBbTLDNBxg0ObO1tYn63rIjq
pDNhEHPH1o2oAjAhN/iVt1Mo8cW77fA7877lk+umYBxQKJCutT5ycISAwTmlVJVh
6NmxoJ4TwQhqsRwU9jM1LB7CHk3g9MO16wXtOnmPq1abucaYJZUfO3XbxE+jusiH
mpIMgyjQbrzFJeRUu5Z55uTwtNH+t9zpXH1VuPMQMqEQkBPmUobHHOglDOSwJKWn
1+nW5Blueen4PlX12dUO1WF/VySy0c4gBZ/lh5W19vYrpeHL2tddEtT5HoBk8VqA
FC9Gbok8aCq+/quX72s390CiNBVlJkvdgyvX3NZr7WEsp8iLY2zuHE4QVEKJ5PlC
MAQrV8IhdvjYFhFaua0qqjF+KqU3To5gXUxZftP3/E0UO+pezjtOlKxgDhXC8ZYt
/Pom9q6UWEk0ksQJT76eyp30Hl4hpmVPoXzV+mpkMlyYeJiywSXozK6Lvt3gr7DQ
YD8mB+kBKEuUJBgqZcIgS+b0wSCk96hH+1bCFhnKfYeXoxY2l0fAtky0tSKGyB91
+AgQttIxYwSSEnZuJSnaj/ifCFDhFUDLT6IlPcZycfEAZHd1bncHTbEiyBF78Ap5
aiAyhhHCXxdCE8j95wbcTUww8XKJZsptr40gn5dG5Wqr2gYkfw/0jydrr9mLqmE4
+HKPNgyRYzf0HqPNbXP6BlCOERatWRkMReJ2YUb8T52boOInoVQ8xNh3xcwLCdwD
v/+MR11k8oYEcX50gXslHfxCVyZJ/RqIUcFtupD3y/rGY+N1a3t7Tjxim6x9eRqI
u+mS4vT13HxZE3GSp4ZSVN8uUJDQ2DlzG/VnROU1P2jJFvf1/f5D9dduPu9R2kU8
6yDRTtNdTunw/szQyH/u5dD66k/B3amVHgwFR6qn1DxFAdeDM5lzkUzrraBPPXWV
y2JkUYNZkfHCw4u/9sjj4yNIqKlHrHO2S3We/b5HR/fZRIeb3hqI5yWdz7MhfUyl
1akrgXJzZsntPNtOv119JTNqPm+9z1ghv36u5Eta96C4K24TBz48aKaL7+41lvHx
vLddDZhrpfdX6w0tMCVAg6XU2CfgSy3hyKcbzWlkVqnEXZt+n/tR8KmVVhryss+F
XTLPxDUORQtmeEUCWbQzzROq7Ridlim10Ksh19iXYqiwUGH5nXnLQkcsOfd8u0lO
+2mzO2ElXWwvK52NuPciizGGTwjoy4EXseUhDuZQBZ6yBXBF7HUgrmL2ds3+buGz
pSd+c2p12I3wZIga2vSpiZtmwianu+QWLW7CY7wt+Yqy5KH00lIcnqCK3NQqpL3L
teL9XNyMWiughI2dmP6DlT8Tj43UBzkvPxVseEG3BYmaSOcw46ymDtMNKGnCYv+b
1mq0OiDG46dBXD/oSiP0GxI1e/A83tv569ZWGrj0U7Z5wEWYX1ksNFqYUHwnl9xh
JyeJvkjsVFsIrxVwvh86yrGkwT35gMni1jjugD8aEZN3cLEg+JCeHqvrxMt1fynE
9t0OfYRnWDHbOrfszhU++WEoMDso18HEPaIxj99brb25XGIkLJgTIjZBEcwxCh1u
ztgBWalBUV+1CqSNF+yKJXtQX5kXpB90P6xJKZi6QWgPt+9q2/y/c08SnSzsl8Gn
VZ9N7wN4XmTfMVYwK91J8Zz3qkYsI9k+kjfte/YCJPUIyFustFdp0s8uV+NOk7TC
fGg/sHs1WMAsldNnstcvsLaOovS+Hy0pPcS2K3Xl+DEu/ubzmUcwUVTDXZQ4Rdv6
6Q+aY2uPfFIAvgPM6dYqLKWQkJrxhb16DZE3QdWsYKNjNtZzrxXtEoucYYM66SQA
DqBm3hzJEc27ojp00pWZAMMgH2d4q+VzA84V9A4bUQpL6d5Y9lTmtS/ub1zDMjoX
jCPOWRXraBC0qL/GfPesRzLfy1Fd6LisTixCnglJEhDJnYXlqPChzJDPhZQ00b+p
Oin8ESK7BpwXpKj0tn4AC2vQtsW9t+h7FMYVf8dfYvKufagXm9is87y1Aojt0baE
LphFA7UL0vYIAAJhwEuja+/mOctw9+TIVOD2DnmdU97ocyde2yg7Nv4zDy8ZJ8gE
4EzWM7JATWHu3ucsXXYq5Lbcj4/zG/nQP0s/RHCmWQZI5mf33LvMrK7OgVif+kSb
T+xcg57b+/ANeziB9K6czf0BnUWFyv0V4O/v7W6f2oBRSoj/GEkMW3eulcv1hBB5
DzwEiFW07Xp1pK7EWTFFKeTgsyPWlbRr2/7pDQlMI3tIlf3ceHMyIchT/sJZl7IQ
e3mVfQHbDoiD3HMzRDp92G2WxZBqnPp4MN1pSXuLIc9tFcJU15mvleMPqRJEeND6
730JEwQBDdsv/0OBWynPQBrK8tSx+ZBzve5bofIa9QU86xVbFdkJwNxmFBTV5fX+
FdPVFm6PGFIzD74pHH8b8sj5+AbVGmsesXFq11wAVjpTV/5Reea2mpjpDQiuzkWG
FJTfHkxiVbKaiNWk2mxHvNMPh5aWkef+Eli7nId1VfuHhIpqrCvt0O2FtVHqB6lZ
HuBjeQdjjFKx2DQpxrvLNsAI3Qph+VCm1CpIn9JOPv+bHP8GKVmsXSEQBFqjQZEj
IJmYXDpo8Tondyp7g6qjeme+D9UbZcl5k2DbKoE1aNe/YXdOnzQ4EsdsosP6T/Qa
kl4B9tMASqOhBYkvdWoEZOfo5JEGLxs1dZxOIfBl3KKXLGE9TxMBwjrWZxWwEs/1
vLBLylqnkLPcVBJAUf2uxfC9jC9Eh7YG8Wjxvm1EMQYEJbfz5feTshR2dTbnbBR6
gxePN4lJTvJR3VlMKV1LBRz83hBHFSvgLugoC2CfNe4jhlxlGLeuzI9Vj1PGzYNA
KsxbojR5L/T2P+fhVNWT8B5q5BD7n2guINNYnJuzDXA1AGM3dB04XDQ/Hgwzop0i
hqy9Pbwz9tY/uhBZbe6FjHUAIWUHMIAh1l0jJnjgTbrQi2Vebm8vSlz14mfnF5/c
kNzTSJ56n3mVoZqiPX+m3g9ZVlKzNUcgfmCFlBjZFLGMhGikPyWGnhi0Rd3NgZcv
3XjxdsYYvp9IbQgOzU/TeRt32Wijn2pK+W+9ugiIPgh4BUR79PJp9v5ss3qzcPsS
ceh+drqqmXwTsUnbvL4kaicTiQwdBtImqevQylV/iFojsx+wXmARWGz6tawtyGPn
O/VuhV32oyC2nRkLi/aoLppXhbr2HKbJYVLsTg5mG5aZGZzO2DUKIUmuO0RKMfu7
VErNGYVYZ+l2Jha5F0R1OPl+Y8Sx8WQct3wDwk+JTxzcrD7HQWV7BH+ks5W8kHH1
34BEafVUfJQGVqx7Jub3JIloUcJ8o1prqEbSSwhKfMLCDQtMhpovbMYKqMNuCkyC
4Vtq/dUzRw0WINlxdMl7qXobJIaA6iU7ELFNjs/b96xRLh/NE1+6K/84nV9OupZ9
WqJL7HaXe+ezdhPMPQ4uX3euqbl+zQqWXlpZ/E46PAiVDWogrRnXdCM5iJ/b4NhS
//3ZyIWMIvTEkaSGSHA+i4sDfcQLUe2nXIMiIMOcfmh1twvI6ViLFIRJ5yrmPgTe
UoEbPXsKGpGX8g5nhF86rCNofjTNaQfqDrk8JjwpnVaNh/P4z+jWcQCcIw+Lf3m7
+45t6cagLYuPCsYalNJkYAQw2elpHs6Yi/UZc6/nt9WCSipwrmiWyqVz6uMBBJou
HG/+2N40m4aT3iFx2j8x/SYxGy7BnpI3GKMa+m2MkmDIJv6jhR+DDAkDXA2aJ2dB
EBQoR5iBAXan8Vctu9+DIFca8F3HacU0zR/yU9DhuCfx5WcZUbc9ONspCmW4VerK
1Ui7lBA+K8/bgJr7rqdhfn5kSxplXjWV2Ie8hYeI/3eZi5U3Bqd7G/HYInAJpfNC
aF7HWZAGcbWkAEFlLx6HwqM0qh5M/XP6G8FJ0UAmJvJpToVjgV1vgKoiO00/dhow
7C7cys/+508kA/H2me2I5MSnTDc6Hcj6A7TIt8Kk3EvyLu3etJ4pufyiiCBoFquz
Y4Q4gqAO4fG1XcBDNSDY+iwueMGv/fyp5R09rxKOHrfXBAFXlPS6aztoD+xmtBJZ
b4khog4w6azC7WKWeZW4KGYGzSlRDl3r+Z2uxdhnNvHr6Dj9xwBTvbxlGeTBhmgF
+kIVRLkJHtwbUH3H5yx4Lo3l+sqlvVVykDpwcKGr4XIwKwZMZeLVrXF+s9Ad8LH7
IfrJiMtGOfZxj/2w9V3W9rcccZwOCnZOdweH2urlEhqRWuTVlz0RORW6B6WiHzHL
t/fHevWe2eSqfT7PyXIMEZ4wVbeE3r3otYThi8md5qcIxfSWhv8LGnhBavDiPreo
k9Nr/AjCdZC4LWdViWwN9jDLY28EJ+KsD2PKYh+OwT1sSbit+AdLboRiUjB5N8U9
SXg6SNB5Noz0JrN0oXg1qCVpqYt8jBzOGF+SO1I2zytSLL/C6rc1/skxjOSrSrbp
E4Vqx5pEE7XvBpYitKVn1q+hRLdu3OmruSSp5NUuhmRRdhM/n/MdJOMsShjuzlq8
t73+mLyIVzcmzocSo6eJg+5p3byV7VYuAHTQ5EFkC8ZnZZD1eJ3uhxkhg5jzWAZI
dZCDNazL9BwW3VwB5exDPQoKruFYQJzbashtSeqERV9pE3cx3N/lUa+jkynm+5T2
pIv2ZvfJlJ/D1IM5spSq3LyVo3dn40t15GUBxfGD7mBqCBJZwdhygkYeBRUTsxG4
gS7bNZMZcU0ItMFauGt2UAqx5wK/Je3uqroZ6wxYqbqSBrg0uz/e53TCIn59A7wB
nsILbEyCmuIZ0Ki9z2yRRzrsoz9fpcxCnTD1JLido5ulJDx9kiwEmWDezyI8kvmw
z/nrfGsCx9qbg49L+2NFVrDeFV4F2rOaFu7RJZyrOnkVM4i/62vvCjooCEPJW6sv
GpeJWee/S0+D9jh8Ukd2vbIUkX8v8osJLkE+U7ZM8H0DXlU06z9mXnqPx4aVJUpt
O4Hi0ffxSBnV63WfafY2is6mrv2Q0H65ijSLUrzvAS5zDaS/X5tuqq987YwkNJS/
NIuS7MX1OMAelSPglbu9yg9wPQA7QgCX8NfR0qw2DpkPxZd3HByfZY+x2JhaZyMJ
cmmYCujPv2MB1uM8rH5RJ6Mw5OG5YRFA7Ijf0hvwE5xfaR4/uk7vb6kgko1MnnaL
qm9iuCs3PAZtdCdN6uvs0xoJXsjLJgRhRK1fT//L4NXaxovWe8hTJJcFIlu3bVsW
UFxamyMXDBrp5rFHFgqG45M1mhQpjW3jn0uMzW6LBxwESjaQ4LonFJqVWYo03gx3
QrchRMZJBUFZRZdvb1HC5Jco+KqFAGxreWfUihM8UV4WlaJZyAmX7Fl4qCUQU+rE
lstgfFDkjmbnlMCtGkcqzOipMGCQtTdlmarYNqvfwz/srq8yJYFJIbWSMaDurVMH
raSsUbfWs44C36rEiljIyEbMksZkJ8uWeG8e3moyZ7guRstZ4fbWYcNWuRUteKho
wm4VIw2qHjCnp+x2VaWSTuOVzHdkEju8YjnLj9u8O5hG24s2vUrfvqvrdAt3UnKT
ikIvwSrYEPkJsa7/iO9JqDtgulkuh96KCY9c+8hZPMHiPM05uP7FTjrVEGwDKXf4
auE0caOyFIBMu1GlnqxWcg/uB+x/eZQXkeMMDkG2niyQRa6BRAVMyiw4Ukat6OR8
QYrY6i/Zhyxh6XHO+vI/00OKaYAx17RUXiKC4xVgAEAw/SD5Flu7RTb23nBrMqeT
jge+mJYEx74PUpNKMXoT6Q4ygKqeJq/3DpPZz9/S076RKnQueWAb3T4vbtXj0VFy
rVFm+8avAuyGbtnWzg8peyTCbXqLhkpEPyurEwVlpFVhN+f0Atk+hpqJ2HFYQ88/
TV8WK1MFQ67QYzvZtEYcWWXVDeaU6sA5IDCTPXeeCbpImakcLk05eG0WEz+pb/Hp
ZBAdlQs8QQa81jkNGoIsez7fpYoWUvsHt4vGbROF1EMoV8aoJegwHMrykXLpDNas
S4L3kZS7ZcNHvLG6YCYW/iWXEILkHhErhRfG2Bxlxtb2xT0+SJkdJzmXuPw9U2mi
G7r7dFgz5zWQLTtgFnVreksfV28vRdmLjsVG0vHYyxjtuKWupHlHerVHnMz2kBwh
T5T6fLLt4WvSvgutXVOTNTa1wKtHWkY1gp0xrnSAOYo1oc3rKyCXD8wCysZ1BbgJ
1y5qNC5WH8QEVkgGZhuXBC4L8NYksNWNxPzvVlAfSPOK5SpAjGFFydp5+OD+QGE3
IPuEL2sgjFlvAHQVj0qcec77bDzHzrKGlsHpc9ee4POHbkJ9Rq+qKaUimXkZWUAQ
Vsz4ZFiV+h2KWzHaDb8Cph/oAvGbBmjID7fqGiGXK2QB2mtVfetnFeXqG3nSCPdd
icjC8Ac67TaOYV3dGt7ekxUiQbvcFtGgNNKLR/uDfqFh6dqGREUnsYprArRUq9sp
u1uKzm4jm3oGdUgov23/KxozBs9hRmX94UWciO+n7LRUrk5zGjWni25Z6AN1tJfi
+REiR8IUIIb6DRmA4U0Vi7B61f6VZ0hD8fJOtIGgAZCS+W0nWj7b1TQGomeMn3og
anAXanYyPO6SUWLi0yQWleOeKYkcR9/LZhGKxYwJoMiqdVc8PPb6oJvk4PT417u7
xzNp4q2tCPpXtnyXOqOe0tHbTJhWWuD1hE5KZ7UBkCQAbxptVt/R+qk3w+wZgB2g
ZCzcc0YvLvqmPv9Qu6GiYgiiuU3FrJFSpX5JUXTQ3r2vrErvyljBVaWETAP+ojzl
zevqnVFGQjYrzhoRqKy+Uw+s0awltQp7z48iWY+0pmZUGj9RPkdFS+1XGbCEisM1
mHBIHntSk6JToBIZlxTT2WcYGzbSTd7esx9PYAmkJ824gbEhn8yo8pY9x1XbxWEU
OIvFWJF+sa3i6yfiQsGcTzIt/Qz+g/g7dEHfINDJAopT8Z153uHjTFgRWcjP5hp+
AbZVD/vttLoKsWJOqTyUAFe6YCGVBYqG92Dsh3vGfkI/hBowy69aW3eTt7Y+M6+a
cIFgrWf8u30e42VakBZRgGo2ZMQal8RTc/8Fjn0fm5CS3zRtKjDiWnLJ6kuotoRX
EZNqLbYGItqm84W2RfAY7eijGuq1/Q20cC+USHSYW/DDBhlwdM27aasB0vCmrDzr
5a2+4clDKVSFupJfwU6QNxJpNEOc4Ke2+h/jtOZgBmR0St/dVuMkORASg5RnyxOx
tn6ciP2n6dahCt1LHPKUVF/XcuDdkhEaZqU/Z2muPwyNnIVL0UJUKiYT1zrmivQk
oTgTZ79k8V3KU/DhhUYngxpVdAvMTc+G68nX7QgR2Wb5UJ3qosBhrMpYbLyjITjv
RFbg4pyqA/e+KxQfCRGAqPVIiPvxdGF+FFaFzBrMRmzM+0hp2BKofDOFHI5+R+tx
NtghXXpdowOB3Mc53iWFBW+qON5vwcQCqYW7gHKzDehtEvoE+Un5bDQ9buOeEIA5
KBpXEtaRjXxKfRxQ/rMJQ44/b6v2mRP7aU2u+yWdOpVs7/tiLtvqkVYw05b4QK71
Ifj4Y9LCE5SrYy4e7hUiiHDwJs3zGxJwxkM8g6Y1KbyPhLpmCH9hBtl7hniw15VB
EoS8L9IyU3pI7zuILff3DhBfLoo9dYFj1Cd923hxTbgwk2Cy1Zbl1cIx3N8P0eq8
ilhkx1p/zi1zq60yqQbIWpa32bkhYuppneFfJIxghBqWdvsoA6lZOvu4xiSwoUSa
`protect end_protected