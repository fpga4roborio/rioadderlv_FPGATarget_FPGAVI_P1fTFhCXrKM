`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
ddtXksX2+yylW5zu6QL2Lhnb2d1sD00763mmSITNX595NcHTEkwn0zB1Dry37fOW
FufOhVzEJp80NC5qZ/+F0Vk7Ik02dIR0elf3clrjeJRK85K4e3Hoo4xn7YbFUIms
l/8VZSb14+JVGURjfswrIyCUotIzlzVYZ6gzoZwDXIi5gQIBf/gI+KxNXPaKV+PQ
Ufys/12rjO6aI/pPlqSm0hCvftmBcnezN2hk1UeXgOIuKZnogjOsf0iJVX2aOOWE
6pD/psybjbnsNB6kH5uFTA5frkzIzkzl5d9+YDm9OyC+k84E83I/7/j+rk4L2dah
QJOvksSIzN867/4Qt8qYTQ==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="MvBXkzurAa5VTw+1JJ70nePUfoQXBvZOku/SMmg4TwQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
oRtzZL4VJ4iwysPsC8SXYCzXS8Fw2gtZTOskLcDV+1B9Nzn1zTyNtlo6lNICRmmK
ZRVu2BmCc2G+fmzynYlNTnSa7C0Cuel6FYpxCBlOuk3OF2tzAmLAuDyOH3Z1Yjzk
a0aHuoCdIRKv7BrZCdALt03JeUmXKPdOmIlkVGFl8yw=
`protect rights_digest_method = "sha256"
`protect end_toolblock="Jn9CQpRhJt4rnzZPRk+dOpzAubz7omckX1MrFd4p81o="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 6752 )
`protect data_block
gD6l00tciPUa6pDNTk/+t0OO0nC/UTtBwLB41d4inuAUA3i/ALrNyoJVcBnAmEQW
ptbcNp5fxEUJjnOxnedyZEuEBxWRieZFQnkRdF269oOuAB7N2N4qZ0uh6kkNSbnv
cmxZvXeeSWVbx3Gznl/0fpjD1PUHUuqs900GTE/prnf5UJZAoRbh1v4befoA//bp
+RVq8CXfFR4lRbqrsoCO/Dn9k8hcwKVNwPDvEScLIAsvpA6KXwJJhU1xb3ayVLBA
VqhzDfKapHHb2DAU7Ae6UMjZVD4dw/QuYfL9kY+o8khGGX+OxRt+qqwr+ykw7yVH
PYy5xIYIONMCn5r2qQehfVXk3tUySs+0Hbix0pf/SpifC328JCyJ+UnsQ5iAUDwy
Ehf3r5GDWDsySFuw+c4rUhB4p61+MUgRE0lZGGzQmRptQIp1rVSVtxO724LADxmN
tPgB2X5ogxurkrlUTi6vnr6DuMyRRqrWfjG1hVRsexwE+remrQt8Ygbi3ym6gcE6
ub8tVW7xup98TM3Tm/b6Afd9IQOMG+RW/N5K6K+HKlm5hYpxS2zWZvWcsAeva4nS
yuVh6+F/FBLi7WFIJ462Q4E/G7L46UJfFeTWFZnVcs3CXs7or5BptLXiielx+z7V
/LBFcNR4JEQqvAO3bpE8C1krpxNqMgYaaIqsndDKIg4wz5xOLATnJxzHI6Zvj8KU
daieSdrlIs3G35k8grEWtqyABZlP6BHiwWImwrD4kP1SPQptsxQZGSgrE3/i7OTT
VHjQ/UG+tJv0OmCqsB8WRbQabrHbgj/QpOgmB/pLP6k1CzCVq5fwaw0flZzYTGIS
pQtjT2jekssSmYEeYfZc1UBwEL3rvYh6mcqsHwK1T/H97VWdxGjxwvOtUA3RN4cP
y6j4MXQ3T28Ifz6L1Tz+V8uIQQ6UdXeO1YU1/u3J9TWZzGBupL9TVY9vRegidPrS
qV2o81wh96dIrSzRP4KtDuJTjLgtbOww5fC3jcyzQCIhwYXDq00tdYKOOmCQTKb7
TnN5xRI05AUxU+8fs11Y3v1XHZdQk0OlCbfDUoIHmwhR6sLg4Ib5NWWiP0/+kMAn
o+bVepFN64GAPnUy6hkXvBRt68aeCkrPrXF3YTLHPz3UxXeDbCjl0k6qB5WVY2F5
KVe1ygxCivNugzQ2ctOWQBRMwEL8F5oE7MzQE7tWBLcu/IVgLvtkhk2qqCN2BcC8
/Y901JuVFMNMDSLENSMwFgUm445oqx7rrNsudmdFXuV38O4Ki1LEyex4u2a3rySO
9JRoqx+/dYCDDwt8Qx6NWTUFtQaP3BL1/9rym0FhuwhMlEL9H4zs0IINrG+v9JlB
nDdrKEwf70VI28dqp08K2xh3fAIMFBXxkBh6bF+ODNc9oQLfCMmOibyNYBMf7TNm
ugiuSkVmvnOVrRZ9dpVmPRn6iZ/ToLKSihc15Bd0p8jtMfjYQGLDpHXpEbN959cl
PUMhUmOrVlD55xXKBlizmz0ZffrMIrQDyz+UfpDo51tV1o3RPM67kejdOVLRqg1T
szkWLCzt8htrvxPkZwKdf/ZBfiKIWLo6+YGJUhZfrpaJ8T9+vWffTKiBcFLUHnCB
DFz0vtqQNTZm6VW5eB6MivsharWF3gGqpos9n30ZYYcA+O/CB6EbA4lVSnsItqfm
ZhJ73K6jhxb+FEMuAhMVcAFQNKeBOuhTRP97G3B8VqpjbJBaIGAp+zfvZq7WAvso
YiLDglKCIFBlZoYXigAYw+PLjLzEWVQheVUKfqsG6YcMm8wvxke10vL638YWmZjt
jpdyhwTpAIHwD8ouF1N2aUUkD96RP+oovlsst44hBwm5cnezsz00PxV1CSD7+9Pv
9Obd7sAyz5ITP2ytu2MgOPOQrXGDbEzVqMMSMDCf64AMU3I7A7pLmro5j3mpjAaj
qR+1rvB/aCA86dugghWyBNiMLgB0SO/5s8KR2vz32XBC1jO6LmfvgdmcriG5xE6F
kK4EUfP+2qWItnNXi/Mt8E7jvbruQ89hRihszQIJWzluoPNGDGvTwOW3BAR0tq8k
3mSISn4R1G+sCvt3BiVyHsOAT3VoibRsJr4leuUpvvAmzNY6DysyqPO0T6jU2QXw
9EOyCWSzZRbZtOzopZojpsq+7nNW0nIi3e+zcBPYcSHaOPvY+1BxYceI2iTKAKOl
qQLRLo3jU276TaeTl4cIuaxneAQuS/5IDPPqVzp489I9/9O27NmDGAm0j/TyBo83
2HVzGbQBaj68bHkB41qpd/X4QymkHmz8Vl/zVhFOnrUyFHlti/cTQNU3Q+W4OzvR
tlCTN75tFD1X5WzK32m/nMQSSdF1LpPl5pyUJaSuGylMuLQoJw3oQMSSW/XbiTDO
jV8Hc/cCEB76lTKVQv7tOL+O/F9JtjbhGs/YD/t7MZHCWxnxHqxOLBe5J3XyHzHi
Jk6+qFXrE835OO/7ZYxrAtofe1WccC1ADHB1mvdADEUzQZHi2RZjZtpJeXRFgpED
OMfulEisH127KUnDwGJuXcqM86HWSTHMK5kHHKAWMoyauTpsZdOn0Kho4aQQjizF
i1VKe9A7FQTkDE/24IDQX+2cyWbrWSL69HVIBV4oYsgsiF5bM1jLgatKhLNVqtS8
7ukc206ZlR/ZLY8lK0ACn5vmDOAnAmDCtGyYo+64Oe1WQA+mu63auNyVDjjRP8z7
KUldCT4Ls5WAxOPRSXJpcz9edznpp3Fmlg74GnZfw62q6CO/oIEbXwfFlPFZFJVs
wWdrZLxSKJLdYNfz/9ley37HeTdS5wGtAsWSGnqw9zYdoOLDTmT7U0XO71+6i9T9
8edQgcoGkvbR6bGUYzoDdoHHRVFZKSZoPvHT38Lwxj23OEKgPQu6TxBnosiyKaK+
DZabGlzUDaCppEOC0CZlx6UsiEMkVL7TksR3+SzueLsmPGwd725RchAV9xXEW+6w
10Ad/4v+TcKBAb8hkQe95XGs6txE68D9kG8JYK8q2VWO5KvfACXRn90kfUgbxK8G
kb38ULGO80ZHbdZxwvl/j1eEYK0jKVjZpzyERqlNWldVJan+1ljYF76eTxiejuMs
b5xyQdzfcDiSxCoUu8b4VFWSp6AeInXUw4ne5VSmseetLY5m+PEyqNbq5ztD53dT
7fbDaJRU+DpE6sj5mLTs1ydx70fVLaflevl69MrdSQtAqn5IbsFDgZHBdApK4IPg
+lDPtlljnx7VtPaugeY/v2lLsEzgS++wonvxaBIJA0y1hnyc/Z90mP5pjUjv7Z7t
aQ55Iitk1takv/mxtzDKFUyQP1+4zgorftihJYHIX4z20TdYvt8NOpfe2isq3GlW
cpHIieYRU2j4CKhVITccizFRMWIeZdcBann0HQ+PoL+VFkfVXFK6juo+2t513Pg5
l9B3ujJ036SlPS1yCNjqlnb3PdUq5982lHtxW08UPTsG386YAGeJ2tNfO902Oqcd
dQfP8rS2lU767yI9jQSUQTvPfF9Wh8pcBC9mq1PUB78o8L9bsmIvzYmk54F4wzIq
9OwnGWzaMTcqGfAdkxZO3DjVeCBLOlv6YIq28vYmO8MR78H5ZXueYtCa/fH9jxyX
BhPPP9DpkO/x21ZJiuX92TnvqkubG64QXLxiLueJaAFpeVg8iWPiPMPDeSOfEeZ2
yVTXt0NMPrN6rZs3RX7CUQeGsYHEPs/untfVC0vGfXODHc2iC09UcX8UisS2agMO
FJbrcTYUDTo1IvnCFNe0Je34bUneWZ4uWC7JB18/XYXQFc4K9vAZmkCiRJ5lPE7I
zmLNqrjuDzju1MTz0CczA2KjJqIZ0373xyLv1n1SLq5OQsF/ehDHzVpzvb+A7OT8
cGs4qw21sJmu6LAQO9ni2btRx5PZrR8ksvzfK/5YagpSVTSZAhsWhJsJpXeWoSKM
p46uyPsC3LczoHfrJKZ1uZS+NX7nYPmZgdfO4Pd0haiI5WXlnrMJaeSNNnOYohl/
WxYRSxH7vD7MAtg8ZVFevVgDoEnBqEQTkeijMNW06fh0nPZdrB3ehra7M56vDQuc
KVzo82SZlspN0pHZvGr0uG0b+wgjpiphVvI2N+SVOxj6y8GuFH4Vr/VpxOcTwf9H
hcN7bJDYuHwUer4NUxdqK0+Dg0gcV8Pjy/gXmczZHTlRn9AkajMfqWhWANuvfCJ9
zfMc7fqxd5aomiZ5eVuf5j+bBn8UuwFx7vI0iE6xr36NXhYmLUZDv9QwikbHHW7x
shClVf4+2UZIH0vP+MV4jQUMZk6XDCEhyVQESwhD1QW3jZDVH1n7EL+hMeCc82+m
eAGLi5n4nLHBrPRllOQ1busStl2EigvKrMLPFmQnkg6ip9s58Rp0KC8J3YOgTu6C
b2c6mj3OBHBbmOdXj/bslBWv175VKiaT+0doegpX+byN2a8tgo+vDtN/cBq29OLG
Y+HdZkzK1VtdH9A7dsqFAYtHTMJYfaHUh2x6NmVukbzgS0fiO/XQoZXKtDXnErhl
KhGsgAMMDn8Tg2xhGR0e2y/X+e742YPkMJFLDZz3KCLwmbUlUUnmt2NNvBmaZhEU
J54S8GGJsp6Jt7mpDGov7TbB4O1gFj+yoWZCQSHh7CsdElWI1juuMeGCz7wbH1sz
h0EIOXP6kB7VXd+BxiyN1OtQTn/1mAsa3QYWYYzZBmuFMMUikbyxs0dLFpfejo7K
3ASpvIa2/NcjnTBgJy9OnE6OcqBdrXMe7GAxhJM1UMQ2CwLBZd4CGAihSAz2ndFY
4lLJsq0JTKn+zr9RnQ8KUolh1RzU1TUYMyK2wKeYzD4z0bgBe7nhJzIQt74j1JCi
+mBvMNy2dmJoNswlCem5/nA9oBX5KCRka1syKjxGZmOtZAzt4UT8EFMUSi+n5xVg
SCoOii6s7zAcgSHoxS2/a5OglQAQsYLkT91/6K0gmxVWK9OsOLyl9X82d3BT2FNj
6W3vB1iJb2L1xDdyuSh/ctRzThBYBcf9IhTxGzDF2ZL+pg+WLFM62y5dHylIPE2E
EjgVRmgI5IpdxOQMQzUm2QAIJv3dG30ZwSsMSlZMjtEY0iUmrqU9aTRzl7qpDUB4
jLa86r6zkL0KEGXc4SjK047hJ0aL7cBwMCGBrghnB8VDzL+/Kk2s16vOaPB5zJe3
IxNElowYMkmFBfrdcaVJGJsfnbxZOsDCJCk7jMHmGBXd9D7ZrT9pzCdgVariymHR
1bRNn19fbuZVsl66trBiT0Bp8elstGa6TW2mONPEisWBJWCAyJJJWSCYSR9fOBYR
aRZR1TMhaNUGgRp/XIF0bQnjdEM2fggazPQSmCM4LNLuXdAffGdauJRRtFoDCudm
6khcRM/fZlbycRcXsBsVUY14yOfi7zgVYJZjKTWpTU9gg134GsVZe5Zcg/jzreFN
Eaup3WaMC4YeM+k2rv1TidUDZIB7nx7UoVRS+8YF4BXIwlZjMYJIdU2/+5NcCPyh
Zg6wcyeuxpjOBlj+hoFh3S/OC8NzfH+O5zGfk7qKkmFCe5LlIzgsISYEfPgMe1GT
4incUlzoJ4uVGfe7OaNoyaaubcHu83jMqemiHLFFRY0jauBZ3VaP4NaU11i1/6U1
LEccoUrQkCQzzxuIFEoaPANgMOtJx7PpopOHmFP7moHPuqA9FJRQXgtLFWz+8322
RFqy46/aPjMc3+9dXZBXTI8Qt7B0QKcbvTmJHrBREYFQExpmB8oncusk48TAZwfq
Yc/lN0QDfre9kwE/HHwFsMjh0ubc2z5SthC7cXRl8rmD8hvZ4S27uBYphFrHEpm5
jW8FpiEWaZYrbjhWzUVsLhj/uZKuyZ+Y/uQA2SF192VnAGHr8w9KGgOhb6cmv+e/
jugkpDpljiQE0TsTapCUtV17G+lqlWc18iF1w/MNw+sXbxkHhy0u4SMEIoAgWKfC
XM6UmKxHXrqC2CdvVN1ccwCpe3OSGZraubOkbJhEg0qjfbrDxNRb8YsLfYfWz6Pg
3R0vMTtR+0zjj9o2OtmATCJ7jG3Lvuc8bClW2DP1ZuMeffQvYLFn3suYw7KJsTV6
/oo6Gq4NZYigEXo+2w5aoUaqvZQm+U+Xes/L2vjuIQTyPmGYWfUmB2WAcELno36O
+qmk0hSVIMwLjENE96WmRiMyRYk6X7rK94WLD4yURLckgMqikgG8vNXccy6lmVSZ
RBgGU7EQ813PrXC8rgF5CWsI9/GHxd2ti7aUugQ9kCCk7NP9ZKRYDuOtmuAmyA2M
oYYhqMKM1JsPi2dZTOprBGF+HxfGw2rVXH0KNNr1I9Hq8K5w6k6kMhLXlkCB3Fj4
wrZIpqT/YbK3kTxu1cFuPVXEz/7RbEPl8ZEhOXAg3gmRcXnzGkHJnpzllVaqTHXq
/4N6+gM0Tr/SNi1beT4vuzSR0mFmfXTBfZbfZaAVtrvYGyRw199OWjVaAd+gefAD
yZ4Fc54GRsh4PjWX7M67cCfMcU0+nv2iKOgo9zlJK/2N45jpOK8gXPYST6a5Hoft
i5VRhlAncAbbkz8sryz1QumlmI1/zFdpw54cU+GEch6xzNJ1S36kb7XZ2Oe/JiEk
dQ55+yWX0KGAFSZFULctrFGqRgtigCA58TqZWpDqkPPCrIkq3SRaA8bvIapAgQbY
tDejvi+KJYtsgEuMjxpsJ6QYMJDwdRIWaaQDgSvz+mVMVUaLOqmwu85cq4QG6v5D
ShMUfyT/AYGx8JhVn221OhmxrW+7f9ezIemL3/3h3T9E4vKz2iRphdmXl5Wi8CpR
i14SboYaxeIi9GDveFud0jldKN3yxGqSKrcT48XFaKyO5g+vf9MQorg1OQdqv1+Y
4rdW3x0Hc8zc6XD6Vbphg95Jb4j4js3SF4OELVg66AdiooZ5WfAwKwlDf5lWaNsX
nhuw7hokYSWJ30P6AHtwx3vI9xyj1Y1VQYs1WlWQdX007l4eImFWIwj4qeRAc3MP
f2Q1fmpbQFLpnsKTLTs/Ohkc4dpyMzluP/vrYo+aqymdeBmCh2AORGk3ou3ZWULO
x2NBnIqcfUt4G419//66h7FChdn7yaWowJ+HTVeSKwl+lBH3LPUUpZ+osjq9r0ws
c6WUlMDhxtRAQmPYvr69qB/bNFiYyEpp2N7SiaolDYM5nGxxwnYY92Letca2btXS
AFuNGzt3HGp31u3zhs8WSP069wnEsnBmx4dRBsGES9/dUoIXvfWPmsivTlTmmIWl
q1xmQLY1lP10kAFKjl6DoUx2TocdeH25YernFatbnfHM4l7zweLIZ4eUp8YjWTlV
qUT352KoklNnYqd8fOvbePfzwqWShPkAgi8zkzsJraUmt0ZL65LNnKF6yFOExFAB
93xT9P9c3boqSfrw2cI9x7kYrEdcMD9lUNzfadXbUJejkAtDvJu/bCisJTvAbBVf
ZMXOJ+b7xyMoEShKeb61G3g7nn24abc7vTVp0wllTCXMybI8lB6WDCbJMoetzyjx
+l4EmmIrWBxQTjJ4oBoOHG2J/xJRiJSv3IZSy1xiFiLWwbMhHWTt+7nE4SuiHuIT
iZihs4lHDXrQjbO3TWl76oWKr072Gj6W6e7O6nm4WmL8wzLfzuEbD/TJs1rR2FTn
+LAAUj23zJ4c4yDOWqs3GCbYn6fct5CeLm/ebaL09JvRoBs9rmM9qvxkrAj9F7rv
GTO/xjyLM2bwpvBSs8RMwu0KJMzToSi6Yu0BGD+jzoOReNkzEUG06mj/XmsDhcSp
dxbbP32zT7GGF6sg1FurAuL4hDGqHJVf0bhKFylNOpDgsLrm7N+cZrtp4ClcpnNI
SNTYdEgkZf8VJJVIYTM/QjFOc+kjAI0L0TRvacqO/UMaApX4IhApL6kP42j6XZik
k6quv5qak6QKIHSp85XuQuv56tvJBQb8BIvaDoe+7Ekh4WLLoX4XJIwCGX8ymHf9
dBnF+6f0MXIcUdEcJOIdyz6W0cUv+An7xVrSt414txLBDcj8f4o3VwEEfdA1S7n5
GD5zSxSh58uBs55JvPIl15NT0cgjDClNFE9LQn4lbgFJFgm0NTUm0H3/YKW5dQpc
oxOcogU5gDM+NVVUPqBonO6+1jvPDBAZUrojTzdCDjmivlSvvH9UH+jLpZGqvvpp
yzYQcLMlCdCwkTcBtZ1S+SjXW12tZS3stwWujC53Gk10sS0mXFF4cL5rk1tIamC4
ZawswEt5pG7bGZD5LIemjJ4Om2p7AVD45qaQY+MpNrnmjv4dVrmfrnTCvsaIC/lX
Q+gp3rwSGIK5e63cCoGv1I0xD+IaQvSNMtj3Vm6/tkazrb1TQ+yLeEz2dzOUPaZs
xd9CXYpCuYWJF1yS/xvz1wWvhrsRuAOGF1S0lJq5sh7P5jljkYljnlXcmSTk34cF
SzwldEBVvKKMRAPnxkxvi7yrM0O6NTmA1dPEqdSl0zl1uyRgZCaO0R6Y6/SsV+Xx
IIN61T0eE/ezIDq6P17q4U3sq2MLg5S27y5CxJhVBMIB6I2kuQnJimJ5+IhTwaGW
jpGbISi+CmzeFoA6JO8ZlumLHejscTSjutLCb72u57YhPzBRlpPfrXSWUHUPB42r
ooRoC0+YkC/x9AjpEA7tLHk1EABCluIiz4Ues31Su5YiNEBSfTMwmuajKsWA7hcR
Ph9peB+GcVEK/ozCv8kmCYq4G24eDV8IC7NXX8Ve0yqLUJ7j/wA404SHAOSCr7ZP
Ks+7yf6zVu41GfNE/cX8nxp7z6m4DXwq4kBcGkY3kSo/jfw4lTs9UzBpcBUj4Unh
ojlLB+h2oPzW1ZBuWbaTOq9OgxPPe9j0hg/0M11GJEsfMZtA0TCNeZcjygMHkHJv
FR78iUyB67/x7K31DQ9kukANlnKDITB4zrbBX9dV0eSuI3P4nN2MMY7lHSwnGO39
4Ggy14AdqYL9OXb3c9d1Qy4VSDeJ/ot9lM91PKNDaQ1/4ngu31r8888fEln9Fg5n
QMSCNa9vCyyt+XA3mJ/xs7RtMBzUqbvjYR9qNefh3kFuXQpU05ZHEP0llA6bUgXZ
gBp/HwyJLwB0MLu626Q2maty8ffHWWXC+WyAVTEjeLo=
`protect end_protected