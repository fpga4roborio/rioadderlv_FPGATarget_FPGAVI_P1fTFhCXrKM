`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
ddtXksX2+yylW5zu6QL2Lhnb2d1sD00763mmSITNX595NcHTEkwn0zB1Dry37fOW
FufOhVzEJp80NC5qZ/+F0Vk7Ik02dIR0elf3clrjeJRK85K4e3Hoo4xn7YbFUIms
l/8VZSb14+JVGURjfswrIyCUotIzlzVYZ6gzoZwDXIi5gQIBf/gI+KxNXPaKV+PQ
Ufys/12rjO6aI/pPlqSm0hCvftmBcnezN2hk1UeXgOIuKZnogjOsf0iJVX2aOOWE
6pD/psybjbnsNB6kH5uFTA5frkzIzkzl5d9+YDm9OyC+k84E83I/7/j+rk4L2dah
QJOvksSIzN867/4Qt8qYTQ==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="MvBXkzurAa5VTw+1JJ70nePUfoQXBvZOku/SMmg4TwQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
oRtzZL4VJ4iwysPsC8SXYCzXS8Fw2gtZTOskLcDV+1B9Nzn1zTyNtlo6lNICRmmK
ZRVu2BmCc2G+fmzynYlNTnSa7C0Cuel6FYpxCBlOuk3OF2tzAmLAuDyOH3Z1Yjzk
a0aHuoCdIRKv7BrZCdALt03JeUmXKPdOmIlkVGFl8yw=
`protect rights_digest_method = "sha256"
`protect end_toolblock="Jn9CQpRhJt4rnzZPRk+dOpzAubz7omckX1MrFd4p81o="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 3456 )
`protect data_block
gD6l00tciPUa6pDNTk/+t0OO0nC/UTtBwLB41d4inuAUA3i/ALrNyoJVcBnAmEQW
ptbcNp5fxEUJjnOxnedyZEuEBxWRieZFQnkRdF269oPK7yijrIkmzs9B8GvIF/P/
qsCdz7gX5n6YlxRILMR+xlLFQfCjkkTAzAdpCZr4857I1EEII21nRUx99eXPB1SX
Tt+iKAHBt3fcPX/3hhQo7E+4mCnMsB4kgmp6zVH8ivuzk2lKelItqI7GylL1aTF8
Lrq01UI8SevRNHmKworxav0JVKqmxmT8cfb15YJUrAw2cAhSsDJTJhCdU4Vx8N8J
cuxyNBadJhuRRpP2ZKBwTHwk7o6lFcyGB5x7JpQ0FHzwDbT0UA8TQGRHsjqyxuKy
M0/ooX8je4hlXCABOWO5Go7daRAp3Lu38wJdYH3RAfcqp/u0VcehqUuwzcop+pxX
JgUYOV3qzT43ZxnBr3M82/UUOamKwEcwL1kxFPJT7yA6pzWPmwZAVt7lY7jT4kWY
hW0IjmRrj29DDRRXrIUgDc5GgJWMsqCR9AMDNT+j/TXqEdlbSNtYUQC3OHYfNOH4
C07XTYi4K+TWq4nEDDpQiFS72ILzYZqQecCRdwxadDnaaNuJjVef1d3c2RJ+5vzw
qyOLApWVviqs7PtGFa84wKIQ0S1MT/RMbFpFfNnBDcUuaqnKhwt9+meQRS/xRD6A
/1hLlL/Tpi+PI8s8gzSZiQWKZLJ5W36dVnShGI44c1P4Mw+CH+2qAE++pRmXl2Ru
3rua1MYsZGT4yr/sH6t/iP5NYn0zeI0w8dYkGy7wvs410TmFc0yrBPE8pSTnTmUV
mRWbYHjjqWGvpMQs0AnYpLFUy1py5MsheBC+7U3gMRchl5kXeC4qiy7Ibk5BF6gP
3ZW5UC90gyDAKFnWGhzhGaKDQIQ1OTpV5oPfee3drSpaT9oHIHVsl6szT6shOMl1
lREQ8jevxwXseWyYOx2VW1/QsxxRK4jShHJcFDqjKvrZCTJxusJQIXwr2L+RwMjJ
PGFuANtYZMRSE9YvYuLPJYKLo6Nge7HoDOcG+zjnnfGwG/rsELwcLEncRA4tS1ru
otKJFJMdT6Lj5nnWLXWDN3Z0lch2fUKXb8hHhvGtzWUKm+OHYdgOP9D64inZK3Zr
s5p2YxZEOKkBgez5p71rKWP5Gfck7nRvH5KE5bO+h2xDH/JIm4zdhRDD8ZCI+rW9
f+FiRlP3ePbbZZYiK53i8gAlDGG9R6dt+/lqnr4EoVOBHAmlFYeOdhfabI9l9jng
ir40EGHAIhpxAIDvUelsShGm22e5EXEmwdI0MwZQA1y2Izd/4m6+Emary+KzCsiA
qzrpMFeVOUcuG90y71LM2TofscP9Y39cOq5qHVoGsv7D1va5/ekmfsIM15dRN8od
YAULCAnmzQk0ePP7OFJ8TTkDhmPioFqFuFFX2Y5e3/Xy2IoxAMImBQ2tmVZUHaeP
Y0Q3XNUjG2rDFN0J7AkDHniz0AOQCii9doHlqHI6wIeM7MN8De2h1s+iup7X1yUa
znwTUgG4w7u5vnhqQZeVy/BxOSTGmcX9aJEdbjtgyNdFQCPRdW5SOiy2sYOEytxd
DYCsuRVyR/yOuHZV6EA3aP1ES1M2hMl3WdRviVqiwHEWb6u8fqIBtfNJ5mvlZE+l
VEg+Ck9vtimVEEsRiKdBlvxo5yAcwhcT55RmA6W/AxcyU/6VO9cduJL+JtmSR4dr
coLkg9pjMpMEtpDtdplx9frjQSzylm1b0kt7QQWVkyiWPnLd3wCVOl2O1k+YRG+A
O6qZQ9Vq6HtMBvWr2hxiqHzf9BvPzv8BcTz0UCHzJYbV7TC7KhiSgQ1XNsRq5CZT
JvBECkd2+ZQjRWug+X0n6oPgBIqYM/LJ6lBkZaBl8ojg5YhXeAXTWivpTyCWjAK2
AJt1sind0d+W4C+X4OhssffM6R1+tyjyGyHliLfYyOX5H7quU2gR2+UPVu9fI4jC
QX0qjFT3BzIHjNQkRrKyS71sQCus60sFGQm+DMsNKY+QHtiPR+AV9439BxssMjfg
c3lwIWTytpoEq+i4R3Z6j4SJC5fWNq5r16X2K6/IA1wCCQ1DtcZs40LMoTN+mual
TyHdTb7bDWrAB+UDDkawOlEWLzfhwSBz6kpY6mbthqea2Ifoywd3ba2qHj6M0bZM
vFyr279/P7DWFqeh4R8XYgVLvhTasdZ6nVflNu3aorTyIhxiRcp3TCm3DNU1cUnF
j5Jcuh0KBBmQN0sZ0M3FqfZ3SI6iuwOwL/p0PWxn1KQ3wB1mokLpa5HMXkDuMl53
omBGSUq4XAzG1NywB33dCo28rBJIrFSYohR3UZbYR6r1wfStEWBhFo8VDnTHcT2+
i8VtJItkhae/pnCUZabmPEvnnIGIens6NHFE2/H3ROlS4zCOK11wogu5FjPw9SPo
S1SH7opUm8ZZ8igU06Ibw2rtVzR21EalXBhCbwof43ZbiXuTlhvYoqaBZZZ3IdGb
aijoykeJSlgLBn5mxsnj9RYJH2H4kncwh3o/MZ5vhG7PTU7q82A5nPUwo6ma/2tt
FiF1ruTpS4aKuJUq8scOYPzXQTehNfWKI1s9ajTKkHvcpdL7N8xtNc2jAi2wCprF
nr6S0tCiy/j+5XZM44lusGTlW5Tvk6Cb3mTuI5bMQ8Di97nVOsBOIiHIR1avmkfA
QH0qbvWaL+2PMUGjaySBNl2r95FSCjH7qoy3MI5XEkZov/FFG0Y39cVrpJKpnjsl
d9zSipy4AEgDQu1C0Vf1r+wJ+x23krlyyFEOBZ8ylRCSaXUa+xtsqj/+88eipcQo
wR4GOauoapiY1jXyX8qfzmhm0VwcVDin5OShgnaKYJXPtYdNaOdqz+Nz9NGndG+1
gQhRv1r6zk+KoT4iNT075/ZQKfMCtGi2eO7heQwsEL/O0IA6BX/7f6VslkqRj7Ex
FMxzMbbqvS+XDMZWFQjVW7MVp94P6pSChaqG/NK1jLfv60kn2/px1DNzO7deRoDj
SGjx6kSOElwrw8J/VlXiGFOdDQ5i5Z4fEucNdR+j0rYnJewYpkzIC+zpRWNzpijM
5NQLJ2Ysw70DnQMCMH8ZuLSwOpOcnw7ZTPM3LxnwK9b4o3qFdX0cfFVT73qWjYzz
0t1W9/0hk1ygzJePiO9MkWqNUIE6YFZa48mAW6j28xwYf74gnDbni8Lo7GNJDnSD
6+CPrTWEB4VDFcD10Absuum6PLFklst/qu72ArI4lZh6IpArFZhFc8ThN0HNnnml
bn0Huz9Lw/LHrVOldCwfqwFdFfiDui1TeF3AIfWGcbVSmNA6jfiy5xPI2Hybhdgv
vXG+F3hSGfIBTzpe2V2msfVtE6TnW/NmxZQQSVsEqQsNhxWpz/1wSYRzJJgws4Kg
f/BERkCMotO/170/GxL7PPgBcj560lJftR2/Ka4CpHHFHj2wOkhPseR8aocj3rFD
YHBx1XdwaNhq7v76YCIMjhM00DBCIm2WudLijosiob5SMUJHWkgr1CPDXBgSB10o
mIMJvsh8uyPvlV99vB33NvgdJZyo4XVe7sf7PgM2fisMlH89T3R97vH6OYFqA4MN
wWk1fM3bcEDQlMKr51FZqAajXDaCtNxalq9XXZcPykt5dx1/KOPSR55evADzkRZc
gyI07u/AERX7PGb/nxlkCkLn2Ewt5i2kwBVCiElpxVOGvczEed4WtkkpZ/gop7QO
75mqQaq7tZ8gZTDQd8vq+0YrvE8AeGTdnQ8Lfe1DeuNqsCRO+hRa7J/TIziyyvew
sugSeZJsqYBNjD0dQ91/mWouV1Vi/ObaK4jogM5nEPBbLLE7fnosv7Yftcp2lnOn
Mj7MnpNpewTTR9HTT2epicjA4mVu1Z7rNRh+AoJHBXIF79rVoyEn3Ns7mYb0lzSn
gAXbmeRfI7IY4i6wR4m1E3Yc7iM3YBnlaMX6UhNoHQGxnmt9hFEjm9DjlkGYIavg
l8q5oG1wZqfAXRD1v9/uSxyvgZC23a6fS07xjF2RJ9LD1fZ7CNw4gOwufVlwDaxz
DIFlHxrPmFmO0I1Dj6B8S4cLog2gloNc09mXnkOLInAYZ5+in7XwfVguUvhPvrYn
sFXwQ6vd+LlTGc8Z+1nYvfFG0ydaS1L4LAe5nC4fQWnLYXIeProNgWsuCJ1lva5g
272XkaM+K96GlP7dNw3kprya5InN9wLYvYvGGQ0M7JmpODEclGbYMy1+zp82HX7g
7uogdCS1WTFuGuOYLm2gfDDDU0K392YKq1o9i04Ghlxi1nHxSwjZBb8QdAlU/ioM
KCvMnAhux9x24lfihWs2UPGCmZjIPf+J4rUbG0pUf8ebwgXF03amYY5evB/QgDEJ
QUKzBP6Qvpj4sqDrdXwzDY/7HHTg0lhSWqn/2L3nbFG6PvZWECfrVejMwFkP+HM4
dHNQE5a9iAxAcPjstxuoEzUWbgm4KCZmKDvxIv/73U3I5o96J2WsLNblTOVn04VK
lNpH5ozfL02Jj8BviM6CSM+g5ZipiFbYnqJPkbsqQsuf85KMtNnS0RXAgHQ1bS/e
gbS/w995BSZFKHB+Bi1+PfjdxxvXm3q7DQgP26ENnCcivMxp4g2L/b+kC3B5thq+
`protect end_protected