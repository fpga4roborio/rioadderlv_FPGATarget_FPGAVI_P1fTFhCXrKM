`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
ddtXksX2+yylW5zu6QL2Lhnb2d1sD00763mmSITNX595NcHTEkwn0zB1Dry37fOW
FufOhVzEJp80NC5qZ/+F0Vk7Ik02dIR0elf3clrjeJRK85K4e3Hoo4xn7YbFUIms
l/8VZSb14+JVGURjfswrIyCUotIzlzVYZ6gzoZwDXIi5gQIBf/gI+KxNXPaKV+PQ
Ufys/12rjO6aI/pPlqSm0hCvftmBcnezN2hk1UeXgOIuKZnogjOsf0iJVX2aOOWE
6pD/psybjbnsNB6kH5uFTA5frkzIzkzl5d9+YDm9OyC+k84E83I/7/j+rk4L2dah
QJOvksSIzN867/4Qt8qYTQ==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="MvBXkzurAa5VTw+1JJ70nePUfoQXBvZOku/SMmg4TwQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
oRtzZL4VJ4iwysPsC8SXYCzXS8Fw2gtZTOskLcDV+1B9Nzn1zTyNtlo6lNICRmmK
ZRVu2BmCc2G+fmzynYlNTnSa7C0Cuel6FYpxCBlOuk3OF2tzAmLAuDyOH3Z1Yjzk
a0aHuoCdIRKv7BrZCdALt03JeUmXKPdOmIlkVGFl8yw=
`protect rights_digest_method = "sha256"
`protect end_toolblock="Jn9CQpRhJt4rnzZPRk+dOpzAubz7omckX1MrFd4p81o="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 42512 )
`protect data_block
gD6l00tciPUa6pDNTk/+t0OO0nC/UTtBwLB41d4inuAUA3i/ALrNyoJVcBnAmEQW
ptbcNp5fxEUJjnOxnedyZEuEBxWRieZFQnkRdF269oOu6Msj9mJuFByYfWSDG3LP
esNKkUv13uA7CJnjn9HelUGop6yrXHD5zmdYRtY551ORZdek+ZZALJd6QgO6SBDe
ltC3MxSBpzZVWTK1M/1HPSL5HQDjfnZWJHnNewwKt+XgWCEhKZVggOVj522L+1CA
xNdcpJVlO1j9tm9kHYwsd66PqPTd4AMGxu8YlFyoXOPkNpqPEhFuFk+gyCkn5pRo
SkP6CTSHHpYM++6RdqLspxEFyG77jcOGIJsg3+RcBlHnP/gRobm/wIgM6ZMOevOj
3PA+nfq16bLc70b4BnCTiWjbiHeDrWi5pEki1bZebjZVrs99+/ha2Tie98eH8Lvl
zOpnZFg4acPlhsgqFTbQ9sQcYEzwUfdSdkdn/vY8YDweW9pxVtH7R4eViWq5UIzH
sWt1fd1aJMis7vWcLPDeUzGvZUbMNo9fuUqTfJXErNn57AtMjFq4/DudU7ZyQTKd
O6dTpa3gcSL6zNEVMADePqaEj8aXLAp2Uwe+LqFJvZaEtTe+8WNlTCFoZuCLX2L4
0SPct+aMwnQQWH0eUaP4yL2k4Hfuj8SoMoITqCM/eQBSVEH3ylvgMT2wR6DFnrnq
IzDQ/wXukUv9VJ4csDfA1JwL7+XJytILjcoJcAVgcuwxrY0YWzrGctS02BTjm8M4
FbdmNWnsz3keiNqeLRfRa+9wf41yhxoNZ8jCQEKtJO8edcqbfT47SUfCPOqiHKCe
d+0ZTvG4dqo/6RzDsvBECQrbU+FSm+s0j5p2QDtlCy/k/sO5FenQoWh7JglMbbvV
D6HQkMyM2kbZMtz2DVpRro3ad68TJCGkbTWApAjJ8bEuyL3IvOUDUig8WLTrvFAw
wNKf9v9mZolvsRWlCyksoWkqwzDFH2E5JshaZygIAk55goTe/f/DxI3+93mBtWUw
frVfEv+uJuXhbZeGxwVXqv489uuCq0F56hr5jz40rMpeHUa5Oc5J+mDKIkKI5O2g
DnUuFWopmIpivHt/kCOG6aAFHnrskM097LU22YAq28RrBfHVmmPZb5LNgRL0+KFz
Ag6xxlw8XZ/Bhhq9KgwZ/QlsyWIGq4IVt7dtc0nVKYdChIiBBFNRJx5uddYoyJGb
4MwCGw9Tn0QnYHemQXYfK/v6fRKutmywGHry+1kUsT1vOEiLgLQOnIfkmRraXQX3
/pTYF4ccU3WZ78VLBYUs92xKHZsFQVT0H92XGELK2rQSAHzC1O8pfQDO9Yhozy2d
XtUoiOqsVA4Lb9deV1oiP/sRUiqh4M2aBG9fXwISREb4wJf32s4p1Q1elug4ZnOg
2H261c1F1poKEz1nWpptkI9c2kgf1vWqxoOihG2eBegfkSPQAohbmdbMORvo4rOZ
jZOviOjXS8d/Tr2Khtn8sZz+sXYKFXJh+/W/zr3kCGAHl4ueU0CsLEjul7EkM7dI
7dvTH4k/SMcm8aNLB45JcfeFsCbG4D4g6e+nbWH2FO9utXxNSdq+SvE4roGDNPJ+
dZSpaDsYTcJUL/6vtdfkrxKLsNm3v/Si9hVl8eKBb0/a13liFnUveTnDC+KD+xFu
OlBZ38CtfAt/3AqU9Vi8y93rCIismCzcOUvXUKlELvADRcf6TeJ9zIniUCV8WLR0
6Hqey6pNtIRDSA09tJkE85oCzF5mNdkqka5NsrqBgdFTbNdJWT69cvHfG5COO6RW
cpsFN2KVBBwzU1m7vA2eUR8Rxpx2PDRnRVTqS0WWLmpMyeXBY4pBTywAk/Yjp4yS
HTeiUzjzBso1Etbs4NxFZAHkzeedpaijA4H0i4J2CRwzvWEmpsyCF+ZzqOJnkOM3
b9psEjLfGogPpTjJEdojtwWqXgDu6tZAyYmfy253/PTZAlIvAK1B7eQowHpPVAnL
wc3xn8sOuR8wXVdBPY6c8I89f6+l/3h4VgX2vL/38aX4e9MvaYBX197Y0tdYB08U
WZwBGv30I/VyakVAWDmzbbKIXvs1qFxU3WnZ+JgAv1pxGd6KsG7Wqxlfu6ghyD2Z
Nlyi02T0nnJ9LxLuTXRf/TzQE+gVlP2Afhro3T4S9ac2YYqNuADLD5FxhHFXE55S
cwCrWFcbGlwBz4/CEZ52Po/jUMDRR3ZLimAMQrCIxfegMsbiMml7x6VhZgi7v8u6
wyizhPDEQm1z6gh68Hi7K8vb+yq3/eU93VEXV5W7RsJrh83XyJ/Sr4I2GBy+qrxt
fuawgyr0C6j0fMgqx1f0WAWO7PzZdpgJS9wwkr7WTpNU6wfKTgvvsu6MGoIHPURT
E33HOifdZvlTAnoTud2fwKOZkvOhW6qbWq4qOOmq715Ml7HfOgaS0GDC8vmTAh3y
3LgCVAUfPzd8PTzhhEe8/XVgEQQu7aXF0K63l0JmKgobyKCv8w/s8dUnwHUAogkg
PSMfXPSXtcyD7XfcLcsmAPMW+bo0Vj7sak5e8IxlV6Dol9W6TFqpa9O3dBDoXJ84
0VD59naDF5y/OlMY7p+FLC4L9FWb38Do9bRXhmzVA2xVA+7uom4YeZCAFSOcXCM5
2benbQVF0Z6qBQYbD3pmhwHJe5pL/zYJHhbNqMqkf0ut1/tAuKy3utTeEaaJmagE
FZ7QDocqKfjUIoK2zAQJPchNyIfqq1dG/1JKn+c0ezQBAT/8adalaDtgH/0KX738
jyRp10mskohyY3vBoO+tIEU5q2tLQ8jy31MmE6YdpbDCGOSSVcroNu/4zSNi6lEb
E6oEWbubja6BSrxEHYDcir/stN9IehD5UOK2Ch15NsZdKtDDW5tuUDnu3WGXfDg1
lA0Wbem2EJYy7IUml5hyJ7g9SbDSaWm7+ZdwTfa82gdmbtAQ31tUlBkU1Kv9xnD1
LVcAGAOneY+3DkC9jN6eWgDCW7uR0jD24jdIHEwhfl8HuwG8BrnE0mOeT8koinQc
wRfn+cMhqBBRXw4Gng1t9Hqvk+SwVF5OUCrOIgxaDMv87HWywYj9Y4TDTb/yKtKd
p80tJyX6MgHzdosU3ZXnbyjmN2qwmykbygiG7H5S1WkDI6ssems8oJGH5BmDYbPi
digvKIBmPqB/XfvzmgZZaBMkLHnpIxIjV+oqfT0vi1yZJOwWP35/vu3D6PqKeFPF
Y7TXRuvxl+ewfISkN6mArVSaoqTQCbQvQ12gQihSfFos3FSpY3VBuFffVTyTSEgA
SpqdI436J+Mp2meEIzZ5NAns/x4GIR8iPadV7r1TESaSRsiiklIUZ5VeFCBtnwZr
JJ+k48JXTp9X7sdERJSy7rtUu5HLazFaZXZOciBwf7MeE5V9CqFIaZCjbBLlYeXF
ClDYB4hwzjJtVNLEB6mumoBv8xrYBcvfD+gkZ8BJshYj5nZlBNYOcnl0A8iny2oJ
cmUjhf/wmsAquzg2rrRbOREgvwbsrwVmRTFYJcJRhISNjq0l27BRvjggdG+FTN6B
c++4lyNFFbFSgMTLUJPlsvRdlaRYemX2syGN06MLa82mOPO+cKdLogG+YYf3oSza
8JBclp7b0yNMI++tSIp0CIPpS7qpatbj3TW3AaT77ZutuZyPWrhufsKT7mm/hf7W
8pzO3bo46k8oNmpuFJ1JvF6dkqYuggZsA+PXLTl4A5oiciNY4lWT9u2G89cfZ8mZ
A7z9fo2L4wtfuvMvaV9eujNhCZCoCCVl8dfcihCNU9ApzhQLJwUtcvtTMRS/RG9j
9yNxlQOm1X1dg2bGO3yEym0qJSjnAZg1sYUtsw7m5VUN0TTgJTGNDw6UcbgYAisA
QQBtnxka8MXFXXqqHWPkre0ytCRVvdW4E06AygOH56XQ2iRm4Iqk8EdoA8kNX4Mk
hMxdwLpw3RQjFnt4nTBDBaVS9JldajLUO0ipBgYy1aAJ/sm515hW8fdo2ajU/wkR
oFMwjs5Nw+fS8IYhkX2pcHjbBf3m5pCSLy6aP/R3WE9DT/hqK4osCUREeyVlefyF
CRYvNDc6hwV9hYaxssPksfaOr5ldTRnJY8c8Nwf5laq0Sp15OiB7CTRpmPAf3mAH
ZqLiSEiSVqR0Jt/kKppEgzdjO747JSYfbEKvxXcwls4tbhObiFFbHGt4AQU/ya56
qrbYo7Ytxa0O7IjXWLob7IxEuzeOJ/HkAioTqMTFmjQu7sQfYQ1nepbCbceLepyd
wjlEwsqLZbdi8aCn1Bg9rAebZM+aF52oPLbm+DK02JUDdjccuT9Q8KIWoWWeBJGE
LsViDMocCbTw0vAxCwOt/LfeWvkkQUEF2zPfNJGQUdMDAfKtCtfD/uPU2kE2BYGy
aKsFv/14786eVaYj04dNnLJsvZXDQTvuT+EghrZj9iGRgblO0zzXGrhZnF2N6YIG
eakysd4RRDsDqQmbZO2tMHEBcVCyt683ginTATXyK9goL7/8VRJIGvjLMBEOMZh7
sMwAGYkOrkO1uihAbqDRcj431P963aPv9oP4xWcHQ8uYlI0oefy+A/M8eVbaAKYc
9/x201zSPCoC+5nWRMVfw+l0aLv3pqS0jJMqBI3Pyy1i0yj9bd3tmBjixGreZKJT
mCbR4JcyZJHzwtkgQnJDiGn7vkA6m5LDRd5fFQnlFcN666os1iokfGO0CvM/0qys
Xaqj1nls+2vCOQECvyIOGMWN3R/Wex7kzqr29OEtFhqh7zUGhKPpRkcWYTMelNBC
zELRM1OgvjAIRaqJDu2GU0HETTEBvO63SQjJWJFN62ZoxAvBperGD+LfxHRowjkr
akCfEplzeN09JjI9v4I5g/WB2ZYLWhncah4a0gWVdRI0Qzh+xQIN25BwnTO4+W4F
MleAaG3byGjGSuHQO15CCOY/W7WaK9xYVNiLlssEzNlurkgaQGAxjRgPtOJiJUMN
atrqY6I8AFU6WgtKh8iFn7nh7optDj1kbWIkWAEcGpJqTkzDMYzr3qRTI5aUYzip
jkF0mQE9mwow8Iy7OGhi5t+NaKnbG7P97kMQhUTVWOcwFKKy+nLlGXfuX40OMv2X
itYWOF/7JK79NlOlmQzMqc+TpEwTHHpv95Qovu35DLlk0x7WXrsIvR+6U59ybHj7
dUpYMGbyNEJ3ij8xccrrM0FRkmjKFXB82e6OaQj45y41KA3UdmOnxVjHkip2Zyhf
Y7pNKxY5qsiQzyidgBzdpkr0yJ+ifDJNVset6rNhZf4jdUh2Fiy+tYdKexQGah5t
OaOhQGoZpMhHE96QOe8XcoszRI1NoA/Mor1nieunhw2QuOBGfXCvbGaUuIYKIFFG
CpcBJAECH7/HlZIUzMdGRJuIWx1Ly4agSc2/kWFalrsjP1zKLNjx/pVjsc+GwBs7
nQO4DvJekAWUyGsyoMZcsn5PLfwtfkjEgdA1FdEhWmOiPkHczqpGeSYpJetuCJWA
1r6aI/s2lj9IS+/HgRbM57ITX8gNo8GElGG41P9AHPVOEmfw0+sGyvKmH6it9xuH
EVIKMVMoHambH+pZ3ojiskuK4e5bz6WhC9lVhNi5j04JneffrG2E49gl3o5mkMAR
Va1MSv3fJ8Tek8RFz/ZXWJc8GUNOFSIAHWVrYhnEmrPrJnj2ujbsjNlc7Duc9O/g
WlLDrMbBzvdcCMHDv0SQH+LCjavIdyoQGEnXxW8tWPA7e9aW+m/OQJGRV1pHLBZF
EogOAhIGkDjffv8boXaq8iZH4aDkYuE6SCdrv7ECBeD8MzzDVgOMUL/8zM7x5GeU
1LVA3LKP6Yl55s5LaiFkUCLGheadZ33iE/OxO+obIrt5CJxhwC/vYzVSJpR+P4uh
uX1pMgiyfI4pNr7mrsa90TAL1vCSmckixNs47uUcqwKYrYvh/y6VX/jrB+doFKAe
h9d9/+iAyc/5phRBP962OwhzI8ee25S3mejZjpgXEB739WksduGdCVguZF4g7LQj
nV0hLc8wrvQk/M3ADkrOEqksdy3fCtKsTjkJ049CFUocyevKB3l9riWJOBpWzQSH
spAvK6gTpp/d0GRDlGOCfobqytCfWHQtCkGZIEoITMXwabNwmumF04Ztd+KfR0Cm
qbz3C416SUgT1zifw29sh6omHNHCIhinJe+rctWFvW1qymRB+eTiV5SDWG4uqK0u
4+Vr2Filfu4nvMyhCSSh6eiVLcF98Ng3GYbBXIwHRgpc9/JLBTvVnzBqxVTcfMVW
ABl3eZzPKfV7m3ddiCQbWFn5FyuezJ0MlXVePNmGGkNgNUfxcwpIRBnf4ebCreym
TM7cFmd+5RlYKUcdhi5FVhYO3DHvHcaJy3o9TjlufQqBCLwwAyQbSRO82Qj2JdcN
HF3t+XO/zZ+m8yCVqaVFjhs1F7NEo612K1yxnPMnJGjeSxv+QsvBmKnQoQd6YCDu
H+jYotJY4765nzqWyrj8v4idxNIoPqbZdv+MuzA+s/P3g8Zsh0xGwwaAblcOaEfG
JNjum2n8Lyk7+eP/snbAgU5/t3FIBSrz627mefn9Lc0mfKw+s8M7UhfhSl5UYjUH
73xyyj/rs2+ER0u27gzIKgsG5Z3kL3pc8vCicOl5ME9WUqqN0sBYSuS9DgU1Xygv
Vo/HnS+VED9KIKB0l+jDdx8XHw7Jlq64UVSp8Dk48iE3wVIxhwrRx1ujSFo83A5P
9IHG+zJB461TMcnQG0z5JmgNjUZ8eDQxLwS7gI+3rECEIECNQ7qUxRt7/M72xLmA
XioRRJ0dQHZLyt8Z+U6FxkBkGucRQ4acFfQLcuLiSw57lnGl+J9JYpSh1ekSFf4r
1yI3HbR3sYYUX1NYSpLYqOiU6DZFoMw9SRzk9mbS8i2sEDFRc1EiruG4LfhRxzgs
41E21buAG3NHV7MxPExodxLUYdC3ougR3Z5FAUgqXg+uSRqB/+deaNKVD1MTPiWr
MtwwqOXGKvH+olqtwO7h4KqYRe5ZhWy8b8xaD1m5J1MBO98aMKAyJiTBp8TGnptn
ETEWhs2Hv4A1Ym5C269fdi812mORswcFdkutG5qFx6lOMXpm1KS/6+nlGHqTomJq
cDrhPxLxcy4aAKka+ZfBpQUe+wzZHALEgVLEZHNuzJE+SrBZpySmQLuY8GHfLa6L
+uQCh046jv9pmETNLCAKF3Y9DqBbJiwuKrV/lqiQUmDFbxF5IVhDzfWnCmu9fpAo
cT/F/QHj0ymcIHLZIvQCQ13bdFvOcUPTCV+7y9+nomXYgBJU5Eibd4KkdnI7peh4
7YWYoqbg2KnzHiWwkgCybh59bHRhyoRgeA43+u2hZuSVEyuW4i8fdky5IG+793E5
tb2HrGmm+PrEbB8IYJVcHHOeUAoqzVjqM/IKExcUSdZs5BVVftZvZQVRR80sLEye
07uyJZ71zeXOCsvFlVQi6hJo2SNgE4+fhspbEMk9EjoOy4m7631EP6wCJsX4ZAua
/1rK3BfiwXjYBxNcTHyT1oulCtL9allkagYJX9emN1Ua7iMLkjkADgLVLn1XtVk0
mTZxo4suA3VfGJ7xEZFa33w4mbsf7czN8lLKFFaeiLHS6mtJqSJ3PHD0xJVNYJsc
qEp8NwsKJPF83/kywar76Kl/KgjTdj2pCyhGwdo4BuPQsjAUo0ZxHw6kPSlbjdop
uc5uRcZwmqzeSVR9cXBXcUxaC5zA4c+tJE51npB1ivW+wX7lNik3FynIITE5VNBh
FYvEzFDeFh78PS7xN+hLw1aVWkGcA3mCFiKVk/tgJu5C6pRKKXeg3pqJXpH/YrsC
mWhvMMMIlx9hz6Iotc4/lt2itxH/0Bjggap6U5e7hkAxkEGq1wr1JenvepouYYR+
1Da5RvgSlNvQ8o1q4WrLh4NHpLMDkJAs0CPXaj0WeibBERtF1C7aRKO3YKwyTaS5
3IV6yCrYln5PI+S2WhGIHsj/0Corvo5830Hiu6DLEUMJnLmlNs1z6vT6lNe1FZ26
u7QoSyB8FSIg86wLr++j6cdCVwm5lV+uUlu0Kz6sPreLqj9tvbJlvBU/eGtKKA62
9mhi21ZSY9vfqmRz4+hWaqS0VQiSiu1NEjYcVFVpVutvy/Pxrx6SPoC+dtfNawj8
ePWGqYOBMMTLyxefTMIK2895rCs6G1yLpLHtMb1jEeGFJWG7CsFQTh55nLHbPwnS
kToyisZn/Pjp9tE/62mt5y0BpBsQMW9ADMNfVcOHzkFXFDnU09Izxql8wB+PZTke
ENXxrQWpC+sUTOxyYsD09MyCZb7AHjDCCuXQS3gMZhp3gWLrxIt/QA2e98ub+M97
pIPl7nLCPGFSR6edEB10TuTWgrDKqlQYiFqrG0v9q/x5DPtvevpHeGTSBn2B2Z7L
mlXp/qlvZSoTt32+q6XI7B9LFP501T2SLZSgMCAsTDoz0y+qFBYmLfkl2E5mGfeZ
njHxnEsOuqdbZ/Drz//4Xa+NMV2nWs0/+FTUO2nGh971SGJmpyoz9raPjcIJWK58
f4KjQPdd9cpcQqczxcHRdSvpIghDijcp0ZuUQxOrTPS/cY4LHYggbK8e6Q50ifyu
O+FpOStvCghpjiwJusT4XJEW80BeUlERuX36N1A8jNJzUukaSGCaPidnxR0fqiv/
NgliY5K27VdNLx8WClCMZvWFtzPwqWR2gKgBAaJh3jPggvQ7Ao/SKOB82LYrJY4h
sX4VWFhKDzQsDzXox37yxCU+mB0pVYeda1PYLqdi1oHlo4P9/uICDVnz3vi7iU0M
JaCEMbuqfcm4qO5wTHlwcB+1xvhHWCt2yZn7WEgzNCdqFxhUmRIOs7oO7XD8dIaF
eCK6X/XWuFRBBhEPEsvN81mz+aE83Vgr0V9jYdjONykLBiaWOB9+yNWLn0T6u7VV
y4jzSdE8aAQqLDUPj4CNhLffW5rVzlnsnm3emp6KDxppcIUdvwKZop8VO0mrsqjW
HxQ3k7q07F0K9CGzHEl+fMNtbbxKTffqrMQctVZpDbBmfyS+rE+oOsiq15TnIN0J
kjwvBZE5cNfoRWSykbUJwb/slG4g55BppK1OSk7iUaXewY7Wncx+BnK72Zu6W6U8
y+hgJA909xRFtLUiL9yCyIDU7W78QuKQ8yzadNFan6xS0Qg1+Zf8m5sbl2y2tn/G
uxszZETYNMGh5aa8MXs92S1Z9n9BK3aDzxfgcWEVxrep+G6lW20gWXmPfrF5brer
iO5KFXFNIxjLDhXpv2KoUyJLzg07JVpIbegbsWSnSW09PJ4D80sSH9m2BpoXVtZ/
WNw9/SXF/7DuYqB7WkoKyF3Dwr4k4RCIpfGDHvbCN89ovU0MtY9vzg0pUupbd4mF
8ga8+/CPB1wIuNlUnCgoja++/3ifgWcV/zXvjn3ae3gHqEfEQT0sBnsQAuRJ/bjH
VGk+zIxBHYdAwuYDkR2nRg4Xprus3aUIUO6O9YMi48xDbcKMHlHgsurssCIkakn9
llxpQyx50IzmohCnHiWvTG+5zGH8KFa6biVttRhIN5Ka0++sMDVdkG9JaR+lp5cf
Na2+uRegQ09AAOhdylGh57GvkPfRtaAv/bhorlBsY+3STAACRgekQtjiyoCx/QzW
L7GM/dojW2mNzPUKyTSUbrM7OvokAPexzfA1lgfTYzoOdFkiRdu96WwZLbGu7P29
Tj5zf4Z9Z3FOY6kJlAl+IeoREggQ1yUQ34fI9BfVYGRlBu01YJ8HIYcOKCuSbNAZ
TfaRopQSOyt7ZTD6Hg+xfdBowaTmrr3Q+aFqGbW95ZUtOFuqvwTW2zH4/ZqO2M+H
Ly+N5moA4FjhlZ25YF528uMk4C5hJG/ER/TNlKLdn7S5ygUSLajEbe/n5ZBI9ZS2
ynckihy6wjMeD90thUAujyhfvZiSe8obPHVVOl32LLjGrvZJ941OX5X1pGMCBaJy
42ftvfok3/PWuv2xn0tbU1+nP8i0aQyhxckdheFK58iPW5QJKZTKSOv9R0WU1Tw0
YA+mpGI6r6NovlSELmYLOJNjlNqDhh0NCAB442xP5/3f0O/kTt2FKNdYi4Xzv6xT
b4ibSqxtpdw8yFpBPwDfwsTNjTiuI8dAJRZXK37xmHpoEHJthEvkwwjjmw8QQjCl
x6iGXU0JJ0vwgQ9JpNznt53lCRj4NfdphzkMCcq+INCFuVXzlm362eN+FJmgf6Qt
0X9CXiRdqhtlonpxDb5HXbpDmzp2VLh/31Uvjy5kddKydgf1UqqphtVBVzCAz3Xz
NZ2lluMg05DsSZ32mYuzOKvSoHzd5YPMZf+/tyB87oV96Metfff85jFFPrCl7GN0
RFx+nBHAc5SsKewwCyuENjv4vY7tLhvPPR2szQQWAbWCVw0kRXe+IHvSXyTS1cgH
Ugy7J786NW0O+dXTr7uD7e6B+KYdKnWXDVG8obJWUByVgGVmPyFldGvoZI/SnWRA
5DcfQXujYYQwdGlT6ZNzs6x3qQKwAPZkEoTJbBlPaMfNxi6i2adewWvX+pOyejlj
tvmcpjPgFA6VHpLtLBdQ8SuYMz5bSQsToW25haJ7sSIaJ5KmhjjLOPNVnBHdsr9Y
rqrAncoc36E2XB4oQP6wvkLEvBE1go6PnIAtWbz9xdPgx/ZoO8GHYE4HSqbTGYj1
FEHENR5QfzKDxf0AC2gBEHujkrE5d9gu9OFoZqDrWr8EVMmkEq+ZceJ8DpinHKTQ
Hz/UqU/gkoNuV3RxUPHHbfGTaZHPR2wZkqElR5NYbn2Vw6ndEjf5Ym16KHh00Q5I
djZvyk9qTOe/dxNiNr+A+s6kNS9lPakP75uKVm/MC2AjLyDuqk942kjpv7gHvfjF
F3ZNttLLVMiqNSsMG5Moqri83CzssNqtUrekvanKvmoCB2QRa2OitNXwYYzTqQXN
X5WqFvzqB0+GiqjEaDycXQa6hLfxN2mOk5zIGniYey2muZTSAewbJ0bNshopMLGk
vHgwdgbCTwdJ8rwX/LAL6te2iWJSoQD+MH81E/m8kfy11lNNOq4Ywdnmp1I8iixB
1FyW1sRZK2pHFF/JO88bf/1F4p6cSqn7LuhuiIk3ENuFtmqC/24K1FtCuBBWoB0r
puTHNFJSK6iys2z+xIs9ttFFYHGRyD5fpuYEHVICfmalN9SaOpzVo6GX7jBCjnOL
sycf6rxNBiAcoiGyJngLTIBgGyPdkT2ehONaN8uEfdXYhm3HHOt5BPy4xisry0o3
OQRUFEurpylYNMhe+0Lb6mwPAJy1oQ9V+o3hqlX1nUetTe59FVlSPovCjArdBxMn
K2/z8YqBfS/zQgb1fzxpaF3biWp9+9YMdPESTy4N4sISw5WNUwetfxkUVhrGUcyL
wUrq0ElViwL/GrbuJ6qFOcU7WksQ8HvesdkZ+yTl+v0PFkk5V/QFRvTdk25BCllr
UMPj3k6OKMAgX9KG2cauFazu5GGOvXBWJSmWIKbtqJFDQbpQRXRfiC0e2trkVXmn
F+sgbWsobkVqDO2mgjgDM7hKqfJ9W0GBhqLyNG8ZrD1p+dKGr7Zb4bGXb9XWUV3P
k2N4QkeEeaiVHGMDOT5DRF50cDmk+Y4FSWPqr2p3iSGraLDBfqni13+ofcem48L2
lzNpLFyf3nw3DaFqcPuKY7w8/WI9iq4/p8PxrtjNk4H4G7BO5sQbsbv0k90Ef4FZ
zIkcO6Zy81cXRJBFfWcjwmf6C6k+37hKwSxKEdtjSGp7+G293XM7ax6lYwRceUlH
nK/KvMu7rLK2HqToudjw4zpjbjsdNUCljI15ccjQb4Gxsvwu6OqXP7q5TGC8hbbu
uwJZp/XHpR7h6MqAfx2/CRaT/AEzEaShFo2LjjvdAjwsmzax70ktXUpyaRvBqhNR
kMlvI2003FWI2F4yP2Tbdt5kzVNbjOxOxd/v+4woPpY6Xb482X/xL38ASPieHRli
jq7OTUc4yvqznASTr4ptOx5tBNBKQH7Ztcm5CDwrw3vAkU2mdQsehdixfm5+xHAd
MlMWZ0DX0kp/m7X56c2wZ/QNsZG3qlsX63NA3IPa+FS7cjfvcPsulzJItFXciSxP
gs0Iw++HBq4n2QBJeXkNH0g+LfpNWlctU7LyfO8FfjIa2eYdVgbfLojqa2d4BOx1
fEjX8ystLEl01g5JgMI5vVYBaTO0fgU3lTbt89ffiPq5KKGLu56yCUzwEA1P+Gxj
O8lX5gI+ccM1wcs4RQ+B5/6Ju3m9aGL6ynnRPWqW/IUoS99yOOWqjmf8bKu1bZwS
xaOZVqO3zo8Dn7OEnM2+bHLlFFZo2AKlaiEoRPoUE6W/siChjHvvLhUqFn7Q8rqj
9U2+I8YSsfGUQgLqImiC/yX1UoeH1d5R/x0Lx/jEv3rpMGrh7blIw8wWuJa2OWKa
tDHcBmsHelWnZE12al28K5SnB/1jONE7femzrJPQ7jqoDrjvfg8IygK++3LGrxVe
GhO543MkWDrhd+Ro8qLgewWMNeMX8fO7EMsCDpa2PvVuPYspl416gdPnGxyPFKCh
ZxlAwJl9vkPjHEyFECN6OcLnreBLETsfiee0JpM6DtWJg7xSl0IGWBCIIGp+gjud
iDQNq0rj2NBqzTsU2jOThw8erxLTKeuKlOfT7qWQzib4t5hoz8uVHEy+bzYn8OPP
cUkf2x6vLnz4kDTkcBJK3oJy576SjbZK8Bsx2eSw6Y3FUEogMYZl5CpL/KL7mi5N
sxePiH02NwIjdg3b/gVoNR21TT2tjQHMlsinHWKV8qbtx0iOVTSfNFCo14Y2pbb9
/jyO/iFHsn8otoGi/JNTUxo2T89OnQ4iSlMTnRtAeNgZHPRfsMlPNosRw6ZQNS78
loVnAifu87d0cmfbQOOmCr6T8yFCC0M8iWcYOmbQ3q/5Hefxdt0UZAsps42TfCyN
G1W51sCCy0AQH9ZieTPrKqrvoYkcIRB+magyZ9qDxD+mW0xEsPTUyx8LGAupKDKR
2JuKxIVuKeRWIRt0TujLFHjJgdYEZQoK/btODtBpdLPeuOpZCupRP5U+M6nThk0u
5SnK378Fc0Z14AGQmJzfFi+7zZGjamB6utBVsweGNXt/sf10JlzlGlYJgxg1ces4
gTvvUsUmuaiNNEZ2lWevdhRJiXxfu3bBV5cftFjx9q+wi2dL8yxkhViLmgCxrrJ6
tM6wOEIWwVnOXIxFMkD7QppmBRis90xMP+siCUgvgMpPILSVO/hvZwsDcJJcWEA3
Oax8kQ9Vxuxw0CiaAbPlNe3UOukRLds8gX/b5BWyU0w2QHkf+6AaADF9fHmD12Ye
hARgN+ruoCF8q5QRBjIJF8uDvd4f90X4HqqTJSxCd2pYufzKQpnMoAqf3ziMSD0i
r4AU0DAzMXcrAfc/jJlW51eTYiH8lThzuI7F7eHqClcZiiqrd6Q0md00FApf255K
yU+2ofXOVCacsb3aJgxkI9le/Wlcb44hevSq9IfFaG/JcDmyUxr4VSIEgN9hbTUL
zaUnq03ywbkzPWXlfTTpjZ9qc/3KZzk6hf2KaPNNFJdm1Kzz5xxYqW6ihgl9mv+j
MczZhLOlllQ4koV8M/dUVSGBk45e4P6EC9j2YHt2xjq/8JI76N7QlWggEA971BHd
6ZFfiSweBwQ28oj3AFNIp7+VWZFSt7yyhCEJS3aQH0xJzSYBbjdD4Bp/GNwFA1IM
krHNUmR1xdaA5QFEOdSFYXSb4Zz3TRhVpId3keWePWm1328o9pj9+HBVMOShznQJ
vFhode3iQovee5w+YFFCOBArncj9Ko/Wh30/IPBpF7whfokTx1pKcBFMBgxvio2k
CGGavlaKuu6VnJi0kXmxWd5zHQGtWMfUrbmJDyp/2B9GQ2/9QD2evF1kg5BA02lT
SwIXh8y3lFFqteZLVQ7CV6VNByKr41VbqPfFB72RxNpwd5aR8IXmaDDhSW57gKht
bS/0SgtOTp3gvYzA2JofumAdscrhCyrFGwhW2wEnaH0JtE0dX+wEEeQVS1bR0xuJ
NObz1h54Kq8YMhkOd3heM7Fh2PHt21T2dzJT8xtKDd8QAMOaNjkp0xwj0O3+qLTp
y7xs4EU1Uos5T7LCcmSvYCXyftSzt/JSv5iYVAJxZV9RjbhbWi2ek1ZFGSVDa07P
hXBCSJRqGldcsinYvmhRkLnYqqhQz8JE59WtrAp3jcUx2hyB/uaQjp1WescGVhSf
vhRIm0400OS7YJdSGEdaNn1MB8fYvYbQExVcj8W2CGoS+QQxdSLzkOJW2QvSD+EA
IQRJQk4k2p6HgWDKlqLFV70oTYYf9HwRqlTLHJijBcUUHK2r3z6oW/iA1jeJhl+i
xAkGW5Ql+CegyKgqdIiwMQqRtq0i2GKAjyPD5ivGnxyXBKe2L9/gZVoP1l7tZv9C
bNnCFLOD/VrKRIaWiCOs4uNLs+qrDoFXg78rVsBHLhsVPf5wSlv3Jk4EU5yPlFnK
QWpi0hN6t0ESCcEL2AjS1wcx0VcGZu3DzpjvHOQENht1ZHVRXV2caBlOZPrO2HnR
lmhhjbiowOpMkJwmor41lbioGC1RI0JWEDyWPenlf7LXsvF1kg0cMHocCA0X4qnQ
bp17bnIzXOb7nHAiix/Bc8sXgY3O9DqT4vkv29cru2ohno/ocntCPyRxQTj+4P/7
68cbmIiHpiDkinkmV9MA0zkfR2AyUODKPqXKxgIU3D5HvnxBaDNz+1jEXCzjESmi
cNMlAGlnbvsCFU7+f2/8fEwEqGuTapSsCHV+xwOhj3D1Iu4Jt63Ov5GHZWdfOnhN
4u8xJjA5DW39epRYz4va3Vg2FXksE0EJU4KGU4tM1x99ofTf7iX2SpNgdAHzUgc9
usZWeozUQK1POKXnb6w3M7O5Fs9TJOgqZ21GlteueRjJ5V5agQYSc9pmOHJS6gtR
3HFAZM+rpaXcQz5CDFZfvZUTnPzpHC3NgAOSzSfQuTTuFqEuQuYfzOHjveg3UUkv
iWCJT14gSCJnZFf+NiZ2CM8NW7PO6PwRfrjO0fBxbWXB9geSNTf5O2vGkoknauhw
4sceBBAeJQ1byJutkkOl6uUWOvZPy2rP4pNs90AzqoQfBhD0qudDdUvBiBpKhddQ
dWtAxtXlRmA7FL6oMITuVJ6Regw1Egj3HliymgL/LHr+A9xC2ZhfytIiJHYNb1Bb
Rvuv8Af2vVMRE/MNjJvjKJfuRt2SJUzQ8Ab/czNEy7mTmSrKlfGKZP4kbg5TTFax
4q6PoX/CzRUnnYnaq8CnD+I42kFVxywxaM0deVD0vntjqS2JOflc2AMc7/joWdB6
Wm6PvOYIQJe06G8EIIAa1Gfrrt+rCZHvzUZ/eBp9xADiBBOkp52u6+YRsMV5YFYt
NjrJhY535yRdZP/0UzuBRz9dwAliTXul5Z4y0HEpRjLaKSkJo4kFKt+atE4XB1jV
KMX2mSUqnZk21Z0HDsQaM/Z0EKKkgWbUnxOFSO23w0O6z6yOCgmhdDstuF41+pxk
0g0JvdrHNZY6oRKYoCxfiXYKlGAEQfld8byGHUGmH1wHy58XZIJZKCCJ9800yylR
SCu9ElKJTV5YE2XoIeni8XstzvMhBxsVrdVnb34zswWJdDr77+5zk31sgIBr5mnp
4w0JfnC6xi6p4KLPASt+XOXmjZzyBzs9MKqQvbW76tfT2z2dlWj/086WVJbF/Yh2
3Pyy3Sxue85jKF/YW/tgm1SzL7CzMzNU2cr4K+njoPA+wG6MB9LddefXmVni3cvU
RUS+XcH0T+Pp9DE2/rtvWM8fmxfh9ZRXqlGG2zlEG7SDwm4TfUWf7ryk22Dmub6S
/kewHvW7kG3D5taiHh5d/6h6m1dgfuAphusUuybEf96EYjAMGfZe3XBizozyOrEV
A+J1JGU9F5lWOvDrew890cmlBqmQ0e8rxlcqlryl98TkZxgJlTtQj7l+1VwY9wdB
CD1KjG4g9wN2+gwhNtEHXyTXzpCW5ktewKcH/vYmXiOdrEHbzK24Xgje3pU8Cjyp
jSYiDVAyrvLTlGsyodwKW7LO7WSM9wskowOV2qEJ4ISN6i00ULyi0A45qdyYDW6g
QmIQLba9dh2+vOeJ9DJ6IuBGy0HJ39XEzMI2IM1Yn1SqSfhgF+eQh07wUKM+LeIq
8MGMUWIuQV8602Ij74lAwkfcdzXCovoJqim0ieZnADvzzXdWokT2THV5e2/TuRrZ
E8mPszHedLw27RCD2k/CT54Dq9BLiTHRgTXw4nL9fY3tBixuYAyi96KSltNA6yzd
lzQBf7WmrD8LDO6XQjr32OlanaptNgMsBcyLjbzT2NrGZutDzHUF/m50MlaoAhD5
bxRHMAMeOGobPDEg/27UNV1JcpsVQ3AP+4I0r6BOcHa+6KsxlRop4P/N5tnEq8l8
QhqX2Pp19EP7tQsMnTdtLB/1aeKl2tgGoy7GdsPD4lfuTfsmbFDQzTe1Mqhd/oTK
yI2cfERmzY/IbZRgd3zifCMFymMpd2yZJPFuNUs5pe9amTxT6GdpjSvQrrUFIL6x
B7bva/IRSeUEeyRNY4R2S+R1HrLyEGlIuzGEoo5cGJEhPzH/63hLD6R1qvEW/F5C
h/h2chfL9/2CT1Kge4nu8QQEvCLiY/i67qAJ9+xnYZ8z90+JPhmOnr3nxxTXazZt
KAXYi59YcBCBSKuif8BACIhrSLKrHtqLsP8jwudQGjj+YMrgtfkduLRYPMAQBCbh
5JBkBW1U107Kw7JzDG2+xwBkvfWBgfY9Rkpbyqx2zzFH0Nm5Cm/DqXGFV0Sc2CU2
D19+/ENdef7/aE7DQGT0LuFP1kv3zfvG1sO2KbpYkvyP+11FQJ5JN0sCzMQgO76q
9mcyYRBZifMgW/GHOxWevpC6CaUbUk2L1Mnt9JqOhkIbPXqM9l37JXcAUT1YXrHb
qrEz14BNDLYTDcqYEpg7ArM0JZscBkiPUsPundEDXcewkTqdaHXl+QJf5XGLlKFt
8pM8Ozqob/2hIRku8PFzyL3kxYTYUGFaQvtIcZzTeYRYFm5D2ij7Qvag6VcVSN3K
kmev16qPWk+aEohpWtzJsX9YbsrfSD21YgfTIwm50pljtMxJQE1ottx6LdXkp9r3
hdoFDAoTRByYCDbnMeCrDuc2r4kdu1YtHoIpaP2IfOn6XldIhlgWL9PuWlnGCRy0
QKlhs1kgm653fA8n627EZr0DSw7i6IGSbtjh+20Eju0cAM6TEP3Q15WoQr+R9RV6
xhccUn7tt4gbovhbWtSVho19TUCC8msXn8SFT9tOSzSlO/BxOrqWvPXz9q+0vBBe
H53BqURb6oX2s8HUo5NFNSVg+WzGzvaQ2dQcaOybPHv74grNDHFUlxzFcF+SNJZU
/Bt7Qg6Zdg/fSO5utUZA3+H2ol36lwwob2JDBxxJpvEDMQIJwqLgk9sUAODkmCMK
ycOqmmLzbT8g0io7ykiBveRFmnm5z0HJW8nmaVjgFK7oFL5aFDbRL7y6nx1IgLgD
9soReE1eEOanxEvpzI0KX9TKhG8rZ2rbw8t3hYMxFqqxAsRgGyzFshjVZ6cKJDnp
wzpi36Ym/uyd9H8LOdHHOUJZPJMf5gYX+McsPPSvuQX1iTWpBup13a4N1S6H1jPr
P55TlzmgQ+28vCMtnIkO0yleu1xDmhJJAMDhDc3XYWwmhTg8dUoOyDESivyBLnSv
upc6bsMaD0ugWGKpG4J1tXZD9S39CQZZH1Fx00oADUWqGvUnQYTfeFJhbXx8cKbR
jIA5xgDiKyldrOjfkOpnLuZN9Btw+oqEvzclrsSMkohrub2gzUSBv2NNvYDzUF0p
sjpKDWmg7pJ0OGGw7IuHb7kKXmI5ihKkCF75/MkFSyHm2Rzxwto9gXiPzFy4hnAV
rR1fqFOB88mWnbuYvfB95sY5k7C+2HxhXrYcpaeYuzQc9jQnntbm8FJsQG5XwQ4W
N5+PTtI5H2gOoAY3YvUve65QdCOGLSnUpSuU+eiepxGhTjbX6qPKFxkpVIdxZ5pM
3Ku4CJ4xh4W4Eu4ll7/OEhIDaEbqdUpbdM56+UkA4E8ZUQYydAVYHnl1Ml79sXIa
LwoODWJCtaAdE4eXUno2IohdNSmANi2lH5x/XogmhSRHykPFx2EiV9iJGlIPXzJb
MS07xgux5zeFtwNCGzbwcSq8y/IvqS5hdmzOoy+9LdsJhmzrHAb3oziNmVXu+dtz
bkBrUdnCFA3q+Twj+x/C942OWiTRE94rMVQD19ycbQzqZOCIWcuJgzqso+2858e7
aYqBwkWGGb65mXakO93hF2wK6QHv91Y5RODZsGIGcEfLpViD2chZ2FvgxdXUwkcP
dCQnxUJzWb1bXL8PEcXZLPU2x/nWVOrJHNFDKKas/Hfh+bYnM1vYbPYckomzjtLO
ufLVhIiaQlm1hiuFsfIaeOF22Qsd/ArJPwSuZmbojf/jgKqGOlNVxG/rEMTroxCu
BDXw4scpemoGn55Pr8f3oXEelIfvEQTwpzTXc5QFgvf4EctG6xhCt60epo9nIKkO
LuAkN/7t+5ZxYNGwaAi10tPk66Dr0Cj78U5aXYNWWG9KhaMp/2qlBX8f6kxuOWTi
1iTwz/XaVSSZJR9DkGHq6yzgn/p5lDTBNbTwHnn6kZ+hEbjK4E1UFyA1f69Sb9On
6Tf065LZ6hwQjYE4RXALV2ShEFGdnUxKdtY3/U4Lwhgbdu6vmPIhiM7QRkzIb2mR
5nCRhGJNJ3kvk4OFVj6I5tTsCaDgYuC05DPHzQKCZRIWcLHdXL4QbT4RO42gE2tR
LXM+Khf3I1tXMU7kCkuG3Ee0+UazoGCvKK3DO7vCepW6CDmXUQ8iP9uSfxosU4jy
+q9znYqbUldfXRdx0EVDlE0y9OwmgyQPWShwdXqtDVPMp7KbosoCla7ioWlIaDnK
ApJAtUthhFf1IA1nV12QK3RDwwizcw0wTZ/dvb2mI4g/O712++fDNDMs377lcxa9
kfHTMPMpnzM0NM5FhAeGl+NUX0bunwVd7TmUp1PdnJ36neuliw92kzQt0xrxF7ZD
PQmUhptOegIuqXWr/eSlRQj/WpCiZA092dWR3iBvzMrxOrIT5oJxI5wquspUk01R
xbJ/q4dtSOFl2y2OYS807ZCTj0a25XnzPopyZA6xvs3IGLfkgjOCld7jqmL+TqmF
Fb63zNSgLDdnSWj4nLuH9QvU97dXwoEI2zKfdr1icdGyiuYXa8UfsPdBj8NfMxJm
Rwj38543nvmYXiP4kLb4Uz70q/hMIvysVH6VPirmBPn4laqN0FomE6sPCsYqLVqM
feJXjpUAh+bkn5CdLUZqlqoMsqVkAqFDRliPV7IEspuPfUB+6g8OeMP+dl8kAup5
ajYYrjKjGIWh1MwJv8LkEOyfvH6u52NOc85vBnfBV4VWphh0LAKiS43wJhln2DwD
pgszkw+swO6ZxsFRxdrNDQJ3q5l5aSO5Zc0HllPo+8mc7+EaqZtDF3Ld6MpnQeEO
oiS9yb+SKLi+Z6E4g1LZQCkL9uJEEMUr9euhPFNjzTRgO33VB7ljyFc7rrlubLk+
fuqUy80d+bXbnfAQwUg1ZtisW1ToP27jq5dY5MQa7G8kjhdaJ5jIyD5aRbeClf+n
VJkD3kJjRfaxM0rBPiTtnNIJXQmtPGS/wOUNNHvGWS6LZ47xCLSNvs6IoRntwseR
xjXPbbAq/7LtB05YmHqR8Fvtd38UzyDCfRcVj9MmtpjL1sCuRY0qHLImK7mIxTUS
bk7Coo/xaLcvNwwaehsD9K3WHblJSaF9aJzd64BLpiCys9iHbDJ6IJgioiEYy4LF
dV1wPU02TnTz2Ziwjm6c7vmI5OdWhtHZ0YUjwQ5BJiH0Cvojvowf8afmmXhHP5NV
3zAxnS3dHag4MUIoEdnQ7NqMDY+mfCDkh6SrSbINHC8vILubPTxnak5cVRbqg95/
C/alNfD+ZVsA+Y/5xN+3oaYP9LKd3RbeeDCf5J6cGFANw+bp7t3NfWdyaphh7yLG
+MbipJXGEIJIgy2t3u9gbsPEWJgMSbUm4KEWoCiknMw9MkYlZnC3g5CWvzn7PVWY
vZbwnp17nFzuLKrDhrNhpsxf1+R4ucwDHAHhC82Kr+HzpaSdJS4zy9od9+uVXtzA
hM6W5PYp27GjTy2fpqeSF+nuFalrkdG2H0A8aLTBNc0FJ5/ckm0RJ8Xu6snOoAnq
+/V1QXoHGw+IEZkXy1lYWAVD68F1d3VIQJZRAqIky/lKeKvcdWNs/XR77zjANwZp
UAgbJSrjZYlpeY8gHMGmy6bXh34o4nq/dSU6GoPkdxbBs7dZKmd+eQb11Ln0LZP/
2YNF3I6uheQGehiAlpMNE35av0HzyhAjp8ngmE2vJAxr7p1CYM5inBvZTZiT8agy
Jf3humeJPaDYnDaBNDKDTe/TdecN1JXWRHxZZH5/ud+T3FF6u+xn9CVB37sgWzyt
iIrr1GJlBYmHILsOX67Al3GlqGYQ+Bs15PhC30ojz8w7ecYlb1O31bDGjRR+6syP
uGDT+E0iz66RBBFlmKggJvtJko9NfgiphV0/9y+Cd1WYZSshvt1aO9gBbPmfnkEM
6TWr/orXXZzrLTcgoJcQsx3IyXPdBEvAZwpmfwuyD3CKt6RaL7HQ59dYDddohQLb
ZwaONmxudT5i9rRaHPaXZ7F8lKzZR4Z4u47qlH5PMF/CH3R8i1jhXeRI/Y0H+pF4
SrefRR2HBtH1r/4whvf3ONbWwuM32J2Q3/Wmn0fGtMQHXnxadHC6NzanLt2As8AH
y5YSmNz0z3cxck4cGKuF4bZ67L5+77W1RzKt3asBVNXWDvmtoAAHKZ2/+k6rTbv2
nqVf4YSyiX6wQMgmL1jDC5p0L+HSuY0iHoCqMBMSkfAg6V54SLqV7dlpPGgCmf/L
Tb/Gu8M7KtnemhZ68izQ2/SPQWluMUpIwjvCZG6SxQMes8XuktIoO3IARDcdzYql
SsrEbTcnju+nE55szKBgAOqi9s3QxVEQhzOWS4GLt/8A13Z1uTxek0b/Y5plkS2v
sSfwNKnNAS/Gj3ymTf7oKL2UN7Awa9zOJlShDuOtHnZCf/Jv8mpnjd6hWQ1a7cUi
nEo455B6B/+OzmNheS8IFc4D8/Blr9r7fZ2mL2l9cbvXWCv2fFnRa8dQpradJGJG
sZs2D7gAG4nvjvVT6ThAD0e3oUuU448Kn8veKYyd/rtnJzNXIQxoQ9r+lt39JTqI
9dgrl38DWCCkUucsIzVOJ0ga+6AU5HhvdHc2iLSYM/uQLi5w7ThMyIOSPjm9ZD04
ctQrwm+QajZz8HyuQR/0sq7pP2qFmdOl6WMj+zVH6QQYZDELkNtFvE2eLjPxl6fd
FEwhP0YFNa1K0J3j09QxOQ72vI+lt7eg48XJ9Zgmj7+T5IHsKk88ohy54KmVtnQr
mmI80n8aTgDU5rEYkc3EOwnO4pQDy8jhSOgE4L95a4O0ifc9dXOo4/RnxJYC5EYq
BEkAQTOWxbbMs3Gyy1FO4oz9zcUbTzgS826NkfCFGGtoh+SA+Q+QXD6wZA91MN6c
G2GPJbm3VLPGdQiRxmcPiPss0pxxZ9ExAgZsRsWGVUbcFXQS8TZBee/jopzdQ2X/
K8QYGIcsc/yrWVl6GT2N6CPIfrjB3tzfQyWFa9YaN0UY+rAz7T43+MU6Y9RndDdG
+YWcAiCaLEQi/uTF5UIwLS8ft3vE7BQA8l/+UpzCPKidgPIi2hIZgTeO5+uG6TU5
MdBywTge0qzaXLHbIvloXIAU1y5uiEnxHmV15rLtSlcCP9qkpwE2BtoOkCMOTvBe
xkfe0S6On4X1BJDfnqg1oOlTs6JGM4pnUpdNvXDatrwbWJWDsKPumGkTQ7tKdCK6
IonNhDRcf5AQEWUi78FjcibKcSfHxQIxpzWwPN2lM8MJwRGAzlQpyflF863M5YhQ
jZWbCL8vlfZIJLhMfQCuwRuetLeBMQgVkmaooTxjDB7VcLm32iacu/TW5v4lb/zz
9vH3NOVyAWqWzDM5erGxnXB0djKMWwCvlVB8/MHOxy6ERB9jrSucOzB+1PVoWhzH
JTZ/x0tGQL0/cFgzMMGeWU1iVX5DCGbKYf9ZgS6LP4B/fqYwY4oJIQRJF1asIxAy
Vb1+ENYDiQan5u9AebCPWItBOGpslN5ut7bjJukoadA8olO5iCgfyzbWnsXBOyft
wuhyC1INq6U4X4i5XoZPNSuxqqsrHZkxt3AADqbko7pXj7WPclVIVFY4z5ZFMPFa
WpFR9GsdS3Zk5TuYXWWJu9M5dg5/dg5Bn/nXCB4xh1fzL7Jt/O0iQSo5NkcfUIWe
mksx1C8mJkYIDTC70u5BmIQyn8Jdl+PBrtFIJa1DxIIKs9DTImVtwWPnlPQmuEho
rr08In4TtWb+9YKXNB5bK27hA8GURwsSOEiXH8mmuq+q46x3ERxhcIF65cuNnMRr
ZLoMgD0eIKYASXyLfdJxV/bsLXwvkZtCN7g4IX371oVlVoDE0z4WQtupUhYsnRqX
OgXgzTWeug3RWXuYdaN1n1L9XRsRsCtBvZH0TQ5usiSCv5ncs+NcPc+EWAK2lu06
JvJj8I9t18oP4FC01wBZXAo7EndY50zLY+Wil27M+SC/1eAb/1v9iMy4EwLA1gJg
sVNlebc+XTgZkRyzdCcx0MmUVvI1g0fjeowISUIRz3begbvTDzRSEhAtpovZCu+G
SPUHgQjFjE0STV64KAy0Y6oAzkJvl+n+vgb/tFmLAPSlmRnNueTf6F1F6pSL90Jd
JkX2gwuTO8MmdNj9Ec0DxtJ2uj8UvHjCR2O5cg4IexLxK0qs3JLqH4oDqOOQhmwB
nX0HqRiwWpU4xswONHbUTImQT18u8Dxepvb2b+q96DK8o4A4DuDTTlsRvDO+GzFR
+m3DIJ6iBnQAI4e0Y3hazJ42HIGDBOMqAXVIBo4lbFs6MkR27l947SCMufI4GhDO
jTf7cZq+Pbf+zcZSerbrWWU/kXdpSOQYu8YCLBS/s0l1aZs88tF5/V1NDaV1v1bo
3qCOoBkru4rEgqMt8mpRq28adDu6aFIqFnYh7sg5tScMvprKOtQQT8hpxZmxrndo
GnCY2nv6FyOLSF3sa4/43m2yuslrQGbNOrIQZpuoqSwkpyBMplyfC+7a97tdVIcc
QdD50gOQuyozNdRp+1fYQq/HzVGQiQb6MeM4cmEdq9iZs0adUmQAOf9bG6+DimdZ
bwc7xUosZ4RGT5+csfH71vAq4ypNXB144mefc6TP+/edLiZ4Yqb5w317YVZDyRAs
z8pUQpkV74+hi9/Apyz9rKAqICKvAxRFKDITGxxdcRIbtphBeh2hTuE5lzDCGgM6
72h7Ug45DFWq4C+aZV+M8a9UnafXO+Qznir02sERmmH4Y4T1kY/uAjjyhygfCsfb
d2COVGpQ6K5gHJPlhaiBSte9lMzLZxAQBDwfQSPJetO6SAUwi6YYXIl/QWcfHaU1
ihrK8r9ouySgJ+83tSx9Dxo7WNbq2ruAd4birOR6QqgcK45VqRK9UEZr2IUFl6pj
tM8k//LR1Ibc//mnxb5DlOjk5FCeJRLtBINoVuUM6+UhBGG2/sX8NaVKCXMEqDn0
9uY3wqW6J7KE3JPdDqh1uML9ibqsJik14iDW7fi0EKZxb9+05zk3NP/sEwUVM/RG
ZvN2Npf6BTdGc6geIdZ2XEpWhUS99I4fTdV8kdncU0aiS2M+PZq5mqnt+CBnefJ7
FL12y4mOaEgoTYZfbdma4oY8lC8VNqhx2RtGugfcpsVlKRg6S53X8e13Zvdx9OD1
PphOYlT0hizneglgFJgYjV7IRd7MCH7SXstH4u/Beqi0ucHEh9xdWbVn7T9AFgiZ
2P17dtGw2nXkuscXIFVGJiR3c37uK6pFpzY3ieVxNV7ecRv0D2YRVYiwWgJfW6nN
NdPdDma8WRRAWOfXE75OWvetB4U2aOpQjk+fbkZQgrWMejcAwXpI03gxnq5ueGhg
eIkZuUDnUqxvb+FBU6NKSDyV/MksdbokukW+dxx+ALq3OMi3Wn00Wez3rEhzMLbF
jFBwUPwIoGJ0QMsO+5UHXwpcpEiT3Qe82m4ociXv8lq0BfcYfpbPmOiAlnZvW2mF
2FbwsET+vm+QTTfpMQWi/5zX8RxWZGCr6mXb3gzjWGRGqhAdthd7NxXAqkVinDpt
m75paD3Hc2yNnbkif9NVS7xG/m19JpJHOaPIyEKU1I28OarLBZMaKkE7lHv+Y0bZ
g7BcFE/ONcORhgcC2A4Hq8r0H+TclL9reVQLzkmGFHjqxA81kLoZkegk55spbPuu
4V70PW92UjsUfbLXPlz2s5d/h8KFJX91esORJ/CeK13i0LNTP4Eyzef528o4/YN6
GhFzn7bC85QvFOZF9xb4+Ube3PH3cGV+Xc7XLj+rqJBJk7BDB3nKnv/NgZtF46Nl
YvJXbAHCBZ31DF2oa/u26BiGwVu3ZHNSUJgYMLFvP7Z7dzs6f7ReFtExZiNnxzNv
wLmT/ksNJ58PgnPp4rjuotz7liA/TbymmH1Zz4zSVta6A2N2GgzhPkuvSSCm2ejP
KIV38RcDOF4i93XIPDajNLd5m6/Jy+K5vdL0pyfDRsQ/YBVF8y2smIWC/tQgknI3
rlXXway4Uv/NhPlda5e8zwJc2WbQH0JBJB5glqCLLgzt5Cl9rpnM8ckzecX2YMtz
XLSdg7h5lu86j8bJrBb1NAXmsaY/TD8lydSVMm3cSjRx4M+xF/FuWcPOuzNia6QY
RZ4elNkDVBkO3/0y25oiwDVUjh8xps+w6XIMIsT0Ugl1ttIItYzrL+drT8ileYpU
xe8Vpq5YPEF5R4vqE+m/HA+bw1Dj3bNRxUFQVuv/LIT4yvvZ91A00OJWSbTRnLRo
ETNREuvo02KbiE/YRZUpGYHdgScBjS09o3RziG3WT7XbDhIUyhsl+Bs25A2ZK/gL
5/mKCSDKElvpYWdqjzTQpU8kHZpu53QVl56R1Y1q3K5jqAM73X94jsbD/OUi/tCk
X3vDK8OfaBF9/LkxSEYfcxCjv/iAdU/gqfu2rC2Pi8Bf6SbmuiLZpq0Dv9o1UIap
qMf5TimMZ2YQGll4uOd4RY/hb38vcaHaePW7s8WidcdEDxged7tSXy/3BrVy2CtS
EQ7ykA5Aycs/8hA+1M8TKtjUeCcLdlSxhFftAIIPKeNCZv7gJUQoYBrqIbpqZV2Y
Ouvp6eW79WNWnJ7/hj60QRPq5uZxApdRPTSUyrp+0IfFCaEHO+KrV9eBHlya27AW
Wl56f6ZYTvPWaYLwfIrUR3swGKRnOzXa600eDrFRRhWrzF0AbsyuTh0J92o4TZac
qBsp4xzkYgplYohB2JTXMImoUyS37GV7k9lYvkEKs5x6ijom/E66ctH70bZwHqzM
zLcMjYQGH2ddCigVz6zHo8xu6wowJkchV9sey4yZMK9hpr5yDBhWdQ+p7eSy5y2R
Yr+yZS5tt/zcOEm7pBNwdKmtUbp9zGH+VxhygPZsLKnqR+Ty0HLU2fjDKGdh7VoA
QMF5cQwGVm9Yp+8iGJeJIdRWT1XwvWnGaI6ktoEtjDLFd5bQQoZfnS2ZIWQXkvj1
SzqCpjSXaynbqSRHTeqYZRvC8ff8x5QIHOBHpyYFlPWx1UbZUwYoVUuQDowhI0Np
1K8mvsPy/Mc+SJFTOKs595ceKU0nyxKk+XajLslacW7qjf04ff/bCQ/1GpCGlAtm
rLJY6FoKl/yXd4vC82/Uzv+uWjNg9CSpRiooalUtnyDuIFcs3uRdfCfodzKCsIu5
sMaoqRpj0RK+QL6qjKMF3gZ2IhJCXZCGkhJtlj2XAr8W5/VI9bKe1D5X8ghnBDAY
aFHea41cbNNmT1pyeXvPxgnEgxkIFcfCqTbcx8EypliP/wQNpE63w5VBzIv0B4H8
ohpH9HVmGKpJpzPi+u7yFq9erPSgsfloR3a5tqQ5YnsdGkQf1WL94RhL6dzYRTYO
+eBLcF/MQnM9Gcozb4jATPsk9gyFkX8vvw4TaCijzF6rT4AgDH6j7A7AbWu1osQr
3Oh11OjaKh7S24ODGVN1+qdW412mzygdA776bminpiGZeasq9ecYn6tAprGYtepv
WeNqAS/KFlmOF1P2nZJJbgJcm1Kl7SVrF9AOYb1i3Lu2eFI1xtVDvXC6eJYWbECS
ZCbtxaOrvwhVECqFdNs03iTE701un3TzuJkeG22rRe35HPHoaZMgMkeOzbJ0DGex
KOaZFQLbI/WmZab/+T0lJJErZ7OQEGqMbGbEXM0fCzLtYE6wvMJcGdEsXaQ9MFGE
dEOVi719Be9YmDQUTRmhWV52dPlZYjG3qtvRzulLIXE+mHArIMnZSUC+wjgP+fTq
jYzJtex5PnzZKjSz2bQ97TPicFQNe5AUWHkfNgDjIcs33tL8podADBcs+2qZJAhB
+wngZJwLXUt/gIDRf7vOplztVA1zrbJm+fHIWY0zAAdEFeok4/NGboke66pUxThi
nMvBWKjBTuva4fgBmwT+Ou+tjR+iWTALAt0Jku1TCn++JCqikx8FWpl+GaN4Po6Q
eT9QgdrukGOufgbOMqUYX39JwSK/LT7r4V3qUBKrVYniRDLeDsTR4rxatHfBg0XB
SEM6uD7e+bczhAvfRONLLtPHh6b2xhaQy+1J9KTbDwCBiSrN1MhtkJep7cKk2uqJ
092DdyuPeQvAXXMKkK/dMUd3tEJIjHk+fNs9+aR4VwvEEWF1R5HACuNngQC2U5fl
ro3BkQp5Ldcjs5d4Eaf5Bk4SU6YycpoUKYhAIis872w4ciR6MF3JW/4JAelkWN5Y
cZg06DptFLOxKnpgKc6PIeQNdrTu/iLbI/wys6OWnk9NcAUD/c5Q/RNcf+qpGyTB
KodM2lyNdl69rnOXGha+MoFfeP2fF+jB+z675ELSSS9rdK16rtcdD9g6Tr3A0sNd
+SelWppCpB0McU32s0BCCEoEWkGY1vbsUrTnk7+8V9OewPlKTcPrFu/E2iEGpgjq
AmBxrt3lYxfOdCyJv/BMNGOEtiH79z4yYvOKVekDKHDZ09pNRUS6KXSWb7Flku9w
VtjVJf0HbD6BYZmV95pnUpN3O1l1KkN+rV57vVfYK4qEgmIG9BNCdWGeeaSTHPUr
4b747t9v8CPC2RGaocLQaRLXQx+8USS907Y3RObf99ne2fH8mYm6UuB/cVI1AV4z
0TN6OfrkKbP0zByBF8NnTgvPUr+gjvlpEBUv9NIW01D6ONYEmlLcceDU/ZJT+aLz
7LCm/8xNetkElWbvsidbSCNZHJK8SKZNnf+T1iuzW+Y5r7QYurywkLec/unI2WEm
M2KR++1wXBBB0Pc+fYU722KQ9SRp9Ok09wyHMRA5wXs9bBijCqwrSo4eY6kDXoyY
k3lIUektzH0CAlO37dGjrjbsN7tiKBfAnunIB8nMpt1MVcShRHkkmTN0jIsAjJiV
qGVWxB+LAczSyNRVCU/S67Mfh5lWZgdlVrt+90QyJRkU9rNtbghyHnltPC4FoKWR
IHnE6RbYzdTkyR0HkjJXS0N4yk3zcS0T3UAVeCPSqGpWmakWXyFOX0DVKHeWqMmB
7FqjifgXDU7/Tn9MNwFd4fIEVUJOGAG75Rz/3Sx1JVZ7Q0aBuL3kpkkZc9MSsggJ
Z5JOMtiLVChIGxjCPvaWpr1/Rb64UefMZarQAlopFYSk4F87XWUvyiafPpK3IQGZ
CxncUBqB3wWD6s6enaT6jEighhwElqWxrnFcdN/pp6sQt+N0ax27tCYN3f10vPqJ
7xqudPT06rokmXbyxr8IZhJl02GGYi2bY9bY2oCFh4QkH00l+xCdu5cdpdN12gjJ
obDLnqoFF5iM6Sokt6I1gWlYFGWQjYKh6r+zATAd6N1/+Z1t7lvHN+PIXD6Wd1MZ
ujGJQ8CUeI6IzWlg2BVKN4Ogk1X9uBrFZFTVsUAdx8m7+AQIz+lkFbrinnF4EWyf
qub6DSyHm151/UbDk/24ukrJ/kosLoEdg1wwoCjfeGP8nhfsesXpg/CY5Ka13xW+
1JBMhrDv3VgPCSerk2BwE+a+P6/iuz2DiaalV5CEt99I5oYgSds3smcWRFVNhPTI
HoijKMYBEXhnraqZSCoh3LrB8xIiL/nivh96+HeqDCZ6CTC5kpRVpmvzcnPRUlhw
G5NqupDQ+VatsIW3ohI274SuCme+IEpVHzMS11kbQ6Sz95P1Xtu7Hle1ONSKMuZc
/pBYsR15uy/wXdsn121dAk1w+yoaL1nsKBc7W8glS8aPEahyo9D4XiJ3AY57v0cd
XWKLuFWIdSrQQNELwjTgZ6HF0VgRHlavyP7VWBuN2hPPMKG9lBZNvtBNpk0PKR0d
FB7PV4jMS6p7jfmQrs1zS23jlfC2q9euunLe/wLAc2ecQ54V5UH2HpS0mMOzpB6W
TYnFzVmXfevyz/bZUbdsEwdBZ6/R9Z3ZAhwhq3/otdtLENG6/aeX+oKWFrY3FCMg
vd4AOpqyLWK07hluXR4x0i81F+8kYu6sJNF5uBJmmOGh9/pH9ePraeX5/wuvICEV
qBexaG08UYxkpbYCcEva9Ie0m8BXzgkqEGgTB3zVi/3qj2osTYUSnpovRGBKxhRq
I156msxzr2xViN9YK/SassJZL2TVG3dDAr20wJ0E1vFgtCYWvDejKz9b4gClLJVY
Br4K6UUnOZeYtWSJTmY7ImUu10YNqeco4vmIMcgh6FxzviKDwcEwz8kvmRrNFxEO
kyrprB092vcwpuCHPv8FT58aXNWl8LIQg8Yajq64fIzKTxmzNj2qwaJcwJRQYO3r
6jFlXAQV69Qdvp3qyLt19rPGTiKOUZ7qLGH/TEUonpb6koZi4PzLmgNSY4zhJJOw
LelXKelTD9RVMnKM3pl48a7AbvpwGNNv8qE16z7OsL4TmSmYr+mrFMbTS3ZMmxU9
fnB+4ETdCoo2GotYsSN1EgiOpNccAXwk1PXUjTvA+FW21dWdi3CsLeiM/hnUUopH
sAglQCSxxAqUZ1G4YLAkFUieXakfBYyxTV3UQE2OPBFRRgMGO3tcfDqLCrDR2Iyd
8bQqyNHI7Iups3FTrl0Nuhnuvvl+3u0Z1k3If5EnAvHiXiqR8FUDX8kChA700bHm
07lpyaIleGOYGoUN1MIvSRUhWqokYYw0H8G9QFT/lOdNKPi9y/7CTjLx3meP4pK9
FbSHltsD1R3RLn/o3rKIAsfdcPyZAfzSHTBtTZAbKS6y50PwwzX1Agd5G2u5D5Nj
0uKiGox/B+jpObZByE9tR2vx/dYTMHD4W1OKKet0eCUgZwy+abqBTFbxG4ySlcj+
eDaADnNUT189jAfumP3J3aj1VWOo3iDcA+wa3OG8YbbV8IK/82zpdqZRcz8rNf4l
7GzBj5nab+CHNoZxuYp4vEGWkNe0pSFWmYBg8ECLSszSm4FNcIMYl1gfOPPtgzak
ub7oKdXNW3h6cSgE1Y4O7/fOukNkvGIiOO0gllZuV16AzER2sFp3kTtem5WflwvP
PUzDUTbGZjiAi51bdJKG4K5H10j2pLzDiT63Ym7NZTKdkEIWTxsZpLSPY/KoRK9S
fv0AzYAe8/wSX2NgNuZtkmHemzYOng19hHkszMs9XPTerSyfOmKrqkYm7g2XCgCj
lk9YrX2X5Aa6GFZIcE84MudXttd5SqVhTPX+Dj5SMJDh/ohe+BOQYqtcS1XGdRrC
uYJmPBNdGqHwhGyjiQEgB6cBtkgdrEDGsd68E+j/QLVEbcqPTLfk1LJ6yKrTNxe5
K3bcE+b5scHPVrakDc+XtPsJ6yugkP5vofl/d5UruOKG+cSILZRycJthE+RB+R4u
BvQwG14hQqD9LZBiI6kcdqUL255y55OoK3gHTxIU2p4OyfBLAwhoTgSw9Iqgvw87
IhCyRgjTJUQjUs6rwkJyvRcKEPpVPL5mq3O6qn8O/Gnnccep5CMDSu//GNwTKLyb
GCoQKiUbNGzYLeGsqBhBM51Dg4v4OcWQPfYzyI+I+WqmJUvBoOmfXNVR73mg9nXB
8eKHQfyql67plIAvhQI0VGYWLfDp/uIrA3gO9VvyypHcXG88lsLhJV6UhBibSi5Q
5qC7hQNdVFnM54iUfiAzxnGw7PA3UnAQzicu5dqE4AE+Xq2xS+Ww6EEjtsGETctu
VgTwR12TAvjuE5XZMYCMhRhpnwqEgSVF/S3mp3uMYiG5oJVmV6s97zl+pyNSf70A
nhvhp2s35gFg8XLv9lLL4GJsbD3UwCkaWah/NaeNW1oVaVpvCzp8mjm2xwF2ANKp
vWLE5QyIJs0X7AOyCAeIwHtLpqSDe1CUa30Fck2FP1pcT2diFBI4MAJgfeSJqnSv
D90DzTh+ExhbNGmNb18XzVyGCBO4kthf2prBIGpogGolw7MiaxlFEtAZDmYsET9v
tVxyRrDMKEII++kxAtLQvpYUbAR2aAmAo2/Q5zhJlQDTSVhlhM0Z+a4Uqzpq7a4u
lmGnMPj+DnnsWnnjn8sMrF2RztJ+hj/633CZFVov3cOTeghkjzOQteuu1rqN1BDw
YAtLOp+97izZQHOZBkVz9+M4x+2b2bMapgfydEXPZP953yMCQYtgz8dYpYDWvjnp
qCZKHfAyq4Bn+qtS44Sk8792U+LD84CIM3KYKLFmIl8TkG9K+cfcZOQIY+87Ioxz
s2RLGx/EjzQksyZ1x6YuHnEDPpRh0R8Wi/tKmKPfYe9pYxGYre8rGscbVTjCJIv/
Jy65Lc27W2i0Q2iCJU69SDLNQlVvze3hSXLpMvL4rL4A4Z3WDuRrLfHgTNI5FzfS
xREwRGGoH+9d0B32UlGAYcMZh//UNN5+OGKiU6ksOuI/54O9pw4mAo90Ub4/xM+N
h33WlFljHS5vfKhgbs4uAl25mvfeeTa/c1/Juln7ya69w6ffnB+JDLtj6Xf1/nND
StorgD0BxgbWnMRrOlpvelnT4cnDbRWhWu67tAce8oCY5FZOMSdYbd6pCXnWLLfY
H74Zib1iTuqNUGMtEE918ry4ppccAv1igeaLp5ioCPYdOx3bXwsqyp+4fq3xw0MK
ns3Fy2ySvmRk1yytwQB6wRXzaoGzyhtSOQ7kaBGB2NO/iG81v2t33N/gmt67G5gI
FBouWxJbi8m6ybS5SJNlKp/k55zSSvuHV8PSApJOJwv/zrcVBYHkf5eDrwrMOJOp
MSDFy7WIQDBGoFGGaf9YQhulYLtsCzOfS6knQi9S1whDBfXBiaE+bymFJYIaeP1F
+GC7CyVPw6dD1GaqvedS1AP6x1L6+CdD1VBi5ik/NaU+qetUeklvKl5JDc/9uO6i
RHjNY/NQl2U7xHioibT1tuJIUpfJFgc1QNpMTVlU4br4B+IoZduBNdPyeWqEhyVr
gngBXWnzkkkYduIWSdhQZ42TszjG7SJVbBxD7zYJ35frWCiTI2LW5ekp4kh4HTIy
xuKmt/m7+9vo3O+hwVnxkw2YuZKdkXaZBedJMapiRQ93XIYdqAO+5hkqIIMoaMFf
rEqJs1Qg6sqQxTO25wCvvsN03vNlWT3UpYRY8l76GfbeD2Zit3wQvfLDl2A1R8QB
mBsccPxqN78JaMVdTAu/Fx99uD+ve6dSBk9guOv17ZXbpGWMRg9EV18lu9bevgo3
+jw4jZoyiKbXNtC7SYnjII/mjKJrpmAeEIJBkBDrERB3vt2WBq5+PlIA7YOXj9F7
O9zQpY9u3PeWYDzOKGCBCV8Ik5PoXyr8h0dkND30V+HtgvA5g+TAWIve5npl26Xb
4Z+5TiB3gEE1mBmczuvoqJnlr/Q4WFvv6wYhWcIoT1DYeUT5T/6xNe9oIEjlKujl
EdjBc6lgr9m9+Ns2vMfQdnpi7AetBoTfA5guYVeBY1jfqpqhnc4/4cC1oxfGPE61
UtxpaVsudjG5qxADPrjGI0wby+E+gDGfNMeiyEN0tgs3BLoxYCQQj+qt+dRutoNw
pHEM2EGs02Y7gjIVG7CSukw9EVR6ly0qqKDCM38IQcwPfL63Jx/qeqyCMv5y2a+m
kaBdIcF78wI7sHlLt1rChkm4sZbzcDRolWRpyyJ70LMCY7UjLdFdXEgtaWoLi+17
LyG0J5hwBtY9rx+9e2axAnkU1iQkdMrG/ONiNuWXvkB9ZMpthya3hlpFjsO3QBwH
GIvlPV9TiW+oJ6qt8DQNdGERrFJaYkdYKvTgHAu0kR4AUz+4p2IPbUbOU1IX88LJ
Rqfqi8ftkM4XGm2ODQIw/vCz3tWzRF6lW7e7FtXUHsvz2ikSHSH2C8FYYgH+UQls
Y4dczuzVodpa/3g70MTPNv+ggn78Tf7WXrzc3NhwsqCXoff8+kH/WyonFHQh53of
0Ady1MTyg4ahAjT1j+cAqJ/9EwoxnoOB1NTcH2A/9aSOgeMs2t/jZzXEjTW7+0jx
+lv4k2ljLVd0nulf54qqKi3+9irom0GE42HsDnCTMfDdncO/j0gyqycR6HCbmUYy
4uOYwZqQ6/1NucTziBq9ufkEeuT+kw/3AXx/ntQwiw7IF/5Le0PEuIT3Bxf6U3zn
6BrCSYXhlnRPXu8KvtTm9x2pAUrSRtUU76Q7r5iD49NX3ON7OUVghjRmv5ISBW4H
nsPZ4Mrw5oro7dgFGSb2U9JimMiAEVeLVxrRHkj1uB/IVWUd2wFoaUjvL++H38Rx
A7Pngw6w0yDbQsBXV2R++l4v9Tv3j9GWpn6r1EPb7L0/eot0Gt9aqgzIxWIg5Yia
cj4ZAZd6xLMjjf3BpLrktoxLT1Dlx3eeCszL7SjHIGnGa+BtfK2WaCaUTcY+5ky5
eK4hOJalZtw7StghYxFKM5V/snk4d9ylx1b+WQF/qiBptNioo3bp/NvqCqmxABaF
T++qkMtqRLS7GTF96rkBDWy0i6jYL7jxyfTZwsNeBrnbM98EoeCocjtdijVjxRGc
m4xwtFno10BktFT3FfpY6JPX8UnoDynolyY0M8I0jy6trdkUJpKVRMXU83M0Vzqm
Tltxl5T+5r0fWllc+mxYerZnbAjPMpbYH0+AybvRvW7n+GD4ObupMDjQOvyIo4WZ
nkHhKgovEA6XeUIAuzkMW1xxhESQnEFCwFRIZA26rTwnxecu++0+ymhm9yUS/tCK
UzYC36nzo0WuEvrQ3PmbcjiAnERoUVDtzfnY3jQTr4lI5t6RySq5oaI9/mk6x5xF
woMzdZwohYEO8m9gXQOxdV5zN97zaxn1JpF2MegVi6m/ILjZkgoCSaXgXErAErCn
3oe0EX2BDxPNO8zfg2G1IpksHuhGHDa3R3tT1gRmE0uGqzCnYhC9qveVDoHBduGI
Nq9vfAYJFXiqpwptEtzLhaT99uulSNlxSuK/XymRdwfE28mb6UJLkb1i1X6moguJ
WUe3y0/Dp7ikPP3zfD8Q7Llg+CUksIuUAasdJY/rdo+04j75+j39YmB32zflo3JV
/9DiAvpmKaxsqgA2RBomSvk9vHzZOn4Wyo/a/umnjeNm65m77lxWTC5KoH2Jv2oD
XOQiQrIYJVINkf3ngwSejQvIadAS2eiq4PCWvsyBMBg19NNWbKy5pEJV8qJj1e9p
PJMOUt5rgpfM49XtA6Vqor2gCuG1eZA+6Q3AS5R18xfWnNqHtO8CaJg7W0yeHOHc
9AcsjlOhZxkjp9REqjhbwY2K9mR/jDD4rqwzh9npxtJdxS3DDWJs8yJb1tPC74+Q
ZUzLdybWrvbePPty1PZzCqzYhsQYtDlaRdlSEhuSn0rMEKGp29kyj5Gn8Oa+OC/q
jn+bOuKUxgk+qqKPWWzHE5u6vxJ/LhQsiaOeiwzzU1pDGYqlcw2tVSf9veOsRyI7
YvqVMB9BqYGaGyOaX+ypqMBllz7Wf0paLcp+oUOZqTUDa12+KFya/34Vo0/Li1gd
6e51YhT4rwHrotozphxQAIWzSBbQ5UuRc0GK/oHl8Xjwu+75IdglRDgKy6/c2S2v
Dm3/doWGQZmYdFt1wusK/G9SkeBSoo8vT11CYR7gIxOHW7/Vzp3RupsLh5Q91FUt
BGCRnXEAeBuUJOJa0UohK0Wan2nzFPJPZWC2qG2+09Zx6lINtCi+rl16OoQGwUFK
VhG1D2ExSuoatHTkZO77FrS44WOwfj9ODjVht46XX4pxDhnCCVcy7tQwAuLYY4vB
QwjZ2ghAYFmw/DmNbRWvpj4eYOTaneBVYaqz+fay+i10CHebjgi+epqnjtORJquj
1PeOhEIzXfP/Hx6Mux4n7suCiOi9wa7OTXovFW51flPqL7w5kWQfWTT64/Y9Cw1u
aQMMZcwDMmY7ViRMdaZ9SX0Vd8Zp1bp8hi5ShvkKjvFgD6zqmbQtoYAMpvJ9vLrI
/0MXoty840qt0m0uPuPF+J7iB4aB6tBrcInFLHpk0N1PM+ln64fuBKcv65fQanZg
IksZNLdnqJtAA/WY0PnVbiFakU5+4jDRuEVOOve2GWJICwLGr3iIsxy+zjfb2IVo
k2biXDd+fPQcxH48ZKhyX4aqx7arcyYXorvYQCIwTYzTffdNq7svlKk6fqT0wk8r
oeSMZBNl0ZTuepP2fcA62kDpl4uf5vaX+fpWCT6VClUtRrESKI2jXuj3k3e3rBmW
0q8LLyi1UtDL4Z+FjNf53EpGY7JDwhvCcaZxU3lAUCqLh4W0kBiplCrKF9n0qHpL
OTmi38YF7j9D6q7qftJTkeozbeIBSmnNfWJICZj7sb6EYZilflixePcpEPaoKvB1
NuFITybKnEAEMMrBOmh9m+LYmoThMIhlfpVghabuYpEDcI9XiEBMl7+hK/tIBeDP
ivRwMWxzEykGJq8/iJiiGNrwwl/KA+95OyIKyVCe0y20fvpYJkMOpjhS/fob5qzn
MZGj8fC9j1kmJ4PfS6MG++AbdLz++gVGDBlcrxs++Un6whxPto28A/TapxuKzXrR
zUinbqyIjpzjSueZrPZ3tt8RnXSXnsvuQ5A+DPnhyklEImDZgQb/HtahynAyG4fF
L6wElqpCYfWEbOElNaNxuthJ/6cQy7Qrv3gOJz9dVbk5TZonQIvQp9uUHTtcL9y6
vV9XYhUSQyiN+MQJR98nNUWsiIaw4p1IG0jjBE8TL4i3p920+SBdzeVZIpCzQrYX
hZTTJiVBTJt7tAxe6VERtofxH+38mkMC4A2SCqr5mMTc98c+k9u2coWaO59GRzvx
5XI3h09QCXWrxyFf3vu+vdOrJey9ZUewzS7ACXdzHTN1PVZNxteyVRSHSebQnPBM
pvODO2GuLDboSheyKT4ckRV6mIiK66CQeem97/MYttpyD5DTh1qR1FPQUGAECK7V
ENQBdlqr4wJyu0EqTmbp7i6NJkowDJfllemjXDQTE9hZovaLfoxXAk3MAMmrOabV
M+y7UzNwJQ2V0SfuSLbqJML4DfIBgm/gE/A+fPspTM5n6k7eS0wsfMFSl72ik6G/
viZ7OS3Ai7vPJXv9UCp84HCqBfJb77HmsGCUFLw7Wtj5gvLVfrj34d7RKv3XNoBN
PaOr7XvhbpABesq5ULsfrciOGfQihkrgz95BjbpPVUXnRjATdb3kiJOSKRtlfSdx
fAsLEXxuuiudEGSaF6jxKVyKH9TONmUplH7be5J1Bpd3PU5SFuvoXQ99gu4jAALW
TgODzaI5gnBMS/JSdkerJOCE2xMoI2GJ1612E1pzhSvvZrTod1qr1HA12YrRZGFe
QURjwEf9CH0GKa3VSr2E/tYAE6GRN0lTozH3iidud6EYJnN7S9VkfzXKJt3s6lne
eRdwRi3ApJ5l0SaChN6biaUG9zlyOkNMOMQten+Wvz43mcGjTTspAJYvqIRt2Z9M
tccm5u01Pon02c9zBg4pnWOqabuELsBWbYl1XkU8rYBPKB3g6G+YrkPfJl0vAn2i
g6tEZw5hQdrq8qvDwP/ZaR4DUKFr+wvzY2RRMJQNRBzpYciWhAF2MAu2Gl4LsBXZ
0ZGTHHGHCzqRBwleLi8kCcJOEm4CxrwIw6oY/2T1DCbOggt2iuVv0MP31BgcM/O7
/bOyFaNlRlwTu+oF/rJv0Bp4zEHblt8SOKu1ABelZCaD/sRnglqeFVM4LQmtN5zv
dhSl0MFAQAZB8d7Fz1fwaR1syuzwnqfPhfhSS1FY6ZJGuAghcMT1AqIk7CCGgEK9
71Il7tLLU3J9bUTpIhjOfxNJVZqDbELNHUnraxbL4zdLsC4P/Vcuxn8v9fhf0BI3
Et/BAu1BaWKWzHN7V9y6GCmvODD84DioyIsCmMbH42eqpixoGVvTgctLzixV7NCk
m9e0Rq7KIup8T+3JmmqmnisPBYdzPCObf14WGNO2bcbEBPvg6Gk389SYxZ0MZ5zO
pbXW3yFJFRYJE1OJAHC/m/E2Q+qTk1kRBYeZ+nvE9TKA7N1a4eGi9HGZWJV+9mq5
6Hkkd5rjHN+V9ZUZqa7ug9NLg6/NIXknJ/xIq4IaPdCFAHsTOokSS0G/PRuX1mzC
sOvDJjzViB3E1y+SRAcY522GwOML86aMH/ZEIzto90jxa+hVY+NQYWnYYCaMU/4B
+gj81vu3KSTkfYKMeHykSETsdn6+HfJQbDS8Zep1wE7zO8RfzLGcVst0930Kp99e
VFXmQPYUraaXGG5Q5kXwE0SQ4VEAVqFcRgn0ftxkLdBYx5L6V05FAKQdJjqYeurU
gh9//heln2M8L3tQuRPbbB1vzxZScl2FH7DlKfz+Mmidyh6n9TO7NfuIQoGsO76G
s5tS814EdSIq6ptTeDOlfBT34SAVBG0XaNZ9+G4gCB6J7iLb01HuDRjWG3DUo3wG
6IOZzOkq75WxMlGn1BLt65PhxOku1IaCPA1ULKlxEKRYWahUQIvp04drHF97n5+q
Wk3PrL0aHJO4cUz3F/XiVUZWkS7NSyZeTMHro8lTEvyXPQMlZEZgfPF8VD3fI8yn
04KJ3rjoMHQ8fkdx9SF5t6xMmso7R2wU2iNxI+z3r+N/mOKNqf7sU4mNnsHxd/R6
3ckzfyMsdFbGHlr+eRNz96APnooou7NBRPNXtptNIv96RIYHjUXYu0OXQSzeDWZe
MBfN/YGswNQ2xjX3IE7z08pYF7qqsy3T/efOO/DgoRUp4s/YAXkuiRYV77gxA7dK
R9TBUknwxSQ9NS8Es5yrq9BKRAGnPrrzjUlDSzPyZ4RQJBGVctHSVwXtdPJOQxrr
Go9e2p4XTXNMnW4TFeUSn7YS5MYCcCJ8ZroEqWk+j3HSEA9ZndxDjsIVdrZQ00+B
tC8Es0tYwU1HqWbtr/w3BpztK4/OztZ4xPkdH70RE/LiQJSPKbIyDofOvdEXyUos
g6ikTydMIvKAqdFJv4VvC7Rh93IS2KG6H2CDKfBDPs6Js1rM+fLGDkXxePgZg+gU
FXES/o+X0o2QIhXq6wki1fPlJURD2Qcrn6L/jsJz/aHEDQ6nv05/hQOECesqpPZi
WFftfXKi6t7ihh85Rlb4/dTpY3BUCok7Ao1tGQrV7ulqw1H6+bw2MtNLa1HTjbrl
1zeMIPwkjaDGIqWe2miMtnSjlvsGeE6es4goYm1dDPgW1Gfd4DAy+DtJ04jIGhYF
iOSRd8aPI/arE1QqpoFEgBeq4abuLl1QwgHMT7DUeMhZr1wcYwbgaOl8RaPZ1paa
PpP9TQWwSC9TBAwOyspCwURHqhTNn/8Nc3urA75hj9dT1uQmi0W3ZrZdyj5cZ6tT
TKd/PRyxh4o0MjxtbmhONqhaPAAyqB0tJtJKU110DqZ6SE1tSRqAtO9U4z24IiDY
c4IPWzldeMqQ70BH4gd/bJl5zua+E70HM3RxQpgBQYBh9pM9AvQopHapUStpjT9e
RRFjlKL2lWMSVLC3ZR8L09eQhU8SZ6v0K7K53MFDn96uZ9ilIc5kdq4j0JXEsAIF
hRLtxMxGfi0V6UURW/WCjtUuiahKSK9gwM+Ai2p66Aa9eRbYQ5ki6tNfdBDMVuAv
xiECohKijMuFUtEA6JP1kx4pygSfuaFzU03iYu/6eMDS1b4wmEli/zJOI31SQhkx
osFwHh/4547aG830DwPtcdr93FEJCFy10VsBrSgzID8+DxL5NuW4OM5/mhGba+im
h7FNfM+p7ucaSpSlQmzBg5QJzYk0/ctDBPP1pc2s6bDb2/vEMCnVk8YFkNUo2hbn
56kUQp1uvwyGK3fjObMeGZDGHUWmWBdOg5ct7mnJNR8J7TWre/Pa1pVn0XhsPMrD
fffTKNqbVbCJpu5yhIph1cuIN2D6zsmXTl/jIlBBY9AwPCJ5loHDbeqQw9DC7Ubt
sRe1y7hGhDYBMA+c35Jam9w16U/4t4CPqWYZgzguiHA1clOCn4gSCI94hu7kTRVL
3qGoSnJj026NLNxOfaprhsYbcnVVuij0u+sEqr7aK08rMbSMHtkplHlni6n8TllZ
0g3BsmKWGGvIhyOYrnIZzDlAtKu5xtrzpf69LbRPesJMCRTYbge/aE1Xge2+tbhJ
z/Gm+oV6QsEmm9EBO4CPCd3TYpkSnRvn5k8KEC5N5U5yCI8leJjhZlBdkDEKN9vJ
knQjYBOVpVOWwkNQ6xduNSZU3u1U1uly/A+p/9EVE3JlpwHY9d2zyX/R6PdD1YhR
cLG8YSD1bR5qx7L5kiWNSDFSIKjAIrX/peLmH8FBRK5Nbb7gwPE7EN5n5QUSgcnP
+JTxKaIP+hZczBlzdZsgYva9ZzrW17IvxYgIJJWzZDe9oQZvBlW0pIFtpukDaOiQ
IK1acYY5sDorXb7ZB2cqoz9Q/Z/eAcpPJa+rOAlcmVLW0OpAlPcRpE8+aLHrd/K4
syxrrC/AQ1FaewCnpgJeicEVYhHEMhg7we7Ma9XmRoGPBgpctZ87QaBG6D7JYxM1
Qlb6NMIGcJVhOavRQr0DG6Sm8R2c8VOyyfeBA3+JfGiPVNXhCt+zLcNMksgfpeNV
UR9fgoS+fc+BSjBzBmXCkScYj+5ff3RAMNLUn6HBn17GS9Y0HIJtw6/lVznyeIKd
l25ri92Z41MdJno+p0hLfG0R9TNvffuHP7/hI2ZWQEpbvBASOFySc9LrBhveK5IX
mOTce2GUI0wZUpLxh9fgyjsr8DiSlIrpXbd56tiE4uui7LuXKR3RjmOZD8/k4KhM
pk7ymdi98sv4XsnJ5MdExv440eIC4vxILs11ByjPvYLjlQjazmb1k+Wc+snwKK22
n7ENU9/rNfFADBAHlasUvZe6lnaepej5UGPuVU/h2YhXBnZnc73wLUeT4WtZwZFz
Ha+5v8GQOAjbKxB9C66f84pY2TLOqkCx+xsws0Of2opyAGa86SlE0UMf5i0maiJ+
d5VC7eeHtcVztqVD3LBp+xdIMMPY2qd4o4Nw8R3cbSr/rIaN6C77kQJYE+Kbm6ca
lB4FQhr45nacoF9rr91qY4ycznuO8hZhFCVZ3mzd6z0RvLhlzXQ5sEDDAZAniaLL
+2IF/abq1MQLoIdfXFIzIsrRZwMiVrD/MDbLdpKnRm8mX/VM3QjYOmCdZbSQvzF8
90JoL2oqDZQjy8ZG5XuKniDMAzAEUFBNPh2gWPoe6EMchVGvBGKj+YEs6QEE1YNe
HjK1CYtJ9YPyQQ06cUH3QUQHKN5j0KzZfblbTiuqCu7RVgQVSyuaovSO+2GLX51n
ESQfQbJ8GfBQm1llSQnKzgZVcIjsIBnuek060btvMMaM/6xCLUx/asXUFleGemQv
LNOytjO57ZaeKKEhzde1agizGF1eZwSNmuO6eLoHAjqwhiCuaEMC+3EZ682iTIbJ
WnVIbrNImXoMUXuo42wgZRjKlZxXfNhMnLW5iqZGWnrzaTLeWMwSxJQDQ1LLlgTe
DzY3wXGMz3j1V9bUCo+mgtjErGf5fq2wsFIdfR3be2neVde08fm1GGrObMpSLPU1
NKSkhX6+CSeQ84uEYCco37oyq8E1E0wPxi0D+zWaNwIy+gS58W0OrIwqUagF9M6H
ZSIl2ND/zLte04CAQXlvSdGw1ZgLFLZadKy9rrMIPUSZhPGk8sJc8zH/EZlg0Jx7
H7GJ1vgErnLnj9fHKSCZeX3Rcpjs/G/hgsfpRN2Z/sT9ECyIXff2p2wRuLlesesB
2i9TR0WxY9kpwqt4m5bO26zOzAagc2axZ2e80HHe4al+5gwmyLF22IkECPpg4Lso
e2fsdCuCArhUc2rNl8Dp02cUxg3CPk9YI841Mgna6YVAn8wZlhvQEbU7eH28+DMq
xoQXEk8U5hAn2AeirR1O5b+qem2z3iWxvBJdtwl92lGuJgZaR1a5h3+WHTvLF+fn
xquNHiO/zFzQGEnCcBJJWVUKISbzV45UftzMg9hsEFkVPFh7LAJOuEm28NHDmXHs
m/y3P0fl2TMUMO6YmRiCTgMdm8llz5uyF5mKwhjBdkIF1KdR6HmrIP6ZKStphz5J
WAlOM7YB0GwiNlKuTzwUBK+vZJhbr6t7/jy3dedbug9n11sYMb1W6YtAoHHVscAi
gmEW0JnqqoCKpVwnoey3I+k37jvZ+XEilAKYyJPAPtIvZoOZfpo+DvSbAGvpgR/B
qgi0u9INkfB+adp+T0di0ijEcTyWacf2tj3yXc+e991F5MVR5dGGdUm0GBpPA1AF
82pwFP+oMp9Koq5UqJB1Nps6yp02J9gIkJFe4y3LoXPEt5BL3NNEI1AkAH7LHjAL
1ZRNqvkdWtYvlKaTnDjQTFqj6ObHGsv604Y+Wcvta6g5xDuyCgxykDmMpxmU5EJj
GXNFuGfVhE4e27GAQu6NU+QH/gQWZkFmTBZHgoB06h31cEaUqGKFBo234i7DXLix
npJ7ekiVvdDvCPuK0Jb+8p266tJgevtsyum+2phr+Pu2q0Xw7dOWBM2kDB5Uz4DO
84RX6Ei36iWMY0akfw9p6tGBo+cfhptemW6QlRcILR+xhPyeNc3DrRwBUNQrO4du
wIRetHIjkZURE407dF+YBHkz1h0CL1INdJ9C28C6u5Pb/z2gM2E7Ox9ojO0Ch8Bb
LtTcBS75Y13f6BRC4GzvTXfitaCHZRqJnkBh2jEhHgu60zOqs/jojr/BfPzaMd+V
vbu/nZmJTDMvZMkwJSnNzqb5yjQsxfaHq2NTHb0M3b7+DLplTkmNavIwK/4xsT0N
wrgQ3zsq7+4HqUPOm5ccWdbsZ0OSUJrXa1mhNJjDOARdOBExHKCIsAQkNI8Hldax
eXJM9hVr63xTOnhw4wufVpuGNUC/B5pVNsCRj85pDZLp3V6x/F/gIex1gsWm/GL5
XxD43zQfgrnBJay1J4E9hX2hC/a4110BsWg+S6s1sxCfCgA5kSXGq8JspFFacHd8
RgLBiit/HIBFHPvsJZOM7i33CBUs9sf+WxiP0FgFY1LTVqi0GMM0hiePms2gMmky
ZNFEPRcKKrhu/QNVU/Bx52nxr5nZO0Ic/ghO4YGhBda3xe4nf56p7BPMWvyzldYE
cKbZXDAxMdr+nKqYujve0SOBJo+EAi9rfdkawFlXimhMnEY7NJIwRWC2sYMCyxl4
AwZ7+LsxEIYQT7i4evtv1GsCv4DKe6kkjnsz9mw+GY7FHvf8XkGlzl7pcNhtK1P8
laEdQJ5b+5xjAaD1XlPHV0PLHuV29WYMOlLoU4ksr6Rlax+8NdAnKQDmhq0MaTQO
ogcT0gylWGlpO8buCbj/fGIGlb+61csyl3L0aRJxB8HQcZRxZkRgXNPHysKXYjtN
FC5qeGgQZ+29FfKGLS4EXGz+LfMRtQ9dcF9K5wKNEU4BIOSWoMHfrr4qrrWSHnPU
YTClQeSK+71W6beb3xlppJAahQJs+s/iY551Uz1ATG2HSGMB/g1PH9cI8oyU3QQz
U+d6lAWJ4LC5boZgCC5f9gznEGz523HlaliExv94zG4ZPVplkEhpwE/a6viLsbS4
Pa+x0VW5Xm75JZ+3Lb7jQgTeYLfbuu9Xa1ordKr8in10BlAohTa6ZIgEKSNVROrA
P7r6bOKIVdS/WVoX6/iM7Zjp8Ybo7QDV6VrFLmnzim37hv87XFdBrCh2VGfOFJuT
0JBbMOtSnqOOD1MJmMnHPy7wI7t/B4gPs6p6RBKSzuICbIpp11lU+a6VfQEJ+obE
dTarU/DEEc/b02l0+n72R026PIUW0/sGrmtGMmQJCBmIIkieVL2rfesFTjaZoVjR
auMayDoNGg/RQlrREKDzJuQzu8V72861Nodmb2nUy/mk3V0C62BAdylSsc07rK4X
rkCyPlBj5p21tHY0S3YsvVZBJYbm42PkqJzwU90+GS7j8jVwNjFuUSWxNeM8pQrk
jyOObGtLA8CCCNH5BuxFeAHErxL/hzqpoDYvIWkzufFA0zGsXSCK5Ub+XROclK2f
NCzhpr3hXX9apXX5ErsBCVFT7+TgfR6WdyjUafRCygeFh+LC97eyZHx3Azh7tE0V
CbMjLT51RLOJy1ouVXVUeKPos7OilSVesHVXmXZM/9mytJCqnNJz6viZ7ASE4+H7
GrBHzALeubjcW/FgullZUUGO4wJl1PO+Yikk2rEDG1MmiyQCkG1GkQ4tw79OLsQI
atLFPN/ZDm84hj1yyaLsJGcIwHJs//WeSNgpldF2LwTMXnF/4cxlZBYGLUkvJen6
D8g11FtlrxrmcN4rkJ1Nl5JU7uURu50AZd1KjTmjGWTC5R99Y8N2gbvqHro9kuLN
7XM0VzJbLAZJVRz5J/kB1XIA8V8YpiDkVd5+aKveFGNrUr9MqIXf0NhdPzxKzPNM
bATzm2yvZud6/MQb55a6wuitZTCcbefTigd/b0Cbhx810x/m6A3j2VKwQj+MmJPE
JIm4aovbnnrk90EDAC6ueXSYd3UcoHK17YqUjNMbN7S66Lzl876AGjbK8vUqs4DN
btADs/kxQdC+hCCdF5PNBy07PKEPnxHr4XrVfjqTEeNX9zRIGzWjXj/Y6UD4Vbvv
9x1yoV3SMyU8JZkSIv9zuE6eKZyxJ586/MQaTy4DsiEGwJGZKe9jXbiwAdsR4XyK
2aeectVO8qm7s39adxbapDpuFncSLN/NwnOZCY101yVndoHaAX5yA7My2JsU1leD
d8oBUtaiiZbspiliWq+W4riHNekPxR39gmqGaE28bjZkVJJBOAfkYPRktveesDkW
Qx7tJwoEWrmjtiOIy6RLS/afiRNA/2qzT6BrJCJBHFXFKHZke1R4odFSg0VE1K98
MuqprJ6b807kyhDeDlPfquV1nUgQaVkLcvfRgLsl9PkGsdDUbtfmNCZ8ylpvHedI
+3o+N+sHWWh1jpLNM4gTP0BydMua7g/bxciAwpzbXCxq/2AbRjl/gnxxegRfXX2p
raf8HoTRqkfWp4H1qsrgyvT0BBMUvg8mS3AZIt1G8GObdTg5iKj9yBoVc90I+l9I
i7E7vqq0cWLdcklWBS9dWy3uWjtZgrlUfhHvIQWmTmCqXHaI03THnPxQ/uUQrc65
HzYbhqiF2K2npVGPrHQS+UkFJ9vKxX3Br89mTo9ZCukyvhchIVvh6vy4S34DKMkj
ri8qq0xc5BOlN1yMYdOGpHMF0khWvdbItYEMHZ86fzKNUr3l5wDYnN2oGRwfXHVp
2zCLFTBYyGT4wobrO2xyAHH73JupNPRxpTauRKOcvZNgpp7tkZLyhq9kcYMYcRWY
R1jIvOxHwj8CXnjFqBG6fjcpIrkVDpe4bjILgtZIc0McsnPmekhGfhoGYGl7p1YI
/T0rLwV3nwcyCcqhC57dwPBdkWbqMJQgwzderVOMGecO5NvaocM7FdZUEBIrhwxF
WZAC9slAy9P83u+1wErlGrE+iv5B9wtUXbOQR+azMsmpoDFe/wlx5aRCpAI0eyw3
W3Gp5Wg5QrZrNH+T08mP+8potIDSHqfKMjPPPHRJF5Q2lpH9uX/wu7EgYethoU+Y
Fjs8y6RJcHpbKThFHcNwuGZUVYGuWWluLmJOQZxUqnNzqIBCsJUaTJHv9Wc1nLwn
zKkWC15sFqO8IDElihcnwg3PQGl0Cls+SX52ZBjYu+4oT3to9Rwxs3ZLnI8c6Vy+
UXL6MEPZITqcUQ1QQn+/pzhMYri5AicIK8mkp3qjpWkBrzPxMKsOXFKWppKrEXIH
9hqW2cja2HsZ6AfZyOvwskaldgqSbsyJH7z/nD/WxrcA+NShdWSb9P5egUJZqJhx
lGOhidoUFPVW78MqzJr1Xkt47fEcCKbVd96bqGeTQjgoz4dHeoQFqvis9y7e7AZf
q+dnJKinHxLN5Qdx7UOPtu3QyMEuHVEX7P4c8h/ksqsimbdVQc5CxQb7u1cGTNVO
fmR5z61LLRArEKGxXSpmtx6Xn8OdreUooGnfwV4lFQVoLg7K1q0SYBmS+uLbFWE+
rFu/qk5xdWiB3SsTYQNeX9cG1G1hjqiH0I5FzAFXp+mQmAa5K7ZDBvWDc5H+oqbJ
IYuQ9clwgBqQ6D1tr2yTD1m2Fa+rOdUmj5tAKvfrCUKpdMpRBrDV3RQAZTtERFpe
H9KPVBU1K6kZeD6J3pS7kFYKzBKWxBw9wJ/h0wQeBku2oDQiYXB3Lw6Og1XiAluY
ykiak4FKwglp81fQo2dgSiLFhUwLMhjkLNfgPrANymvFZ0I3qWqoQm9p7JjKt/AS
VgP+e30gC2Q8VKj1jf63YIDFxImc7WkMOLlsqkxQ8ro4E4D4Nr+H/rK1JEdF4xXz
gUoioU7xyrLwnIdh2cRjTTkIBKn49Pc05I+0EgDwG6JdKJfOR3SP38hKbWSNP/sR
im4jVFMEMUU572e1lMqjP3n3biXJaKnDdN/cHBRdK+2bYn7hbwJbeY0goPmXpkOe
qEKQ5eLEja1wb8QhQRasNY8o2Ud1tvLV4Es+ZrzzCk4WzEGVQjzpLlghtqv1rjO+
BDAkAFjZwpnC+sBm/UfBNaRcB6HMILkn0UrtXCaOCnN/NbCgmWUufVG1w/JNxkxk
vHPqaBm1p69AnCeQe+A6MvWBu1TsGOrrBicKSljxZfbZhONe8uAo6aIhRJOjgduD
9D8nwjX4dqRoVZ2V9pqSHHyynICJqy8xn1JAYVQ2xz4LvAuNIfVKKPWI+Yw93p5L
r/Sm+EtX2YHCYk204P4pZ3KsZOHempzmQSWoll4rxZPGyNOB3nDMQsHLVxS9J++V
9jr2iK8t3ShLuPU3fWsD/8QRcyueRLwtXSoKqIcq8QR9J36GSYrDr8KVPkY+mFKv
dvQmH1tXtygWT80ME+AFVQz0zosVKhWfGIhsVKaDhzJXkJQwSlajDUTGE+JD8X3+
L+guLalZJwVT7oe3P3vQ1TfbcwinGr/SQt2rbpE3JbGQucT1/iLwVqeXR3jViYex
FZuMKsDfVAloEfqvZB10ABsiFku7evyDDJfq4wcZoHt9BvlbPGYfQYyLoLGKHRdS
2E5NVhtS5juKM4FyW1J/cb478W0orqwh9WZFm89rngQUI0tvfGLhnkVk3WhPBubn
tBcPQ8O18tRDJaMDXc4Bs/I2LujH72seARTRyhvb7CTvixpLhr51w+HKdqevbWqx
Yg0NrvpnXK9Ec0qJNny/x97LpAR9Upg/U9uRf2ZdYjnulCeHH5DHhgmtpi7aG+Bh
NxRzDmmnwYDOb+4CouircdR85GrggxAoaog3T7igUEadxyNxgwTJNRtCrOIi/m54
i/EPT4Oe9XFQhRMsI7Yj9/U5YAE/mEPENSMk4/EGBGd9gZ3SamxVVAEk/n3gSwMf
KSrLuFA6ecDd1Vt0RGES2oAqklNLUpMU4zjl7/eHhyhqvVxGev01wikp2EfL/G84
7olEIohEWd7bnK3Qvmx0GCYI0UyuKnnK0oDoMZJFYlwbfrom6Eu/iP9gtVLkaEzd
r7BbUORc3SMcTaPFWzoNZYeBD3dPYRjEksLmmNccM1yapj9ZMGdSKUUSPi1AnZdC
1AtCwLVJay5r24Wrqm8UQgikqMy4I7HTLYbtaAEhJCPT6ESYPwDt1ngpM3QefhKX
uJSPUKWmnTH/C+x5P914f1+PU1iiF+fglKSa/E0XGywwXROt0lqiTAOjdm4Det9b
cJtK5Zhwua14hKQVxSmkp8oARgOVhqtvvsrVojHAk8ocFx5szCZq+fkUZK+VqxG1
SOdsyUp3IHA6K/plPDobmzrmhoUaQKVJfjV2MRJqjmPdd1zxol4MLLXa3eZ9SDwd
Q7tKA2h3BqNCuYPHpGHhAxmbCkwoBk6iOOwtMQSRVD/0un3v9Z0l7Jm9ouV8HwZv
pHaI/7hBgbv5X2jipxrZCSYqRbVqkt1HpQsx2CQoR2Eo+pInDAOVyOvIZPRGt3ib
H/MHvLkA5e57V7Gq/f98npoy65tQfS+t+XAJrfWzgMspeOuD2nXdDmUVGtOVdLjC
28M1rh3uK+WPpewLojAwgWdqBtjwy5zRfgBHWhk9Ho+NqjMBPVcsTQG1ro2DWjMu
WTw1yIRU1sCIxQO/cDan8HeGSbh/RGAP2N2C3HwF6EmtEp8wf+a6chlSNiQlVzte
odS6pk6ko4KluB91O6dsEq9pS8N6Wb089c+NdSHRUNXnwd1qHA4X0kesJQKDmfIk
Sz7ClMZEMZ0leyHdKSlsF3FBWIUIePJakkQ9TUg9+IaeDynlyQ492oB9s/3L+CwQ
II1WjU1XmYQuCFCC9kLWKiMIJPXaoeucmYyXd7U+NgefMoq7q/6NYT/r9F8OsvZ6
5UKE3czVYZM0uFlm0bWcd5/sCrn/Kvk2H2FBkyUubSuwNO9npF0knozaAvYOpBp7
bN+pzTFxOmevK3NBYZLMUvy5mT0Ws9UVZdEblax1nHbZoXWEV0qD6Yw+UgfC+YxS
lFHcpRrzr2Z1Wom1n1wRmDMFOauRCMzi/gmU52uAnhMvD8H0GwQHK0vCqsGVa5Td
okAb8KnqRnIVYgP2m4r2+Vz3L9TdaF0qjCJIvousEPyK9xQZsbnxYS6AA9Z7YRmm
+1MAXSpz/RzBHpQCjvU1RJRur550YqUiZW/hmzCypO8PM3vBvzHzrMQGEj21WJVQ
X4uKTfxyI4B/mTk+z2s/KMQFC733OsfxErgLnxAjJ1T3knOYcAB2ACkVScLtlln0
q3IHHoyH1a1gA8APBYFkOZiAKxvagWxHkvHGroiXz6cMVNUKJbero4YhQ473UiwJ
ahjTyhDmzSE5bDwOry9hvxmrAFTNFKWwxH0Ubvm0ESaJ/lv7BzJd55O+C619uy4t
Ch1tOidNh+RFmYjnrMEToAbAY0a7ChZRetRp7sWo5ulMTsQW5XDeEzsNyeXODouM
/X2AelpcN/6fMwNHiSPeJ7LPBPAkOhDDaykO2mSKMAaOMM1QHHC4FvQydWm5gIxt
GSxFZBNPPrztr5NLnLavYwuxVYG/LHQBCxYATohax2jKXiOpQap6ncD+3FrXCZqh
3o1e34QIF4hPondxgs/BeVqGMCNRlCnjPP/OxFw0DRAgRqzMmGChqmvrMDzIl6G6
wOsHFhQf2v8fP7Jc2JPMukbuf9r/9qqIoWsd7ne+wdeE76vrNZDvr/JWsp/LSGS/
vv2GyRJq6rjP8Y+TYomIWD0kzm1GXtEMIAV2uVd+2kPGKsoAQqbZMBXmjsnUaSSk
4dYQYA5DII+4tZtac0TuKILpS5GkbTsvhQBxJ4T2GzHPEupXgcZDXcky8DEjMgjh
p0stwwUshEyso4A21RI7P6CbKZEWqQXn6EezvuMsnYSdO5NOh48Izpn7nQXsQT1h
ByBXpt8YIaZ0PRZHxkXhiHLPsg8R5Rus8Sv8pjLUi4vqqniDcZh/kGyu1QDy7esF
+y4W1k/yLEAA5E6FyYVfuNCbZYYU3PF+YySHcID5y8zRGLkCBD8bVrCpvbtbRqKl
gqEctojhTguyQ4znzfahOHqzjDRlUXSJWKtXw3vwUj7hhoRV2IKrKnIFNNejU2XK
gzYRdr53WjnhmW8F+0QOygkdUMpf2zvmzn4PmjrS3ZPtcg/nX261cEuMJjdiNdto
lSydz1+g9KZDKSyKygVPyX7mRkdzk6qoZ43SCjzHxHKMjIwKtqxrHAS1fR3uoBo8
nssyQ6KZDgRRj/m07zuloUTh5t6CFvXA8brMCRRwqAtoueAYLXWfN23yTyQac6lW
lSyLJjnmlRlyuLMhQb5OGlKXppK/bhWPa+Ga3YAoyjj+/Gc2WUoFjQZX6FLDwV6h
8wHtDHoha9UFKIdA7Dq/uOypkvTisJCXyJ2+bX8iYRlPNnfAPJ6qIs3YohmdZ+h5
TX3HSjbgSXfbmjZGV0WKlsDnFZTsWHZ0A1dSG5+wEZMJwqn1wmiiETvOIr3TLVQZ
MqzXrfSq2YscNlNXBciqds5Yy9bLAJt4VFgFfCIc9jBdRbk6S07aELjaMR5XOyyw
VIp/u9JlRhNILPC9cZ3Ywe9+okC6sIl3eiTurq1IoOFXHPeS/BY2bxtkTSSwjIih
gpCyl4ViJQIjDLkS1TQNAgyeg56kopKhzrJtpgXM/mwe5T8oAjyQJI95MhBiFCaW
Y3inYn3hR5w6kniyvurZkLDD0jjx6gZYTJce2f7RDj9xR7A6dCVohC4jc8ESTolp
Ixn+qbn25nWdGSgXbcTXt57mjoqetMd0lKf7wbOR+MXW5hOnuxQTHDFwKjJcxYAu
llsJIyaceZyqZvGomf06UT9dusZFDtTAyOn/+9dETCRHQRmfsPY7rBPSlUQgbwW/
A7KWAUIAJDQJV/zoZpdDQQLHxJjxz2hLJNXFuE9kY7hBj7rrfc0yXIo59UgofMqa
6CmgmSoC5vllZNadZ3Tv/DboCkAmX0nwcuQVqQR+1FOPmWdI5wDEvlRg1HrWODFd
QOyqX/SYIUIRGzOa3jdn/mALtrq2wUMsGk4v46uQvSM0D5OCElsM1q/nDNfybpLC
Lnp7zLShXBFfsN0X7wZDLi8xsPddFyCPR2k1EdLPySVdzTjklbvgSougX10B+p5b
+2H92o5WHB+5mWpt36XCbz1k864YTDXqBOGQFd1S5jf2vdep/W5Vu116MpRkjEUm
eg0H3LF7c2xW44JCsnW2Lur6deHc5wiO+xLhV5Y81IlYT493KTvpTU3VCOKYIq37
gk5b/HpUMVyPbaPn7JMqS+ENvjmu2ylHrrkUoJpCO9kIVQWxF2Ox2F2p26+JPzn4
NyR4/IDIqniVSt4rvcBkkIW7e05J/zBrLAsysMG0EmmTGlRkznyJREUIatnKhjXc
sWriv6C/po60n6HsBhBKcRbQkv3wUTKpEQO/UYuo2VDSxhMzAH0hUYp/KM/AUclp
UGm0BnAwrFutVkkyOWwwogJY9P4I/97gDvB+912ZgzbK4YSxntVGi1FoW3h2JSel
KYro/jXaAOhAEQkJ2iLjtheLfMw8LAowGgeFSPZf0k+jSb13wdyNZApnJ2qgj46e
sfJIphbKbRi+aoEA9xw4Jtc/+qQf7PeN1TiFYCJ7R995NHA/q3yPzms/mxrDmmwU
kyRtgo+ec7eMPY6H/IbFhMVhrtdrb/HtZT8FvVXYM2vq8j4nYbsQY2r2FNeUlcTt
w983sn5pyAmBnpl2CCHh0FCoCPnJY/neg0qCSvNPEXJamKAsP/0LWy+Ly8e+u/hA
VPKKDz36XnUKd0Y02lVjalctdVTWi97dy6V5lWEe9Nxug4W+KNX88WbgOMjwIOqg
Kv3yB3z+w8obAjCiFq8wpBC7H49LoywohCVMcZea/p5rgcqb4YWTTTGaxKJBrT2G
5zLqpMVL+SlMuYb3/GXKN3KjTYN5FKPUf/J6xigFLAH+CSiyt17KTExVji1s4jR4
Lk20y1q3wATsfm7qR/zhPHoXNr88b7NoTI8qJjpOY/HtG/mhyGyp57idgow9/rg6
JIhnl8TsMUOs4XW4vNlTm6fmmtqMAB+deeMF6EiCuznHfxgBnjLxTScR6+HDUt//
W1QMowJlofvE5/WSin+ATiD7ibXnEaaNYbwTobKcsgEPtvg7oSQS4EpDGnD9mDV6
Eqqxb7psV9R+75IeV9DNl9jeCbVtLkregaqmTizmsRjFh6NztUlsFDSAI1DsZW1b
JtUUyG0jY0r2AKXawidWxhVUnuaxeQhKF63Dc/bpv3BXTU1vy/ytT8045OZVVWqM
EvASZ9HtzLiI1kLLZpr3G1Stwl0yELZCVeb0/kVVYO3yIHKjZv+iY3DW/jUUmFcY
jphCAzYD8ImpFxPv7R0Nwz7TPErl0JtDcy9+fcWzEm77RMtfaebaYUegdcuCmmQZ
mgQYq7vk9NsNS1q5Q5tbXZYox9ZR40d4UMAukHgJzebu5Mi7lL7t+o/Gt1Pn7R9f
uDdYAF9bqV8dVLn8EEmq1ubGA6QEp+kaspT6L1U5qSHneuFMYR7s1rJGtXp/RcNV
JILkfW6X6q+2i9pxKY4awYeP3LUmRxxIi9y6N5ci8Qx+EPjBWlvtKHC+v1pBl11M
axLfDpp6NVyqTRk/tqYJOtlulOqksGmJPfcvzuBpoOsP6oAB6VguCnk1bX6v0QfR
Dtxi0FIIQRd+gcsgXmeSRlM8Pz7Kk2rRl1kETACNKs47rD88rLN8maHPoBOJZVGM
EcFC1NAuqQxSPdTBPBr1VT9b888lqa/9Yu4fo+GRdZ7bomc1rLwzpbgMPQLGjsBW
+/cFz7Kcy4wZhI2WLY72pUCk2peVPvo7M7HPwmWaL2zKicRiNjP2J6TV5jvg3DvO
gJRQl5sYCeYUyhgHrrUWxF3sZ2Gj0XROT0xAcyfRdcKNNGk1KBlalkktM4PrjPNJ
RgMlzaaE2DvJg6x/WBNm9MKDlTRpijhVVo13HFBYE8PDMCTOIbSteYG9t43BIRys
LKKHhcQx2UjmlAayN0PK1fW4FFRq2v5z6WwzNl914Ey37k+MFhn9q2klOr6lkPLR
RZ7AI/BLSI8XNRImaZaFjHPwuAyfLlLM35XlWROF8KSnArFC2l0l6NbARFQXYNdn
GsMeDtMNMSeX4QWQdIUPHlw+3xUb2ne42Hx9/0vT7HrCPTlieB2sxQiozjawap8w
glwfiH/gZRQ5l7mKei0hhj79NUxojvtfGOmor1I1KctwtYqGlKRp+xF5keh2q1ss
w2JTs3keq1jMfyZJdW9EV5GD9yHgx39DR0MUZ52p0uclJfrRP1klfcxBNHYBuzjp
wEHsr7Owi2/4ikQ95gQZgM+9g0BtLxB+LPJD54u55IFk8J+LP1CrGeN5t4tbQXYc
vn9ifJFV/snUTCNMJfXx8KuIbD5e40bM/Bib6AmuIumFMGLEQ/HFeVcS0gT2AKMB
RmYeeZvj5HgwD3rlhY/LtyyBVrQF9ZklZRvvmSeHSsQ5bPH0TZd4sFgPmYg2XFhH
me0xm0u3RHb9pFzF9htFidPbV8idWvCTXcvadiW9IpulNCQVGAnAFmB8qg5yWw5m
Ah+BNGWx3wTzJwZ4kXTuqJeEk2iEXpaLLt1jLL5tm+W17hng+SZxZodjFqGrlTUT
FWWZ9mQk4mjvnLKrPCawMOP8KH3H1Xwj8pS6YGvmACt/3mYJTrN05YFETCWuOyZQ
j89DPi7Q+OCBnhbIoU67xITHldpt+I2PAvz3U8DSA1+tZsVZtpqwCy+Kmq3vECql
nmqpcSvcrqQuYQ+dsT/GwvtplHlFH+b6j63RZdsQ0juZ0ilpSeQinVg7TCxeuHOu
4yZUK70td6cubxY0g2O10GT0jN/MqO83dB33LBAWhB+IKWowW40kWQK2/kSrrMAf
yYFyvE8JHrYpFPJSYgIhi2vRZc1wqZPpj5LKem9Z8IJGraHKurKEpp+qpnROuHdF
Bf7XJOp6RxeBP2JEmrlYXVzRfRFcTr88ke18X9xzcU7FvxNYMcoJ2rZcnXoyHPEC
8mhgmulNsBlYBgW7zCD+JeLvvYcDQ6RYGMw7sIa7nvnndfTa3PYLkIVBaCVkLQjB
OrDcC+JY+DN2Ub0YBY4xZzveRteb0FZg0EhfeQe8AR3rcFRUGUC6+kWKdugKBi7A
YvqV21xS/z62OeRfDaVRjJRiUKTTw07/GZDL8AZ6YExHQpluHyTebmsX6pdJl6Zp
2AKg651taxso6fVmUY5rB7CbDX6vU2FGofrknAPQJCibDLglztDVcHHgrKNJI43W
hAB+YKbJszCMJTPlDRuzb8gZ32moBXvnmhmPax11y0EiNoxG2DUBkPW7cTLX/yyD
CnjywNvWdoglskt2q6PpjiYfqx4EK3Q54JiPvEcR/fmGWZ4pb+DdPkX2TXmN08In
LAFXMLJoGflKHVnWu0VQ28xsks4PzdKhgsNfGN5Au8rp5tZtZoSZB/ZE3W2ta6so
pbC4iV8gUPa7yyYGY1bZWjqL70hDYJwZjrE37Aw22CxG70FzaYqzULw/ugxOQwyE
hVPmhIXBbdiEZFiPCdwn5LBMsueVn/okuApDeKQB5yhznv7KWD/ArIpQNd+/jJND
BD80jxXhb9mglj40DnnS2EIVgLKl/7xofMc5lOec3J96yZ014tkuKATM1PZUwbw6
IK28PDGq2KkeE22jy/+pa94Xm5OY1Q7E1TJeLwwW3kxnwAUVBx/jMkb0W8uNJ9wz
ZYRbUCMQE9nqaXB0DumHdJ2L/utS9X/C43P+Q5wMTpM/Mkc9dEfnzTSNpDPKscX4
+KehqHl2J5rsodRJEiTdXhzQsE8XICXWGn8sm+ybUN6U0WRjSsannrDmEr97mEMW
K2DM1G63I8DkQ0B4307zx5HFYx74twWX77rvxZYQCWahHR0cK7TueuKyPBgI4wKd
wor5DV3dglwOBHeb2hI5GHajcHIoQeffkXrdXa2eq2KoUVi0wQus69B8W2gsaE7H
u4qmv0BVpS5wfRzUy+eLUnbYEmwp6auQTLZFNSAVYnOP0sH4RSI8ijykeE5jlF8k
4FendMlJTmhxAMsSMZcNwt34n3EGpPloF7SoEMVxBqKtieoS1Lwkn8QeKm7abjgP
lzAGSmUhBICWV8IfCGGG4iiIiOb9CCbmrfDPIaZhmjemFN4WA7pbnh36iK9epBOK
1JPd9Womaqyrtg63n60A2b0/eToRzXmHmYBbwzDgteCLvauWFPNFcC5/2pA8q5zB
P3zC1qI6G52Uw1uCR3MlF75th73fYeIG/xDKRu3GLOj9q8Ln52R5MtVcG229aLv6
tiWLYWE6N6a76Hbjx6jVxjnDofhuWm/qg3OXTE9/l7929nKwwdYFXABmHjR7HXT7
KTShaEd7/eIGTKnszoQcqc5ahUP357tEBXLhypOg5oy7m4RbWVUmAodemxQMCelf
mjDwcQygYAguyViaWgyRfWXqsKoBwQkhCGi4jW6QdX98o+JkUi6gtf0H00HCOyyy
hdw+NtwM4br2kxkNeShagCMBJDKDBW94lJjMG34A2b2ANcQc0UrQbWkXjehOnar8
0ip4qm7oQMZMG7FXfw3b5rR0Wj//5t8HGuQbc3cKKZ35ZIt5XzYUucT4fP79r8Fz
j+x/nSQQ8Kh7kT8vl0S1MRwacMqUS8/cmeJIxXQUKtdSef2VKN8i7Wok0lJbagNH
CXoQTRTGk00t5ixXkS8AovhFtYEXqON7U8CQa01pIfwYypQA1rG75h95SjoLPBha
A5u+grpiSFLP2ViYx/P6rSGquCgZ2adxL2zJKLzsPiKGuxqBXgVidXf2M59+Uy+z
M0czSmiCgBKLZyQLymzy0YD/vJcWa07fhhgniH9t7fUrM+JLqh/10PzCmQmESGue
vhMO6SY/friirhgZl41pMOL581DNQAchdJPwewSEGMrPrBoE62k8wDdU6f4y5UZo
0cHIRzbKLWm8mC6+llyANQhsB6XuyeSxXq0GlRdPO9WwzGChWf1UHpJunBv+3lXC
+a3oWXiGLX6076nwdXPqjf2q2LAI1ENYyBI+70avZrGH0qPXIr/6p2YAdcyJCIg7
4jM4G4XnLWqvPtNqfq+7b1fhJhE4oi2fRyFdLRxw6sabq317n6YMjlelFtgIxH9l
YPYYyt6pRxOp0RvQu+hocyTViw4eJkr0IW0QpraXF93vAC/ZXIS6VEDrd0l7AJlU
g8NAOWkJRjzEIUnkTAUfj7MhX3xu1hT7ZEixW7VNr7nwPW9NqO457PJG2VXiG1GC
O0QIAI0WUKBQ6vQqKCp1wZAqMEyT9Bspb5h81O27Ji+t/WwptBiHM84QTK4TihmP
ME9M2997UNlH1Fn5UCUqebPUl5rON0tiOYCeVnSf0H7hE8dmjiuu4hgQ1aVOdWrn
WhNbrDKZKQWfZ6/ymrFVwtdAokfUA/T0TfIepY75rZWDfi0971s7py300P9q0/gU
/ly5XeJGGddgxq1fa1CFL8nEfh9n9IKbR2nZbOYsaGEr5o373p6LodbnunnrEGkJ
re4M9FWEUJxj6uzSFC9J9G03OCzYCxkLAunHH19/bosVZgx83Bg6B/rl23TSMA2B
wims5AJpqouxAIqsnVeBJNLaJpqobuWJ9K/4r3VOEXEsPSp9MglZLV+EB0try9TQ
fr3KkFpnohsgttngDypxlCIr441RDXr6TYfT39+Q56oXXUFfDe8E4f4OirJDHLZW
0yuukNgSuhQW3ruRY6j5kfiNL7I3UHgDt8B9p8mf5fX68O7+62iEg0evkojPavAM
grA4hXXuedNUGiPmn7hk13V48hVPAM2h9Zf7/Gr0h2RPyPtdVdISn9DfmqJkmBwb
546dqmxxNhzYoG74Z8jh3lAX7kGwF5HPT9ZWobaRUSZy/PpQ3a1+tdFFiHGQzbGy
KpQ9TF32CKAqdhw2c9vp3hx6bZg6N1e/KdIZ6xJILh6Vkf0mxCDPMC4KSDAJ6TGo
TXWMv5x3VZBB9a3N2y3RgZjp31dD3HrVAPkSacVNykkt03a02UtEYGZcoF88DLGl
/iFDj4rZweSV4VSv0OaCyi84lFA98SrcroMkGqLjGFWSMugI66FfnUBWlfl5qyU7
E1rtt0TFH7JhcJZOVCzjllrYpg51M/7WKASwcGEDvAn7rzOOwYfCPOf0bf2dgh8p
Bp/PNPBZF00wABQYcG8njxoy1MrgHKu4n3/uxQ732NBdsjK79kFDwRDDcEiUFKbE
+v+xSfGPLZW1E2r3hwlGrbxLEOG4nt6X8mj/f8rTXlFPN4DcMeKKdOnsSkckwCHI
BO5xfk1ZT+v6WbisGPxUGH/o2vRmPv2p8CP9G+OUPdZfDd7bfMBux4O1PWrJEyNa
tn0r/Gi/nfzAUjKCR06N17PodZmgBNZXBHE3rSjB8NABfF+LHTzeYgTdY2nI4R7y
PJcGqgM3WFE4QvYUMSpYgwtrMXvgIxaHWGn1gipqzpUDZ/PtYKS1xqPVyrChMwMo
PYDKzEN5R9CGULwKcB2mvHqlAoBX0cEoZKVks/BtN2E+vNETMPunzuRbPO+Ersrr
BdybxOhgYUFXmfLKedlX8AWgO8lMFOPDgYc27YymA3YXL86mk5WtkgauRQ/QiBIS
6muy4oJv/cjIMWy6vbrgNHV8n1pojJLghUsM0OPD6rvYZ/ZF0Ar89mxZo6uoqbA8
ibDgb7v1vwZu3zyQq+lPA3aCqsyUD8KoqzSDDJLIvI7ChGpOItI69z0a+YdVh2zP
HDIDXoAmAu19S7QA52JLtI4OQAPUlwp+Dcjb3j8vu8cc2dWb1erfDJDe2ECOLdCH
FwHs8k7CIyuwvaT98lQt6OsrY6kzTbK6g7JUD0hIUY+N0var90iKr1ShKj2JQ3tq
WpEWg4v1I19GeVOb/KDNopz8Io4LW3ijE7rUuYfV0wUVWjTGaLQZGHPsoSGtfvpK
SLfO6FmNRwuBcvcoWcJ/iRUz6qxvZvKkt4F75O0BZCdMJtf9mx6tu++N56EzVLjY
wVJ8mZhxVazN/vS92e8WV04rVXTeSN29qKAkC5U4KA6ecH/VrJoFn/rcx5UutmpE
BYKTrxpqpxseSzkFvcW/e5QtUrx1Q6B1iC9RnaAwVGsRj9nHSYjPohaUh8LmC9SQ
0wY6RzlhY4RS23PQUtB/HAvkt9dXTFTvnJJZSeJ4FEqy2XShk+uVmmjnJe8mtLF+
0lc1FB+W6ztW0YilMOwpUW6xhmII6LnEZ8ygnWnZhzabmhMVYRPL7AmUQTxFVire
QQumkT/HIbG8J7SO3wyluzimvXJjhytUgRq+kzF6zaXjjSQdQ9F59fui0X+l/uUo
S4ghjpC5ZpcYBJnKZ1uCB6YMjKP4Q1+jGDFBxFS7igIueyn+np1tfrsupocnhB7Q
OeMU1vO/wJNhgUltLj4ogALuio8W+KcBxmTwuToCCJukm0GDAunTtZoUmfb/PJa/
X1GH5OkJiugb67tAnQSAmnyM2jh+lF2mDSzw2JT7kRQEA3RRy4gdc2Nwpnbk5DLg
UmKPYK6NAXJi5RgCNrpMZoikfY0b3EtDwmjVPBAhiOboZEDQeG3dQ9jV2TzqdlwJ
levaPHxHcO71n6J/ecCGbqp7FFSNw9N3RZTWWfVx1U+R0Qf9B7CyBy/qxp15dY2o
Hx4nrYkryH3JgFRuOk6EM+luX6yc+oZRaqoIkLymwUGP0CVArXEQdid7Ei6kNbxk
S6Pi7X1OZ+k4JTh9p43i/IQvmmKhzj2iqKmWvJRXVjdEiwHlZv3zl82LHX2Z0P7v
ZI8vHCq31nnnH3vJI7qQRGmTWpD8sLTFUJDsPyB1KdVnlOyHCjHN2jNRKs/lfylE
5AG/Ek2jV6dqmutdXs1qeVUB96j/E8CGH/pp7cldkIMLt/IeKtkNY6M/AWLXyDuj
sw4elmhYixllNUEPRKn3JwKDoyIQEJZ+CLiISInBtQ1trshTBEJ7QxNoc5wdv3AT
SU2a7oJo8otCkT8xDKLz7kkr85HqGriLw9+5ez7kLqgC0Kk2GDiIfxHaEnyIaEvx
sBwBj0UTO8yUJ3e636MbvjB7ioauIGfpOBsFWFxmKh8RhfQ1kPAxQltx5PgX+xun
F1GN18+BPiErGWhEH0iL5x6Xj/nLXKIStxY41FvMhT5o1Txm7mp2iTnGyT6GzsWn
W96KAZJllAONxh7JkTxvIChd8rlw90VRhcoKQ/ViX0xiqnxae2akINNcNkmZg76b
RxYUYBoxBcegt+fbvidR/SmOv6/dqwSSHGjGJp46JAw=
`protect end_protected