`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
ddtXksX2+yylW5zu6QL2Lhnb2d1sD00763mmSITNX595NcHTEkwn0zB1Dry37fOW
FufOhVzEJp80NC5qZ/+F0Vk7Ik02dIR0elf3clrjeJRK85K4e3Hoo4xn7YbFUIms
l/8VZSb14+JVGURjfswrIyCUotIzlzVYZ6gzoZwDXIi5gQIBf/gI+KxNXPaKV+PQ
Ufys/12rjO6aI/pPlqSm0hCvftmBcnezN2hk1UeXgOIuKZnogjOsf0iJVX2aOOWE
6pD/psybjbnsNB6kH5uFTA5frkzIzkzl5d9+YDm9OyC+k84E83I/7/j+rk4L2dah
QJOvksSIzN867/4Qt8qYTQ==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="MvBXkzurAa5VTw+1JJ70nePUfoQXBvZOku/SMmg4TwQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
oRtzZL4VJ4iwysPsC8SXYCzXS8Fw2gtZTOskLcDV+1B9Nzn1zTyNtlo6lNICRmmK
ZRVu2BmCc2G+fmzynYlNTnSa7C0Cuel6FYpxCBlOuk3OF2tzAmLAuDyOH3Z1Yjzk
a0aHuoCdIRKv7BrZCdALt03JeUmXKPdOmIlkVGFl8yw=
`protect rights_digest_method = "sha256"
`protect end_toolblock="Jn9CQpRhJt4rnzZPRk+dOpzAubz7omckX1MrFd4p81o="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 39680 )
`protect data_block
gD6l00tciPUa6pDNTk/+t1gcgy1iCdpjTkA/bOvU9JA+cpFEv5u/7dp25hHk7lLT
6tYtR8HgwcLXTcx68BnPlzdPHkVIv0lwXo6yhFVkYlDWBcqD9ubowgKij0UjlXmV
p4anbpVt/gKvAYRDYe8Q5F2CQ8AIsxOuOcJ2vhCPchS4QF3n7+oG0MKU5ZyzxTu6
4sibWTVQTTYAB/sg1MLPrtXaZ/HbLYmSa9XT3n70aJlqofFi7JtlzwZzdpCiq9aP
0xR8h6CgL8RjsaFZUkoR2NtFBqIUR9HWJv1IMihbruYk/8LIX97zN2tWl9/uEXyy
INJErQNQy8wQ13B8Hhg2Z8sqBJMcICtzeTjXeVYIc3h4DSb8TcevXu0KhxTHAsCX
qpHhq1AonscyOHSd7K/srxY+1Ktng9d+KDEhvO7R+t9RKj2G3kH3i1i/uPjnzzle
KOacFSuMdZqf/skTSW0J7DTv9JDoo8Vubi6r3MwIIXksYL1LKmLpzREpnd5367wJ
EgzFlWLDwHZ2FkCsx/qF0qvxm2rdprxvpquPSFi+PDOGCesULpdgiASRoIWYRPM3
Or8LIuL7rC19OueUHWMRcybAN3fhy+81sKOkk/lGnUaL2lyogU/ynGg6rifqaXyK
t7NmqWV3O3I+m6cM43CqB8AiVeUI3VFaU+eqAoE+6Bh2pSsLkOERPc5+y1dYnPzz
u6y5sTXRUBVfLN5klNXa42+gjMXJGK1mJrjGll+xcWsr5u0JCDxpNlXkbAjYHaEH
kM2ModPZnmYR/E/CdUTo+IMopH71uJ1/29jbZiB5UsFYUY4aXT3wQsyT9e81ha0s
ZDtFoei+t9tCBG16MVSnYvRjGJBDod7mJ9Y/onXJuDNP2xSZkOYKSewgV3Dayi6g
GgBCF16217evlMod2ea6std9NA/vORBem+e+3ram85o/3flpXpKUenaN33vvNEWm
6dEpDj2P0JVT2nmwRcyb3i3hd/utfW7J/Hgj2ilzG/ULWUQqdwJAJZEXHcX0rskz
jTEFr++lxFLr62bpFAdrKOpcXnMg/XSY0lIUVRyxU/ilebJvGUDkxv0F5sckgfaJ
tODSzwNcJSyxLisd64GcoUBgnpRvkFO7bzc2gkdn5oM19yukrqtbvw90wHvp2GNO
owlH+Ua0VErtQikeMrScviD+eahuhnggSxq5b15SR0zg1snaH6MJeWKB8DhhSzXo
CxlTp8piv+8qIiM6HbFx3qSZZNgaXrgUTMh/s0u2MPC6zXUtNlU5fvk0tQQstpdw
qOhUlfkRf2JSaJwPT+KXgp97wdzvzSfSDDzO4VkejeRgsP+nHcKIEApF5m0fRWgf
J0XMoS9GSIHg4PvJazld54BwsxVgAaxAUAc/QTsrjXa6d+utsO0c6KB8xcXST04V
dG9tu8EEHVM0Qlgr/+9L3qU0rv5DG5IYqOtgW++vfHT9g9LGwspl7A3V2eOku1Bu
Y7P9q3ECBOXREyq0bctd7/ZPBdZTW35wOFgylkoMm0ncNZrF3YwCqls2puxOHHi+
UgLQ6LTqcezij1bpNqjVrWkS7crX5cUzfZ+iirmraWuLaYVJeNxlnvS1kSSj/Yrc
LBqqXt2UYLzwIqCeTGFyrn2WauzPt9Ig+tPa0TktbEdURB2sRBMLlpWwlvQo2r7h
PAIF4JnFuv9PaTR/6Jpc3C51Tcj5P5a46z5e9bFQYkmMbU0Dhhfpj0S2rh6PoXio
jjv6fHvMVjO8Gz6dWHHI6m8bE4ENfX9qLf0FUwYiXMnS1UVkF8XUZR8koHeVnWkA
Lz9TnPqzjLgEBNumQrbYxDvIiGQYk3aIR4zjLOH2XDKb3fE689lbN3ikcQAdsh/e
Lk6HLitOB/KWpTuJGKBroHofBMdkC0ascKSmYsCvYekGRrljNsg1JWIyTxFvPYTg
T0iDtKYoXPap0pN2Y0GRA7YJs1Q53/90cOpbmB3oxG+406TwEZQt0cNbCTA5sT82
AIRBFMscrmgieAAaamfdV6Luq9ZF/HrYd9RVqceIijkx47Ub81cC/MxrnmwjB3zD
tHa/IjneS/B9OsAv68xty4ijfNgKU6enCOE4YCZh0XWTvdgOF8WFJdeG/HHIuPNd
oMx5+btFrdd3nZdKlCLRpNX8+9cNK+kqbsUN4SaJOScwJcStpImOhJXfBTxxFr0S
+kfs4e8hmPV87JxQrlr08GHKauSheL9a4Q/p8G6lWwp9DJhVQfpQyVb2hBsiTrJ1
SbyfO3VWRbnaVf37+bY4Ikq1tvxzx/SWzBjhfqtYzv1ADn6YbzIMfgFcS7jYKEMk
CM6/7f8kDmnKFFEENmCbw/2wm3xIq1EtuGGm8rdXReVyNwcmpaZLYX0JohF6fSCB
Ii5R1GUS15Z71Fzn8YU6feKnnlpU6R3/ENNY0h5MAUzUkQscI9b80v2/Psw6MhmW
dMqyDU9/OdDFLW7kK+60YMGkkB6BIq7nS6avPuWRXiDQ9evEq3k3ZM+pq3gRrJGp
+/pBRSyKjWybxX3HZyFB3YPi3b7NoWYiZOzFpQaalJQlkkr6wHlZnCQXLUO/4i8s
30SKSOBDT6gMwr55kbkSiVIgOh4QX4Rz2h+7LuaYmhvx+30YgPcckbLy0IE2WYEs
NORH9s4AUMyQKO+eCtK96B2EHDKg27uVJ5jL+vGtPM11bic/V3vvTav+pWT/jf4h
LoNOdQe59bfpTPRADMwp5Z7/IFDhiAwXERUdr73NLh9cmvXbrd71iomO3kte8wpN
Y24YEBOct1a9Fo/eY7mvT0n+ijfJjcxwfvryQ4MCJlVJm9LZosALAVFqVp7Zge26
yZNO0y/eS7QtwYsxtV13jLjR9V+3+gIzJV7P87TgOhfU7n1btMv6UD4d7p8et4KZ
7AcowkrpLiWDRGiyMd7CJ3+yWH7Y6OAd4sWNcSn30brFS7iOrRdINPRCU2XzzVZ9
kMJ6fEF+qX9yHFHQ/9s5JtsiQaWEw1jlxPufp6Jt2iOLWVvuLCL6tJkROhzpBvra
xDimiVcHjpOPApVNgDZgF7y01wYNILmp8DaBryN2RjYxORD38Hzu8xVDIYE2tn5R
WIVLWL92A7+E9s1Zcjs8gR3K2jcx3XcBRdHZ56UYTzLdqs8EK1ob05sKLVcovqkH
3xdgdOsRrI0yQCNIqK5GcUDeSZ7SPv2brKbRaTa/pt9sslZxg+DGts9U7JIMNZZi
w9OvWmSBwagDTuoHU8J7LP2m5CbRezf6PSNYE8LZnj4Qw+jcKqDrJHdGrt4BXTQz
YAYSC1PKbAHLRK+csVbhg1I78iE/Ep8v6SIwWv5ZGSBrGddmZliJG/VhRnJ2q5tM
L/VG7LY674+eBpgT3Onswm3lgslbmMRp01Dsj2Yk0KCotlBhrUh/dH79dbT29qYL
BYzM7wU1I7o31m4UlKTRs+wi/I1LR9PlSAXXZUG6CXn55yt+Y8lZ/FSmkeYMV9Kx
AojMCtvp9+7QkZx5umHzjt4M+sIrNlEPqSoabo+h4B/qf4rB5ntT9PJRllpGY+8u
tH7TyU4I8y6FcKup1JHBaCJIp9IpR8FReU8GOF/kKiJmchZKW43OGQp19o/MuS5H
KTmyTGB4P/vorQALaw/BhHWFJS2dYLs4u8KzjlqqWzI5g515tG0+PoKn40JqcJf+
l9jOnLJPJsE/mSAIcEypusCfHcx/k01tivSDg3Ph7VR6bmVrW73ubqbU/b48LfSj
lgnyft/sHfYlcdddCoF2uQEleMwNoDnfPftBdx/cDsJXs6RGNAUTOerZtBhFVumA
qj+owC7WZ4KLgjb27xiIhywECm8Mb999KAFhiEp/p0zr5qEqTcIAqAyUpKyRrY5/
pEK/45Qfp4eK21rDtPO+v/as3ZTCEuyIDzkKjOMRso0EgHy16Lc2dh2F+EYBs6Dt
K6Q5cHap9s14iMu6Sjh8GaJFRLnCt6jkNiaa1fywNGNmubRp7M6sFymW1GPJTaBA
59hZL+XiHxjoeevphCPQg0GZQSzNJmIIeElX8/QZrRkzMGjIOqsEbIruNI6sjl2+
WGFGu0o5Pj/PKOU0iR6HctncOLhYtHmjwCKueoG5hc1+TMhflSfZcWpTdmWwIEdZ
78g+rvBYYASSQV51MjSFN4vcK4SZSq8wq1lb/S6736dvUv4ly3Gy9nLhjlekcRYX
L0C18NQympPjAOzvokLnSJPnOvx1ncfz//jdyHrh8FmsU6fvhQhcoTJkepQt3Ddc
z1o6DjOVKByzCDETK5N0tQg15pyEeynX5a6QarCJBvvL5vdfO66LsC3Aq0/pJWud
M7F342HCOvSb7lVVefPi9oB2z1C7t1mCkd7NP19TKiaXEfor92k7FDXwDHQPFQdt
2b/Of8BY/ZUHJqsxeNimSaVU2sosT+YJwJvOOon+jMW5zXFMRpHbKWBO2dAeascs
Sw5n48ee0nqRv4lieRYCpwzZ4M92V7C8vWGNiuC65Krww83YSDSpqdA3UEyZOjBY
Nv4lkI52yVe4/KdORIrx+Om07fqJz+Iqcz6TyeOgL7aeyIROg6IZNb9yVA+fhCXA
cXV+57Pkxlsi1SGc5nZIX1t/C35Shl1CdiwIx6axR/Z/H8jcxSgbPwyXvT8jfOlP
PYk7Lhra++3/3lzCsWZVdzAqUoqmVYWSAqYcqV6YzA1Dxxp98RpjD+MIoD2S8kT5
MgqWPgDYRkvE0qG5BZ/GR1CN4buJiWXflTTfvrGWM7juMDOUp2huLX1XIBdxJ1d9
sIJOMkvgsxVVtIs/UgvDKLJ/lgz8fS3+mtP9me9enniRGa1PFK8Hn8+M9VumVp9r
avx6LcQs44b3tyWzdx5XePw1icRRxD7dSLIfayuqlq9Gwmpaf8F4MjX6qJNlxx39
Xdzqw8eFOiWissaUQGpAi7ivCRbG1hFmqQlOfk8Fqm8Z7cIEiA1Ab7aFWWocMC3u
2Mtc7yh9kw9lhc/U5vy6RB8j+hg4WnCh4Iwfkv59LB3gQJzTH7aj1nV0CKzbS0hf
hNWlE2Kd77tgn7XQoJHbyb37Jflob3XZv1SvuM816yg00NjSjDCJM4wnHqJmDaxM
+WLRTGYuJFU4yC4NavExxB3vH0v+bmZE2SeaCvcEMka1bcaaZQolEeLQDQxl5z2k
Yah2ISVASxrVUhOLO9C5wNz5iurseQVooRC3O/rEDsA3hFqWjh+JZL7MQ87Qj1CC
9m1J7DOBz9y+SZ0LnqQv57jLYBzlbp/BwrX/QPqtsEcmOJFxti4X4eoNZPZhu/LZ
a/RerijAq0A64y8cuKjYsSLJdl6LzZWYAWB9hMsoxTrPalGs/l2gbvYPI4TShwLi
XKdQum6NLX+XauDRhDECVZt8yibZ+GMosLSJP+I8SoIzaZt0aV94U774yEXKgB6g
spr/W5vANKAh8QaTA7crHDD/8WLXMSkD4MUpE79z79MyQxzXs1J/72Dob3Q0oQQR
DWeaLMUjKj7v4h5sWNReMKUqePfqGI/wYozu7OaGq/DvrXTGATviC32Hl6BsX/J0
YIdzDXGjfYmdNUI8H1/3/GH1JbudK0XLlIS1HTdKa8YKQEJG7ENhBM6fj9sq9miX
HrnFvgwwjnG++nQ4k4ulkkXy0p28of1Fe4VHY1d7VyeiYVpRk5Ljso6MrVSdskP6
xT+RzmfFQxmcoe/sMob8GsMOadgOqWYCFG1nJ05fsjV1C8Kxak5Esi/FNf5GBZtA
cVzrVvrymBQZ30gmnTjWg7AZX0qHebCsu0p018aYp2WJtxJvYLYSM0/HDldiNS9S
4MaY6rprzN78jtgITl10HZfj3zYhKje3hd3jJP6yQWYCvYAlRl9xZXIKnLIzIswT
uPGVCx8roz4a/D4+eYKZpUMkTHmNgJ6X6/WXjbGWIVn360zXAZy/ppaOi3Gn+8kI
tvpouo4Enx5RwA1FLE9xWze1jvLkk5bGQv8xSIn5ShOfoTjO3bGadTnlcQHeXKo8
zJ+4rKoyNsyr7OIVg+p/SDAslzmWOtMewtkl6hhQlJvd1BPpk6FC4JlZgTFGnAdY
r2WDuKbUI8M51D/XbqWPmwi0zhux7DytT6y3Z+gJstZYBdtI7wxiArocXbzxCpKF
s15l8Z+GSfkCkw5IG2jMF/hMuj8UOvn/Qdh3CHQbVDb+Mh4qoZQc1ahqmIbW/x0m
9jicdrHO9Ndj7I76Cyy4Nt26x8StdXTX+7C4eK/sGzk3to9o95+pPJ8Sp7Jxjvbc
TtpcrXJN1GfmN4QfvkjZg+oRPyqmBWTqfONt29soh+huhYobFlAtT1N6J7nRUlka
JlnHCfwcLzlIQR7a49soc8YaqTAz3uOLr/DJ7/6KmcuiVE7X98U8VxEKb/KnQW+H
fJMMo46ji2drIYz/u/wk/EAQPtUbxumNce91ogrH7CHMp8UJCbrXv/gS9Coa3Zlu
Rf2tHMWgtgkFW9KlmIbjb4503aG3X27ze1cA92HN00hJbQ9rbFZNPyyfU78XsXbY
GngX4gJnigv1tXpP7PS48qmtR7Mr9srK+1NwnuRPwgu2DaDNNihKq+FbArlX0ukv
Io7MUa77SEnLtFTHCPAR7cteY17Ds6xLSqkk8g1b+eUQmeL/ZT8L0R79RhrJCe1x
Eshokikvecn0RtL/dePHQmkk32lQ/vr1mLxzFAsSNxtCK1vIKv9jv3xgaKhaL3eh
bQDTYr7tEfVL2Krll3o+jA40B6Zb/rw0iltYbBw5465x1NMm5QMUJJDppZ6JfMbl
mnr+rES3WGGb5mho3HhPw3XN3E/StN1fj4qitmJbBuI4LWhZmQDxHgQxqTnbXt4Y
msnT25tsf/7UX+6TAo01pk35b6dZ7kOwIopIaUWHSkpZWR2zdj3WWJLfD185e/dU
cyyDzKpzlClNRqd+KRt5dgVFOQmKFdzTGqqgh8L4Eq67FMSSSYBdS5AEb5MvIN8t
6yAlo9IJM5IafNC7SnTGRXe4ZoWRZf9K4dTRkNwkiXYuz3yeBajTgOb1BQxVWojR
VIiEI9JW1yxStm5G22AIYGGyKOsn5KwMcOoSyk3sDSFbAjPPQXyyfVow5pZSpm6E
H8RKkwcmIhZXO2UU9h57wG0n9QVFkWr38H3NjBJnr3ZKyOjDwgva1yKZMAxC6ob0
07bxD6hQ2i8oOl0i4/csEl4z7RVlXkxyznlg7XNdirqb98Jtyu1zrQ5ZIfbi958S
eoCJxNy5TNt+7FWcV7g/kBUb/92MVLjZVMmPcYzHxIIQaTgmCDN/nXK2hAtS8TAZ
SrcuufKR9Qi2ozmkXTLPzAtgfQmGga7DZJE4uxUvDXIDilA/jglTIP4FKWp5FMKw
ippIwTS8LbaqlKfun4++flVZFUCLBGBuqVUSltjnAbevzvdNNkSgJGRIA/G+V06f
wtTIYAp2IdnQ9KslQAWZ4cgqdzDc+CJ/zkTCkKdkSwys3LJXx5veZcHXyeqss/9N
dSZdgILvVlfLLiCQCwNGh6C73GOhmv0VPc1ll7EyyNP/weA6+m7L2CGLX2lgf8dO
jhOq9NfPeICKc7XNvxVrf0z2FVgaI3qipCHTH6JThq7uiKREmhI1KYidDfIxG1+5
jVYkjH76W1b4GEJsViRVEBbltzcNObAKidSmluQ5E/LUR35q+wJQabDyr1SF5aH5
XHTqe2tgfGoe31F3sJ+Y3P2N8u+1HgFqnm7pzdB3i3qQef0d4RKwIqtRyUuSJqZb
3J7U1fNzbPCIod7Yra/pX73Gne5SWZo0uSII9GZm4U0N1ByWzbTHZfyH1IsNLH8u
1VMLtLTZ56pdCLWhV+ZOVicssJvN9rOQ2ckdyjydFMLTcyQcaf4/AAyBS3HjThJL
gYB6v7G95W5jwsu4TzELVegA+UiXatQUUUTCiYgZCXUc1isJpFYAfmPoidEHS+jT
lmsidZDd4K/TNYK/gY0g1fnQhE288pE3fSzsgIZmHAZenT0lAWMLuOVwE5qj6Sej
B/ovuXgzAoa07dPHeYFpJDcY313SNBCtgAKKvdynQXkteh8o6CYfxa/QMZb2q1tM
aro4TVKs/4HUDstO2Vjxf6SoaadedWqDD5poVC+LRpb4ZGEar+LY9GLa2XzbnRzR
AiW9MYA4zuWRPnIGKjMO5VBAYL5t/7kIkWsvYc8HmFecYFl2VenKnwzXomYxRdxP
CVBcd68BiWXp/74DKDgAvOQaZEM9+Lj+3rk8SoALObqltmHSAklxrb78Afqmv7Ka
Cadnrq5i4mbaLRV4Xmw4uiMZ4XZHL0FClIw5IRdgKuuRdIGDygB7KYTae2mfAqHA
4mh0Nj50JVawpEg0ep5k21BGEmjRhNVHQXaC1tfMVNvI+i5q8fW9esgZG41Cih1P
ybcLy9Q61Ttw/SRL8uCzOUIyMqNgjVA4Jb7WzhHxx5nTeSSM3zHPs0H4l2h2az6k
h/uAUvERzuEBFG7qjPx1dwJ0GvBgFYHQrkoPLSL06HxHQhnkQlt8NLmPN7OyrtcH
yxWhBrhbAmeldQCgz63/EL0TTmuM+aTv9y+AxqI8tu5/Zw+wMMNrH31zcMRkyMOL
tY854Dcq4LyValNntX4wTyonDNTmWoVRBadmmXgOo1KwoVcxX25PR3oKCrRj8YC2
wFIsU9SN6VwXnPuyQBUs6MEW9taAYRssn/JOfSBpV1Yh+JrOfiEOihFSYdqx/kHI
zPn7+FqxWA3PAo4sI77oCOxeN+9RLj8wibBA6kIl+nP1y7prt+056ZHEYYadTZlr
koSNBbUZyPsYJEKLJ8YAby9RyBYDWI7h8zXg4YZ1Bgk79di5aa+BrWhFGQR8Q83v
4/P7Igq0IKtfFoyzhmaW1PNhckMBo7vJc8ZNftlCsUmzaWBb3Vvip+YhUspV6I5O
IvpaiMmvWOibOEH/u0gkK44Fx22K0SZk61ozRlczddARKNQu1/v3gXKCme+8N4CV
TdPydpEJEiUGms8XRfSvNmV9qpXbYowCXBD4eYLlWntB0IxMecpoPana479cvsAq
Ru7mDun8iSZUc/fxV8dzUtZMlMUUTnv5A7wvuzHpUsmNoV974VbYbpJjYZhOySQb
X7NRXndzDXat3R755SZoWcQCoVnWqQ+AQu9fuMi0xx9QvfJ7MtftixIw8ace13Zw
I6/8FXmiiEtrjDhGi6gSLIFVWNDohDvy3Qo0GuhnOF+xr5z9GmGgpWWGNBgxX/3t
vS07pPj31V9cafjvgPJIaiJD82u7/GI4tJh5xmpRLp0ii0WSmb0gbP5N88PiqXU1
2LBdZiT3bB5bAUW6hBzBMNKlIFZnqE+6HOmwnUmhOwy0f+QsRD9hg1JOBwuzgAwf
J/7DL6t6w00bsbLG3qY9ZdKq+a8nwWAEA9cFMBKQo/pequWvamEfZ6WT0B0kioDd
5XZLUsxsew1l22xYcebpWQCe8vlKbnrveNkfySeXbF1xmRVSVLRNDMKxRUrGQYtR
CxjBTRxZxJ8fvzKuB7I1M3LnNDfx6O4rYOqfmIVqT7wTm+3XMCOQ6PvHaUUnmh6G
IO8rk/I8Z2FqSXf2vlEL8smBG3AU12V0R9v5OagH6/PAKsN+8jIhqf4VSrtaqFOI
RDFdTqL3rSHc0TPDU2IQT2Ow9KkOufOGiSCIcPPc7c/tpIukzHds6McNw4kYlm7H
zz54hEJXv/9tEI/CGMl1tNgKaC2OY5e/ua2dExhbIs4RWmoPaR0VZlRa5384sLiQ
KDaoEblpeU9wVAk6yqtrIfk89p92pmLXNT5qVdo+5XEHMuqvtwbTjECXhHEqNC5/
jTySHP4A1fyZUNc8ncEce3yik/lVVbP7sgQsp8Y+qQ8ZNic6VCzVP6qlCzDnOOg0
cTuSwS4abWimN6R5upddNEu7IKNds9oK8+H5MZd0ADP5GtF4OaFmOI1FskwP2jd7
vCoMd5fsn7cAuleodxngdRb6C+MiJnKP4zMQQ57xT7a8nAT8zQshRGFzdM1XB91c
v5pS7z659CO1uuXyJip/ar1kIF7z+UI2TWheZ1CEjZW4tWcOF5HmxILZbvrLWeam
Jl5DdcJP2+fdW+322WiEQItr/dZ4e61bBgWrn40wzCcOZSsBHgBgRsuDj2p3LYQe
JK/J0ltPNCFXUd5+20qal3VpmGJyleCcloySJFZ/J+PDF85xpc83PWARrgz9THvk
pdynienVn6Pw7+L8AQP/Hm9YJ4rsJhXkFnOtdnOii/uERWo3/6arhD5YCacd3K+w
PYM/sMvNqgzuoLBT8UZfZEZnW6Khmi5/xN1gaPmGwuUa35eQFSDnTEV0j2kPYa/r
rJw2kwVbkwaOtX89XJFaA1rB7Wzga3OIERrAQHz+Br9T3qEq1Nh+JtaQezLq6Z9Y
uDN4HGe5fbJ1I3qkHR7RQ9YhBAN2ub5pGQwo8guxShfsCVCNxINCsyI3aUJh7o2w
BdfZt2SHRbhd4KpK28JT5kPevFJyuIwSjKLq4wOzxIe8zfTjT8v5E4D2fA4RK5pK
YY0/6ewaxo7rZjoGtJsGlFxkMk4vriWtP+C1fBMmB23Vb/nw/A/lbdbovj2H0yWe
DnuzbmyH70y8g+BE9X27V6jtJ7P3puJdvmxrCScSgOzYkj9a43Odz6x36hjKOHWk
WhCZ0ETnDW6ViVF2OBvX7HAY5ePcs2Hk2wM20AvaSNTYQQPml9Z8RfX5CuX9ukee
aW2JHBdcaud1VFUeqtsNI4Z6tTiGMAnVFTxgLOMBepO5Wqw4wEurHsyNcvoTVlfB
SPbN48ckO7FdDbndFv9hrX1SGUHKWEzABABBMVcxisG16QF5Buxr9Eyny1hEJzUZ
VxQtjGRHgd8NS/KyZBXcy3MR72CCP41J68XvPAeswigNNKfJtuk6EtF7zIxRYqOm
Hr72FIafXrDMGVxdiJ3sEPmwnJEUVmHvoUEB3bNUKtHM15a/ZjvBgvb2WxUqeNzd
YMwCTvkJyD4aQG1oAsESRcdykogY7i19MlIg+WETgEcNAPSTfC5U4Nm5jUdJVmBu
KfbE4klpbbU32fnDy1wrh7B4S4RDZeFgP1AiI/gbapv72xaJfrRG5hS4Vv7lBTFL
5a5ftx9kdqsDbnl+CBAUssSdLMK1gHjQU/BYJqWIbMVc9mURwmSjc9mIV1CykqEA
Ua84XznTlLT1ydZvTHWK/XCmevFM43pXyqfQzP1NHep2XCeUBCw+tg3VmD6YBh06
2ugqWSBGqKiK8/Mm5YRYyhGi956IIaltNqJ+3uqvFuyPbAcL/i/74NpJvCrBPpdG
G+IqdTE2PO70WAnKBUWtkV4C/cKU1F02ciIJhOBkcrmT4C0rbdjbq/x0vEqbe+EC
QG78Yo67wywoiHIYiMKPMtYLU5OLj4EAYTSEOurMSEWyqBOGvxENuFKaR/8KBqrp
gfSzqAfgByPbp0jXazgQWh4tulOWjuHjkM5E4iMm7a0CdBgjOK+j3Rdmsa5yniq7
cD4RHcSJiZ15z/Em5JrFOGVNJ539/1bpF+x9Wc6exKYR2UMkeW+6xTk1wmduy6Hy
UDdOrU2oKjrmoOqRzFtOkJAxCS40cVt4SH+ms7MuupQrrYIxjeWnj5ua9/CitUaN
ueFI3WeTp9P4kIezG4JI61GIXKZIun/uXBUjKGGtuOKsWh6vslsg8NCxX0dqxgrq
O598MNT1lIBjDPeCrQ/lweTSWOqDdaZpVnqbG0JCHPOuyzYc4R2Ce/4fzUrRPik9
4LqQzpY4aKxAaD9mGuXj/QGEo6UBVB71Jz6fEzFjFJMXA0Ua5+dfcAQyfSRhcGyu
GVutI7qTDZVoVE4Jmmj2WaqgSJgGkbOQ5WvFZtVs0dT6fmhDEzwZpsQQORA2LWcV
o+cGxHM/nJ+SzHvIbQjFE0/rkBF3S04tVQwcEZypcCVOuFJcC7dHKxVjo7yrg49a
22SzbKMyIpazxPeUkbXp+ETFcdaI0NSdUyCRbN3LHxo96YRPntC/Bf/QW9rq6mzS
t26sZPUzvjJaIPiS7iOm/IOH/m5j1EhT3Z2vVVPR+yYutfu3AkxD0Do4jgd/ltyu
dBEzf7UuXxSG3HZ1CrUqGqAGHPos9HFbF7UsqofjSxRDlbRcVznUXIzch2ivaGcc
eO0cpwRUdijRdg/Wp8HnG8mhDIDAWNekpPe5M93sYNkkwuaj8+wXdXJMkQhfZzzF
HGz49dsA05nlbGj3OWVfN+AN/pK32pQfzHtV06FuCSH5Bt2Kf89DZwhIo2AycCFO
VOslZp/aRuCbRliljaNXKEzReZpSoVirDfLARZPcjDY9/G/R5rIM/xdSPNg37PTm
w3kymZwqk0lVifvO5G0A63cvRRLDXmbbDbAQHhKSJJvwlBtQEgERrLqMJ8S6lywW
L58c13GIHjG+ZwzYkDo9R3lR3eoB8FF+ewYLYAFmoKiPsUTapyWkSMP2or+7lTFv
k5xkMOCinNd7zNTspfe1qmA7t/2bt3gbZlDlHdmS896pccwt8VCr5WuheqMjGcAh
Eh2LTY9hxsqmiPXmN/kTGFPWS4xq5gEGbuUesSFBcfOzHQfV7c5F1aZXRfffXYfZ
DxahNmoAx+oQcrRc/niRcUJMhYFVofsXAg7/CpMaJrQi8v2vhXgPWWrhsD/QXQQg
g8kqvwKcp0fdagtGCEdJEhcVixNM3UQ4TlMpc9VCcrxjkPWxUHdy9yV44nuvRNcA
h82DWJWid8JAPbXplwH6TIRf5R2E1h+ugyB9M97XHjzDn94+Ec/XS8eQAxkbajEk
3Yr24NtJYhjiand293zEToBQLltoSQ8rO9fuT5fRBZ38JLoSS5VvKH+CT5XmRmg0
CuZBiLl1mHhI1r7YYDEpuXQ2IJML9+ac+fQF6PD0b3JIFxzDhTWoECSI/cgl3U9f
OYyzOToUJ+hvU5jOKRVGFM/NBAN0QVGycUerNi13c/Ml+bhxOBCWN2Huxsb7AcM8
quL0J+EB5Hror/yct1G7IEnocdUoTH/IcQySMVt4a6KjV54XP6F/erViZExk4W2C
16TYWb5yfRjQ8JIm70/5doIajPYmrVtLyCA3IXaB1ftk4JLat3LLCTLjNNyYrRmO
HQbLjRYtk2SRyinftEeNKWYs/m7jqk6GcxE6k0U4gaw+wa5bCk5jnZU4dPh+qlc9
0YOJ1lCSS1aIksvOhVw/vj5uqSg8yBQpRQ64HXLQrL/DvSiK7Af6Yx7zn7atTpCo
QzSXyiaXSRI6DrtnQmcHHguEoYdggZIVNAizr/ey1hlmxkSqJiJCiA67yv9uFqY4
zdQ1QUxKEuX0WgRzx2jFisA2UNyG3tc7mQyTx2t1EchXoampFhqWTVo0T4zb/LMm
tZjnierwUtN0ydoj7bsL3Q6g2djkKNA5/iz3PHTJWiH36Z7DPJ9LXTOf+NbH+ER+
m3WwpVdQOIi5uEwMXc4yuac1Gea9Ol7F2tO7idHZW2TiJMp3QqpSbX0iCW/PL4TQ
dzxSbqR9S5qcaSNX07hyKT/OWr7mfhTd/aibwAiVF7SHMSxl35FgZUBgH2GI2fDO
dAMOO7MEzez/NceaRstcm9rnebBaCYena2odlHilwNN1oo5ycykZok6OLYeek0yp
j/nBBPnXjPad1WUyMtnF5xtePCECZ17VkRK/cmyAePMi1lpFgBgqFvRG7jAHPXEG
3FTeDRfQ34eXzKZQQxXiisKGGa634NFXYtE9sNqSviuB7FqwSeps79WCpc+4jzJm
azOD1FRAVmVeImU7q48GcY39oRQgjr4sPfV3vzs11Gn2eMBU1lsADQGqhm8OWVV9
6U2E3mt1knD1wDfzl/kA668RYGIhJWEDTS7H+Mizd8+JlvbJC1mgSZ39Vs4ECRoP
JKWJLsXQ2yqsPyqzkdYixvu5mPGB8XgnN1ACXbtXaerusn+6Kj1PV/S/YifxkSlT
y4lnPFhWNDmOsgpgUjX45IkS916WPtC102bWOfisCEWyq/0aOxW8RZBvDcX+USBM
+5fF4Xv4hrO/uRH8PG8gGzm3kW7ZnYr7oSGX3m0Xuvgu4ielhuz72H2najDTokfm
+6C6lIsoXocxUS9SpcIP4O1BNO7yZoHkvJXgMvh1g+assQhYBYMPCFZSuN5HnKyT
H3vYkZypOXrYDOCx8+yYpcmbhdWLHe1j3dbZbXiP190ET+83/v2sF7OVmcEbk+yX
7yoQhTsI4Zfo1UCps0HKui1OO+0vVaNLcOTjg/QCORA087gjjidPRl6WuEymmGEf
LZOlEtGchKvDguH4xP77ZEvUzLVkj5Ci+h3hxTxbXKcj0H9K/cOBh45iwBDHESH+
i0+nQWgm5t42JcNmWOaIHSiPyoSA29fWouc6mh618sR0YRa0Q2CYhrbvbqYyEdNc
oReKtWidf4wIte6xXM/wFX0JKIS/GKZMMNRQocalpK5AWAJZyw832aAzpx51/x0i
fBflUE+mPzgNiX/embonlBXVTOxAjwtYIwN+091s9WWvERwua2fbO9lzG5z/445P
tkBPKeuzNhrisPRAtn/G585/4xWldgWIs20iiU3nUnljSBOlbjpJj2rIXfdHoCUQ
HYryTUfLgHGI8X29idEKLz7hw0YP0nzGLBGUn9Ghe4Mtqtr9lRHrMmq0trV+9fiW
A/Q9bpp9HXtUapNJjQaaP4I2Wr9fZ10X0SP/2u6odG/Pilm26hsBG5boK75Sh1tj
TkWkGRFjVh4LumdAwAB3yTDCD65AxsI9Y3BQ4Q74CaY27y7jt/0+JgQfv52QVAxI
cqYBI3tF+lv27VRGWUGjMYy8/cqmUpIefUaPmsipxLh32BBHZdtIfzzPuf0cflEl
umsMlvkJ3OzoILArfTqex91vnNeBhHISDYffQdUbcZH1WGKTX+8ZZ84C+78Y4FCH
Lsh9JvhYkKd1JWFjsNt/s0bbfHuGd1cvaLVtNufJHUwh9kt9a/dad2S896ltfhxl
LyiKHICiT7pgRkFlMD5K7KPCo+9EADUtfBmI+MXQ6X7MCVYdDwY57G6N3HJJyBOh
goTpotZn9c6xB/lbMjH5rAzTvXraCKXrWaHQZZUebW4WxHoXLxcsaEtI8kXhhjVt
k9f4U0ys9gP6WUdNTWz+p2b6V77jCbTWgLXNEcw4kY3tVjo0LFFT5YL+HFFnTu5S
k5hIpK5AIVIimEFGy+W1xfP8Y3BVN+WKewjbd79uTsL7u/KBVJfjfTS2l4WHlA+P
ms2g4B9nene4ZNIhmCyaPR5KDVho5P6frLFM1HEiN8TWL4D1fF06WBwMHZkTFoBv
wDT+8A0R48VmBXgYYv6dUDauRNPrqCFpLheUXTk/sTpeWyaNuM2sHW2m5+KSglom
w6k4ZqCymOX38wjTq3fllajR8vXhRseK6pNCaYyHJsy9HcjbIiS4MN8mKgc5sIIE
HoCDo6Oiz2B69KgdVYXwLp5E9vNbLL/JucGF1bloyMrpyVmDzd9Ti/SnsGwm/HBE
G7qZiM8iBdVBo3XpJu1wnBOTn/w16DcjUTMcq3ceQ8nJBTkYxeBPvJ64YaWoPAIy
+fUPwAq8IY+1RWNrNVJPBlHGP6uQ1OE2x6rhpLUibnHTuZceFACWB4IE4AfMDUwX
3+qSbXrOpcomJI3xZn1PYbM0aE06uhi5CHovGfBcT/q9WtEM3cIQtzriZsVJii7Y
X9PNQ3aymKikLJ7pPzNwxsvcjq4iMK/s8eFJemlKrJYS/ACLjo/AmGUC9SS5os+1
1/gEESfN8cEXPrO5pnNtJ+25gaQ7ilqAiu7qLQRCJ7FqhN1Yen+6K6niHEXEE1dR
h8Y4tRvPgVP4vS+cXvRsvGFNGPjFM+NEqk5+JxFQa/Qx6On9Y9C5k3MvnIchgMPe
dmV3q5ZSbmR5k7/5fPRegUlkMFTg574YdLtWno+RBD89Eeu9iXOyB49xSGvf9PeH
uVZ5qOHdmaDPZzj4pVQHqArlvSdBwMn8D3llNfBzT8VdB1kNvnEcEK5fwcAYQJuv
cqwA47qX8xqffE22tC+jqN2PKDHw1ll5CVnx9T7Ep4MdHldsWLPo6epDl47jkPRG
QfwS4JBy1PMJ1zP6mjBMbwbxpPknPTkee3gSlBQqA1Ts7A613eTJHj9JHBXD2LkM
RWeeZ+ibAi1F2QUunhjfJzuxPbAjRQZu2p7VIXjTDf9jx337LxBsjQroyDUOmV6a
JRiP1ypYo4XhErc+/NKExC90SDffDhFMVNVGUxmNHhahM8XSOiNCCodoJoEmqanK
EF5W2KvM+/ZCV0N6Z2ATKNacor5eK4zmnp+8K4RIAIWeKDDpLNH/0kznXNn1+LnW
6q5VW2oDEoUEwC5pe3wPxqUPzln//is9nnhxFB1/ufE89QxR3TtJzZ0e4tQ7Q9Nz
DfYU7yPIoRsPkeWwJf0IRZWT/f0gghomYwLJVihfoc2b1x3beaOUYGYlRegJ40RJ
dqplNTJ1X2nzAI8fn32pgUsmeGZBpEtgHqNmex+ainCw8eJuFLszR1WGZtSFpssZ
3ZPvw6Ks1VY+XDfd+4zLVrXoW//TsqPTdcXmdj7UklDlzlZVOdYbs8QNJq8JbVUD
vQzVzWC1GYg3CUMQvCNmKJnQRUsKakI2jDbf+9LMr0I8AX7FmZUOWwTQf4QFajnG
035rrGazLj5Cci0wnyjjiT+ykU4uawTFrLMjmI8L1ieQHWwJMuZPFWG9kXgnVPBl
lhSYFVt0fP2WaScEwE3AnQfG0UXeATcJbvMKZ0m3MrvCJ2X425wBbVyFmLjXZR2M
fzeXlVdn2RnvvsmMWvPplp98beKf1EUaQQFes5K/AVytZXzZDXztHUp3m2an/t8V
eWIEkbMvMZkFA+2t98mmTvlWtE0XpNpGxeStsGxZjr+5SUFOn0kcIaH0mCrRS/pb
5PtIrt+wf1NARQriTio5pv+vPNWu/C7Cvcwn4iGRTL1PqBqEclUK5b13/TQ5sBqs
ylqWWfUwFAydeMi8vgTkSxf03FKiOXtoK/2J8UkAl4ArbFPxoATr17hP3wSIDQ4v
DB6Q0Fu92bVEPvR8oaRsJLr5ntdhISxi05kFeiTeGFvLlX4+x0GKL2BCMrYrdRc3
q/DHBLlcdp0wZXJFnPYMpoqih1phiRluQPOIuUknFpaXuTpj5C5WgEesAEoKjV9i
WKUJaldMLsBS3qFBB6sNqHoXC8zmXztozsd9UyV+rD6F5vV9McZfHnhH21LoIA4R
xR29AyMa2+q7SJOGmNyV6HM3lz49UO9HF1t5xTwA6glAN3SgRV02otO+NgZ/61ZI
e8O1NE0mVX218+wtoix3p3xWNlxr2HHny1lv6uHJgliDji+PYX+8H3PGOorCisT8
lYWDIRAAY0iCBiQDf1OIKV2QwmaaGIWoW3lElkQygu7SHnhs0KkCkBA2DyNuFeep
/Iiq3KG0xodaHCg2eHWcWOfzcVHSXoQcI+CfyNj8B1YzcF9mwUolCktD87RJGyHk
VNZ/YgIKSTplmC/0/LHiim4AfUHNldPTqgy/d3czOgPTi89CrtDo+42zBtjx2EGx
0wd0YoXvXvvrttCoxfgT+L9Iq9ubeUFbw5tlrFtjlb3qevHRW55gCH8koHGQUsp6
a5WSwnIUtwnH4L9duHPMVSRZGDGF97Z4wS/l3qstDsexlathMIAMhOw5N5mzWj9m
VBdyckh7dvZvFX5RB3cDp4lEnTD2sNmxKW6pv07WMUkrokNRnWuNcc9ooH6rrX9r
NGFXQtHWU/cS4gcNBpNwjjD14Tz9IxaapxAcimbfnJv43+BK1TSdnXYqMvGlw2fD
55UE6n3XzkpMIvmM7eE/wpmktnuqSrumpz6wzd9nYe5OArtO09pssk9yHaqq3Ouy
2Zs4LphqppASSdjR4sxw9v6MUNRRrXns/kZoboW7XA3sAYP0FL+oIAL1SwjYBiLv
P/KV3MZsOY5j0Mv5dfrbhRqgl+c/wyteQ0txOaRgM+pEbIOzOkyLyeHa5J+XBrKq
vwtyYFM9MyQCRKF2jsoExQcxJnnvDCG1NdaYCR5+oFoFrIfpOFzVaEtw8msWlYsG
yl8JiuhPVTP5EDDmK8yKrfK2Nikhxlzdory1/Bfy3r2tAwXM/DEH+Ho3PRXy1AWS
4eTRebTeW5r6UkoQNKYUO3hSPx8RqiKcoEeRvvn3hHnbl7TsPDpcEjxOzhWoQ4p8
trT5vcadAbq/j576OpyolfFG5eB5HuOxcFBSM+UfhuLGVoe8xkM3Cg/bgDyNCvO0
DxwH1Lrg9KaKw/oW3Wm/NsR1SmB4WGNn5uVSBD4B3bJ9+Zf8Lr9rze43+tSoRNFm
iLGs1jX9+jkWKSvImp4N5JeRwrimPAMX4Hc/Pi8p0iUHP01bWAfQCbz+W88v82tx
nLvxmY3n3/zPGBfB8FCw9V1AnM2thsIZCxE85pZbtdqIrPMiUgrtPg47mZeidFBP
vD6Zp8Em8w9CtL4GJNIKbVdG+I3l9OQXotycoxI8XlMsislPMWUm4EdknVf2SRzg
IFVsX/Z/ndx8dqrfEla+KuPtP9rzXf7iKe1UIDMKkbbngSWC3+1TopWWWwAmjhBr
217aQXrhCATDFRLg/i20PKKfQPbg+f22kVxcM4g278PxuhqoGKfTridZeTpFKFs8
9FpYg3rS9oZTqQhdoIrmDf1iQKR/XMmETGtOOAZXDZLJXr6hfBTSWutushyJG2Jk
l0RfUP9qe3KkxppDOK8Ykek8G+tcP9SpytrkXkELsVeUzNPogOYMAaQQGJme0f3Y
CBSw2WCNh7aUtDS4k3YnhyWDYPORmdmnIk/izE1Lzdwa+W+jSWaJg2Kq+9VOSh0q
Wjy/JinNiwNTJ5GSzJhHIyk1mPIciOtrBg1ajkfWd5V7+QkX/+nxgtAlTQcTSCjX
hzNuVmRgHBWNqYvxAjAk5GAC7hIYYTQ+Wa1KfkbclhgKVfbRroc3gIAe7xtCCo/6
O6tvA2zj9fPEFUfwtaZUfulx2MX0rwZT76N9nixvavwIJAnm6AeHUxiE2ZEDLkmJ
T3JixTNhpwe+xXqraJwL7QkIxyLBfBJRDUL4+U5sHEKYA3+SEGBm1HlbA3pcHCAv
D1RFuPIOpGulZP+eOYcLd4ekPJkUWctaFPPHYu6d5p52yfdq8ApgKtkoiAHNXJhF
/PQq9Kdfm6hO/JVUzpioxZt+qd8AwUmvLczg+t+LLN33CjGdkILioBM9/I2X87X3
ge9L4GkFAuEWGglMj30H8TdlXmzZjFlhVCD1F7PIoZdBrtMm3YbcbkvRbYrJVces
XltVv0IvIUvYphsGsb3CEW83/Zv2GihjyJMokdw0zvkW/VP0K+C1kgcsTLkOm0CP
BGA8E8vgFf3SXjQudUkQROHfl87xmij4qrGNZXpfI10LlZJQvXZj85b9M6991WT2
8UnPFBb+S1aTa/NIQ3MhMD4ZcUyjP/Lam/jQoe24nqgnEqYQ3riP9xJ98KgKy3xi
zYgFOtnldrUn7LTOeLmeUSrxihK/Ktvjjp3DJRyxttk7jyGszTpquxFWzdctlaGI
RAjXefOlqOP0Cl4eLBbQiZ6Qfi0bxjfXlirdoApzuleGDNgAa1vOCxRRkjfA4MpD
GJ29VpkhA9QvYYVh3x6zkqcK4KEvjkiEY/BGLK/wNJowNRPG8frUQZ7geGu5j4HB
Lj46gEMjX4jX7RgBOL/g3kvRqzwTtQTuuXkHBMDSjwQuq8MCROOijA7A9QT4Grg1
H7eMOvAZmX7RzywnL35h608B3DH+XmdElf7Xw5wyX2OHpYvoDlP+yBb/TyM1Jt0M
eSx80uPhTIAq8U7muifAWib99lVtQyaT4JAXfHe0gR1ab81Y/rMWcRkFD37/S0cI
AYgRJvNWbH9/MJC1MTkWELMrf9aBhmGXB89cbSB+z4r/NgrGhuAPFDSeKVXGPAfz
T+Lk3/FyYIxEsIv6jq9v1RGy0MhK6QooY2bzF8ORCSdN9ROSxGZZZcLfLI7F5n9F
3+v5Mw4ntqh1jMwwHYV6TN2mEU88EC8AlpIRTTUdyA77dZY6RkCk1x4+mVz0SCpa
GxWdtylR4oMwKq6xI4yni/hm98kYkzI9zkW9DJ955tHqptkuc6SC21DPqobtjPfE
9qMXZDWmP/Bln0f+WkooMCj0qX3RN8rId0YM6kdG2+p6e4nuDaJVWKU1yvMAIUje
bF1YB5Y4O7MooW+9CaaZsUCLsJ7AEjsCr2uweW6CeVHoFrwJfEb3CUDi94d7sItN
DLwjLN72LUhVk0KYLVQdD1IyHUQp6ppD4L5CR/p8qAJQ49MlmlZZI0DqPcMTts2D
IFF4sKejenhZ/fzn16HgP3Wl2IcSEXeK3VYxnge/ZQSue0fYXMlsPr2Fl3A8IVpY
qwedASSzxtEWVIaoISqMslsuS8B9SaNlm8blPuoZsRFmglKCCjNvq04zC0q+OQmK
8M/K9xs9YA1ue1LPwUVfckN88V41qHQl7twSGxcpeTkJW9koA7V182AfqsPqC8U2
46YrILzArIf3pZZhG3qvhIUZwO4I95t6tY/Pqk/OXDRSPw+YL4v65tO2ZnlwdBAx
dnpj8diMDiEQjLbg04JUA7bj2ZMEfZUtEZ8k1RVAcYUxc21ndLwPiXxpNVPiQfc5
yRYJpLhkVh5gvZoQvfWQIubijD22QLHt14PaR5REUpRRYPY8Ciw5MvBh2mug1549
3P/nsq8oE080WdbmmcqlmsaJL2/Q9yiappNvYv/MTMV4clQSEUfdx4lV6wuOYY5Z
auGs0fb9q73/vPMmgFrjD1FiNiCKF3o4qWjI8jw2QokGYZYfkbecnevsV17yRvOi
vM4VXlsw8X5B63WlWIcU4pM5oVP0J+z9oTlx7JTjexKjada6G9T9lwt6oaaW77Sz
1pNWeXk5jab6hfBuDzL/jf2u5fdx8MVCUq6dNyTMr22QphhSfYixEEj64y/c+PBQ
qo+4qrOe/I2pPNpObHYOAnWyOHcEXF+RgRtpTZ5F3we/lrOMY5aehHW8RpRCqNHm
lBmIegpe4ketwMl3H6ZXWhIlUBYkq2bLd9zDe8OYk11nYOXnu0KACosZ8Ma+jiRc
zjrjDz0aZUX4NK17540XqvJ944edsB5Ix+fnyZgjPIdvCUXQkc5oSyht0Uu0cmwB
3AorosxFjpUDyWC8d1ixgLLGCAEfzhKCS/eCzfH7SVwslViWzhBe1HLUaMkvsd65
a8ym0h/7ehfhOCBbGBE+DuyyYVWy/VEUq1k3mydjjSnKs5PZSUfVodcC1YamzaCg
tsaZIGWmc5vhb2gcp2dDJkhBjsZk5J5f58prlr0i1sx42K+D+Zu1Y5aaJUUSQ4aJ
uSdDybZ0QfFCIJ49uJqLPKL0ez9/oqPg99VZ8BXfeihYs01aLHIPdrbgxiIw/Sap
2Pxvzd2DBsEJRSJNO7wwa97W0oB3xaKFdW6WHBjwo5cpoqScAv7wPFmuMgig+ER7
QI9du8EbeztmCIKwrTBcnUZiADBI6odKUuoAPpdUT1b6oZs9/crIIS8aZ6NVfa5J
DJkVQaAQ7JqZTP04ClH4Wuc/HVSuHhfwQwyLD+6KQjdfZdDHR2o4cwctk4924Tdn
6Um7lG0Vk33Vtw9htadAxAZSfPwDYJ9+S3M62ZI9VcEpNR2OLOZlQRGVSnDWHwmi
O2dKCmL8P7chTxqNmrMGDF2JWRGLOHYYgck8k+DtwI77hCfe1hPCD5bJMYnM8CjT
9HV5oc7xPxrVBDSlT4kgdJOWmItVfNnyJ/HDB56LHaR08SftxJCCVb7OgbMYFEkq
7O5v8QOdVX6vjeT9tDEzcfh4I9yU6xVZjAq+2Mjp2TpWvXIAFbl6Bn0AqQVsp7oh
I26wrkiK80HampxoA8AQt9oMz9DsyIDptuwYC6OKgccl+oqPuPG+ZI+ZZsu2yx9S
KWFw7TJ0aaBbmCfz1iwuvT1l9zaVObDojHeS9TsyGcRG0feF6qQazvcb9V9QygX9
mi0lzJ1cW/HH/6jiw2oIBNtbcfUN+h6bzPhXjQu6vyQtQh8sGMrIZSe+gJQQh2qr
zLY+aAHBSWODR/67CFga0gIjET/ujuMixr2q2O1T22u8r5/xuoNOo1TFQAivVSvL
9HeBUdZPAIftdgSEhY84VTQ4IBNTExtOExP+fl+FTsXv2I8VeaYe9FWs6IwkA6NH
qZvZRnMwpPVvQequeU72GIm2X4BjTxqh9i5LWrHWRubanjPRjr3PlY/RwXbn8CP+
h32GRIi/MU8sTFqMPxSZGoEmkssHWl++4K6C8kQoKjWg+WjY0H1cJvsc8En/XRVe
sZbazp/plFYguKAG9oZj0vB3l092MMM9lCoB+gmvPrS1dDdg91ReEJySDSIWs/G6
03jJxeHxJpxCiLmcUYMaOwY67I7Vrk7DpG9mSPDo9FSNQBFqi6ZDL4kOxW/v0PaI
RuMFqUYMHq1AOgmcowkwBzOSTxB+1gMKcNAAkqAPDDf7FzFHEyhcA+N91smK1wdt
Z14gTqgRYXJIW/TogtDo/qCFih2I9S0YqMdTeMm8RHKWTJnHSSSD76eS9RgAhTca
2vqylC5av3w5nB4NvCvdG7h0h5Hf+hWMbeDm0Cm/xRtpjZ0+sLMSJxKfhwngGani
mamYgY8Pv2dyh8R02caGtMUefI2Tbiv8oJNnsZr7BLZlLSJAnihRFruF2QFMKYMv
nUTdSZ0SKo/3Nn+7jDQ1RhwCRyVAW2qTfy/AtFNSgaV1ybaNIn9WhxGV6e+oKU8n
PBX2rgPjNm6V0uIwA1d3lhLcGYIBTa86DdopI2WpZkdTmi6OYXUewQzlSHkarqvp
Iqq9sXpchQ5bWZWGn6NbF25fqPAqQzLMNsRBHL5MXZxdUvg0cP/TpplS5hEh4r6S
JGcbtOa3WslY8s5fc8418tswWlWmlsF3DJjSmo7XpedTLNng8LtPlZbDVT9llH+U
oppMWimahorvUelqV8U0Lr98f89y7JVNA/WV/1XvZ1cXwp2tRMwuMdOcn1t8+w35
loC0TOTV4fMZDy0txVlDJJnjHzIciiGtNlQqzs0OWyu5bCF6KrmlwGme6O7Jqlvw
UBwRKXjMucrxHroUl0T0xdLSDaShlGYnsLlXzqtvNC4W/aRBc7WiMSHBWeTWZ5z5
G3/978T64L1tHb+sQsxT5uNqiXITqi+kuB54jl1F0esXd8d7olvryLyBr0Drw7S7
HN7YGrbL1cU6b8esi21wv9W46LXWuYQgKvjsoZbkLu8H9vk+bFNuGIcymn9aGkga
mLdKM7Cn73NGHimt3VH7pKkHHh+Vk7hFiCv2xl7IbKVBY2HqAzOO7v4NnaxoI6/T
vAY6jVyDQMnCmzJY5D/uEjFKwcRvK/0Cc10YIh8vsw8Zk/oPpyeCPGinanvsQwCo
7FZ671IobNPfFHF+s8tZnlciVenvaR9oCrWl+z7oHHlxOS/U0HUYqUKTX+YC6dIE
NspTHReXiqUxFwFe93uxoP8SVqnFR4rCLjPUIZJTUw6D9GvcWnC+MYZeNIin2c+a
jCFpqQZFN6WsQRDQO6RnMiEG4S0I9WGu69c4JuVbR9IvTexkHcK5TOTRMf9TmrHl
+9ixKpLQoDefgdX/VfxNe2qhoLWH2qdlNB/k+xYh3N/Q7mMeXc2BsJQrfHdEv/bV
dpxnfwDuXGVEWf48++x0WXfvAGlEuYr3WDANs1XMP2zDdPNbxgZ3rf7Qwfn5NJ0R
2kf+m6w5QHtHB4KcDAV9ueggohdg3wt75G6QMKpMuMQ9PlnV3viGBLfKN06HDJMx
JpCCObhTNzwMr7YS0aGQQdz2UDy0d2rz8sEzjwbbEhs3AjZ2IUN+kxPNenh5vm2K
97HpByM9bC7fJL9dqgdkyvAVNiwU+9O+Ycc8atC35TPwWfHE9tYfeu4A/wO3f8Zl
cB6XOXHWcALowtrR5vvAAbcH4abh5Zy+t2ZD9xykdmGCdMg9tRV6AqTgfE1ZiHMC
Sx2CrHhgXb3p5eUPwFz+04IiZ7Ybt7h3VXQKnZA7M9pMglz76BmagPoDpu4go0bb
lHD0RSV9/+VMnMmhFdJWP748KkCUzppIhlAT0SKC77qQ3jMiiqITFPyg6fQkTvOI
MSLsMihvVwbdmKKWdr3EGQrsXf6z8N9POIzngVKQC1WLzF2ll0d+Lq23ErlA7AKu
/RFzG0RN1ZFFvEpR00bdO982U/XeedYAZf+uHZRkLnaKA1m4/j8mdArJ6jutUapy
uy3zF/D63K42HrTM0bqlzObiXW4W1eWXD6AsjlrVYhJajrB2X6YRZv8OWY4yngFg
9UN+i/514z/WL+8pw7HzhJGaQSDEVdKSHMQAWM0U47rHy+eboACzkUE1XEF6ds3x
xcuv4bX909rE5INKyTBxWhIiZSEZZ/tuQGHxUxFrpyRqrJgCYfm/+DX8O7jPk34S
yNF4W0TRDSQ/T5axlQLFoz5tWcRwwbejnAdb29Kyddwk7pNlDKn6Hn9BJqGhE2ft
JibCCoEE7F+wrMn3XfrbTC1u4BbH73abuBwRfbfP0VCE2YrjIMT7/3aca2PaqSZ3
lKv6YOjozHqzNVj/PYGU28FdLcRxyiyX8/uMUK/+vrIc/qmiD/XuIg0KKpdnkKJ3
RNKIhgjaC9ubwCYp62fjouZuy2LsQRjl9yK0fBywwVwMgenynqcsJlFakNs3EtQW
avAMD+HbFA3qIP5PTiKlEjOLbeFVEiy/sqyywsGP2Vbe1cUGQIh/0lrJrZyoYA3j
/mKjoRsBV6xwtRYPMEsqh+hszrjEXC5ACzzB8gpxvc7hzVzspQUPTfextGk235yC
WSS553iSqTYiasNA+GLevZiBt/WiayuTLVoYT8oL+NcwSEyXRBEP7qXlr2O55QpM
hDrJ2Zd6MPVHT3QiLV2+5FOaQhQdFpMQtZPy07Se3VkI6OzyXVIm+p7dttok9vk/
0InQabjAvPiMkiag6qgahK5OrKBN1wL2HCIuhSzJNExN51NSbfvshirwYs7dzUqt
y+K1pIwX9ecGyXn7iyuIGj5Kc+1uckE2cDCoVVcsqRHJdAv0I58TXYlOSaN7U2c6
AtlN7GRIYjnC33YKxTmlN1mtIUVq/H0R7UkBbIAn62fqskXfnKSdCFQbmH7y63PE
cejaQD5/b22qZ8Zo6g0ye250kkKwerrzysPbkM2h1/56jZPkxlG24xl0+Dl9042P
TsAKRP89ttF4pEIldPA0mOSR6p0zsdrI2dI9GzzMkAmLVTVPbJX/Zphy2ETKhAb9
EaDtmJZ5YUVAt9mYa5RA2O4fvpc4WESZguw440tvrNRaCLU/0taD80AM/x48XJJW
yJEPOc2PmqPXDi9HuW/vxDCKBJaWRIkGYonQ5e1bgMY8uKiqJM6QmGQASJqsyxya
RL/KwSQivfb/dUUcK9wSN/A5WLKjrtu3+tUeP4mI0a/LSKCz7ivzvk6SW4wRVLXH
xV5vAQmqI8OnyUz4HBlEHkQuuV8UUG5hR+0INp50RLx/J4GbZe1Ml7Ya/uDbh7s+
m+OYAXawO8Ia+1MqKiLRJWx+gx1jN0ti/rGpmFO5EWwowPMYJ42eu3iAt6EotbcF
5JsdqyURmvAfuVH6VboAPDMmx89wt8RuIlgKpKjHM7hHYgeToZP1oJpPpntsCJvK
vCP4FwqAhdB0X0lgqmwLezC2VN1oF33h/2xo7OKmgYepzHW14b1aZHoYjek14T3o
WbHvItV8KvrlUl6QBSuntvMZf0XsnDZjfVgPPUOOkFQ8wWmiHsOq2hrUD/sHjqxQ
j++qVyftKynTlNfGfHYjQ96ZsUz83AbXXIfnUdStcUNX4jAnb5lGTOjQMUvlKhqL
HI5ohfiYKK6QYC/LORBr6XxU0rUQf+cxqWUpwnvQ/6s+yQIA8Ko4uCF5wnyOw3FY
83YWXZzsU6TmsKdcE89fsTO8DPzgawBPFsXwYOfmMViCeeynWMGv+o+uHc2RNt1O
AE5P7rvsr0Irpq/M7XDW2VRiXyFBw1NIuNKIDw+xBJ6tSGNLpbH0KeBuuu8kjs7U
Om+mUY3wV3Lj4tZtMpJ+8k4e1YkRxddfUY+VpnAkubDVF/LxERRhhcD66ulKa+RW
FydJuCEy7ESFf+7hPdduWO6ol/WOGDnbcaQ5bYxRQz2SJOsvecoAr4ULnHcPT+vz
Uv2RuUv+d2+v3t66Wn0FxYuSA2A2I136NoflOzqkP2/bVx34Jd1vbSeptQjA1y0d
/gFO3LBFdZk74Zw9ARIiJQ7FDSv1gbsMdi7N/BzzhoCK9K0pJbFHeQ2GT8tdCFKP
jxb68edaKQKdduuNYCwlzFCF8+v7Z5mTVQ40EEC2Zv4dBSVoMTL4Uk5pvxNj3ajq
Q03X84nLtNC84dDbISeJIpfDwcBNug1DdIlZXEXjhhKTv5HVSmRBd0S4uBM919wj
Hop8ahwnTHMpFmhA0XWgSoFfKRkzsQoeUoOEAyV6/BJOiWoAz0sEwTDakxE5EIUN
ImBVScge8sSpj3i/wbPwIvdEYvaGndbypb/OgVzkmYbm34hKxoTlkG2U/d9GXMf2
oT1eOpJV1P4Sn8Aj7YKyZpKl+LCBDP/5jKTeM0yzVcgXHGhGnCBZYYlJJxBBamBP
FYzGlcW0ODNG5FHqXYYOKQUCDWXVoCBahd0eDGchd3SY9zN/xYe9taHktHWzzBTZ
4iDzQtdlZ6ezGsboGHt2EFIT6ni+pnWTNqOnjceh40Tfj7NmQcWjHEPDRn7Cglu2
ER6yjmK3zw+QgG/HNj88h8OXW2LtrM7W8Sa/y1GfEDQtASuDqMSjYpZXjRC31Df6
zH1Iu2jpWM+UuLb2ycxFjw6H/A3LXhPNMvyFdEWWqp66p4HUP0AydpAGay3Ynd7U
8VnPkq4+dcl8vZgnejky3dvqALcFPENpA4ocUha3/VYBcmOU8u/k9siFU6nCUZor
aRqrN/5KS0XkWqieupJKv19U12QQBafr2q8VqJZv8LuFpuaFc2xpb5Ek2KDAgpDI
FDIF1qwHiaTPYY2xSx/jK2KPZIJrECfuAZ962/2w0L6wFpeiVTtf1Nr6gVAaV7BI
qJESOdrvcBp8wNbYRsIyu0wCxHtZL9yXT6CZprvBVn4vwTDI7D7X1fTTWUzGu5kv
bheRBuNzqevrpMT9gx+S9zTO8nhIV+R4cMPVIxIw8ZmftVWJGoBDuOElI2nrsHhI
fC52MWO0u2ZRJGr8l9bE9K6G0zwjk19VstD7vFInpd8Lvko0QMWYRveNeF5TEAMZ
IOFhPP8fDwpObFC1S9DqQqiXo7uU5VICTdMLpLucZ2AyUGxSeYENymzh/KyHMsnu
e/5vXTSlAgIsioiFG9q/u2/V3lOvzn1Hy4ve7AzRCNXio6iXEbwZ6C0C5Hg+sCoy
JYYTEd0ZOZ/+o+NRga+Zzs6onEbotkEyCUwG2O97ahumT3LIUhEv+P/EaBDh9/25
VN8Vw6N3anRQmNNSMd7RTJlbkpEIZ7BF+N8DU1PsBrzhsqOjoRoJZ8oly4pJPTGk
fvhoI97dRN4zqtzNoDtQ9MLsiOfalvcyMisH18bjtZdrFsGRcKBkMitBOAycH5BX
FH5KgeytDxvUOvh3W9QwNr4z+Zj7EB+2vfBAWNKHHxxEICvNEt4I+w/weDi36jNG
/iFUGHL166ULXr2EVAJz0za1SbsebRRTXf7n7SjBsVuQdLx2x+0qgCsTbuXqtvrf
UnvLaVvIbOi58OtaCKbtdvKnF8X+yyg9AArYNVWgnnB8ze5rkEk+EOlgz8PKXrJb
4K9boJo+AkVbQj8OSlKYG9euQTqlKV0OTZ1RMu+61NLvKy+IqNmwGFtxZoyYtTVf
pondkz5bcBKuRYpTKJNMZhUZstWrXO2kvccizZDthAB5+xBi2K7vu+U/ttb7233V
SriJbb0v8RETSoGLrkdAwUym0x5YW1sm1KSmpQ8Mi5ndrHc1RCGtTuMJqudgsr2P
O97yi2CbqB1ZLWcRMMQBnxYabqxNa2qTL8IViGwnbYJElq6vnK75tiBFP9yKs/yJ
KhahAaNTcB99jzw5BOmuFlZnLJUGjEcEnBL099duPC0D9c9TLGGKli3JHEgkJ0Pg
VQSoNBVyb709HMVV8hY32FYxn6DlWdcACZJJa806AW9dHnjp2og0rOSiiMpE7dvw
687v8LZ6P3slo1k3zqrpEaPhvAUa8Gf8S+FnzlM8fe8NNz80J2i52Gtvz2v9dVpb
W1M1IretGW9psqquDR1TC6kmANeumxYGNQ7XOgCtc0m/N1kcfUiql6NbBcCxXGnl
dbwA1jj85ep/2WMmmJkAmyWXHRuC5wFc99+xfbMdBWqiWPB5vY3BSCGqkcRIklu+
MUPuG8DA6dl3snnL/isg9pdat5AQHuFgTFH9aq2vuf8ObHTOAEBjAcQmB2KuhigH
bmfpmsVSV+mh5JEt19Pes80P8QWr42l+4msR3A2YYj54XVjthUKsLDL9TbkmEgJO
CBmooERscelgYw/M9W9ORIcwzEq5zZDiyrdLP3LkvDyn5vWGAy7TGAPZ0FIgesFF
FiAD1pLJyA1AgSfwDEHoyUBgcnZ2q6TEcHbla6wd5vJAFkjt0RjlRFaUzZRcmAB2
L236AIH25Vkaxtm7JDReuU/5LLPQAELbiGTxA23z4lEX5FwZbTmmvC0daiLUEfo9
u4kI7EMAspaUEEaLav9YHof6Yab6dpObuT6PaMe5r5VdB98/ZPpzdBbNNTMJKal0
W88xKaEl+pRLZXslP7MIR6R4DNiCpM0mz//KxegTowYwnW9ErlXDtYMTT0kPnUnM
YzlytDIEU47D9mBFKl2I53mlaaox5jLGFj0JJkxXV2voZNzxNQq9nlaeRABy0/wb
+ocq0KYNCz8W4stJTapvehvnFriRFdXDF6OBYv8asJ3tzGtxVxq/Ikvhl44ji+Vd
rqSmScTIXzEKbAiuXAOtRPxgZ3W+mvNvhOhaX6gnoNhs6zg7FqvDhcOpdQtXdA1o
rHL/H/D5eMXfLJS14tcC6evBC+k/qwZwn1FokwrUAK/d457d19pK2T7VGKi74dbu
EZUEcRJQUyH5ofOsLZbO8SiG+GEBFev7y5txV/AablDUnO9PXltlZOsi9HriC1Rn
3Z0crhjqFeC8hg5h9LeW76RGwgK5hgSbqEDEO44KBKaUzp3AZqU5sRPByGvT3BFJ
p+NEZ+m+2kXJ1eGZc/LkTysEeVodsRp0zPalyDkwRttSnFxihb+SGU9ETg+2bo33
bpkUcKoyW/jumSPa6SxyZCYG2PLvrHSxULEjTrDWGjalctcSa1Z0IyPyXb0QIPOO
/DuiYDzstcn5nepO3RmNqaiSKLtHZ7+AKcQNIeALDNSAtrkc83HNTXS7lZJj5f1h
3Giaey3pZRew2y4gxTTDe+J3djh4a93teNXMwKAY+ZXafxNQzoIl58eQ81KGGGXr
yY3n8qQlOp4VD7QQjYBpXvJSLahnmD/K+FG4tfs+bHDsAkz3J/XD9vIG/vpuLeSQ
izCLnMVpDC/UPqRIcbexAWuVkENnSlZEoHEVDHxhbqw/+iJSD2U1YIzYYKLDljan
etbzp+CQi4JT7cewAK3jVtAGcPvhfXdUP/X8C3Q7bxIiDjFYb+A67NRQbPYxHWSw
t1f/Ut4AAlyD9ZVfb4j1bFnDrfLJQkFcbvIXS0j6ElPezz1qoVhZ5og4PYD1yOmC
JmkjLBVOsMtvGsr9J+VX+uhFlbXYF8dFFrkUGLCuCajkcJ5r17tuF9KCWeil0JZp
KuF1f8c6EtWR4/KDy9jT2eRNH6eDk4iuWqM7mf7f9cSz3KXVNQHNIQldsMqlt/ys
HHMEyADyC3AIlSLvVB5LA5dv72W5aUPuVU2HLiKFEyiPbetBjqmlCiAwErMKjmzV
e6Z+7lUsuBiQh3++C6w64/LmkpfdB67kWqm9KPQupkyL5/z/J27D5lEUCiqSadBV
ZC6MFEewcNRWxQKQS1USvIe9VtPAlxjLr+YPoFkbq3tMhUUSaZRqDmvbBwoUW6Sj
0rAwChHvM9PLqFCNLO/yjt6XQ6eI4HxPQJZ40PspC4ViNMbOtYHOazvkYiUEIbtw
LDJ/WstRQgdgMV6yGnvMkOuu/I8L8uc1bSsw37lXbNLhE2A0JZSUiSquX+C9+PFf
VauyscNX3rXjeQbgbUtRRk6WhBz+GFN/Tyl/M6PrxBlO2KlFLRVH2tsJ0Co07REX
bZZ4yE82PbRD4MmK34O8slT4kXudO3KcvNWIoYD+PUQPkWeGQZnfBFWo97vzcQPd
3awkpFzJjbqRx3dwMcnBEHOejWxmFrebaGb/YmX567pOCmdQoV0zcFyxp9KyXH8s
JIeddr+pL0sROReF9rPMYit1//S+sAFZCQgkH9XJLJ38XzPZAI0ISS6Kd1DqtSN1
1hJZahMbCwxdpoZcA0GF+lRxFWbSVi6I6VDc9qIX2sXTNPnSWV3Vt8I01HIJZd03
RjCXIjWngipT8x30d09KrdC9LvjbixksfRi+5r3Z7yUP6MHka+bbwo8nmSqa2jZ0
dKmXBS92fF6hefh5IaIzHiQOxdIrEmfDU2saC+JfDcmKbHIf5AfI0cM+6QVwMhwz
2h3H0xDCGS7xHs/6mtUuxVKiXa+jt4/uyxopdJhYrucVjqwUHZ+f7PMbJWpOZSQx
AMd9eCjl4RJxQN9VR94ZEJDA5wfrH2ucp8pVuoSTNV66pvCGz7QjDRkrd+q3m7Uf
X/2p1W6XjW/2e9PFNh7DWJmLVGUGMvV/qr6Us77PucJgAC6r3DahvQ/1ef4d5xgC
8GzVnFJETp//2CtODVKgaFB+JI68CAprz2ICGfHPgCALHI0psAVRK4yhRaS8zVUO
YHLHZDkq0Guf6fJJY27lGfbvS2YeiBnLaovE8zk3Nk4yliBCZv2I8a+SwET06Ek5
Qx1h2LP59f3kUojtYZsMbzmcPVXRtNqYbtNplPyGRTlkuBBb+Gsm5xuhpnkAp/jU
aGQCVZfSpbz/Eh39fcyUwx2LMwapUm89j4yK0VQSxXaTJwM1bv45alegLk0/GpNR
UUIfJeWgyfoDcGDyFg/2n7cFaGABJnS61if3xTx5tcXbUHwb+zVfxmP3YIKjw7Z6
lrvOW5A06chKIMM6I0nDFb7tpgiBB7IgKW1vokneDnmTzrygcUe4kI8RjXkSRgz/
SUcjajKLECILoH8aVamxMtYYTGxeTjAML8ByO7peiFpAj3TMGpZZYd3cv852IvUU
K6NFb+cXvYWw+iRXXUxbPb05XWViHGZ4L7HGhqXVvS0A3j/bders3sP0bAyHRGCg
vseYDzLXUp7A71eit5pssohqgGQfEBOeddRkuVkZY+Gdi9pkgSDO3YUo6zJvl0g0
JwEIjoll9Pg43YU2H26EhS+0MuiE5AKLMwbUh8Iqefyx6+Qa79fhliqi6+X/SO1t
Q7q8dU3yyljE8iu8Ur58cn2AA1Myag69Z9YK6ZnxgBrZRU2W0dFz/bvmOIrc6l82
p/V7a37rWZWqhLXRHWpuhiKLFhlzK8CrMKAj/iJxwzvwYG1X1ZpEhMhTEkwqZkhm
WdptNKWmagKnVcxGSDYj3iwwti8A4SvA2Rr1Av56yaVl1H1CP2RTFHEyUpfOOM5d
eodAkvxvhDOTAauvDCDLtDTmb+3HT3QlVPx17MQm88iGDd+bWV3HhOFpIekidL/j
TsgyMBKGiCgOgVztdljj66zCZC78WILa6Lvkg8P4sa13INQznIr+etPai+YrPU4N
enexe+zwJwUNqxWz2Ehs+x2azNyfRD40jpER+HgAIL2EYT2w7qiQAf5mTaqTVLWW
FVy+Q/a1RzjMX2RNWP/WX2sbEcSCvTYupSW6Yq8KxCP9fgk4jOQCEbrjA0rJvHWW
XIVGCn654zsEupIL7IFXbptxJiik3C0y4UuJos9gl8y9a4L1OU3BagHito0lHxdl
u/J3Sif2WtKnwZ/6EN6ut5PWmGqzYWlc08kI15W2HFo3ZrdwVBsdm5ay7+altmPa
OyX50Lwcd7v5SrEiTEmojUKeAeK+Nyp/cLA4sPbmOt+BRX798oLfJDYVYjVbrVlu
bi2OthCq3HsD8a+85f5j8si3UocBhOLb5Ij/nlvoc1L6Oe5LUicbwTpEYgGSqkdk
+izjKIx0nu+FUOqLKUoemjdNtFewMQzrjAGVWwvhPDs6auQOgp2+cdQwVKkJsP+1
w4UbaPmjySjYjMCD83A8pl0fN754FKdmrTau8usfMcNiLb7uLzBpxe/nBWn6YLJ8
HBfbzoeD+bhWVXmE7Grbv9RKFuQYRJG8WBEc0ZSh60byXt0v3Vn3/9bgrzGu2wQF
gGPqVjFMx6y/KEkGlVo0GqyJR6BR9QSu3PGNoQXH/7NbRbWab58jyr9bktBL1SSy
NnIt1V2GhkUFPF9VJKL2UAEjxUDswXzict4pSO/WHaXT92/EEGbVGjw0vyFA/12B
f1u9Gwzee3C2eAQhztIhc/QmUgRyYdWq3DHN7UcA4m4mch2hDvFva9KDk9zLhXh1
7MdZ9i/6H3aovTopyjjiJ4W7O8koqo5vNWjE8u9F6kxkeEkf89WjYnNTpfP0kGgU
FDMzlBHLhIQ2qPrNU6M+rjy25yUXu9YMBTW5mDmHT8hOyC0AMJvmH3dzQqTna0Ry
7FMgdA7NnXG5DAFfHgPkfSO6VsWq+hjgxxZrluIPqh0kje468Rpfcp2Va+u6TQxE
txIJJ6iqqp5fiNrcNGGqdPbm3Luyi4NCNBpV7Cx+9OQ+2j6qVESqigOzP5Gg7V/d
yo11SrAapPSyE1xFit6Z7LUxFmN99OJpwAgalxsrlml8PLbeW27go9FAIR5sNztr
C18nT1F+HgYYZmbGMb5dfe5PHrgbncaNrVXm6WrLkD6ePy3v/8ZlVIrvm0mi0E0S
j4d204ttL1shUUc+NP9k/6y/KgJZeT2sxmkQPOvKLJADfXvco+n22nUO8e1np/hg
WRk/tyhkGo7vGNMAsZJeVsV0sakDIVjA0UFFwWK5fwVWGTPMpqyYk6kaw5TX4jpO
Fg/7eSeoNnxq8dfNswWpTR/ilE8WHxpo/hkdy1Sbll71ql7wBritIk2BUq93bgct
vNZtGocaqcwF/wkQZqYWkTUyhpPcw4MULx/4w8ngEQ8eocgEyk6Bzo6Sc4y3/gtt
6a2ucYUF9YqLtEOWQXGsMt6EmLfvF35+yaSru0EafEz8EskQMxxcXSdz6IdsUK+s
JAVqauQ0dbv8UGqTi/gMjbscyQlky4ujYR/yRaFlbmKS26LP6TDXBY0G1uWdhRKz
m7NZH20Rw2GJjvDzsThW8xTUgN7Fdc902hmT/ywJ1Jwc/DCu33mSNb30V/paW3ZP
1xyNs2qfOAV5sbCUn1v8sV3XZsTED+qdrYehpHVlxmE5fmIlwKyn6OVZGv451+Pl
KVY5v99TL+MOHW9tAvKBVkUDv42ddAjyMfHVXPT7u4CnEvYXT8R7Kx+pmln0OdVI
kGL8RGsYyJAO7czxJejGwsmILFUDQ8qljFiHAvD8TKs6pUzOF58OCUXNWcerHEnO
X1Eb4TJCcvTpeKBbxbtB3MJWPYUWkvtRi4obZpVAGHoRcAGSqatokyKYOJ6oeOSJ
bTm0/HDgx2o9YXmO9ruA5fbKoKZ+OglfjnPD4P4NkkZtOgP+nHozleWqkQ6xZtd0
QOsnr9NpWkwwaqCk/NGHGBZKWrAdOTL6bWUR0aUEMB/3JL0w8V7aES5FQv4Kaxv3
7GKMLmoENmAYl9LOlReey+A9lhGE0AzmLNOj09PQqdBwzor4U5TAf2WfT41oH6qX
35jkT32XNWn/FwVyMfaYMdPUZk2A43RYNWz09thP4KI80pAPFo6q7EdlF9SxXd26
Yy32Ho7sU7YTvSMIAl15xi7m4UWZyz/3Y1kqdLjLsT4vCn6ZLofKx/tkQLa9Wjc2
SMaSQiw5mig9PJ0zMWEFOREIMupO+VroxPevj+XvYBqWFta8fumGwkI6MlKmo2iu
vju+M2gLvpDL9LwbNHkc+PaeQp5MyelR97wqKtvW74nv7GXNBo2dGkpIOu/ZtPmr
gM4YE6ia/URhZenPmbBFqP0RSJp3deGVIThA0yqBwDuOfzBD648a07X5gQLyGHvc
AKWJVauJOzeeP8DpK6sqRnRIdyo5ciwlLLuGdk6C5A1SQkyw4mzcAZnyrFWVUwND
XnqHbUzqt4OHYjTEtdArSvY0wbb1PIaFB9mv0Sg3ub6+JfZMACszFHHlIEKD3LVz
+BdpnO3aHoD5yEc8q17yxBVn0RIupt2V8OAfZpqKY3VYkBwlyeN7CxGg19JMrHnc
Oj5ngSqv/3AHVRv3CFgU5a6e7rKz50RUmGJL9uXyuMEYH2k5ANJEQObuxojxKzbg
UxWu8bDH1I/aeA5Eo4qflBi3BcRMRuE8Sv/5A7Nk1XP91EAVSTV+xy40NnFbHGG/
ENsLrJMZmjLhv0XRQyBDHVRNI9in+FoK4eDbur6/png1qcx/xi3aqzQTykJBdKf1
fd+EOlj5mYU1aLGfh0St9Nen6ZTtB5mhNMJht4M5tKtxrWliJGWdzclR7qaVIPG2
UxN6q9pMuUBIt5ai6TTG/IevhNAY5AjGIy9GuOnh73oHB8nQmuxXUyXKvKfO9MLe
lfaiYxrzWYcGOQNHrPCA+XFlN0HK4oFrpoVNybz2/kAMRuWCiCdyLfe2Jb/h2ugz
eRzowTX4cCOebpfGhiLRxTljDBcIvV+F5BjGNFh+5lX4jN21hh9Ek3rfSq0Kluwx
SNW6xueA3EXqKUlO8OVBC685Y5VhVyQzkbTKAhyAAtooojbSucE+QNKgZgV1ngX2
aDMQGwns723zQe1m/j7gVLSRWyf7zV8LR90X6O5mG3fdC8mVawJXjRPL6iikQGU8
iqH/H1b+0dw2PN2B5MQkYTlYIRGMqm+yce4BcczFrgHtoK6QVcs41u1D7jVWErcE
c0pgVVODkWxBDHLlxj0o1kVVo/GiHaP4YBhnJ5hoZKP2enawut63L1XDKKxnALqI
fLT/Ex/iRG4Jyv+u6/0GuHLS1pmmurdOsSgtmPmKiYJmMmTQwR92b29JflXH6pob
3Q4TBNBAB+N/C98V6aQEHaCoRMBrmG1kxjleuWBOM0rApDz2/MDH+Wogo8jCePux
jdXqidkwkLD9pkh37ha4qsl7q+p9/sPXj5Pj+ENxf9pS70PDnxi7CQAReQ6wx3TQ
Ph0EhnnifI8SHDTQGaaU1Z86MThVTlhzC5OtPwqOKP3eexzNgrGUTYeLMXVwTKFf
mwY+JjlSq+TvMR+S8ej8AGxvC2GWX9r/DInkS1FW82HYHzdipG8bDBGGFYqQNzdG
ScqMocP6qnbQ1ccLe0P1LglG40lxche5BjjQ64bsfji2jCS1oXyA4W4YKsjvZMKZ
smnRtTXuj/EsOChRZ2Y8MIfiuaZzRji5W+7kBTfhBlN1iTEChWatYbsyUe71sD18
bbpr4ZD5ESZNWXmu8aoQLwFzFX83Lm1GqiWxHHmNhsG95KV0RFjEg1lCgqHxNMEo
lrY/pZ8Od4Ak9v266UEWwbCJP52PeDxl2qRNIo1WVhp378F7fC6AzLHULD1Qt3MA
O0i4Rr8J/eE79X7T65zkrtqv0MAMdf7lxmiaRtU9cki5s5seIolGCPAXBUSDZ3Uv
muM86QVbfaa4jjC7oKdVzcoMAQ7X5ua5VhdpKfwyJoNNmqfH5WjeQ1N2xq5fG4dC
DTBDQxBIWP9bLzdIKjGkYzJ4VbAOMdQnlpCmS4dRw1zQkjPMl9LZZEhQbMCGUHbm
yLp1BWvyuXH5ICNQarb8xcBeTICNSqpUoCM8KJ/x0jRcdPkzerGKb89H6Coehl5t
+qjChqVEbeCqSqYVFK4kB7O2b1P//EdTcd+//t8bNtRdmtmKyXRZEmA9eCc9YWg4
N2F/SzwA4ld726e1wBsX85t7KbL9d9yjG739fHaPZYhk/dx516vaM5n7JQiYJ9Wq
yr1390+/KikDO1uWMpJJzJsZYfWXVu1P4f6O6o+vVSjBqqkXBy2RSjPzaIQANWdZ
id/R2HU6nDtNgcQK3Iw7/lZCLhNwmHLZvsFyXv6CkiDsooyAZoSyqZdADDLR2YU/
E5TTpFzMDAp9RCnl4PgVDcG/lQUxIHHlk5ITAp8321s8FfQuxaag8ag0HDn00gXg
8jUb6bhD4VK7DMz2n+h6oMOZDpxvI5U+r6YIv4cm6eoxUPFLXcwY4oR+joaCYjZl
70OQ6eP7+4XGm/jLNxt83e1awQ4nV5wpQ7BNbJIMLGo2UhOgFMuazYBvjJrJnkVV
IkAwYw4zIg7dXREM1hWPAefF37ZCZR5x8LWS365dgMzltvOeU2kVj7vyf4n9siiX
vCGWGOQXpTrdMCy0XLxMacTcMwjxxXJ66aDbbiWXDTr1/dsqv63y/FllGlm665mu
9LonC3CYsPoSUg57Qvc23vNp8e807rOU27XgYgI6P1aFI3fjze8gPYyMGF4LYxB7
owzDeEQjL4kfQRKRbJfr7B4Gkb6qxUueD1FCZkTXIejbKnt62L6OyZJlK4fFkH6n
O2bGUeCwEi0PvSxCoy0TRq5Z+vhBdTu5knRzH/PLZrivA8HSfuGmtXPGnFaegylw
+bBCaZi9zTU/KQw5kjjm4fOfdtdyzF5sY726atpztYkSjq/Pf95CzwAPvZPmcCxs
5NDftxb6uSnMQixc2F2yK/3vVJMc9mPYArl++KzpPwSpaH3PAKAseH3gKz427kCC
YdLCNkEW8bVVTfGtTXoG0zJ5Wd1xYI5h6D80/blxLrMfXANJ/kgQHhPgvneFh6/C
00sG+S/Z+d8Ksu4C8kynZmqqLP9RMPah/XRmwauoC+pKSH6oaK+9t1Lpg9U/NPZy
yeozJAkO6ugdP6OYavw8SIR6oSkZNr32GgXyPQc0yEx27rKB69Bh2Z0NhwP4143B
RLLdyfBRYp5UYHSOt0nGFdFl0zzIa3M1PNCfgxzMhWb0T9v3RvXuV2Uk6kBw4ROd
LxPG4yh1rZxj0fogNeKn/T7cuAHT72c1VVrlkab/3ho8TG21h8nsDgWsJf1gUlqN
yatt3oZ3hpFNlT9uS6TZo3hjj8S5UtemYy4pQuFORCJfVGud2i+OQLXdAzjJE61P
QQvAT1e2ajScd/nbIqt0Q6w3mevf9i97hdqmbW42dHfBI68rhlgb98Lmkj/gHtvG
KuR1zkwzZH+nHfGLvTHGkh0aYJ/kcz1bCyxl0cX1nLWya+tFxKQWL7nh5dEoxejG
WyGoZfdsIYahrzM2JQFBmGzzjEFI2VT1XUXDDzWjhZX3fEbM+xk9Vz5fZasQP2Sc
PQIUdehFV8mEkYtc4eTSDy9M2wxXYig5bc6eEP+6Et9O+gg5NDyFPMzpknR8NCfI
MF+s+7mPEO+Fli8wZ0OeGRyqDwweSToMol5o+S7sy7/vzjZWRftIACI3Yg46Vbpn
2uoEz7d66LLS2GDdjRWt6iH1vvNs9t6xvLDuZI61YvIVBiIw/Nl2ZZ3RNN/cxhYJ
96qczEQ90ukVI/3StiyyY1ypPyccIm/9tvO+9lDbeZ67C5P/csRzWJvQM5cBGy4I
8i3BKW96C9YW7sY49RY6wS9l8JTJfmiBv/0JXGjjd+3daPoiLHZns/0ADDrd85nU
4i4QVpPxZQ8fgl6QQfNVcDOKz28b87Ml8hGioaWEWAFbDtum8Nif2/ZM9E3fHyp4
BraMURkBkqbLm2lz6jilGwi1wiQJMY8AG1MeRNEGsx/ThGRWlzWN5Ho0uSCmx069
3lFCIh+ghE+6W/iw6LKICLS7zQ92aL/5i2mz2oCprXks+9+pkGg3PDJqbb3ToBgE
XAXlReMIj5WwqPmDUpvOw8R8fQNHQJOy1A7hqgKQh0diBAnFLjrsXDo6DYvfPVOL
7kSfdZkcdhuUCP8uBdvmwpMdpBXdp+8lL3hu9EbwFIr4x1vmz+sfkUNQB2nGydoL
ByM0u4MZPDBwiXrW0WJ3jN9jViTj8Y+28xjRupgI2j3x84tf+ttLWsVvgKJZjp0l
eZloTaytBq4/6wcVDGj70pyQpmg4+uTc+KJdbLJmPW2j5KmmorN9XpKfoRn4tt7/
mMmBCyxQ3Tr2ItIidyjALmAmyM7yESUA06xr4bMr2V6kbThjDUiYgxE8GFBSDNSC
9+x4P7FhMNvxOkpJBpddRl+ZlhPjkkz1oLEa8k7GJcyIiHicvzZkBO65GKFIGTB4
162K9N1bEsPHdQ8GOQV6ABu012xdTBblza4kbAsaqkYAGtZG7ZVGASCUbO8M2KbC
I9eND7RStQtj1hL0qanJznLHx9t54THvoEs5/XL0ygmQNsvtQO/gVmGU1T9kdtF1
I75LaHe+YUlJ7WwMRjG4g+bKUPGsML3HgRMja7jTGieHpY+Rafzjpe1bQx+vz1jE
8TIX7AMFIGtLlpVX0EhnBk1LWS0ag8i+JekFohv/Dr+5EvOG9+a1Km9UCfTY0eGx
BDMnE5iTIQwofzLhHGJN7zXOrg3tN9kgJyw3s3M5WPgDrR5F0kxslZ1K5NwvFAg4
cBDVjyoqCVZlVUR9pnKJhdY3Kek866l5WTQp8gqniqPZgs7Rhhja/74eO7hWDgoF
hcZAjVw0AsR08pBRLwhCLq/MM/nDvjAKuC0nbLgYfTP2f8HLb7luALEoLr07hsYi
1j4f8Sh1s3NPN5L+40WoWcorhEu4WaN3eghUiamKnPCCT6EynkgzPR4OCYsK/z0X
v0GjKMn+eLMe477JngklqBBtQ44HV7BhXUnK/DtIpyo/zY73q4JmDIMVP5me5Hbc
saAM9flT52PypjOlxsr0/gyJgVOXv0h1KfvxiJpyBV9vyk+rNlUg58Ug4r53Ua07
VefxmQlHKA/gXZFbLSLam+2rabdUtavJ5sM0KTypi0ezVI+K6uTzfJMdZh6k6MFn
bqPghhrIIHjXSGeMBCYRp03xqcjaDHv8/A5V42bqUviUF/vbGoKh7IkS/oi+/a0S
/2phVIGEe8ILQU8TBwrJHTX/HBuROs9gjkwR/rza3zA53V9fAeh4BhuY4H/lJGhD
BBT7cgoZb0qio4SlEhG3x2FMu0hU4XmOiNLE6GfGeP0ewiQf0Z57TyjN0LgDccQh
DK7xXGkM/A4TpeXl1nfBH3Ah8JlalPuPQ7SUsfvXYlhx9mOe/ZAQBxXuBi4Sndn/
Mm5YZ0nrpJ1L9GfUaVHoBxivDnams/CpVPfc8u1Et2DZlE4BExr5K2c6BMPmeXnu
2NtoU27zIHkgNzeBV2QVk+sUQyMqdNipbnbL7HPl9dwVpg70i04pKSB2NroCb/Gg
uBrS06ec0Jgx+S25yt8GQZEp2qArlF26eXmF1Gv6Ms1tcva9+VDcQodLvmQtbzBC
4ZKuFp7wApcED40HavXS1hytzdekjaBRzIz7VjX2yDOnHW3xuFz9Z6QajX2h4BKN
a3GHf4kfKyYBqP+56QWcdNMyjt502bHgGOr9/XZghUpZ6qoGBsPAW7+KDYwkFS+Z
RHH/fcoJIpkvwn/oQ5Kzwqru2HR69H+wVtTXmiijjPlyHCm4cg5XsMKTITkwggdD
aZ3i+uSEiyyyTPNOXiyc3mdzAx3VBNGWqrglbKwvrUGLEbettJ6+LlReyOH09VaG
DJgO2GBf/Fx3RPUWKh8SEn5mbSHq1PJsGRhTf3Zm34q6QiyJLSrIBTsvjAZ40c5L
18b+5sur1xTT09NWrncyGDD9wsqBrZtCOgdHqbvJfIT9mk6qGU3kzNEg/sEp1WM0
XPcaBn4hz4I6eN5/dDfaRaSgo2cN/eXDPJ8wJyIjZI8qVSgCDFU976OQfcq1feXF
5y9ahcoIqYvUCrBPGXWsreKIwr/NGiam2ZF99i+L7WO/hmBD3PWntLmm3zgPBwmQ
As7M0SEVzQg5M7KCayX/GETneV+rijh6/T9NnZqm0iYYMz/iGoA0DxNvMhY94PL/
lCSLHQ12tw9HCR5Jxr8bAFpIdrDUQKtNHDHbG8vw28SYTkx2zjlEoO/T2lybk1zt
jaspvDrTi+kF8K4iJshjaU8BQcbwcYhcgML7xSed4AbqesgwlHZ4RZdcxnosoDgn
tgQHpOAoXWRno1ylr+OoXDITbeJl5nhcuY0TXJjtOPEgzjlxPcOjVWBxAE4kHPqj
aMQnqCazXPvaFMwv+FaDYzyDA/EXi2mMs8/CfdI679phrf8N8tqBE+4nFznD/DiT
ykMZWg+48CIxb0CDk0MpLKsS8bOYJReiq7PwgITJCLx6WZAkH2ChPvKKoHKwqHnY
ZCEgcUqUeBjBFlQ6NfTJaZYqfaZNQw6NUGY+RVnOlGSLONUy3ulFhkLamlfJqpJR
vW2ZqfiFqjVEyLCB7zbgjYbExNbwruVGoUlpELGRS4Orbm3LRZuULILLPya9UYDD
+v5Z9XiD4bcCdna7FRoxe1lo8MywCYC73G5pnwmQZ4DOA3ylBkB2qGoMjLeK9Ind
xCDtswUllii3mfNCx+L1LtQ4F/jkt6imP8Ku+fTRoKl3oR+e3+Bxtd8IqgJ5Z3J/
3Rdkpzj2MsBi8ZRb0A1SqhEz4Br9z2+2lslpbe5fJt7t0l4ioQvTq2coYihR3jL0
x+swTJsh3RxXNTHTAeXXZyOLr43HbAsPaVfiazZ3q+e/YlE5wdZbvVJ1idAOjDam
FVBqiwdnqfm0ZNnqQnxCUTSReLQOABQdjTT67xjT/nR44dxe+v/L/UzVcDHVJhPg
4lju9sXTmYr57KkV1czHAyaf6FMBk9Q+iIuVVJoj5R1gUwt+w5Z2pOUQPW/kFLCY
QZuUvedCgsvnMcKPDTUZgdDpvRl3RJLh0YkrvFhz+/TtzDVVRWqUjdSOq0wl7+rw
XeGKeaZamabjwW0Q9iNzHmIbUR3BXpY11SvFMYB39yOvAikZ6cZj5F/8k0zDBzFv
otVt1KUzRI/nEEGGmUo3IPGBWz/TvDzlCaJLzlJcO59jTYKUNVWf6ty/w9owk9+Q
4d44pxiC6bOKawRxCDApLxH74CuVQsEqZXO/bAfLmGPyj5z+Y6axtbxipEj7FPr4
r2Jb2OYxnrMeDrYqRTpTGiU8Gs4Gu5uxBGacR7wK8lLTckDmO+vSzHtnJI9d1B7l
sVU6dnzWbE7q3m5NbHQBNeKUjBxzgy5R32lfqcPX9YRXb0KymkNw/ghnpW6qvMzf
+rebv1xQsmrRNT0awWFCAnI21Vxj/Oli2WEV9RqmL47Y9+PcaHpViHmKe8MHR9Ca
svWKgogjsY3xzrh1pIb6+PY6CUgQDhaJN+28ZW6JVwadVS5TxtxZaQZFtLPtGVrJ
DRzqmvryOoAuLUi5LLs1WyEMEQ4N5e0gviloBqphKRYWfJFq2QDxSnmQyM6HcPyG
pES9Df+SUIIM8LQ+QWnF8g0zTCV/cb/TQR3pmhnp5ZOfCjSWYKj/S5hJkopdOzOe
6E0XnfOQ2qJ+zn1HBaL25PogLmTw54FABtXPm7W7aKRAozxWZd6tYHWLqXjMVVVo
ssXtpMYN8nIcscJ9RKKjKLAINbALjl1qnF1EE7HRdYYBm23KM6vpDCOwVCXliI+H
rtVhxMLHnuPfblCUh5dIzQ2he+0llKwLq4MtlrNxcf8KDNnrHNAAf0RrBWoccof/
UxjndZ3d7eUfWvOq4KDigdDgsfANzud0T6kc0Jp46UBYq1jgWBEXQJ3088xrvt/5
7HJkaX3uLPDR6genuKSkW3Uibdp/CwdvyfUK0wTLYhujLRh6Fbq/SaUMovV0b8Bl
rxpi5KwnMgUsd+3Bo01Wzs8mE+VFbX+HAiLR9YAjJITm+KHojr3WQUrpLfaE2rPL
feaJrWmZ14Emo6+QczwoCSQ1Z9MW2BSBdIEyNCkvky8AK8XJjeqdC2iG1HWYkP2H
sjQtToYDQL9N6urLsMNpnsw5kN5SQTqGhR7Dy4nt45FNsoaNVWK8cug807PwR4ql
ZJHVeg9prFAhjbMRFLiex+g14HwN7hlR3gjJm74Cu5w7ABa2u+ru0EqxwlyuCFyQ
viDOxBKmNWTv2LuO88orPgQqSTDgh8/Xd7K7yHMIuE05ScF5KIK+ml127EPd/bb/
Ert7MmWO47X3810hKbx6DRaeF4a+GCDP6vxKFcMoLGo5IIUU7fot48hcPG9s9hxE
G+fyFZXHk1266r2hPs3DJma2pL6uwX5/gFZiuD84G5z/baJ5g5GBhzhDZLJpk1kk
BRCK3S/ofa4l4QDxNi4toaJ3jY9q5OHmOzCaGNwHbnwqavHL6oBfhzQNWJOAAYrb
eABJdIw/Z2esvVKFLNXe9GSc0SkhpKsk29mxu53WZ9CZIxfmVPvH492luHV3GQ6E
yO3mFBtI1Z1cd3++ZVPlWDbJz1wVe1fjjUYLcBssGoJCvu/iHFKDV6ce7Wtgw6Rn
ip3jKJcQkyaYcb/Nq05RcQfyLDh6MyZfrIOVuAtGbxHxroOl20tHeT3IF+oitNgH
Becxw4zLFnLr4P1Ofue2l+a05isjtP1Xc2Dy+cXpKZv6vXj5unw1vmYVFenG4o09
ZNa82DIOY6s+BtFSrObSHm0gdeeKCBFAexB8vzKTdzUHTK5Y/WCx3u6d9inqCVHg
QpQIJT+DASh4G7IufavA3sUKyi9ClGHZK4WA8cFTCXmzIynFDLRzQxotOqRydWd3
uV+of+AESOlWVMIK7M7IP9gnH+39NzmGph+Fa37j182rafkfwzMa1Dsmth5kJ3c1
zkbr/Jqrf9QUqg4DTPyDTUTefbJN3rUjA9I6Z46Bx11XQFUS0SwYt/yI4DIaI9M1
0GR00+cQx/A7Zp7a8ISWcJ/P1Cq6l5od6QdkFC0ZcqA9nqrv2FP00YRHmzH+A0pL
8xfZst7jw1UNeF9RV0d9v3UD08B8NTGsvmGIsYzls9+u0y7nYaqLZA+LFV1jGcge
WBMYk4fvq8lus8T14LTMjhi3OjFWCsdzkM7/K++gEQlGs6Puly0S/McfQxvXeJvP
AQXWZTPNRhrfmuddQej8NIpQcWCkBgoCkHcmvGgVFHmerz4VQO6bd2+g9eYpaSmu
IWN6WLLYDWyXZxzFq4Ed/DENcRmFnESvTvuv2RlWdkAEKwrSNL0crLSX8QC3Bxve
41ilOT5CRI6RXZ/Bj++pxPpyS4sXemk9TP2lxHbaesOAad/GFywgJCMcAuOHEAkd
6r+wfbLUnElNUFEHeNp7/zY34ekmLuttsXxURGU4TuJWfvBUetht2kigSc1PTlxt
C8kq+Sj9H1mZ6jd1Po5Z6bB4nR4NVpvHDcWYTf2MXH0l/9cVRrBnTT/Ms4M1GNLN
KJFoAAxtv/W+i+rMbyP0E08s96mVEA55r0R8fraQImksVMjo8OkOSqEZpvVfjCPk
OrTlSrmj+iof1npqc6neZmBVELLbTlCy7by1cIaA9FyurN3fkLjCEaYGTa0Scw0k
OZfdA4/JoBTkLkDtDtYvki5D0g+NS8lTnA40snlwU2ZCwHiRhmmO18QXkUD1gt9/
6EMxklW/09mFWKBQGkchK4r+Iv3y7XFudJ2f0XfcdM3wZoMQFj/Ng7DwligyddbQ
Oi9L4k0MTcHuWrrSs/ttBrvRnxJCQWYGagAjsIUnUnxiiob6Xi7IzRAYZj3eamNh
pr98rdyPr8KuoqQ0VYSUcsOKAF7tD/twIrYPel1XA+j6AFX+vfNQx3Cf485rlh2Z
h/dFsoBpypvDXStHMvX14EnwZqKsJ3Xr19Of5oF5rHxv8T8HnUWCk9YYgdQeBYkn
TFnAdLHxlnJAVGrUKuZ3sQMNv6j33LigUASL4bc85z8DbhtV1PdWM39xTdMctWwx
HFolW7DIcZn+VhAi4SZ6Or2MfXkqPn5CEo7KPAn/bROcwBrcUqA0Y173yTQwjwpG
2Uw/v5B1HowKOEhTXdv/wA6KEHc0ZlJcuXgsfdT59+F0AXDogsILA0OWHPHvDEhQ
MSnET33ItdQOvhRQG7Jun+uzSpCeCHYqHgeAa8TxcCVQSyVYzZmHFlyaYWy0W/M3
gqbgnE+7BVNORd+XK0RM6YBFdlP5qyYTIVs0OiarlSY8jfqt20KXShlJ8TYXYCqz
6dhMZJ9FryIYL3UEoAQgS+v4mdSUGXO+RYLHlCIvZhCDF5qleloataAjxQ7V3Mn/
u2xY0Hgt0iHNcgzN47mqg3OgQJjjbjBqFe+Unk9ZSw56GPBUm/EI5iJ7kodLPvXt
WZJetV5KPcRISg0YZlBi+tM2NUnzxuVu8xWKPSPX8y6yXDhe64kKbteJlx02yCPI
sxc2li1H06o7p7I1nUeXqE4A2ZaZwxm5/bK56AnMmN2MXTdT31h70CLvAelmJKu4
j++/GLskcsMZQLjc9ClKdInd3FmL5g+G1/AyCrj365NeniF+7Dst0H+btsbG0tCQ
4aEfhxo1GGAFCsycPS8IW6JfARONobYu1dOWcVaqPn+RFGQdC2UZXN2HxmpYETBy
VvW0KkWsTRVwAPqKMWjT1P47FOhvcF0+M/LlpNofe/fjOi2QU5FuJtTiroBaB/dI
pcFFKIDbQbry06B5j50drGLcNsUOCjTRYg9K+6noK1xiGaKiSNesPr1sXQD5mnLb
GOT5p7HbkSCdVi7aLGPwuNgvxOQD/Fxa5AnKV1JPWjFfv43xTkuvNGN5VAuJm3C+
9n8QRTE+N2EJNyyFDwk95wJR8igV80+OtNonNEL5yDSy8q8/u/kuTDZjXob1KQWJ
P20LvOjFOsyltP063sXAbIj0DvjK9R2kYOgR+tDEOkSGuTt/0qMQyef7RL2Hf64Y
Gqf1bea4xOGX0Y1yX+0G94YsU3gzTi+9FSwZZ0K0wR8MB9xAX++Y0sjZKzS+aYG3
G3ZfP54XBCm5zGOovoeNrDLOfC5SfeHVZKknMTuyvl2FiAj2UE4sfwu263A+9o76
fJdBIvxrK5kphblCUSlb3gqCoe4CKKRAfn057mXZDUeCGezGmAKUSuIxSOhN2K0Q
am/URwIYSEEfPbnfDAFGmf3vdyCtx/PhU4iwXpNK7L6QlCUoBG5r9bZgQ21yw9Kq
BJYqANwAKQ9Jjfvm+2iLC+gUACzLtFZRTNezml8h6OnpSZ7l+iKXo7txiOHJXort
zPXHRRu2OMaSM0bA0EFecseibkv066XwfMm3wEHXDnFjDvqHsOd0F6TO/TtU/Nj9
ryr6LSsaCEdDRsezA0WkGrJ58wF4ey9ZRPObB9zyjpx4PuiXQ31HOzGTPf8Xl5/u
HFBzSmvVY2ybvdEqAGCBDEp5q1Aee3GNMBwldwjXhBjdyMMb5+aHct2q8een7fDf
2W3GYHPLGUSDL8gLvZtPKSQhwUKZMunmi1BBLOB4fFGv9sVLqjWAOOnh8y32pqyE
5n3cXH7mKjT0KNjccaIdI4WI9lzCpESQ2TR7/AjHzKhnaYzdz9+bkzN8FYHEM1Zl
WUFxlWnqNK+miM/L0QlFqgIhynyISFcb8GcwwYaUy0PjAyz6/UFe2XSPU0yEjw9D
2xZAykCiXrigpWXDlJ8RgJJ6gJKs46MHS2iPTVYtzyUi+6a2M8j5aA4Hm0dFc7FP
UC7TAHf+xOHSK4mFlHLidPplhOcBzL2PuwYxIfJswJLucarhUJ9dAajGNSjNLHF5
mXQQojhJHNDbMglZpG4Vr5cV5V9wnkvoZrKKy1AJE4nxBImc9gEeg+l09kTzgMl0
zg34clMyjZeXIKW2f6imUJCsw3N9SM5a0Pr4gNC5zS8ZLENxaLo8mvZ8Ki/sFW2M
MEPJZuPijvDCUc+djoAmZJy3c0wrvz927apqeeCeRhVH+qCVvjaYT90gQ+l8bk8K
L8njBdXuZ1L32eFpxaTa4+oz64WGFQK/jh4zogzRkGBAdCegFkmp5mrEoEqRKdWF
YvSZjTiKVJIQrjBDUQZ4XKsNKCG19i6+ASr4TW5OlzrEpf1fxEK6PaIXK8d78evG
wFUlNocBvqduWXlhaGrkdMwGrcM+69WdgvifpNuOt1u9N7iX9PRpPhy/kN0jg4C9
dI9fXM45+IHXb22iKoOcW4uIZ3dUNly4W9iaaN/t8ufEDO9aj9OBL2huuZfeUSZe
Z0gDvIqD4DDecc43iwV7cUTrvHHB76ykevbB2oRrKm2vg3nQv8i1SSGZL/igtw2s
QeG1TtaU6aQIPPJqC3iEegXkd2kKDiBYgn+THWMMisiEtXIiHGpOXECMv1iWlZ45
8N49xBS1CR+Vz4PCkwRfXTCoQtlHcP96PeUkHzCIcgK4RSA5HxRNmtoVmmbNjCSU
fl7uM+iOICu9OA0ZbCHjZ+RbqfSK383OhKENCTHL16cp3NURqkeVf0eYc6ql6s+w
ACs0l0xPZMXkB7h0jI5oAVbYnLELMfBFnFapuHDaVRPJPB31udZOwCt9TflKiGIg
5EOGuwxcYdFtF7TMYNwg7Tz3sKe+OXkNhOJSxPezLIrS2LGMnBxeORQHb7sk+unM
3Gvr5uAwTJc+KXO/ogMmpyVvgqJOHjcIT8oDpkoaPNoN657u68YEmkUfQxkJRbtL
g7hSTZodFKL9ilAiXlQr4ARw6roNdlFigwwvwAgNUqPvIdit5OwKYk794hb1W34U
yAaIWllWh9SNuh5hJ7d2A2kDxAjIjz12KvV+IEaOmXLmAbGhTayQeJBvCF6lMHjz
rWN5mVT1s+4q+t+J6aepVbJ/6Esog9AY2HtK8TRZdoVkHGhD3ftljIIX7I2tRtD4
hpEsP04Y4y6KbrC4MlwMZPnci648mRKawxTrl5AyAvM37nweNL7tEFYI/KAJuRmT
gnn0gKigXK2T2+1rJqQ6c+kFJbsMejrfMBlj0AyZ/doszTPdndMU7aRxzor6es9U
zAmz1oOMW6raHX1VECw6Ve3HdXVkdGUYyTETVwyGfQk2JH6P4Cs+sx3DSdxSOp+X
l4yLm7cYPSzYluW8YvgJRTxXbO9bN0niJ9jsmnqO9E1Vp6WkhwwWRTE99GP2N4no
6LJlf+SDBJR6NKhfrm1eRCNa7boTSZs+EgQ6Skx2lCu8S/J7oVfx3Z9lxGFHhdn7
1hp7MJS+h3RSc8SgkVZ0mHu7140PvF6RPjCAL0ht98ctk3p9L1LleqjBtOKov6aA
529rBEdH0K3jt2LHqkHQc0LpqQyZieNwjSJSTj3NxJkbEZf2efml7cBwqcRtYMVZ
ZZTx7HWtdli1XE7sU0QzhGAmVyonTEx9X7Mfy9RccSZYOMzXSCq/1rh1KXk4B4s2
g2xY1pDkvgcHkf//zHYqwZDWVw42quVX8gDxAfEsGkTxgal42BuKYdJXg4lMoVu3
YvRPFIyH3UpPgB9oVNYlmyW6lC6k4kQBlRAtHwOP2NA0dCz5PxBfIrk+t3hTO+YB
wIo8Pu4IPVGjvDlLJVdpXcJg8iwlhlF1wyEmZqmKmjRRBeN1pUJJc66UXCxJIFSQ
EUUGG2Agzp17DuKNa1FFFYHpZ1dlGRUxnIqyuEebshJIXxEvf30aPRPbnAkKOeNJ
5miTUxIZyZnnmVV0OSq1/VfICSo3q7j34VslZuZEQuiLaikxDR9uHFyR5kdK6bV0
Y2bmiF89jCrCAm4iP2ddYXV/7DtC42JeDGhvi35XQV/bjPXtA1FxQkM4oClN/AmO
SCx9Ht4qmn7aLg1f4yuBDbb08bFb2Vrjj3rWFWTE07egApbRHk7eDUDHcV3PmGLr
bI02F7UoprHpqoG3pa1CVc6CkChKh+Jx261yp+O/nrLgKYp1Ys45s1ESlPkN76ro
TtWbbSMWvaSh/fS71wQ54Xdj92IPtP/UHMpQPVSXVtuYL9/MQ0mjzUk4jSspq9y9
E7Be/HN2k/0aCgGLSc37LhYzaqV3jWOBTtGUwIQbT2jUUphcz8syq9gaebmJRXCO
XUb7Ng0sAQpKNpisNU9NvaUm2jCRwraKb1WS0mNWqPoa0tfV1YwQBJiL1oYENL+t
z9nPt2TX5LfhS97iBGqHOSrMlJJucS7lEYe1GRy24un/kCudMla5R7PlApTkH71t
nwtgerpIqwFe138wdZ9CbRYkP8E9BvWrmKfqsIWVhGQ86fI86iDaFvfGWwBwx37j
XnrHgFISGPX3E0qZXJA66VmB5moYZWJPEB7oNNxc/Y5bIw2Ir1NqD7H1haP3Yv+p
PHsIsDBUgH2wLPONJLHlQDhUYH2xBT8Rrbc0CU8p6DPk+njda1qkQjRVTMQYGV57
vrEXTs6RI+hA3ss+z+9rF17a5qqPnwl73ClEvEJF09GBztQYlxFbiTCZ7/ZvE+Nj
Mc9uh7nfhOF50wf/bT9OWu3XQbYcYpVx9Nx1dLXDgEUQoypgh4KVEbCSEW5p7oiL
2zC8qj1TTKHmQrYPkneiiROVcMLAvw79S0a/KUg47pOVZ/5XlU2tbTVrPjRSSJJf
eaHRTTkry9yHfL+My6l8sV6UnCul9wKdM4iwJmvwrX/X+DAGmxQYQdYPKlUmy7wT
Br64Z8JLyfszHza2btrmimjFzRxGcCANvhIM5wPK7hH7JY881LHCM/3dkAOYoJWR
Y/KaO38DUUOfbh6gDW9tmWWQheCMBsWvTBgKBqV8CL+J3y4AIOxcTY5v0kaPjRTo
Q0vtKaFhUjUVfAPwWpPatoU8EctY9PBTCbhZGNGYX6177zU6O/O7GCkq45R92E+2
ZLIEtmeAY/nYaJ3dayeumvZPloUXOc/aq4r6w/ZqoLeNvWQS/rdvFaArZ4dx866j
gVf7PmkInG8MNecqAUr9bjVhMrF0QyCCxUUbhTdJpTZK8hYZ6of/nuYRKgizwQ/t
VzkNEjT8Fse77oDPrHD3v5ZVJGh6WHjAwJEKYyoOzyoNwpmrsHdJLe8W/wBS0J91
8ygsG6EDcEEPTBNjVS5NiLR6AWCcaLwJUXez2pBoDuE9qpTPZvtqF/eCi5MwwxYD
YoSaL7dz5fMnPa8I0oBmawiDSdk3eHF2UjG75hXuwBgPua84Pq+6qw89DrmXR5UE
xUTIQwJoP07DojgBxR4Vaj3fa0/NoBPTCGHtCjC2uxCNVYOUL548HvE5nlAwbWs5
0palmDmrwnp3y7VLabINrw9OHHVyMGHM4hQ7KDJa4kWXYTIU3Isg/cEkV26QrJ/i
t5gLjTkBlXRVPIlWaab83g6g3K94w3OCy7noNX4Abmzl7lvsOegtF+vktbyDb10g
Zr8/EZpo77u3RDhVhqJTJu+kT1WiqmPFoIijw6o6PXa39gWRrBRufqCIxKUlHk6u
p1aLJILPhehkZciErpJSH0nGlgvbb4gdvZlxLEC3R5xnUjs6gLT7gSOWiTAG/GWW
v1Uwtvx5AX5X537miDqoRLcnDsRrc7RNIMcI/DLA9uBGY/qO9z4tTx98NWqH0/41
zkhkl0itWVzZXeG6nz4U0Mgfszh6NrPaQzB7qD9kulU8zgDiLd25jetPs1gEApYn
Ip58Mjgo0h7X/KFp0JKiSh8e4kemzma9AIAZzKyZl02RMQYkOANf0t3yjSlAUhqo
Wkka1zG2MFHXxYNSAtlbo5QFjyRP2iuTUItQMmBo11oCCYgNv6VXvv8jJuNyBj4L
3uj12pUL7uJHduYzVviY9y6KcS1CFv1nsHo6Tfx+eVqFmKWZD4CoCnIsijC5lvU4
ZbOtdaxryb3gm68+fzcxUksFVHVDbd2yaYF+otvd1D8o2O3MFYItWcGCNJrNfjzR
FiS+PB2NZKu9Z+zxuIMlHHFYKZ9hGhAfbn9E52rW10gjPVTxUp/UncPjErpoQLMi
VUKWJIC15OKr8oNgrPYY0mjUUzNhJ1EewJR6jskat0yd2Ccxkp+z3Jf5eY414ZnS
LUTBtRTOS6Y3e60fcpcl54/1bK+Bf+SiDz3MXl2t3DWLTtW0hhZX+oMQrqa3iFNg
PM/6uh9lypcjGfaI+CIPyx7hBMUFWV/ZzNXS5w2CziCZqOd3DLA5ng+M4gDmOR+z
jgttD0xhJlb+o1L9NhLFrLfZyiG4olxI9MgmZ0c3n1oe4OKNXlqm7tY/lYeUnZXA
Rr9rQBHy0WDP+56gdu0ViCOYU90hXwbq+8bnk+a03PvppHB3sBDWOb/eyERymA8f
RW6x4PXQJ6O8YkOinOWKvGXWltIT/FNx4C+xuHk/Tj1atkTXmYKk0l7SPoG3q6sn
2Pg2EbLLQVcx1GT754YL4f9vTBif2ae7h4HXJiaF5sf/OckznwvYo32mLWTxalL/
xQI3Xhvjwe93Dwl4g0fmb2j3JdWJeu+ROeIx/wKaLRgfsd9TCbPki5eB81yVXwur
lX1drFkVgumiWhr2cN0QR1FbLrkwvEdsgi8FgAiuiHo2HdXtIPxjP6tlAadf0YsO
3lNzg3mkhvwbC/NK7evDUFAGGtFPjbkWS5PMBWB8nsDD7a1lVzRRo3+Z4lYA/fLz
/UEDsWi2UWUH5COES2D30PBZ64My+5IrVpBF0wsdb/3C4JyW6Q6g4rkrPqcIA74L
AduGUcinu+CE8u61+vdoWNyr/ozbtdlpy0j2tM8x9ncLkS80W+WOZa6fW0VcGm8l
MjBxVn+fijzEKfpSWo8XnaTI/uFwEQUbYIycTwCemFufuoj8kFmE4Os85fG1byWb
El1FBJYyQc8dqx6CS/wzUehjjhj3vutZpWonf4bINtfbnG/44oqkOjBepVPxXToP
iieE1LgLnjvTDmfZV++CCL+2D9dHFhCUprZvjHwIVnDPmOnWCc5zU3ieS/71Hf1O
O4QmjIlPAzjhitINjLd6CtkjL6rQHkMOMdWA5NJxJU7R6uD6fvcoavzWlDIgzpiz
Wij1KS7UpHFMPPOtxkAGgDhmUVMGy6A4e3tglJlXL2xpGPNUzJFX2bIZ1fhm2mvD
/5uZnhh9r6y7LZjWLS7xcNfEC9UrvI5z4oF+DN23hGC5U1dtv9Io9Y9f2NblpXf7
elKjz3IXuhFKPzAaiPlcZortcq7WrlT4b1v7I/wsLSg0gFZKGHbLXcr7rwGZx1VF
xEX9IAEa78EesCzsmZtpRpADPN9unozKsGe0Uf73sqVYwkVwbznIgNSlx+BdQnP6
aQoeMwvQSrfkIiAGDc9VyelKyhZwlDP7U/uFu/0MCJuGYCjjdjITL3fO4vx94C6c
OXHIxCYzSCOSerqBPtCAVIWgKKiXfP7cZZ8mpKDeQhBij+uOTWHu5yWnCyT1vo/y
dAX8r9kpnJzEtu/q+jMr7SQnzv0S1NPLQyCw7BzYVK0PX2X546OHibmANq2Ac9o1
CGSJppcE9+AtJ9QSu8sbD4/8UoYw/uw2GhnGJzzGAAH6GumJ0avgmozCKTn5Z+LD
eNlSAet2tlV0iwOmCJ1d/rz1TAbYnyIkzzfvEV7SHF+xQVZ4ASXntZIW7Hljd8Do
xxMvYGD081E0XxeTQF9Uo//Lqsio5vkY5FamXTP3crmF574jAUnRVpjTb0xqwxCF
7FfND4WADHAlSYFvDLaQbr6JmG5oTFhccwB5LJieX4zWq+90jSmjP72+fquUvMUt
2zuLIK9SdORF8Tg5/DxP2C/7rpYHnfl05uxSgVGfwuPyH4yFddXF0JOeJOxg/epr
XFopaCwuLvZFby+XazY+YwKQiFO8viEEPbzCsEo811g9T/x2oHHe0ea1zke3SDtG
cImswO4fztP+ekBwayA/XEJqvmuo0Cguvxobw04AhSkZ2xtsKFLIH4EKTxt6VcQh
An5hIbtic37mFv24Jw6WP3BB3etZoAV7OtvnYIWHDHRNdi7z33L+LKrUljaL8gxK
Ota8F9HCy8BdBu3yGtZUyh4V8wquU/1Ai0YsoQGpyo3vYY4EdOahL8KO61OOgkde
30xjX8C0P/GJUiNHoP77Mw8P0uGZdvTAPt203vD9XigOadgFcZLj8i9Pe2ZRZqwA
kpMasQM1FGIhXqgh4Gy0lRUhp1iYp0H8pqklEYV9JoOsl01KsSL54/Rq+4QoO9gx
ACTQRtyMId1sM6tJte2sFUNr7a7ZDl/GGKJIt0CqtiaF66Q6GMzcVedC3O1b+x6i
PXWp5sJUCeyHKi0fK6g9UTp8ppnu4jWOYMOEq5QA9/CUYbDCgPZC4QJRZXdgk1C/
Nj/e1i3Y3/TI24Fl1uFbJAL+FEdlZBCW6YSuXNDB8p6flejpL/ngwzkhw+Ae1ayS
PEGrDSPw5nb5fb/b7v5jlEXJBbg9eoo4Okbdsfb/kEw1QlPy+ayMZVCZYmK15h1k
wt58CHbsDpncgUPvHlTWIrHl7pFhYoRtCRU8zLrWouwqnn1dzOurRB3bOzn9il90
YZPCZmiNdfrRv7fkzMmPxN7IYzpvqWOtwjMNieHV4bXH+LEwoZJgTIB5G9l1jfur
wUXlFxwg3irqjhqCXT0WxvNISyCM59hJs/Zt2vPR7zz8pYobFVL4z6jDgPquirk8
/NbBdq/bQwcyPTVeh+BQVKruDa8le039j0D78jn2tNqXylCh5cGkb6LpcN2N+wtv
JA26KfMevuiz3y20r8ySOV1Zz4qccu5r3b+aVfhf9KDXj3vhBb8fR6/8Ao8uugmk
dXJj8ukoQMUNrvF+CWES977+RsnrEcejQMgFv0piniNaOluZ09EsMgkQryS44jjk
40QHlYGWPqQz++VsMLxH7mAYysZVRCIPGqURh2cndNCC+EQr6ga2KFiv6vQSd8Jm
E8J8dUqXekL/4jl9axVo69z1STC2r7AoLrlmMnfSuYDnqxd7FC05XyW/0UMbHQ/a
CCsUQ9/0iqeYwss7WSqst/xWoRQgzKSbQQe5S2iuHj2cZFCWg7wzCXqTO96HmqKb
y4UFogYQNM2gkg2bLwtiap6pD1hX/bWdwN0+pt/GwujftxXi3mdcE6voVBzqmEUe
m8mh+pQEai4pTuOFdLeuEuXWfMOWMnLtqkBfl/7W4a5Vczwj8S2v+GA73HYZ7XHF
Ix01qsOAcKEo7zSXongMRHsbzjoByTQm8YNAiwLcrfyH5CYMlm4kXTqJWnGq9Xsq
CNH3UyPzSh78VrjhX9lWFyNF2/lKB2AosxlEdQ+OmQ0wUAks7koREWV1LhcfCwao
/LjaJqaVWigImnr4nNJpJQr7CWD6RjVeWrb5Mi/wl71XaLaWZ1V0/wnEs8Wp5Zql
iH3mfvu3bPzDCee+pmpLPo8Dm3xjzqX/VbJn51JPh2XGttnhbiJnkrra4gYebsJo
3j+m6l0xi2sVhiIqCZEd0sRq+vrm4Pnj0frGk0n73uE=
`protect end_protected