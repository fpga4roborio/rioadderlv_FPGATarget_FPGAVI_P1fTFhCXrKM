`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
ddtXksX2+yylW5zu6QL2Lhnb2d1sD00763mmSITNX595NcHTEkwn0zB1Dry37fOW
FufOhVzEJp80NC5qZ/+F0Vk7Ik02dIR0elf3clrjeJRK85K4e3Hoo4xn7YbFUIms
l/8VZSb14+JVGURjfswrIyCUotIzlzVYZ6gzoZwDXIi5gQIBf/gI+KxNXPaKV+PQ
Ufys/12rjO6aI/pPlqSm0hCvftmBcnezN2hk1UeXgOIuKZnogjOsf0iJVX2aOOWE
6pD/psybjbnsNB6kH5uFTA5frkzIzkzl5d9+YDm9OyC+k84E83I/7/j+rk4L2dah
QJOvksSIzN867/4Qt8qYTQ==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="MvBXkzurAa5VTw+1JJ70nePUfoQXBvZOku/SMmg4TwQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
oRtzZL4VJ4iwysPsC8SXYCzXS8Fw2gtZTOskLcDV+1B9Nzn1zTyNtlo6lNICRmmK
ZRVu2BmCc2G+fmzynYlNTnSa7C0Cuel6FYpxCBlOuk3OF2tzAmLAuDyOH3Z1Yjzk
a0aHuoCdIRKv7BrZCdALt03JeUmXKPdOmIlkVGFl8yw=
`protect rights_digest_method = "sha256"
`protect end_toolblock="Jn9CQpRhJt4rnzZPRk+dOpzAubz7omckX1MrFd4p81o="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 50608 )
`protect data_block
gD6l00tciPUa6pDNTk/+tzLxvdHE2s3DQL3/JqqujQBC/Ei+vcAB8wM3doqg5vTg
mdfn9XB1bLOis2CVSfu295W2DNwHfMSTc/8BhCDRnTlLIX0UCJs9Za0+LoM0rMrV
T7EjVWppbP+Em6PkVKCwlmIQ7JKaifJ+Y+kjw9HCGboYo5074hY+K/CBbfsBQY86
AyoN0MKhsIx+eViNgnWjAw/QlPdiPAswm27LDiDhPtMGx1Pg6FkXy5lpRv3pjI1f
f8I6W0yuzP8Xg3I7wP0LryJf8HgL/4LXWK/a4jJurivib/gX/NJsCMij2pmwBY7I
28azS+dL0Q0j7LKrecwZCEhX8zhMBLqa5m5kc2Xac29e/ZYLN74ddtdTD8y29ayU
iKlXUottOGZjJeMIHFvWacVBpOQkrJ5fxEL0b4GRtOBzxv7UqF7oBeKqNEptFXCA
76cPDG69mEkedDe0yzhYp76QNjNwUaK8YDcRMN08qmkb+v0NQPQFS4hLkBiBxxwT
f4XUC20jAA0TH1BHLe5ZbFVvZrEWkvwnLk+zbYevD6i/UabCU6lapv6O2sBudsWp
tBHltJJb2mlBZdjrX/mZbpQNHeZQwieV+YOtrok6ZnjSMLRkDpYfpue7vKt023ua
WUwNGg/SwQOkuPMNEKftVX3UeSJUfSqSH6RZ0Z+LlPp5mU+ZcDXKDTcSCFZzIPAZ
Qfp80gnqXRrG6MK0LB9IOdTHXEI/uNP1RZG6CEotQUzEiBPV2Gm8e2TUrRBpsEiH
wegOYd1UIDdr+iOhpDg1Ow3tggu3Atw0JKChM9kLMCkMvZL7wnNla/kSTf0+N9TV
rFWVlwgqKDlX/EYkVCNF7uCnL4iRkhtiIzBo4c3+T/SAM+a5LvIe7y2dAkquUSRt
P3cZrZV5/oa4L8NLX1fkAkjNBj0ZYTakl8+GJgj00xwvxoLXbIBWSbLZAOJIkNVi
PS3rRD0cMQjj3xqnZbxGqqv8Ttuk9kG8VTQapkUq9NzVWzhvAXXMWndTQd0DDJwq
8TrwYwPiYTKozMwMIEru/3zOUB/47aD4fHTaIcQPRP+YyVmOqACdYuWW8xQ3gVze
+EUJxmxqF8iUlHBYRyni8QepQEx024HTxjEH/YPV6jcXGmM9PtBH6szEJZ9qACwD
kerTlaTAPNDtWlAOwBugttWEMLjeeNDHd1dDfDeuv8jlGL8i6fWJAJvNN4Bu8Vp8
GqcDzNGFECb/X2/MkCUk2PxuItngGVXRnXXEeyLj7VotQUqsWPMLtxkKg1T/gkuf
EDBukH2K+kS32+N0nJaLWaODx0hI/i8DhugYaIsGOSTnLHxKU9tlcRyxNiqdaXMO
Zd7xOjAnZceD3cjN6ce6XcJNNX0VwwLNqCRrzxL62NCPw1HkNP1120AhKGPsMFsH
bGAx9Ydq1iTGgOYhu5GXoOFp72xuWkaq3vt2HWpu74PfgA7rZwSMufE0o3UVNbuq
ROFjy/+ZXxTff7uO2BLhHyPywy95zzc4h8tvOdCYDHMhgthAJG1TUXmbshemgjDC
xpEmHw4iJqghSozG20BIHKCcOoYTfosI5ts7XxPWTSGpzMvPHaRteR4egIDbfWuN
VOpX07A/ackeq9cnItQcaEEeQM6wYDMgoFfiiQ/Ox5fTurU6yF9LX+DcleCClM6T
8/x3G5TisKZdoPReljP7lHcBpTBO2dLz7i1Tac9GLK/byUHlttzbdpmFjPwjXJP4
BHeKa1px/Nj7FqUVPwSLCHAepDoSEHEWdFyOeN7mxyBpoE/jl2pgWACYcP4KBxLt
3zqOw3wyX2s/tC3Gd9M3bVISbcODiq2qKGY48F/GGd+Nenx5HJ3PijLm2BqF3R2V
Invq7J12MLHPoru/ultkQ4sB+rpaz8MDchG+XCJmQh/D1ZEWgKHr9b0kPv5mLXey
jxkv39oCbriqd9VIuTySTf6tSwejgBvkYd3xw5GBGtbgqthcHclnajv96qUHtSB0
1RNyotcVPm/utJLiEsrZEDBftY4XPjT2bHbiEcrN8/vkj97AKaCYPm7TunPgREQO
CBjxvLZta6OMY4gCYhM+zrG2tdANQaMTK4sNjIqCgTccaNMRyUPcMdujAofJVJR7
GGVf0pT1A4FZFdKIcMESH89KTu8EopnpXNlUOdM0c/gguFM2RpW1F8HxJmEphEso
jPXraIyPbIcwsVd4U6VIv0hZyI+HXLdFdnpGRYKwcK6u5yjBs2SV2n2GdyfTNHTM
lLur8Q22Yt8FG10sFI+thlFcFjJ+l7hgM/o10rTGLSWv2Uk1LPDdizm36bR8Ji4X
WqJeNPnyTKewy+vy8O5anb6f1mx2WG/GvlcMwKSdUhPek38vy8giFKQyGO/78bsu
QqsWAcASLZ+HjIkGydggdWjwXqV36GpyDV5mtBqQSF/QvG9WdNhzV/qfY/FY4kPe
MrAzI6jXyh87oEQSOZ2vlh9IuY926WQVD6WtCADdLtvVeNCEJXsmGUPkumXwhFTe
3WwLmattFFDUp6imPHT+ldkJHiwMT3MOm3ekdJbzPJ65lL4orzeC61gAMEpO17z+
KuVkcYsgETqZwg88UQbaW6nXxcRrV9/3xn8BW49kAmy49dIOmgUht4evmo9Eo7zB
DRm+bd5hYtxwTXqvkUq8M05gWLhhs7MJQSrkjT+vkZCS2QXcGw245Y7xQ25EUHH2
GPL+HKbzRi/fDb9kixNWeb3/rrgChtiGeh95/Dob91ZqDEPvKlWfqLS3r9cRFhCk
XYjp8RmQD61p+cNUsAkJEZXLaloiH2Acon7qRlLC1WEDXKZoDBTRtSFKJZRaG+NL
ZEElaIrmcfNvsjhzyhlynSv2w/EeyMjLdthq0nzwgnS/pyI7Xgb9R+vLAm83ZJhJ
k1Tw6dC7pp+lFAh9n0wTcKiVozo4+A0N5tmqfLWAnOPQLTZXgaYQ3+k0hrkY5+bB
dEkSBZRTm7taatmsl2//D7KXiTGffxREPm+gIWQFDY4X/DGTYx5vybLcz7zhKKZE
BFqMmo7NRyK1sZHd0p42LVdHqjD3p1S/L7GG9ViMkKXY5mZlYKVxmNQ+TZYS3kg7
LFsckBZZ3pi2ddsvFJiax7sc/V/qEfUflWNdPmfrQ3k+4gJuS2tzRSuoqpvt6iTL
JB2jhtjsYeKL2Qr4oP6P+ryDLObVWQxywjsgR4bF5W+sLn3R8lkONY47f0dZE/gf
DYN/vLMYKeA3ndvzt1IBN9bc+o2JDNYKK42cEp8p7Mif7FTVGJ5yc7Ausk2q0R5k
CzVknNwkxLwq/T/rXFiCSmB5RsD/Qw7ji+DkzQPb8LFeqgw7bO2h9k+M8RJYFT+Q
k25/KF8dCXEzAWPWayVU9+xrDvC1yOjkJouXAdoIxIr+t2WgD/3u3OjTWeJlShI5
QbjJLWIuSGN+2S48TQNuNX5DQ3eBHQ8WVrvhbHjQilbHfS6XAFDRJP8toZ3tYkQ1
vYNZj1bvObm7gVBwAVe2pjH27JPoDza/4yJ/PLub7m5gQusFxaOP9Z9pg0Jnx/05
u1pcrvRxVRXCcngBmLbHjUcMdhRkkfZNjVNmd/gnCz9Q1w1hM8FobEUOu6lk/O5o
LFeBoBYoCXD9aZZ/MD7Kc71qPsQKQG042vuiKuopIcnLinzr7Nhx5GW1pUODhgPB
go/fwt1PEz7ZUvZLH0WcU9A8KalITTVRbw+Q9je9AMTOX0CREUhWgN4kh33liZNT
q3nF9g87exyIO+FI7xB8A7+yRmigMUtpy8nHrAX8W06PEeAYqGKolkf/ZIhiXtpI
Zr0jhoCUrEFXOhZewPgLj/a+Fgk+CdRouSRs7fInLJr3quhhE96NAmO7ocb7hqyh
rnSKArjBfTt/WjFh7TjY5xlBElW7fjcip3duugTclFaYO4Lno5Pe/YrFbypBH8ZI
rUaVmz4G7YzGtp8zmGAiU3r3f0McOk5/eRd5NlRt4nAAKfb4b+iRjy879Q7fI6Xo
dbJg+hwxqajBpBfl0Vm+dty88PKIg/fWL9ME1h3p3Ho9sndWMTRJclbi/2HL4XyS
pAYrDtrLaAXhhGcok67OOZ3IPR8breX0BXgIwdTUa1haE9Qw3RNOxl4qCk5PbkqF
j0K/HF5ur4DIFfX26/SR3N8E3+qt+xoyBjoNFn86jhzOhA/7gRqEUTj7OAHDU7SN
o+dxpyNDX19V+Lf4whvCnb0VPxSJekZRXm7uY2Ls6lXYNVwBiVkaLHTTqBk12xD8
m45AK3K71c1Y1u5DOXr1a3y2W0sC4lW/H9h0txhrPep87PmsDtsNDB/ZjPNn3ncA
5S+mNuf5THJ4GFyAjORFJyTbjo+MU3IbzZJIdddMG/PFd6FuBNfLVjBiyyHmeFO8
o1MuLFRwogjuGK6GB8gPtBrzoKJI/f4+D3Id76ka5AlB9kA/nsoTQZpSanpy15ud
x8zAjuz6LuOB+rFGxafruVOLeKEIsLoclxTQVohvNH4MJcUGaCwqANbZ6xP2zuUZ
5jVFtktLB4X/rAD+PS+o9J1eoD2vFdugiEKM5jymP6AoMDnq7Is3cokAf/Q07gzi
a/uWnNSCmc+TceSZdqjBvnVOBXk9YRLGe9dOyRudvNQ6POq2uRtdTRHZCqaT1iK4
MFxMKYZR1VbClMPCnolUTu+jW69e4Ma3h2teZCYpnrFg4Jf1cDd8QH7D7EoPQX19
3sd3Qv+hlix2yTDv3zKzNE62hzSbAAqkHn9Z/NoWbww+96DeKbudDYDSo98yoGUy
l0P1xMleZ2HPYXzoqY/Df0JvNCPocPKpHkekm5Pzvim884ZfC4rNfz8U7go0PbWA
Qa3397ih/+x8nFbyLr+yu3flTiSqbZx+Em5vXF7C0hpmqoHPdY8Ilgx6iglE38ga
z1jK0v2K4OE/Wjr220UfcNXWucjgGIzfwYn2L4OPa2VrFFHq9ZRLseQCmyOwHVvg
4MCyA+nXnZBO3bGwjcOdWZxJKc/7mSraVXSoqqw7md/tzZu8GN/Vn+mnIMulxAG8
05ShGIjrDT9T0vDNDNMehBjeO1+Zt98l+3WuQ/z78g9fn5Kn1C4oJ4m/QDS3BMjD
M3xAFanLpGROCQ6qcPGEllABO5JlFSfA2PJ/BNWLK+cHgvqG/TpaCvnOyguLBBoD
tU4pBx/q1vqz8Gqit6uX3l1HRLncwEMFqAcOx6npHOvT7OB5cDXcA81zrtLPdtmQ
iiI0wf6QCI4nbH7MSdShovUSgkXnjbcsbQzkjLsA1bbRz3G4U6GBpZRenlR/hHjM
BPQebnt3h5Xt0rhBbttSSS/GedvRwsdyuvHOytqfVg2nItb7Y12E7g+OsnKvHXyY
7ad+vR5m+0fpH9BhXiF9jKvYwXp2M+ASa6xJFjlmoI88yfLuYJJLYxZ2VAIJUUpk
aawp+ZTovmGcbXF+BWeYZNX5zvAjHVYBcAk/bAWJZK2uAPcdzvwkvrkLcrl5Lzs4
ajScxwjn6tb8QGK/yvzoaRML6SU57kCElnYA5bDQ9C9Y3Y9pLKXetT5JPJMltmzW
uwYvlT6Uv6mI3TDtyLF+1jNHVQtg4CZmsOVhAwN4JwdZEag2i4RZ8dq/ubSrB0gR
Qq3zJkmiWl4VgxzrXY/8xAGJOmH2jyIPvftFr1adeDLj71THxTY2dfXwaK1eTqof
KSMtZnQkR++tkgKUgLelnXTH2pAp/v+9hOR8x3KZb6Iwpr4FfKk8/UT79zrdM1kz
ZHUSAEiPBBNyRXMaltIQneCgNl9rf9Kx0bdpFxticdbOo0peGT1KaQgFZPwJC4i3
eH+DKZFkxIOCcWM1T+OSHwlQ/642knO1c+9MuwyRTazyIQlJmbOwEU8NhWZ+Pr77
o/c97IPHJSZ5tU1+K23EFp0jbLcRPvkcNElqmUb88uzQCDMXMtr1zr3I50MioS3K
iJjtoHFB/f+MmQSKR24ymZ3HO8vo5Adi+DiLs6B3RjM1GWriZjQCzEcocFn5i0X6
L46qjPoed0JHMRsUHmGCqVU/PqRclS2qRNVjKoib4Lr7qHxbFrcEGfAwYQczxiHq
50vmKhuuCU+QWhT7lh9iSyFObzAercO5ZRZMP62SG+8frKIfhBgFgtjNBVBjZS9C
/F3Z4MkHzOO4X8Qxk+FSPXDy8LIjlMUOF7/1CDu757naRmZOh8xmO62tVqISVHAc
Zzeb1raGSgShZAqRE3IIXTby1UGDOs+VvM5B7ITJ1XfC48xdENFlgMcDox/rnb84
Oke5icFnT19qF4dnThfxrcQpW8fUf8YXc3+hcwJExjP0rmREerTHLyHajBadfkuF
x0SxCojX7gll/gsPmzpqh6MIwXBQZkuYqfcMp3LA1+Erdba9HMI9o/N1c6BcgbKO
LLtRf2uwwQbsT7eKvLfDl6/18d5vJoC+CvxVbAAQ/OV7k7R7WrIEjKq6vBR54vT8
ar0vsggfX4CGusPF8f37vyEqDWueub/aaOTLMCURPZ/Q+TZ6dPfjjCmOZ4znNqUk
dn/q0qt1H2NYtP1qZb/n7Z52aroK2qqTG3NMz5kXLotCeTzn+dr9vIGFuH4c9ZPM
jev1bM+Tuq+7geAW9/yKWER/q2fPk2a7hEr07plth3jd5iNxkaF+ZVEzcfwPpCI2
MwDlJLnVyi2coZs6JV5g1itAXo/UNNDdyuy2RDTs8Typ2iG1L4gxo6NHpV7XnqOo
uHfzrNOHvwQpFAxsPzwcNzVSjaiU8acPKY+MVFWF6lggb9UYSr2oPC20Fdwq1UPn
GLR3J9OYJ+AXSOjGWry7s22CtDW1qCbDa1wuUSSJsTAIrNVSAingvUfrfpS1F1LS
qFVgmuBhPjRzKhjLnxyvmlgWXfcFGzSOhkdRwR/poeiTSS7kI4BWvfQ31vHEHb7z
ybkzb77w+bvOzVTjoYkOSH8Lbq+gYFlzH7bpK+cZ4UpYlUaa01T5S00/XwPf3ISL
OYt6wc0a0iq3bEw4uaVjuJ5pYsY7FlfHUPF8MUWKe7473fzN3r3KKU7hs1ElyVoq
FxORJ4DotKURsolGD8HS2t+mOascLR2/go31jX+HfJl2xSwHwuJXZMQ6Dg7odLmW
M0Gtt8crYxo8BndrLh2xaI3b/O0sK962qNBniYANIceYDcnxq1CNDRr/YIOWhWsi
lyh00zJnqjqvqsmCxWkxuWFGUU+h6lwZGsj4LfPwg3+1KwwcT0ZyikDtJo1f30HV
fuW2CPT1j155omCVRy00t3afcmVuP6s2aeQpRntDtwAln4/obBKS+Szn3Im9/PqM
zLmVg/uMGlp22pEWvlsbcXT0QsJNPSKhyi7fvDdE8h41woHuVfe5xXSrnJJQ3km1
VnCL+UxxqYjtmne8bQoEsFxuFsG58XEImoJ7TISm/fcYNzvhI5LfC/u+A6AJqbJ4
dKsMSQVOujZXYe25dMEmGv/OBuNeD4suL5mYxx0nIOelLFoQvl9aNN7QQ7NEzP/0
RuBtCDWFeW8y9Zj6yGkn10dK+EQ3/0aX24nSN4EADc6L1TG9R3z7cRWCfrqPQRvX
Tzvn2g14rpL/TCsASQiXJEjhsMUIwwY1HTWnvZYBmGEaCmTtZlg/NpbHx7RJO5Uk
/3AKGOgJNmOPmcvFIvQ0DNRqbzzjOJZGWPVBGZVe517AkiszRwoonTrZqx+JYsEG
T0IW6RDCyCfnXgOfFvhkM3KeQONPsp9eWbopuxhdDoG7IjAzVK17Arbke5HE/wml
MLyRh2IAd9Ckg1qiHAebWN9PwZE8nVnev7JDUOJHh/Q2JpiwLMk4O2+A9RX3/LdK
3J7YAdIERMD3cfUwnI62KjIQBIOurFWTgxgQnWXR374AsHYK6SIkb5tePRL+Hq9Q
abzafCaMJ7v2o1c+1sDNnz2aDLItfUhWUn792N7MkynqKAiyfsytGxzsxbfS+5wH
f/DdNQa/Y6xhr2T5pVqUnin4AYvW7CiB4vdtoBsedtY6tO/c22ArwpDmx00wOH8F
UHBbG4SdYyxH7t/wn7ljxY5ZAuPZdmn4mDiq2lxs7aHH2Tu2jGqiyQaGoXI1zgXQ
DinuCGMBtHgSQlGhWSmxodkGUti3/H4iwtUxaHdNcg2siPUJjLZKJTiFMaCod4Rl
jBf/78o9dB3ozZcv5nYz7F50WNoyfX4tD9dVmGo39oh61bP/dXfFiQ7JK92/DAl4
8JMOvYY9diM7uLzyuKIIEpsrptipmEO0D7VcFaqXCtpZaOj2UnXdGDrW8UHg+cjN
B+UoMZSChEF03Y/LPs2c4S7XRgwPPan5qLrWUUUFP0I+MPmCr9Y2Zn8q402GkPjw
9Wwwx5C66cHOhr4YsFGsJX4g6tyVCdIqidh00xkE9WbIbXwb7DbNsNlcEs48C00r
nAtcdXD6isNEQr0PErQMXgvwB2z659k+M1s86ZQlwd7IanNvW/f1kfxuqZbPkipr
U1JrCmw3qHb+iRt7S0r9a0IuIVv9r7RgL51iR9kJ8tt7yg/o6gyPqEgkLldBg+g4
3Q9LppeqvR1aZdLZ4r1ZQHzn7th8pj1McdJJfGXUK6nYk8AeoMU+QDmApEsWHFmz
5VEk1aqaQ0j7t8g884l1eeCOZoPHW15oZS1yzxy8q0pDjij17vSSNaTCOeiHBhv/
1Q5JqWNUKfNclWh0yYW155IYHGFY8/nfUPzA1ztVhcYGFKWTsbMgXi1Gc0DR2fjc
MK3FY05T+PBNmbyAFmxa+eEmftBBJu9WHl2L2TTiToYN0ey6o6b15ytrusx9wPh8
qmTn+SK9Nr1HBhiyK53mVU0gbsbBr8EKgw3KtHRunUUy2ZSFD6+Yy8dr+QENb4kg
OEZjcj+KEUhJ6BVND3s/9DKZWPRAtiK6iZVmLbqj9cBMGzRExBM+gYG6P2D1AINs
fYam/uG6uEehzGdfQek0DevX/SysK6dzBpfx7nHUEcOfmGQlBaN5cLov9WTNggq0
reQBrH3n/P3bTR6hQXAOputcweiQeRyVz9YSCXtaFch6x+wBqdPjECucq+Ij2tmo
TS2lvSY3fG0Hb7gJ4lA+uwpYp6GpkI0iOTVB2Rs8j3YDCFNz1F3uLuHoz2Ydjhn+
aheafaF9uhXlZ0KiVcsOJjkdaOxXjfHHKdsgcH2IEa6BiHrWsX1BqNryZ3SpZSVc
RA94H4nXKvRtROCFfoQvJQHBsCVK3dNN0uCycu5s52sxrG2cHI25ttD6cU8V+Ikk
LWDhWI0xPlzLgEFoN5A3n8sqNZXuFijPlYIazjVjcBeKH2MpyV2aETg1XLsUT1we
XB9ntcf+lkqdZct0I0tyNxwGX4bO8B4miWeFivH+0N1OOLdtn1YLyDp0H2eQ1TwU
oT8PVz6RmkgnjNxmYWVX1Jd1zuQ5ngUeQkAir/qRTcLnJdy5txgfArXDp/aYgZ+9
RXPlXJcJESelxUABBfwbN3/yijdSs1nwmMsRObNW+Do+dQYkkyQ/000Paayyra5h
btgpzT5T1FMxsFvrUVYVr1sDj35pGuyS1QOSujbQFOIu6a7LTAajAX3oCMkmatM1
58x46LngqsDRabaGTSTVINhNwK3krbCTAOk+hvTke8Nep2waXn7bZqyEB/oikbrz
1NQ2bFqBtRneBAQxdk7Pe0VXqdopkgaLjh2rLdu6nAeUypoc0lnSlXCoG9ohHbpg
AcwYgyCaPg0yJ+JWndPn5ge3nOK9SUFN5bkJdUfaB1EFJbR++ZS1MXwL/dE/NehY
zwqhPokDzFQCye+FbqAzy7qcQ3a97p77y2rlzCFt1gTmKupIZEv4kjRLkWg0EIV/
NYl7ZTNGgRxDqdo/3RmPnilUw42B5X3kOERAgeV+4xoeX3Nh3n1dQuTHjvfCbPPJ
5iqOYxdgN5JJmzDnfajb2H7eBrdBaw6s+Zq26FbGwQbdNtn8qdNgYFKjtH3UVVrJ
qbh+o+XVPj05YXEcaUcgEVAHYIAmNYRqVt/vubt0kjEHZsqBlMXvqxAM1F92up3g
wzA/6Z0KbZaIkPcF8cO8yT/ox7AJLmy6uKZgRRxRhaHFA7SZrKCgOK1GU16LJx1N
hRlfIyQg0bmsoQjHFw2s0YkEv+vlm3ZT/jYR7g3hkaseOn/LhDOxA/PUW4Pclp9K
aI+r6I1vfC8VTD1MiT5Tw/At///wYv1Chm/Dj5ht5IFTVAlWWAZ9f0pPNuUTcaB+
FJPH+21pB2+1k1aQEP9F7GBfUGLeEdvmIiq23Agnw32M0cZRHkHoMwMFVrWVw2kD
obZZDy5BC/fMuu750AP9F1wwkydo2dFkLejam9gzQljOYV5uvuqVlSUxgVQ/FucJ
Z9przBh0htHBnF4lBSxcokmYUAUHc0364VHL9QqaN43cjugp0DixUoyXaUdJtHUq
eAKN7HXmNi+g1FMO+Njkh7XDwfB/xhBjxRUxvlj6dnBsY7UkQH5itsU/UYzaG0rj
PtMajoExr8OAe1XGp/PDcpFC4x8P7GNpmXnhn7H+OTQJ+UaWPTW7y6yoCy3o0QEa
QLw5IiNJ3NADDErBtTp8yJ8T6X0xvraPnuRRiz9bIbckU8k5H0LhtBE2ktqcx9jz
F89+CrWouxZekfLiNplwmh7hqRFej6NL++Ale8wGSJy4Nyga8Q9Ts9n2kQImbkQa
LNLS0AdC2onBhBoFf5dlgtD+KH2DYbc1grlsO+CHI91ThQqoj3v4K4nM+TgLceYP
T76yMHpj8y3WY6f4vhk0PxIeP2hG79V9uabR7QxeHvafHOsTVYSOpDi5bADpLSZo
5KBnyHjknnJL+bANjDfXpIue0muhJIv3+9ZLivAdYFxg9+S7aU8ysiHwKCTzkZ66
mpqxMXFxnc+NsiPXtaEvW7hg0CHrXZeChHC42QC/eQLPP5DU3cnLhEd0z8CCVqog
SW3RJQsIzsJe5BZ/tWqovDkSt70l4nN4+AijECqfAMrJiTFGwU2gRYLwOXYyTg4t
q2ji0Pp4Lpox33hdPpHizowiBVcIvduPx6iu1FoHhIzRPjAB+mq1wSRkHpLhCQkh
4m0jUpe6IIbcAOqwpPkrtJlkb/ibI3yQpOoHjTe7GTqYs/h1JQswRq3vE0gvmfpt
h2Gm0fOJjLwTdm2HrXmq5u2+zd6WzweULY29tUqXIOTy8c8hAPm87lIs+MIAmYnh
NR1CYVXOIdVEhB6GeQIQahGxXXa4RlqqjQsodWpSF1e4C7MEWpLhxvxF1LrWKTDg
yd+Xd/Le19ug5XVwLajZGLMAfVpUViXu2M04uGYGZd0m4hdD0J2SUpjSsTDpoWip
qWETIGXoJgXp2tasWm036H2KA+pQHtuPrM3HlDRaxG88Eo4eDBPQL7zew7mGCY/8
grsB0xBDBLYLZHUQx8X2Z6SClxztN85dunO1Bp7RFF0zw2BiChFsRnivdSy8owwP
jixBbIuILC0b9+UJtpyEuuQaRLbT0Z+Lh+OzNUn/fzws0i7X7qNtqZRzBdP0pZiJ
qCBRz56HoMsB6zR6dbrS21qqXNspNiG0cUR7bjRNsjZgsE9zazLGrYJ4pstpqBgh
lAjcyymT4egm9qrh8jTOKi6Pi4GnSPuf5QgJSFx+qQmMxMtQmB3ysMTo/96kJrEo
QFdaAth/TCsmKyDKtpr6uPS9AHba7hDvUFPtOyqkXgP9nUggas9R438t9MR/jagm
rzmKdXEMI5yIrmBXgRv8AOHSgySmuLQwj5Wk5jngrEH1atWlNRyti45VVunDlaiJ
l7OJE+09r3nASGqpdfgh3R+pSe8Mhpypp5BDdhmGGSv7lEojMUz2N78UYark3op3
OOOCQIzJhohKI2KLmMDkJC1fqPEa71bW1ixLWtwKm60bbhJ0OaARJoPMAAFX1Ru3
bBzENvxjlUvxLXkuHymZ8X8fDZIGFaTGlKw0VHxFpRWiefAo3MbUoF+nvIVvchJe
+7ORrLxh5UE2QoedQBFDFhhoLuYcW6o3KMcywBMKMk/t1gLyKGZhjPb2Y/PL1CXk
E1UuVdCx21D0Dj+K/P8LiB6lTxFWzKcaKHAhF6qoyMnrjLKpBW0lgrJQHIMChyqv
olANNBXIqlXOlP0OoTzy1I038EtoYk7hm41q7qIy6mjl8aBY54wo7p6CW5kQSGOg
gXoadP3EMapVXP8kajb1uj3x3iBYsjTQAJoD6B10mYpIVRpLWFKkTNCExJkXYtT7
BDfpLsseto54Ic5+6x5HkvZF/C+dNjIKHDieKZ7xNvBLOtdeYZd9iQSvS0INwkMv
p3tyaIGPV5mizC7mR8eDoJSHqcYcK8ZoyrPNQubwFsg85J/mQfTkGk75COF/hSYm
vJs7RPLzfKge5qOP46hAf0nClHwyd8YbWtVqbqjCG44InPwv4HTL/ltbYVcB20tG
j0f2d9FZcv8Va9GJCCWA0aQqyYZxoLrO5AIbRbjP4rpOu8iz//SPhDAvP8dVXSSe
1ix14zshDCBiiZRIcIM6vo+wleKPiUxcegKSCtUe0GqeEwuaCqo1B0uR3BpyZ49J
J7tEr7BqptOLF+uL4hopsstxaWp/9UlWpc3GjXvQUCIEMipSXj5FiU9gu9YIFtIZ
KvPt09md7GWkdTzVU25T2sypK+oq+wzOGr5z2h/JEHNP3waVOVZWPgUcy4aZ2hut
3hlWwZt5zstBqI1Qs9to9BdssR1Ni6VqI4/x4hYVHUQIGlXxl9jvX+cwgRTBSpUf
J5yNvxFhuBcNp5cS7o2YVRKJD7G7fT8oSQ5kuFnH4vvMnrR3b4VTYVC9JKsjGUUB
GtZkQ3nVRnXeTwNd67rC0C2bakbsiPx6hcfrmLQYpe5SKAiA0C38jcjxnwhWzTvC
thlvd4JDP/EM8k9fLjCszz9xb8/hm7U1kwk095DYfgOJuNOikjR3Ojol1ss8iZee
Ty/fAxzAnPHsIRKIXvPKFlQc4julnDPlAtL/kGMPBDX5rxf2LOWSbFjistoBhngP
vSRHh61SIhVYr7GLztpHlQOjRrRwLu1bpGchWwtIXVt0wH7u7hwtsErHAufCXEHv
Q6n862O3XR6GInC4Jq+5T1gZs4i3JjIh40eSvg7HPV025r9PCIgK85vZuDTKp7Z0
OvIwuAadoTfr3yfmWQVJz1Q3WVXtvF/PeUMxNEHPhSf0J/ApqbsmGBVZBv9FIZOs
cwbcjiPfoteFWc8yOFnN6oTNU2BxJ+8c6+iZpdkxaJ+FARYbk1966/wZY06WPG4U
bidrB2cMKBypiDB3zTQfmqdfpZaANJMvNbcDCJrXgVlofPX+BCKTLHOsA/CxbbTF
IaOU0U4hIVtm50yDjpLFRTB+R9oCwpPscH4x395DskKtw9janz3WEM+Zplvr9Cky
bvp5cC8l0Yx9fn55bC21ghpndSumXHb9DOwROJO+QWlLklcHo52+7CO6izz839GY
zxoaIRVLC+T3bT74RSaP4NqwOm7QnT8uUwXOOduEs/yvpkKIMRwL71Tropzncdh0
pOh0eozi5sLFakFat7TMbVgmGhn9rOfULv6mWB5a2NoFanaM/QyBf3/BPuZF+M6U
+81vGll+JxeUpzkonitq/LIHC5e8o4CwlexZlJuNEZqEhKywx/znr0h6oyTKSjdH
aP+ruoNOX4Xe18EMljEhfIcoSde5TIPFH67+iatjfviqfOte6wr8RjSliKUTT+4+
hQ25bWkmKyV60RXC848EerkwdQ3petygLCu2Kl2Zp6j6CLn5AKu+zbdGzujq0/A7
jna//NqEEBmy7j3/8KvZodYRD5xt7rRIUEihoAOI8DJng8Geef5yxEYgS8HyPt4l
yCxzbm1hit37K0teRHvaSJAaTsddfpD1MrmSsv1Qv0tpfSG1IX9INKA1A1jRyEdJ
vTsPqF5m4pFX0jedqSId34Dx2VS3qWoxNRTCdvUxpq4SntofNANbva123rGdK5Nf
e4MMSHmOg3uaEjwVi4IsJwNxJsWFgXQB1ELnkBsDrAzwbA3Xdf8D6V8dm54s7z/c
36/P2SKcowVx+d/LO15iMfLhGQncgMbSVt532m9dJqSgFm4CbrvyROKTGGX2n/pB
8SPPAHlXXx2D6i3mzAXsirE7wopU78uH3pizNQjwN9E6/wENQtESsQZo/YdsO0C+
AsoGCBdBo/og6DdLAgzrBPEfqRgLJT5FLxTnCJR6FfjObruyAq1sjj894gjk0xgJ
3X75FQSqXisLuxDKrVQICOR003MR6fHljbilqDB07HNXbuOin9ch9SvAukiWJxrG
uaeGohSiXbuBAkhxCngD3Yn0QeSyjDDBmv0TeJbOp4AJKzG5MhmdEasAYO8Peidi
52DOut8MH0W634AkDZAy3RuSeWPK9MvIeGwOjtblNQ6fhx0Sl4PvmntJBVKTUKZ8
7ZnGFDPrhADt4vO31PCMG2bB/ZtzDLp0+Rk5wExBJ1QKpZSOEptvi/s1ut9K3glP
7LI6GjaHHfexcGYgJtKnILi/GjLyBBFSnwlqoDVumBB2rWXZhjH9cEwSkkWJFkx8
j0HHK6/m8ZstJvXLpG69a1wbPWPahQaloREKPjixyCrEQ/s9MtVP+Lyd3Xxwnce5
RburDp6TVOPHYXbqf+SJfErINo9ZZFpM0oD93F5Oa8d3uMejeGABrxR5THg/IrSf
QOABbTizBv7SgQcGRk4faKXBOC+ub6Qhukf+SebT+nGSXJ8asA05AsJeFTzRu3bd
OEbcA2CrkaP/AWcvborp9Ub3kPe5X/uFIflR+d5f8pNPIOXY/6gW8LNcFG3ETk/Q
qgHcThZNxD55TnhLScMHr++U4jRj1XxsHp7tE7oETulgIWrs4SAn5c9Mfpb53aYM
LHu5CpQQN5yFa23OP483+LF1G/wAXFpBfwKsTgdkHXtKIICfpiIPC5m+jdUO5Nv7
RZYkR97dDJIWH/hluG30ROutqU6T0KlPvjj/qYmMQe0ibn4woaZCV5NCE7MRDH2A
AfNVJrF040o3Ns2PaGNcuWvOE0+vSfczR/XIp+qMl158aKdPaqyL/PZOlZoaOJ+p
ESVKNh1536IupEC92ulevXPjt4/1erCWXWVMObed6rdbyUQ4VOukS/bQJ0lwxERo
LQ06ufJMHDYJZ46bmzM3ZCpRL+DgCRTq/T7GmnGunSoFZ6Bk2X43umNOZ+WorPBn
CSCj0B5oTadWUPkLNnai3urf5BpPEU1ejYiEWpQLZg8Sz8wWpG1OBaZP7iGLHmLa
6qWRZ/lc02i/Lzh7AavXdCyXn7DpdgowTbD4t9laXoMGE6UKdNy0KnVjI9H2wE2L
m363Eq0+ivcnbyjRAKNAbegrnz8krZ+Dn/l7WW3JTjF62sDjCIId420JnOm4Pj9o
srExFMOv0xV33080uDZT+2E7NAWYIzBeS9Le8kRUrx6TEeHghnBZqrWJblCyDEHf
WR4vuJdKCvSz7M3S7t0Cfr2U7lBz01SStjucr0aYHS4FklVdfYVpMhheNMXhLRdp
8EdAvDVS71uNbW1BedS6FrGmo1ESHNsvwXjy0FVPIz+FR3rh8EPPVvxOly99F5HD
/l0xeXnldx4qgQYYwD5VR+FpvAbMGILFlOy5yiMWhnyaN9Rf+9qebiwp1rvPtzOa
P8Hq3D0Q8HWugL0KSwj0Mpre+oTY1d/H7uA/1kyhzBqTgGX7V9bKXAuL8zAlr/IA
pV2r4VvPvrrJBfuiBU2F+bVk3AebEwZKOoO4rD07FCG8bQ7DbgK1sPGV+lLTPbOF
rPKpVOZFn3KCiSSXz1DFygUc4fMtVBstXIMMRX6iJ6dDx4DvOyndv5VFQDxiOXsp
PE7v+T3IRZKmGcj/ZPvRjXU8XrZIbqQvoGEV7JL+kqVozcaRbMWM5HaRsDedmd9P
lWN1AeuX+JZClAL6P+TBd/U9NHwDcAmwyPWbUANbd5la9/v4V8IMOXcZxbAsWUEE
3CG/bVEHCsjl3xChRRLMzjuZE2ZRCVcVKMDillkJc4MIVHbMv4VK+lBT7JGRrkmt
mPhBDL9al9KrhQEtEXnsKzYJjxnNRm7jQRulSpEVeR7luL3Hluu0/YuHQUeRBYH2
PDPuHvKlZaoA3wtQ46+uFNiPUXZefFdazlUj0PRoqlLb7XM0IDfRhwqVpxlwc09S
wvY5Q3tgbAeH0REPh6rqzEqNyW4DbFRMkr2JO0vhAx1Xw+EhpQ7TcTb11sQqg3vJ
mRyovX295AO8lrUWe/7bHbrVCPs89Mos/nSRTaSFcYJsvBnSzplrRx/4rMMpQZge
Sw297JxQHOc2naj7u3Kx+27dIU6H4AjE39ztDLRXfrV3yRnwJWCZySg18ExTgN/e
u7arUETad2ojCC9cbKljBfLkphiaINWSQFMPajVhGPrusSUNdu3IHFoAeZJGX0co
+uocF3gBSBGHMmDzXqF/gfv0oBUhEmxed58kZoJvV9XV6BdrVpel89T1qNCy5VRV
1+wZ4cwiUhxZR1P1RTqVvMbiKmPapF5v/uX09Nec+JvFunsV+ktNvMLhsQ1RFvsJ
lMPoTvBNskTVGX7RuUv6haVnbfMXMfbQLHt+UW6sxZqhUqAAy4ySqMpnVzM7x3h3
0ovO7KDsq1PW/+SCkxHGt7x7yzfNhckuIlH01uqBe7wnOblBckEXA1PI3oatEm74
wKASOq2s5sO7g41gEw1NKBkIQwAmARQYM5Cz+/fSTjUe8z9SEBi90gIzMEeMhcYI
nzlY4+Wp9qPbpXEqgoeC6KABQZ/9hBuKxEkqBuIeJYPhGI9b4LRJqgOcE3gMu5hF
sfGepGb8+FZenxd1blueomyJG2e+S3i0LgpvEn+Bg3Kqwn0NJAPj9UPLpJjV8gXQ
hQ2qtGUOEGg3WQTvwRYypJ50ZbmKZNB9DQymT73ZfOmWjvJnhVXYP7lOQxni9zKD
4Yy7eKm71n9yp4SC7HgadX5gcBhogobUMKrwjexxMMzLaxvi/7uN+5HmUeDHEn42
xhTFeO6h9N6mZ0lfCiNXqRY5yimyYM/hRsZNsP7nClCcbcB/eAA4XIN4t21vfSAf
sWCg1nRQJLLYgiFHxNl/dQSl4uPElxwyPCDZ3pIRztWdNeV5R7hDV6rqnsFXZC8j
nDC2bzrnU/5ZXOSkiiIoAgAGrVqgT8e3eE6F34scQNRHb5XASt21l6ebbo3CXyaQ
XB7io+haTmvNYhgocLMYa6T2CM64zNkbBr/QSO8Y06UJ0FLbyDuIamcN/GJ4ydgo
K+tD17hTjU9xs3+xnfrT8EP5ce7kEaiF61CQfBxdUngWmcMx1okIHLdnzZo9J4hk
L3gc/yvmAu0HzSd9nlScCAFTGaZUN5pNBFhZ3qrPDE3PA8LfK8V9JnVQUaPVW65t
9FMYnHUGIoHLk8oEAm1ve3RtM1IEK69sqf8Vc+2wQ6qloSU4Z+YoDcxuGCquESi8
AFsa3uJ8BWwHuLTNe5yQ1DY3cCwmm/JGP/wNNQjB9HXbP8o2NKChgFDS0dY6o6+f
yi9ZTZeZUL0bWsih60pwnjUv26ffem+82oq6l4LfkyjWVS6w47znDbjJxqXDcIb8
NUeU37+0N1PhbYezVhJ60fLM7UgV+Yg4e0qONW9ojxeMDraS9QvbcplAV18MCtm6
YszNywk2R0pRIQjG7hjza3DKBLxYXjBeBRXjk4jkiCdV3NtRxr/2K2p9UrhmYLa4
cv9SJI23Saz+ejETQw8GaAoFtJz1u3AfvP30gbIbA1RL4WDKItd22po0IM8Djq1i
jzlHL6XcjHk5UeOYMCGsqdtegWnapmI3mTOR7W8k1h102/MEda3mlXU6xiJo6aRo
rHSgPl6DHKX7L/ZlB7pjNkTCEn3oRDUsI4BY/NAkCQTKzmt9f5Mi16yqdH1VboPq
BCHJCnwuzRt1l3Sz1DIP+axy5pnnEfuYTfKFQdu/dPlGz7MhVx+rUsirvZGlIpKV
XjmMGrf7gpqGq4gDWTzL/yVjeo6U4Mn4ssRLcLoCyVhSGcas90XfOrI5S65InpNr
YPmRloUeAsIg4+rPjlAtL+NiQdPcxdEFrbgIb06VZS8Zfr8wBItPgejtvriP3+my
aoSDGhj+BUSFq+WPh1L8dioPeo6uAOzvIQ5D34NqTHmQs07sBxsze4mNGYCl2pRy
o0T8unYYv6iSwr4FS5msWn8uCvTr/q0pNOUC92FoSycQMAOs4KJwryIyRLxLbAge
+KxMyvfy24DX8lkvVFkRczKk+XLHNHqFmUTMKzV93kpBE5MFySPbuue12brb6D5R
+OpRFkHOijkyaNqNXRosgHd1AUsP4a5g/VUETm402Uvgcu1SqDCfbEHval3ViV6q
OVBP1VQeD7UuTi95A40U2G8CCPRXo7Lo6puCUE3ouVjs4wEaErzlRUkfyDRwVp5p
ALk/1ARQyUgJpR9KeAlYyHKnSI22Is9/VTrVaqKXbGgmUl4FiqToCCjCoQjwCiAr
EiYJckOaR9wrcfhFs5QMSVOaCqfnTIi3/IkNrFYQWDYAVTb/ynGWJtPktace4uME
FZPEj5kkOfbiJtKna/Niz6HzUfV0MyePw8UKWj1Hwzl2Qh+d2SgYwyFZFdJ/sp+N
kUUTcGDVxu88Vu8w7ZqxiC4g6iQte6Zseg5SVY8jOUGgth2IVUpeERLo26iT9Q7L
WG6FiXvQcr9agH14iZUpYnDRpneWrXNPm6KSv5P6OgsKFzVjI/qdxxQFciu3e4z7
Wk+quRSlQEJoEC3HqHtuGi/Z+pE3QoYrQkOf2vsJDzM8XMvD84jzg/hQMOtGYFML
vBD/5TqSVJppWh+u7WkjOTfzKVoovaWK9g6LMQbGtfawOo/85s6VF6PqMh7mfQEt
YRD1rM6vGh2hV3n7RWg0gYv3RPt15D/dmKKzmEGHq02/mRGqIPmPY7kupkpqYFU8
TBdbTn31oSynO21xCGC1dS6fOn4SSlmpJTHQlqmfaGf1+/U7O8Sbs6kKiO6COP4Z
RQw6gl63AuO731x1sG0jX+V6CrmvO2U3vaL6xG/JYYorwiM9gST+Ti+KXxf5hcDm
2rMUDjsYs2F0pk7Wm1znGlaIbBYxiJdxix94KvOY+tfUDpyUJgbWRw1JVM2Y0ElV
5mUKYf+3CxT2p8/YqdOX43eV9y4uzeKEDgiaBkyZ/Vqa3JuXKbYpfQyNsQz2Y29w
oMIauEYpyvT9gIXmNTvqQoEWfpafOcbuDoXG6FX8gL2JajTOfqJLcqjiH9+qgqrt
B+eFD8sppJMhoVkvSU/EtnJFqZH7rzh4+ewyoSm5YEt5QJZgx1V3hHMbckkcLHUa
nqitlaKI31v29zs+f6l/cZfvm+EGlL5UwgoDFnxtdkxT02Kr9a6NlmUzhxZ617G5
+Sp5OWKI5KUU5wLoLv9ydSOoWzc2im0GI58YSVen1B6cFPvIqmLUQ9N+mNh2/xG9
3UeMGZ8zdcLTfLpEKjLo7YFPrHZjp5qbjhVLpQM5+pbQp8QJjfIB/Tje/usdOjpS
00R+DgoflK2chCTONH3vNE4lN2CczF2sful9Gjqoi5aaJV2azQgwzsDrL/oxX0cJ
7XBXRs/4sS9qiNsDeNg13LxfVP7kWBXou3HMIuSbhtQ3UWRmwweXHx3iMquaWvjs
psmWqgilIw++x7GMbo2kXeoCD7CmKbd0a9fAZqXlo7kItTUAZh4PfQDdtH3KdoFP
3M6O33kJ4zQ7kyBgMgTCdtoH0MY4GXTzCnf4ij66BrXVHdYlXfBqm6JiY+bxzO4Z
SbmoUPBuFNoYKqD1A/ogN/mBoy7VTVNL5w2Kxn7hgI9mr39bd9t/QJTzoXY1rar0
vNUBR2uNbM5YND4ihbBH6rsvuEzq5aNqd4PfBKFSNeSWBtULbQJcm4jUQ/I6IaDd
sxUipklBEle6VS841QerkOtsEvQnBqytTgwrNFETMa0SPqTMFWWnn62c2Qc3PHz5
UQFgshNUkBiAIIAs1XjhjKJWtr8RTZ2y6GJihNcRp1DYDtGzKfTfmFkjv6trMuah
auhSXZI3c0RfZu8MhDNM2brvzqxiHdIGedqfqGgQQabrKdyGNwJ4BKrHfnatrIjA
uLwfIzqS66ARVdelcAHqu40A84CnJ3IYPMkwUGSC8RCdzkyefTGmVzuVhU1cBofn
XldhluTSJUPBkBh56SjkoUVLH+e7Ud50AwlSwbMNjJibaLR1/BREwv3WI8oO2eTa
v4El5G8XoQUi9w9frIiCl8qnV+fuJPaxzOB3IHUqZbTrXyVtkvfgIeBzkT9+jIYo
59oU9pcyZRkO/3skdRHCf5vIo4A7L5qpss88k4YT4oDHdOZKPRkq+Eaos2nD4Ioz
C4aVRJZaMyvPtU85b8fvV/7uzWXbG3tpdAupIVuI3wtWrxlNKWLkyGKGKJHCBNEs
c9MJkHs6OVVN4EZ+0Spjg4Jv44zxqfjfeGIh89i3f75pKitMkNjdF7rC05yLhLSL
dmcUdMVopRzIgRLup6G+7ZrsjLRWqk2VIY8eIfCKOibeoY4dY/ZVkCGNJPnGQX6j
R6+AxUc4PFnJ1foMwbsPH1ca6cDXL29uCjVhZ46EHMHeQL9cqn3l0+WjMgdONGrD
s/0rGHDvvcZdLXfHmNktZtr6QutbSUnt4dbRAkN12e7/azEnsFC40E69SSXc1a0g
DdOlv7ad8VgJYKK5PToKZvNNED6d9WvYPdsztLHxDil8eiyUZg8omXYJBwmvAo8B
PTrtuNG48ydqvO7FnakAaMLWM3Ot67OHXuIVtkET5CVjkghmY9llK9HZ7v3VzDaU
+U5p3qmeG9QvG1ZUcRfT9wCKlT4vYLfn6bQW6vY2qKt5IPwfEcL7mtynITXAxemB
lx8pTuN+idun2V1iA37Mi8vu8FJ5pc8Mt79s6U9+L1vMP8RkYJP51DU0VufZKZX6
Pe6R0NW145MUwuFZsPPRdnjLgTX0TToKSlCR8Kxhx8w6+fMg3yzj+T2fJkTXoVIX
Fp+yY5C7gphIpOfalpMUAe47sM+HWZraSOjwUAe2STZ5MYetc6i6VaOP+ez3nRgE
aNLldcHMDPdwSeMTKKyhxPQdMkpBOpN9HDWqjeTa+0vsA6eddobCuO/kjD4ArFw+
fBVr/opGMEi96iwFzeBK2zVeVL+53L+zi0Oeuuiy5Uy8Jb8WK9HXR7XeJR27D0WY
35qWn0vPtKkxA+ovkGnR0MMJw/0+rEc+goLYdzEEEUsKNCJELp9vgeGM1nNFBFH9
zUphBfmPGxNAS4ocC8rPGmbQIWElEegi3p4fqDzaMqqdOD7YIc6L1VbWKtdzTbMh
JMcDLrUW6B+LRc52HhL1d+yOxnGxaC84Tju9BhL2xpOxgDn3d5E4v1vCbdDVsAoX
BjYKM7oar53k6PfA6fUoDctwduEF+FdMn8H18mw5UUxBTDlWQ/VScCHYxhsqN4Yy
PmXwVdBJViVsxtyOG/QGHq3TLB5+UARjkdekSSyKZ9skEglXpcrGtKuqxM455erO
SevPHl+6ZpWjWgrBiNdKJ4LIKcRHfWHNegJsBwR1iy77UVGb0M5I3NVxltIRMxQQ
Xu9S6MJrb9NkzGJJtvRxzOBWfoGPPZ6AdDS09iFUUXdJhi/6zyolf5FCayiYqsUP
JYAhVSqTERKWFvlyyr/FaUymE/h0H6Fmf7V5J/891w3OHSeRxpHqQ9QJmURRbxWm
WpZ/Tir/M0ZmPBqYqWIersg20Rs/06TVz9qPGOATkkk8yBK2FOrXpTBgTCyVHhVM
aIVdJ0uPWOA9Iv2zpXeEuXBHQKeA4Gb/iJ3FSEm2IeFSAujuA/l1wQ0u4+mI73kc
2FWScV3l6fbTEWBHDTbzdDdaKyEniwQQ6a+o+GBuuOwQqnKB3tpy3NK9JuG2WASK
0LLqt2DEgoKgiRhizP8UyVn3XWnC+Lu+UiXRLBq2WlTc2VNWVOs+PqjUbR2ABOLg
8LRj9qu4uTaTqo8AQGVg28+qsauyQVODRI3vfGlGVBnxVr0fA9dUOSMkmMoi0DCQ
5ysKE3nw4vhJsJiG+qTJJ3KGeIvv2fHrTVMtkPHdc+bt0qlQlJtK1VtCf8AUCKJy
eaCQ11uGvCGzOVZccWZ0cdEbh5rueimhwmArhEyLy8eDCdqhzB1YH2XB0qWYcPpI
FUPwPzteDurhj4ljurrCBnR7MTVZ8qsVGm5csK5SVrA0TFhzQGdsxgHPr/dJVcIU
XJC287RLuSoW/wV5wZOKg3keqQ7FFML8tz9xIyCZfZVUzxRzOTP2juEZTSOY4LBK
ss29AZ17IcWmiaXbLA0wwxLiGt1UUeAhfk90NI2KOQlqX3UQkY6Qxo2OxM76X6Ux
XjRYEoE1EBDYV6fbUYkYTXOgUlttofYWZgxOkaFRr2VB+1vS9v+3GYcS897xe8t0
8HYA9oixtlFXxkpVLvnrWlgRL6QOClUIaNtyRmxvYcgj2nxZV0zAyXKO9MsgBFuH
foeYWXO3g6pSxO5dpqEDWXTtZq7IylCRhmWuP+Apa7BANm72S9VgBCgTadYquSmH
wPY1vr2GrPb2sdLtvdTybEhdqNHe9V5iCre3SiKOGWgsPATvLwZx+Wm60fl86WVa
x02Pk73pzV2MbcDbh0WEVhFsu18DImPIebU4GbtuohVqdy1/gzaoicAH3w3g0seX
FK8MLZmm2MGgvrRxAFjnf1TPmMKtKwxwa20lC5dJ4h/jQrFMPd2yjmBU/ami+fs7
MnDtA00WGIter16rZmEe3yKyNL+jIOdGw/fzsDhCfqIXDGNMWRx5dQU67Ugly6M9
1RsTd5+JbAlzcjVGtvbOUogNmvVO4S37Z4+QiIakQgUD27nbu69wfEaJcQzckJnP
Cl1mwFfPELlXrGSBcn/+7zFnfFsQoOXA5O2fKfRMFUgzm70mYffCw+b28uc1m8cS
ZyBfW+cr/6vimiSWPony77/WnQlu0DOv59M0Ko8dqjZuElX8xqznjl0+TD/9It2r
kxaYnAaAP8NfDg4xKm3sgDcyVvrRC/o7XOLtjjq55bS1+KfBQ06aPEYAO2Mf2aWp
9Oq3UjJtchB0/SmE5ehUGtn0SObgvQpk3NfjD4JeypuOg4xli+fgXcQIShsCVkHb
rXvciDUKVGcd5idEZQ6pLdHUL/2uAKoPElS9MmKnwpRUbiIOmK9hl8jOGgqI/8aW
AqEjw4bqO+QwECdZIgpkkn+RdB4cUyXsfxmCKVnL77jAZLzHjVfGXPiO0IiyczXE
Dm2AqgRnQYcAlfB/c5+4Mi8fC1KuMxq4xijIzeEybiJL4HRVpGB/yU8Vx8RGPuLm
o5vJioXCsJH/7IsmTQVsAssciUSrKuwlhxWY6TmudCmV6gH8K2ZQlO9QnjH/hLp8
E7N2faAfdwRh/ZFJBuiY36vaPkb82CZVAzCaMtYR+2lJAKsrnUYkhJ8dC9+xgpEV
YbT4QpeKK5KheThoy9/vklBzUOJMm3lO3RVd8ouK3hdSpAVgShq38lfIJdPcm4sO
pf09Zzfi2FTtWAF/Cd50k9RmJk0uIWSlnjuerio2rE3y6T0x3ang62yLp+uUS2+/
+Eb7aQJO3UbrwjWegR6yMFF+1CSUafLHr+baylSdPanGxLb2emng9Wpf/9pYQGxV
7fgfbYK83t2LWVdinHHjtuwfeQPWxH2SyFDlRS3ctp/8ezSBI/o5WCw/A2LLO6Vq
pf+oK7PX6lDrvrs925cXue0faBp63x+HfaECjs8gu5CMK/MOlqIXyFxBvcQbGGmX
ZQ80Z66hyTtXJ8AEShNu8v384yWi3nNHCo8zNbPPTa3J7ookcV02eiEE+I93ecc+
FiMcl1sDIuzFXInQOAs2ENNa93lfFngnL78gU06xF6XjMouP+f9Upr4y5CtDzmi3
lIGrjIua+rinrI7eRcZqTmxmbwm4e6V3j2bkeT9vveP+hxRSGDrtEFNJbTArJ3Mz
oUbx8BahlBgdl6GZHqhByW0RSLi3QnF7jy3762yxpag3qtBfVR9ve0/GFPBVjk8J
o4nonVx8IrsYPMFZ8X54EIDeVDu357qRa26wSDSlr/OGqiu+2zHD5P8wqnYhKt9a
5SKala65oFBQQG+afo+ArGUmb0DGZNZ+sY6TokMmN9D9LNOpkvwICBDHi/6kblhx
3abkfhy1TXs5wPBUelBidti6eWotiCJwFIrfFell3wTlGin40HGqQmTN0N9Vckx1
Sw+hxiXKQASCMM0KqshYW7KPkh5YbNpDVXkSKI6ZoFwIM0naamZ1NkSss52wRLe+
PPsmztUqQr/iRukIQZEBi00jKlKtQiO6I/nR4BczioCbPwyPOjMdzlrBzyoLIQjm
qtl8laE+uDxTca7SpRhK+i0b/iNkIrV3ecvZT3EoiLK9HoUfwyQNXzEydCtzrJBu
cVg2nxC3zECGZhRF7hU5UbkZxNJPr7MRXfhmHsFqgZaeW9ksH2xTnIcudvCXv5ao
BQJxAI4NSMvnn6utQo4jdCGBKi9vjq02faY3Z6k+dGQt8Kai+Q0Tu6dnn0D0Hx1F
TdF4QpoCqehn0xhrTY+94QFVBkTT1HnZxnfID/rVEyyYztb1aTOqY1KUwudDPC8c
IduEF2CwmfF7b9JqTt+nyUVzhVAqrBbkUtL4zAfRZfREjZu9mFCVO6K/earUILqe
C+aywKJVHdM91zTcRgTv5rubZHi/7slYvMe4wARiWB3do+/W7S1wlaf4usGIj8dz
6T4Sn0qxm0Fd4Dpk668B3mL9XCV+l4zk8pYTB8cfag+fsGk57ewGrlJ/J+2/QGE/
pEm6E0OgsAuNfq+RBO3zJIKB+XtrXHKJHvJXjmC5zVD2FtjvVNmqvCjHW9OWLZ2f
86xQnTwy8CzIKnv52TlpB0UH05Cn/6mzqPPd7Bqu0kEyNUj312ZLEMkB19MKxgrV
HpxAy0sXiwGNhhPWZ4Zamv3Hn+l0Pld6KwHodpu7DGQJGmiTzWMdsIejYeAye68Q
F120npgWRbqDf0CsjVV0rXp1I+EtrioTsYiQhneptCfOY2Hx5DlgH6LjhZVBnQbb
Te+8FUgK3qS9QJYqLspz3EWuUDrWMJR+EOv//FeXZ5P+3GyQBRuFp5usJ+fht4sc
/kdshdEd6nvdqUR9EihVKXroEzlm/muD0sgh6ckczGUDD+vpVY/XOrshQ2vss0ac
qU+E9Rqrw6yxJ8SrOvzVrkikKjXlRxhwcYM7G4SIsW3VmxvH2M8gQJWXRHh1tRcI
gDTypretZdG04fpICu3nvPAo1H74gZhm3/9e1736WZ4KorTmS4EujizLAYBdJoig
ULqwht8bEQIlYtfwa7upl4Apg3+W3EXQRhuSr6SDsiedqfYw4EW/wyA/n149oM1C
wonb8QwXqTcqj0iIrX99I03ES6sMhkie2zt4JpNjs3G9c/U8DI35MHh+Z/h71yVr
F7nGc7WfXg1tnfKN3dtxUhpcTD7CiX5SRBx5GCY/XEiFdniXXgkmWI0FjYSXUad5
EmFAZ2UVnyXX5NiD3wJYmuQNrOqtLE4/7nwNbVOgpft/vr1ayof4ZYwvcf62o7xw
CdUTcU+Rij6sz50w3HVyvGYLf5tHlmL0LQaFCXyLdxP9NNX9En5Yb/9rnzqUQOSd
YLhEXB62q3CpWeCgnK4QJF8FbmXhe/muQiKc2KRKq3bOjb3lIbAbMYmRNnsarspO
VIYhIVSwOj6cE+oeg2mKAXlSiMb1aG3CpijPJeC6yrUv5DEziAH0HZYhThzKAwRO
wpBgqFkgOGx69HisOcswwWkDK16WW31nvQfq3bOswtKmDb5dAgADrpJVYO5rDOTw
o88mcmxdpe0lsk44W+QHAUe0L5eFlkNaiOaJFsNT5v0cjD5qb2aZWEDG8GOOGjRz
Hv96Gw97V/0uKC/Bx9hatnmvKnTgLdLLmJsg+CbS4NreRHOdgFzxm35GPeQxYmep
/LN9ANNhVL/AQYHpUCwTh+0/0RONU5XfSQ2N0O+cst8avHLevozBQojRLIswhtXp
A0q0bfmnqh4dG9lHnRjnMUWeqOynpMeJTLyy4I9YAPnRlUAcZxF0p1D0BoA4+hkR
WK1c5hDZF4o7AKIWI4AWHtSCatoyIpIdSGUsFqyCDY6VaQan6Hi5i+gMMyyNDD/X
nJwt4a8oUB2e2ZkP/jnC85cChagon25/x1zZerR2L2lsPYFuPUmMsWXb5Rk/oQCC
hsnKysCiK5Wx+/ibaxLcfAbgmZZWjDrqr0wjdPH1C9U1vO8Ug7yhYnxikWKErI5r
dgQIoFiwCb8g39AHEkkNU8IgUVhaAowUSo2xYADTOP32jrD6Vma8i9A6nQplzxUU
kCsxmYwxG1kfsvtvHOeLUA0NoiDtPuCHiWjw8hwXm78k0GNX2XAR7DaPG0sxDKsJ
ZhhI+6vZ111rWHXVEpteT2NvFZeQmu9Jn2DUbYxfKCWbQ4AKDszIo8CoGubj4czj
duSF1Ixx553dq6GcRDdOb9CAusAVl0UJABm+knoijzN2iy+QZbay3Yc9GYqo/f2G
/xMTAAArU9RKWEgTLD4GV4Pdlfp6S5tofrSZbhS8YYAAe2R8ojqKGfW52oRzBLz8
XqkJPlisHcDepU2djbQ/iDwOIVMPqMoSgPYITfYzAY3I/ELSeEAI6YWbXgMgDlmF
C9dP+KHMN4aejW/xVgiNMkDESgAB4pOstnh57FfYNAjwTP0wRE923efyNattYk/F
Q4Y/YIrFWYJMIqPF7muuzEu8WlDFg59Ea4lQS2+BK33CWlkT/hSiLWcKSFls+v87
YNOUMMiy8h+w6pxlXtd17XemVUXoLbO5Qnc3uSQ7Bg+8fQx0jad+rJyrPcUZePAU
P8XNmyloCD1n1btSNO6yX2R+8tprttX19GMARn1JWQIYZoYat+R36wcBo28z++kL
YRqGIldxbgWVODiVqPjdgVhqDVrCIi+6IXxcN+0xAWeTLKlQuAb7E3tJGjE3PT4s
VLtDOonI1QhxM0bfexGgDhSJm7QUbeKhS7ki2TYuRysNbY9Y+pMaTmgS92+pcool
fCnFkKsCtIe8DkjRTRmL4DJE7vMp8A/UtHk2wIIwAg9pEs+TwO9tlGj6Lm3fZ6GS
siRcrUEEoQ3WEZvmKwM7rADLnKLNmotsVhe02fIEW2RsOyjdlCrBNKNNeRzPVl39
vdrXkgRH0IKxQOGbP+M3O6p60kx2wD8oeKOGCfVwBOTZnJWbRGz5noB16B5thrmA
qKWgTLEtEPDWRI21c5LzKy4Beq9Aju/oHEqdS4X2+NOOKjLLX9bzoZ75aTXWMuin
ERbH4D7Ncb1SPbeVI12PpKmvGfOwKWpivRNoeuEUc+rUKAJ8bcGdPuyzcnA32i2G
IEg0E2T2TzZWAzsYsxTvsGGUXA3Adfw4AM18XWOtEK8mNiGLGVyGKrlo+CpFZbJ3
G3ZONYo3UYb5iYln3dQFQJlFjXrVws2jJVVTfbv2A8Jej6yLAGqIj3x4DKz6wdRn
BoA8zdWjMKsdMvAXgQ8tulF8KP0YGiHQ07/PWUGoiQ3btDn/GG3JrRmlTw/bQdiP
oIpXC1AX3Z55rlban/+BsIBlf4vZFwuoC4tP4wxi7xbpl4xyTAnbBoF0gaeZ/6t3
Wu9r5C+Sma6SH2Y7KCb3nI898XjoJ5pjq8bwKnyCGtXX6zzQhcsTkLhtkRfwp/3z
o9+K4SfLAwLTSXLcmTbLZcnu5je4kqRKGR3dXX/5FIvkFmmnoV/Nv3GTJaXqaxqd
FSNfgiuz6D9SDid97Xv+s7wbVg4pk5m8fQM2l0fXXh9sAFodguyYmk89RlIKF9Fb
TAbAwafMtJw9gIHAN5p+Cl0cGcQ4hbP5rdIHLw79vUBA3pplU4UBxzNmaR12gKYh
FH8dWNtyn+aQwAM9CHSzhRnl6c/lARd7N4kaQ9bIywQpvQ0ume6R8Cr5ITtsoP9w
4CBUAkt7nKs0kuakMVQqxQpCHp2dXICSSul5g27Frnkz38NyYZ/f9gnKfVKTYbM1
TIZDT7Re4khmzbg5dKaltWAUSSK7+A9e09nyJqp5INZytTqv3wcoGyBC3NvswwiB
RCah2OC70nA0sxLVirJFcZtp1HC4BG4o2nfnDPFXf1plf+EIpi67xftWlPrYHSVG
EvLgmjpatpM584bXDuXEThMZ/eaBLmab7o5HSBVj9PSeMIvzU2qHPHBUR/VGnlCC
7JrezpKkCQcy62hVBKlF3xTLnOhhZ/Wdxjw30s4PsY0KEEs5XvHwzzxjvPw57a1s
1Y5l1NTymPT3xnliXbV5aGWMy5n2cK6+ag4uOLOKYKhhOwxFWw9U5ZLzudo0rWi7
UAWyXlNebVSQ6WX70/U4NM/Jl3tKUpX5UmY5Ycej/CqIL39liTOXV6dJzKquldD9
a0105yu3rskLRfT68u51rS3RelrS74+YbdELHaSH2Xb4bKDTQ0Il8/oD82djz5s4
8KU4qFPy2GkymiloArDhsbkHzxRjdN6oufNj9NBVOrEsCx5nUcqP25n/tVdajV2B
+gbnKSvV/gdnfIyfkCL9qlmYNChhz0+NAmUFRKvLA0/As/1+DOWt7uMKtrfQHWM5
D46uT9FTT3xIN6L0TBq7wtZEb2dfsk7y9DBQF3Rfqitt2V4oIcErX1IIlgiuNUxP
WOOyHye3JBj6q8axJBU+o7SX3chm3i/M1r4tVfjhv73cK4mlRwHaEwGFGppTwoE8
Qmh2cqm/vFkM0h90r7Lwc5kILjwbSnbDL9JNPcinCyBOFL8zagzmVne2r2mxv1Yb
chsgYO+R/OrCPJCQD8RcazjFNITPegAHMmXWpcnfgrfMgYVQ//UnTnVbUVi2VsPo
2J0pGdxVgNIlvZLFJNb1ZhXUdGJT9lfuZxMsJzvSXS8ctThyaxCHGoqTsPX1i52L
G1Q+MQiB+mPkTvLR9DLMn5VjBYcWAGuxhkwsVMZCBQETgLRmYvFS3hxbTW4jrMnE
1GsRgncpsl1yc7pKuJEawd9+g35iV0TpZT1k7y0sFr5FJqBsWPbvnJEljVzPALrT
oCvdc3d/zg2n1vMerzbGThFYKAp4W6pcZwamfluppN7YaIOP9bKGCDiaYMGbSbl6
h3HrAkm/kEpcGu+4EP9nGuc+KEo9hrbIxcoUPRm28ErQOA2/NGnQInWAHNV2LsOr
eouuqqca/WNpSLYlFZ4nv0VgxrP0DG6WJXnpFMe1CZgrGnQtwyUmOGE1tHR3U7N/
yFl4RBdQv3yJtmc1bKvGfR85G4hLvV77hKQ69QG+ECh4UmbifI4ZBNXzhD0lOr/W
BUrIm1Mlj6Zdj5/3RLhpl/QkyJfeLKLf0/ylQ4g9rJxUOZbOWwH+4ZWnnZ39Jj9C
JXoRrkM65AB2YfcFF2VjO5StCo17WZK5atw00MoWCnBePoXbGiDRS7C0wpUFehfs
cBBJoY4alerDYWO+PB8RtBLT9bDApmnZOVgpdaoqkoWGOxCahSEwHg8B+jMhvkLP
5t86JStBHRjh+FfGK3rPPvlGC1ZZbfYaBMfylT6kOxE3M8va2uKhAIwjVlVq+Mrj
jPSd3jAa3TvZOliUFxFjhW/XXFQlIDllf03hqFm0mX/hOS+lE/OFqyTR+Z3KSh4T
WkKuHH3oTdE59YNRMMqWek8xBzQtC4dPqQB9YtXptvq9EsiEttgGvKiR67rXR7/A
ybz5xerzR26G95hANdhVWW7b+6Q4mWLv88mOuRgm/iMFgdamnfID/GIS/n0mtv+/
GP2f7uJRJ4eqeX7RXWf1cWAOrCN9BR25iplMlSI3dYtgmv7eWSyx+xoIQQiO2RTz
kW4HuVYBKMnjWVCGC5DCsNHzq6qwxRZcICfCudoTcTRrpVF0iSi7teTckVDiUhdq
+SLAhqsH80AIM1W8Y4VaMvCvO2o629+MfdVXafdVq3HdAg9eQPh+AteWFhRQSrsV
SFtzdqDbbdHsJ7FieAobpwIhB9CvzhXqZeDJNTzCwiwPsjo4P2ATbvGgJ1tKuZLQ
fHhy8nAcvzcFoh5Er0yAbVvpkzy52s5tR27h4AHWP6BpgtIm9lrmG0WBVHiCroNJ
3o2WoxjVIJRhtAbzWFSrN7glAo8hI9ZWgzIvHCe64LbtXkn5Vd/VnwIVbDYbFtzo
KiFzJby96c0RydjdTkZyAQGdONcCXyjlL6IosuAAJtNbw85eLchyYkpyFYKwjcg8
db5O06uqnkiHrRlmkb8fYH9fplnEGdtMllHl/7TziJ6j+v4ynoqaf5O73HQaxtBk
055iPulDaaxqLKaQSTG1nXm0rTHX8LhQ9n5bsClDkh6XQLOAKPJ25PJR16t+bL/j
LqWhIawvehbkKj+UuttVP9Ri/CqtYZ2EBWXjEVsAnIdUJB8dT7tjJFVNIAmxefno
oUAEOQ+kR69CMKOzlUzrm0ChB268I+P5GCRL1GXqlKjWHzWxfC3X9pqJwjWe4Emw
EHAIBFC3pP/v2ydgcOlvQodv9YLlb3vY6KJHFlaMwc5RqhbfybmF2P0a9e3YdZWw
LG6lhTPCPgK/2SQZwLJPf7tr3iKsKnaX1IZ6xdmcymj42RD9DGRzUPB6v6C9tE4m
z0NUcB7maOGI4xwIA7cy5L8TTylMEwR7Z/xK4xWxmIMg2CtNrsTG4kRmTH6Zq0wG
xpCZPi0UriQdk1HJj7fATNTbYbsZsDQTblo2QiLAm5bamSkGOaUyji7pp+qXGck3
jYEhqjV6xr0hCvpeYnGRukNC19M1DL8rPUsKfzaFDzQU/GsTyUY6rwJVUqMKchN4
ssVHkcgjiCVXTgI7k7iV8GOXeY9CQ8ZUfGv1GBROxNHITmzV5bnpsSFcR6yOKADP
1Rq3EnnVWFvSvvVmEuRrTXQtT0xUd0/goxX6IlhHtCOkB8XRtFnOdaEgwF1+1tRx
OAP5nOmAmyTwQJ2PQli/HzlB2Y7YPADDb5v4n5BLGs1i8xcGP7kmHIDP550NisPP
K+Lg4bpeyccauXfCB9cXup6hkseCI9OO4DoiOUYWgLz4RcdQrVqIx1oPTBCWqrEY
up64s+Fgw3HSnA3b01LwT+Zdz+/ttQsvyJzHs3cEoPxuynyFoUI1OY+LRk06FdBu
dDCF6X9QYzjNhvLi5jSETJvig9Bhs91D3ygUZUUN3o4w+vzPnYMRtUq5QWYBormb
o0Zr3pacaDcro6t7zqb70DReUazu342jrYVWJpyxij5W0wNzYcFR5aosTpzJtnJQ
MUfQjaYXf/oC8rt5V+zLTBeoOZV0RO79kOio8Jft5iYGPju1QQ7L31J4RH86ocuQ
y9S13PtBWOKKGnhsVQzPTEBKAez3cZuZYAvIdJQa7KraXK6WBR8KQEPRKQGthHQj
GfjK2rNAsnuaq3A4WfLGHQDpgGyWQUzXkTsiDqc4MaBZod1Q8d0L2LbR0EGxEBun
4nHQfP08Q6v+lwSUtEAY56O/5Rf7j6fgwP0qOoPLMg/J/ur4A6Eb5CkMiqBm/If4
nwoEuArKS/8+QMeeER//nv7OGp8m+88XxXTsQI1JHENjDGUuZ5bUcX9AA2YahtQ9
8Z9OcCm7DhFyFUY5ckCo3TUPv9P1XCH0BBWwyVFxfRFt5ROvF+okEgHhat1w1mjD
Oa+QsAPP9Gm7ItJk0dO8vnODIunoL18v+fwxZb20/ak2YFxP/ivXg6Q/BUgfiu1D
d36ilRxuzHxUPPNNZE6MgDJIfJ9ddr3ZGrFfJUQO+5jF4eRv0X3bVfVi1p4eeU9s
k+za3zydI4iWvbrA5eztoFP4vKJGjhIl1jA+FpxySzokPDWEMqCk2BV8HWb2gm9j
UdALcoe0KlJg5QhRDRgiDL5idaD/V3cg+0kkNgKqJR7K3265o49M5YBV4Lhx/0O9
c28guqafQK8Mzwd+/FjzY8TKgIn7JOzW9fmW841PNw/tTkfWi7fyCXlREGjZ8gUo
H/ourh12R88aekmWbVvZSKtq1fkqMhYWTdPg+MJhB/XRzZiUiama6IofxzA42wW6
t6/MjeQink7KUhEHR1zX/Z/VaFyJRgLmm/UCqhHmyVhvMjsQpq3GI2Fa0+BSUj1k
vfXszylXFIHFk/2Cwv/SiQP5Ur2XSqNAUUHYKEQ3P6pspCwTAqFBTehTq/AaEEx/
C/kSIfAYubP5y8rDHskL3KxLK+3IJyjdadqw4Q4oY8Jk1I/PuTeqmGiq850r1Y/d
8EAXE59OZYYk+c04N3ZZpAeQtMyyaJeP1izj0P4DAQfKe64CyL55ksgKIEqoeOH0
rE5S+lohGQBdecujJdMKnAsnQ+YNOXM7jUBu+55OezpUSkDRT8dija9ymUEM0ZiV
Jmya4uVvjMMvDqKTHCFu+XN3MI/I4BVqqfHN51DeuVXFtVuPba4tv5RN9UhGIJ6Q
duBzMxjRYxK7FTiLLJTletkqfE40iE69guTr0DUjMNbl3qY6VU2guGE61gCkmi0O
Ucb7lKr+zVGAKMJTMbVBtUVLQSF0FJqA9X3bgepEzTM6BaO8RHTIozZjXxEeEASZ
qtibfA/z5Job36PTxmmsTp3AQ4sp0niMst/tUUsmTqQl9uKFwtF+tKVtSRns4HKP
JLbCMlFKEtZEzGNawRd6hBDZ6wFWWRBoxIXMehPpTi24hWgvnZKDYyDXFC0leRrm
zyUiICGk7X8iUa7bDPue6TSxIhXQO9IiWqVpk4ht2FteYhcMc09bThrouEHSlmJz
kFTuap/ykHndC627Ky4w7H/CRSKsDVEMaHtku5DRoUk5wNPnxMbbZvDC3vY3PtFw
ZrkAVU5thx2RhrmMeMCEFyOK2jA581O0FhUnsVRoCvKoTbaH1oM5uDpvtTbKQRhP
uWuu78A+DM8JbD+bZ++jBRouHrdttTfwBI7W5XEFlPvie18wySnugbreMqCASTDZ
XPel07e/tOmktVHx/lS+SaxXqI1o5get3B8likducMxjGjLPBbhdvQSifyex49+a
hFZwCgPWiMc8fINfNV1/qrnS1bA9ipeRVbadbSwbw56mWKKlVJtCZiQXnxrNWm6t
ng2fGC2vcDtF7XPBQriEh5q3eYcFOQ+3K2dmM6dna4gJK8Pv7AdSpIcqhb+B6SRY
lbyShk+J1eGy5w4TxYcfox5FhRfe32v1RCGq4EFtF+dDqU31PA3tZ6LFhs7AHqqd
tBd8fNlArpvxmvLvSpn51aHvIbBY3LCWbYDRJY53WPWKb4g84nBKyaEwBue92qYQ
frGig4QmGMjkQFySK3TDKogFyH2/bSF4yWIHo7KgaCPT7z9XfQGuIHR9zMMroipb
xGOAQPe7voh7+kyC7hTvEN7mnAwLYWUEvB13Q7m74/yXfMOClG8YkuLHOYKprfmD
BpQ6ilHPWUH7uU1aLowsiXpitlGoKbix+ffG1QUHZFkQQfNH1F1/UNBlxaKA69JD
2FGy8qP+mhndgRAOBzBsoY/P//nDqHKwMM17PqVIBsaHzXE3KSSiJyAewk7EuGL5
UV+bSiD68BPA8Pl6nE24cSightYyfPnA2dsSmUSrVZMcQNV1h3VrO2odsB8nBj6y
GqE3mvqK8GQx+jqGhmxzvcJsP0u/AEtBpuwGF4MtJHhO0DefJbRzrS4dHyLeF94a
UsXhHy8umTb44t3Y3w1igo45Rk4joy6FkWmpb/uvPjzYItM3dPe/3jHOMGJWJZec
GR2nQyMsQsmx1GBspJAwV8smCDFRIcExGfrE2oItUPueatQww69sAKYw3dCVAuaT
MtrUnOiMcPEnrzKlmho5b7yjuRe7d5ufqYcr/t883Xqo7BATM9caCQUSk76UczP+
5z9N6YZpw7YyNlPYniXFXUtFBfN+afV79vzAFZXDjzzt69sxr1NPxtllTX7BW2wq
wwAsGVeI3yJRHF45ZZdj2CYEJ20B1LDU66+rLPtfmrJBzdfS9Xy0BLmYSD64fBEJ
NwOxoIAjBj5j0PivTYVHXKmakZafJKF/zgMVcfPZfxLpn8adVs1g2ZJShM7fZeVx
oQZnl/sPj3krfHk1Uznpe4BwRHPek9EN8aVu/DbQ8ULOEZ43Ljg6/S3U3xoH5hI+
IVVm9pcphqgSVKtmlIpQv8Z9NTcdwm7p8z+PYqw+3dvUL0j5vAzIV7WAWIx1RGFE
ag7LwmoodshUpBd67S1zNeYeS+V2Fx3zJ2bnZcZdXJG2blw2Jgl5VG7TwPys6ju7
DjzXS9bp5vGANRXuwlTaT71G+/7Gutu1IpkjrXP/Nrz3V6nJaguKfODjUkxHO7H2
8a5Ip3W7kZ3g3ARKpMYfbUnKIiveH5uNJpT2ANdYHiJnjrSNc2o/zBIYzsVgNmRX
D+yYm82b4YvXaBxrm8uXl6Gm0cBkdsS+Tlnea+K0VxwepAxrYSptuBcvIRIcfs7P
35PzOVd7AeLVw2Sj1gtMO/7vOofdzgCCv6dNsAVNiQcBNLwdvrrxS5zkQC9fOIhV
GdheCjsL0j7Su6/wxISPI+CTAIz/OrTA8R6F0kK7E7b2pp7m/t5N+poHJDQ2UMHu
KPmgBcIi98Zi5TF2j35vG6YnyVTh2n3l1IP7MExLjRnF9dzY3HhE8pLqoTMbirwG
c5ULCT8UOHesYNQPpBlOB5Ljmpj7CqXtraifqgQCHlYhck9Gao/mYFEPFzcXXcRL
UzvOMvHI6NqWR29Rz1XJ1LGYRlp2Xt42nUalY58HqNG4XSPQeoqmqoDjb1qzT8s/
Nwf/pzO1zOpE6/cPMCld5zOvn1X0TsNkE7yNomAf3WNwur2Pmarbvosa4avprCB3
8X+V4mv0xMPhyXPU3PMHBJs6ate4BwI2EUpHIF0uGCXtEurS8aZxrulkPX7suMyH
lfVaNKU8yxUHDs2SG25l3E5vKuSozAMyOG0PrlSic0QArHMfGADgNQye5P11rGsH
zGUjbnYIBD4/po3nyP8KIAv8mPLB9KNtBPwPbuFa8jIhhg2ihi1fEWE0YT3jHIPa
EIg0Jd7lqy7gtE/JjunSZmsHA5KekukTyhlZqIdVcyiFqQd2EzqpZmCVR8Y/Vj9X
3M0Ak+idhwT86VLieYefaFStjPvB32bJDMsI7kCy8BJsD7sWANCAy5zbHLpn6Scm
20oJ6bPelhrvDFCYuomyoMkhtKbSik9keUCj9A73OHtKik0upPxA6pAKMUFFa7BQ
NQVtaFQR853SS3jBQd9CLg6D/Mut4dXwMe0kYVaNXuNa3reseUQKHEW7Sq/Mz9eA
ecYXMrx6lHg7GquhgAealvdR2RJkW2yT84R4AzxXP71zIPW5Dk3K7VGcEA24U+yG
wSB0Onqsbu9U85+ejWZVtnkNNtdkFlhgGle7I7BWqXRJOaqu7312oVZPMyOi7Lvy
YoQTkI6RHIRoayLWm3OOInvERB/1m3mzj6GSk6sNDb/qWUTRg4J+iO6494pTQ65S
eewAcGBbgcWWUJpiiUE+w0ZN9rOMoexWS+QQBv7cLAPzBWckOY5F19musYzGNlgZ
r7IMMK9rgnH/8+GlEXkdHzxp4OYAKIc9G7WPMCjbfvoLjNSzkDJ6Tk+XzkqafNW/
adjn1B/7NetTQZkZbSlvy9mMMhFCvmtc5CxgAlTRCjrb2jUfzgI9QoXxy8YrtVUl
cZ5RZ0rnt9ca4zFga/8dA/If9yD8Y/zTa5m3Hp41PHQH7CuJiOYXovGljJWfjVxl
VlvEhMlhgS1OQOQ2r/QCcZ7ZsXHIT0BqWRkTlyQqXjAp804eGMQLCQckQeKQxxEC
XYVByO/oSXShuWOVzes8APpKkC4noQFZ+9g/Cntl8hI1e3wBVIiflv8Du7a56uN8
A0E+/90ObH3ajGC+JGylt2FkDqS95FnlMjbzoG41Uo8H+8Sh6znoQv/5A2yk9kSQ
SEtlWL1eqSVat8cMbBfjI4gBFZWxHah7a6Yk1K/O7HOSbRIFKFF/lFfAmprz8i6v
4bTgTRUYH9FrACCmhLFJUQJjVPt1aPfOJKUaL2lb7lb+PoDUloRxyeZmiJ8N3iRK
+pURaewv+x53DT1kXJ0IZ5UwtJuyMwBAsZBiIgh96CcuCLzJe8sxICaZCPSbpda5
vF89P1CTbsOmTOr7RYODINunUM8dl84sjq7kqQA024SBOjm1w5xdlCavcZuasxXr
Ru/Gc/R60l7IINb4BFOS0rGPh2QSpK81k48BPFZ6nN2sentGsnnzby5UOBJ9iwks
2AMHaIYWjfzi1d7fiiUmYPj4VrmX9gIrliE6GEBQPQRwju57329IEW6/0Q5jKxk6
5kS0Oy3Ck4BygsTa3R5j0EZQcmkTBm6H+VnKzrLkImD06udildYRRNsOBXu7Sgrs
NmqJvP0zvAD847br1JwgmQA01Z97XUQMsuRMJYET124XevhfHHLJ/+GI/NPbyKip
V/KniCBvdNoxbODpXObu3ViE3QoRVfDpuak0veojl5ijv6BNDT+8JHmWg0dG5r4N
QeeA/dwU48LPVaT7H6/mpGPUgeD1rj1RGOHosZh4bAZQh5axe6/6eAcZQNkDDzzU
IMFgffFzUO+S3i1MoA2NB/tS5aiexJ/XfJv11SxaeEINSSLVEIl69rDR9hlAO4wL
+lYRJT2ehxeA2XUv7EgjY3vNRMGQzpM6BhNVhwUrdrSspfHwN4/BU8J725G6Xy2n
NPX36/XNzZ3YU3xjF+b9fqxMuWU762FimkwxtwQNWnpIJQOL/9k9KSwih88axnVz
7qB6Cw37spRWQ/uWZaCAye++O6lnsR6OwQmeKdJ8CUGtfWNnZKf+U4iRwyXHyxaG
wQbQ8LdSQjaOW8ChRfrs4geIM6Ad1/6s2TbrqLnFoRMDFgTU/YzOuCfI2Mn71Yqq
Fnsbmthvh5QVp2pTPqrL7LreCA5JFale5XtHkqKvhtR7XgESBPZbAngF0HF58OgM
4Llv04MvFVRpP89YjRLpnTCsOO+T4BOAx389omHe0SOmbbJTi1j02vro2Sx69B6s
GMa7G5k+7h+NSSIkdTZdTQk0rknhvcAdsR2RaPSL2UvGBmB15pk4yhCNTaeTBtNr
Zrf89sqj74gJNk+OpToOSRbtJja264iosmRGPaUxwB8P7xp68mIdw4/Y6Wflrd44
A/uH18GJmh1bpuO+HWJ+A1AG+c39q0IB3KEP2reeLBYD/i1bQFgndVgOVcg1IVev
p3jQhODqyRb7AMIASGlQVC10C+a+kRgCcHcPzyajySwtbzaz6qs7Lw5uEoACfH4l
iRSa+Kt0oXVEOm4XGLU2Q1ot1wHlIO0B4t4mLwEhhVBGVnMN+Y9jJGf33ExgyOUu
nY+78pXTPXbpsooFLpQhDK917AAWAVXBB7MN6GCiAYs9gWfbmMGt8U7WjRhYcDbX
b7b2jM5GVE7L5dm7Q3BO3RcWrrPp9418S7F22TaH1Y3k3fYf+TCckYdCMNL+DVNp
wvGuHqcCG+h+1MXO6a2/IVxRsD8ZFJCVGbRsi9zpsSNeSZieEFlH9/D/isckYm/1
oC3pp83uI5+dJ+RaLbomfSvmRA2g1VDryZhQNOXbQZQCAU+1zukdyPecZthhYr/9
Gc5n1qVzqnBh+NSZN4VqNNRnMB89ShXEti5Vd1www9tjTw1DMPh2H017NI+YIrgK
2HpXIwkvQpIjzBtT6veveVoVnt/XUv8PtYTf6knhHYA6KiB+37QPh+6D5pFfkonh
nFDyOyAFkaaQ2EH8arqpex2L2AHZv/r3VR3SM4SqB/9LgjG181W/GtwXekkBNm6K
Hq7g24AEzeZ75b5FDNlENUwoUiHnWZ26ZjavRaKsLPLx7OQssvjf/S4AE9zoGxHk
0v7G1wYjAD7LaxvPzDLgqFewTk34QVOggCMcZKA29EzGCnbaCjj7DrfoQvp0gwlv
j1CF89OecBEzGaXI/RuF2PUUike/dPL1OlYVVhYa263hjLvFxZpC7xs2HrEhTi2E
TQZdlY8WTbQmCYKyPFPCNs1ZK9GDvj+lE5lJDaBYfk+4OXoRCzmgjgKRlYEvZ2UD
3bD89CtFOL5p0RtJGN7Uk/DhqsU8MVPurPvX6NY4hL/vRRgNAwEpjF76lSk4/uLf
ZN16M+JBd3aV1KuKHLJSpxv/TOJknbVwmpsi+RfDZ++si40yKjJgewhAz5qAKeLh
QFUm8zFW7cXjNC0EXQak68V37S1uMsnK4LlFs5Mo+RRoa3jSbyMQwsUUerma2Ii1
O48diqW0+0BWZhgo71/qmP87bJANxX/6RPjDWLoas7oK6vqAvF5gMVgmNWuc3XaB
ke/h0EKHM9WPITVKCAo6qwDw2BZwN02aEl+RJ+7anbe4B2MTq/qlZyxvVRukAxus
GIg6O+YHXitx2drcgwRaMOa9ERNksKtM2UnBBSnZEf/XSlO9htNc9Mb6KjQv3w3t
ObZOYadVx8VHxw+B8CTeDx4k6UJM09rf1XkXfCzm1GNDABwre9O0uzlgiz0J0D9o
er0HpBUpRPIjIWuxpEyCqZBAbFTarqpuaEx9aFKBOe5acJ3n8yEkXdLs8D8lIw1d
bxN8AOugWLRHQrOKFxqk7BfpvyKTWS0cEjtWRRRau9ApuI0nR3MzvjFTzkOoMN0s
wwB2quIxaVzcXNYfQt/aNuEI6GD0Hue9kRPPapX8jwmG07f9RhUbo+CZAb5YIKoX
LSfUMamXu6lvdtX+z3BMV7VyGBSqipFc424ioSlwDPuvtidL4kfLoBFtB4VT5Sg2
0zR0O7jUo8PTyGkCu/azvDvJt3ErW0w+J+g0ths+5xSwWqVU3DMoTA672C9WlKif
17UDXK2VIHbWYHJHaLMYHuhlTpJMRQknxtOiQ5cu6IH0gSW0nlLIpSZeGy/EPj71
iQjM/15j+r+cs5dQbTIXXbRvllCu2480J+faxdhC5yZHA8G1i3brv4DOYceAwAZS
Um5Lr88XRa0IybiWZeFJZkJDENX24el+GXZpBSBKGDVcPKUniOb2INUWFrvgz6mc
p5z4L549VG/Z1b9XxuYMCwK3742a0+tH67otKBMIPX7oS2LZqTQu8WXPQ5Kh5zES
Quwz+T9FaEek6RwLgqQKoiREyTwb5AJwmg/aO+QIY84O8gv3YeyzqTch6ONwwE2L
uipzP+uTTCVWwxODz+dG/fkaQ1zY0MTI89S1ojPGxcwA7PLkiQr8tSgUzNBnbOr/
E/F5F/aks34BNC8bnxdNBLI8vB29k6EuNhnLDst3lPp4B9l0/m7mEgqzjERVL5a/
4NUqUztDgrv1aLk8N6APrErcH+G8hyXEvzlBPnpJyYPm/cKH+tISbDuC/WhHQCq3
stEHO351GQSe7TtvtAHJRVYN9pqezF9X8qeIxLyKZQoxwd7HQwkvbXPKvkr2rbRy
7VAG2zqqsQtMhk41E7/8UpsJQ1y8+psEztC5loFOTDBP9tvFAcsjOU/uMotqYYrD
n2pcRgnMcInZa5qFzkx5S/V0sua05wOoo0oYzB3kYzjEC1eDpNC9HAgu90KSIJXR
fswLDB//AaLZCnTJU/zhBtC605u7XWU+lSODFM8LZU6nAPo61IwJxtJej1gsE8jx
lvnjDu705uw+o8dNCmHCDU5QDhM8pQnVc16+NdROTkLVpQGMak2VRTUqgQAF8nUT
ML/0qHN7D9Tg10KGVIlJfarQbkVqc68GC1Q3d31e3gCwjPQgIQ2IIs5mlZ/XwPL3
5hKRi8o2DfIHH7OOo9ICLjTOFp1mL8bVdFwLTaJjvh3ikeMDakMqNJs4avlz1kCK
rt2Jv1G2j20dTURNcA3g64ws4nHKpyqQFDhmCH8mbsuHPwmAENb6BIvX3/2koqPC
4NZ36UTpkoRGjZRY0b8BOvlSk7avQOHJU4wmvPDceN/ca6qBGhMKmrdgQAaIU0Nc
Jt95nWyUVYgRMp7OHvMgaD69eHmVJoDjNB+lyUTwaFAw8NevbD5LAO9IziyVEq0n
5/ukteQpbRS9nxofQUpzQac4wt2wACRy77kXdSEKG7SJEmhyCKmWJSsIkFHwyD2t
YL9UWA80zLY79l6XEt31Tev7gqepa4JdkFCUPRFIXy7oojc4pLUuT+lU/WAHHGL0
q26rdN9bPUPK99rjT5oAn2+KtcjQX5bqXmTgXTEgkFOci3CS934JOP5HGgI7hSVp
i9h7AmCW51tqMN6lF5Z8pPkTWz8PL9kKGVg9jDGlLVhgwhL/clA3wwHQj3tqN7Ze
3kx/3kqgnpN0GhF3DmDR17GiqKyc6eRVRyDpBx78rkGoBN58W6r9CUvavUp/oodg
qsuRutwxO+2hr3cOSQ36aLNWy6sq7zOm4pHote3v9dUNRzpR/+1QiSodnzDwxsgd
qv6nHe6xs3tsQCnX+fIH/w/xRKgTmWs4kZHBZzgq2H2d+QihTL17pWROHlkRTHqG
tjZQi5cyZTJUlgnYNIARl2PA17ZtHSfKYaBcSs1vKIuvcGLbiU8iOj0q+mI3fNFq
8+erjLXl1XR0hwkhserm5/4Kb1/gFTyvgpE3ePGeNUmwfXU8wf9Z9MP37naxRKp4
A3VY+uadhSan8q2jvuLzH38G+cKK0GSVjH4T8k+QnwEIovD7faEUepM8NXR//C9B
Pkjx/Lue7Hc/01DWv8bKRj3LcBY85qqYM75mpLWjHdikOe+WDXT6I1ao2JP/dAhV
FemopujCCoQZ6mCuUsiuSqS1IbbKpqmO/REr7m3TNgtOVvzEZ2EWB0bzQ49t8c6S
vIbSAqYOqp5+zjJqYIfQ1+sDwgkqfnq328ZDbVeEvPGgnSnnB30syGgyhk5nvuWc
f40aRmxnTntnoOy4cwlzE1bhBnntZghlCJHMD68QXz8wg6as3Wppu1A1SOXhpBYu
HCYHVyauXNsdfFK0Cw/mPPsG42XH8uiAYLYDsFPdOjx8wIyyJ31/+q4NuMrCG3DS
gbpqkVebSH1pehBbUp3VJ54RGYzHsNsEGFVZFwWVMxKgc+z/s4mOGBtXjt/IQNnd
CLkeNQ7QpXbOeujRbXb4jjRwGGIDCLrb2EyXBCjUxBhDaThvRUoBDyicSfYnuJDI
seVhTr1iD8K0GPfSpqdlz5s9sOKPCh0vc0Ps3YLNv4Tny1MYJwpBcI8+NxEIvy4m
tlqrlvEXEbsdGma/YErQVb1hgrMAb1fhISuoU7At3gqOlLrofDaHOTM45bMacW4t
Q3nyFSvcP68rBtUvF81LQhZPyVdZhuy8yLoo1vcFZolukjGJgxHa+mR3N84xr24Q
LJaroGIgxkiDbn+EtNWOAupBcniSclmlUYTYWdo27a3kNi4dR3mk9YY6WREN0/fC
WZYiGFS81HhJyWho9OBl4ZOFF0rhMoZ8yugYs7lW9Tf63hHxrgbA0OPK/eL8zcgs
Zw64+nY5jEXehenWJ/KTcZ+bbjBQjcVqE6DRUqfJUfuJ9Oq9YTTzuBMNsQ7AgOad
jT7oCsXyXbA8I2uVCKmbmeJHQnFIcXgT7aGVeh/82OewnDYbzyDDq67iQxA/6Jvn
ni45Rk7ExB0ItJuDIHR447Wh5yohOqOjuUd6EueUxWK8td0I3q+cEsGt5VQZ9kml
L9b7LHlOEz7bmW/Y1bSOQ7+fi26t6jvNMPbAco0+dfyKtJU/pd9AiZ9P1pxEqDsL
7KnQ63d1zPmmQGhqUfRCsLH3Ku+vN60mtl8eqWx2aSD2m+A222yNoed9qT4IDifg
9BP/TPKYVrdbWfXk31mcXL48WfBX0K0uxYuvjb8NM1n/HNCkfiWhYXSA4GlbIXdJ
GcRQT8+GpPc5O9AFJUPkVsoROXSyXnYufDzGYCsUQNwZ6ad56fvxV4g5eIFXHYz4
8QLcUyRIPgaXyr4qzKpra/ZSsI72FCgU7pRXwGnk3FfXHUBnwDxKXhT7GRfnNYV/
dyi9Wo7lweKDUEgZnie+MryTyaa3SQnnA3WtMhVwTBg2Y+RhazYoXvnp4nqIDEW2
rxJ+AozkLy6M4pl9Ggb8JnUQSlG34WL8Ozqn5nLlUi/N8v2AdMcB/Mhhiq/qThwV
Q8Cw1VaRrhYndZvP7uM5FQD8TxNr7bcZFiezYBrdtPH0ekSGWRLaItsdgTnatTzH
NeWyOPkYYndIlTaAb76Vh1YV+a+IPYrcrFtVHbBWswN0OTwpsSHHDRMz3Q7o+5io
7K8MRuEkuf7wEx1qt8V1TZqYZDf4XFeaKgsXHEQT5CIN4HRiowlEi+LFRwboFc5C
T0K1NMEJiIWBkaZiEv5Yu076A5gtCzXPGu4T34A6peHO16UFcM8wJ6FJpp77I+I2
ugW6+JKQmnR1xoxf3tdzglatqaLPWAg+2GGXEikzpiRvVjStt6203ylqeMPMgYIP
sKphIJwXwy8t/zw9UGwrTDASClXzW82r/0gFh2jbQbI5KNo3YMbmEHncjSd9yxAB
Sg3hSm4ncL2ZK3+P7VEtDGjpicWKysQP2X9x5+D2vMcBOleI/W/Ymc0mUjsg/GZg
NZzVMFskf7NDwsBLcTMaCH+mc/ZCFMPpU8oyrplB0RxSALQnQRn9WFerlvRpOzYD
4QWA/yAXMxt3X8x0g9gMfBbOii7ZMG/gEc6BKGu2OrPPboMjiTUYIRXTd/US951D
k+zhxP+/IjZpo2wWw7CRIz2GtzkjaJawVF7wEj0FZ+PYaXI9SNC8Ex+y8gfyBYnT
58YGNBy+HwdOUA++3EhPM9SfCKO7DNRzBgzERIlClJq6fc+qYSi4RM7wa3V7JLf7
YWzzjIJ64Frnv5Fx/I2m1wv4b1DLdSxz+Ncs1a5/LJb30AI6IV+dWedYuW8k3U1X
Ei8DiOHnj5JCsgqjIEgnK1M3VYo683XZdwf3eZ1mhBmyy24e41WyONJG3rxrkKVl
okW6mGuRwlxKc5ZaeoQP/n9HVehDcHIhy/VY+6HSWEUL3IEfi9vgO6M2yn8Y74aA
pkV3mglSUbeCGB1rdv7kAQgOhoDPoWBty+ajLVcqgqt4yr7NW3M24SPGI0ZXJWF+
C7h9eo9kD+WagMnm0xKGsfO+B/d0YfQlnngLz8e7ewTeFsxKg6fkb5NXfKOTW2jW
qXyIp6QiO2UEuRHNLMqn+f1y1fhIdrIjVX2X0VCI1v2MPQ+EHfZP5hmcAY1v5FzH
jDXFvFWBKUfrsPhTey1EThA+FiSEpWftWNsyUOxEJUYSpcgQicW1pZRS1vSXOfRV
72qfMQp5JyMRs8wY4M5m+u33grCq1lmAD0/EBrpf72HM43+vC2eL9cIAklFg0kfr
IfiA8iyf2l2RBAqyhYpGGvgTaNWhlrqwKcCKHWZbWamhNMYpZh0LSij2ZRi5Y8VV
9XAtTlqGvFiKIFNFFtgJjixO35Wf9B4ccQKUWwMtPlLl8ROm4AWbOHmmfnM2Pc3Z
MDSA32q3k//QIa9NXWN0ce0HisUrCLSms2hYz86KveckfU0CwhZ2zAzh50QGek5O
XXKuKdhCBkwUBb62arnR6HxhS5xIduwxSDgAALoovWWzxQ4RaZxSHGF9FEByZaoI
sEzu10SGQAqaWzA57TZkaNxUbIlER2wOWnmtX7gFnGDrE0tlUa3vGSZdO0jDrggX
D4GvyXJE0fYDKCt5tGSAGeTFHZDJ5W7B3rAMykAdtjxvfMmEQPY6Bygp+I6+PXas
dlcXlY3JWv4QsPO+ITFc6got1h495q4JZNMo1G7YwDBqeDfOTty9NFufvZSq3lKh
NKNeBZL8x1zjYHwxf5b51zSB950XWvNRbJGBFk+6PWvzklRMhgIJvYQ9ILPSkxMC
IGGgvC1u9oYbuJh70HYM3lXlt/1MjudiSVYsTCnEjRaXmETh96uMZ9CTqs9/Yubd
oi/p6ir/K8/Aqb2IKHQeIgzZm6GrmahZyuSDaafJOk+XKC6IVsVbB644RbRUAMSX
dugFVn1kjSlu4HOu4dyrroUgUyPXh+P2DVqKpTsmEHyIJBKIk3Qs6WW4DHjCEDYH
cjeOMCj49eNhYkSTAZSxuFkAOxm1JEHXMJ3j9Q7wi0lVflkublhunGmxNpzqMMCw
lr0NguoVmxZPtrftMBprbwQvNhkmkHw/HiYVPS6AbwBI5a0sWHvFgk+kGCUEQNAm
Z8rggearEhnXE+TX4wLJDrcrEs/nBfbmMQWUfNaznVhtjQr1lpXT9CFTdQWcciSU
7RSIkTYqt1A5BdKexrzttYwtryWvxRtirfrpFDwljlELtTGMkOuqmgrm9UAVWLEk
lLSaK4qWJFROZ9Au7S+lz5xVkpu+RBhD1bWcoKFXWKwWBf5kjj/KcIgOkaNoJ3hm
52M/MeoRSR4+Z7WCgNMBaSeSOuCm+6StB9e1xn9HAV9lzr9XXJtsBMOR0ZORSVvI
Vm99+UH6YPA0riEQXvirIvNjWAmIHTc3XsT91aDKgMzku4MEH3GbWPxHjapFuBu0
2ijlMMB7Kp9+ocmQ+UDizOFhI01+vdtqe1307ObH93avycTvlNOvpSXFnSaZKwjg
7+a/B4LGd9+Pl7g9BSJdHa7w1ZqA73y2q7J+MbnuW9mKhon+PLJOMg61Gj4ju1M7
rz2E7NVVLI7Cvuoe4nKG8s2AxHeoPk1PWgL6RjH2pcxdtCRywwgtQk9rng7r04Za
IxzhyppnGFYppkg+9RfJJochmp6PoVnQ/vvNKUS0CC5YuQIBAcnKfy5i5wq0l3Mw
L6M0qCrkNbKZK/0bWYnTOaM83U1PU2pIkvywjv9RMJC0JbG2IRN+qvXYRjzIDJTm
Ygw5bqaTc8UwHJNH9+Ztk+3OqA4vlIT+En1ZoDMXHSjy3kNbk209iHKmigZJekvz
pfqNQTPVl1PFV2trosibUqkFyX91BfmAgPjkWCvy93JV3t9p7Ip3Pq28EMjxZYqf
xwtggD144jH0PFdbZbFMSqUEnvmz5yR0/ssNDBmhu4Iq6cSOlwgoS6kHwad2tije
He4Ru2nLh/QutQvJRaXvjd3uM4WGWUzJIY0mUKpx+zxGRHt5pXJiOMyQDauMDvNf
nykZft6mS8I82/7VsehPI62KJ3Nwgv8lcurktEBL2l8vMZ0IA/caXeJ1ik9u2iz3
u8eweFL6vq/9z7RWcH4kI8KSNSez5zmCr4orcsI1aLJurB3X/sAm7IifUiWoO0G1
jw4DB3NNxaKHTZ2BE6s+yKAXS4kCUBwiiP+SDjk1VE/lhq/Ck2Ni2+b5Yam1lovG
7R8Fd0F1YsgNZ1aW7yGoRTdprTbjDhxiu7330IMJDIyycMzzLqP3Iv11qsyrh4l/
0JYtktkEoask+UWwvY9x/LuZlNpSqGvAA6GF7zv5KXowezaT1WKBXjcaN9/DGYbO
eTVlZGTbjhCs2fgU6xs0zoSmo5xtvoYYgHqWEhVNzUkzSC3S7wMWUAc27E8yjgmY
iNkTK2BBZsW2ZqR3tgSvhQCvigWa6sH/5sLnpqH4Lx+53R0GO7fUymvvHse/JTMo
dA553Be7EtiHOF2cuZwivN+T++5Zv+URl25CTv9Ge4xeje3J25Tbrt3NF+QZN7DR
7q7Es5OiQ8I+UdbB2igEgLWm3z9+TxqLwaCmja1S4Mvh9iBB94mw918ALHWzOzCu
1Y8jXcWQrvDFDJWy4wzXD76WaOYuZUoqGwz319XnH2SOKyngYIaKn3G+Do7CZhrV
jZ7zJ3zU6ccGbjqWlVekODg4aXwdvLDMjqHVhMzZxYReVpbW4XnSdN/MdKPQXMYp
gC2VgYzn7EStt6Nhb2dKnvrrQ96+J/UUWaJp6IRmRDopXp0ti3lU6z2RM7en301m
1nLVG1TmOxBGinmCLYVq18saXPmucbDkRqYC1cnqTE3wZ2CBF2QQB9VxFIA03qc7
uZvCse9qqVqgOrOQHTCfEQrLm6xodmDe+C+NndcrejkqIlNlm24X+0fawkdiKPFU
9kDdpd21MrBc9L5mylzUiLiWw93NUl6NuYClCSdI2EeAP7qaXr65mLfQyNT1zSk7
DeG8FRZBFAcqAQdkU3+zBgOsOuNuvtsmCtey5EcXjr0z1n9/Kt9TVe5zV3Tzt8+V
Zf52R69Y7UnjSHBzzFCHWhbpo28bejBmVboII6dYwBca5EgWDNvLSrH6bjcgJMEH
BWvSjgCuUjfUbVvOyiJVG/W+nCeOyZ3tO5TBmUJOOT/zYHwVtInNCpoRIAL783I+
XHbc59D6V8I3eUKtHMYOZF2B+DfZFzkHHyB+9/Ra6s8cEuIhFBUROOcDM+EMUtBj
FFf+0ObOFVm8/5oQz0vfRbi6OIQagZOWMdoa0y3G4T3k42jjuXhOUzDnTGSfALR1
pUYWQpMzzaxBp9b35vfIqQfFvQBwmtuk66ZdUBK5pi47TCWmMrkCUE/o7S2Sn2WS
TIdVyXAGBFIb/jadj+sd9U98TutEtR2SDdDTrDtU3scA9HF2ZBHug1fKwbIwaH5t
Y8ydg8h4+mz0U4nHbh4hPc/TJENE30jqXvmeckxycWtRG1ZuEEClDwaY1bwTwPmI
kr1msdKsReYqvq9flE5T2U8muqiFeCfSVT2gamY32Nu/X4B0zU02HEFhY/9GZ14V
TwzdnEKhXo/5dKQki+812N926/U2WKzkpBKb7uYF4sT6wABYdjOtrqt5RKzj79QG
DSHQAMInyftvrMLwQyfgaRGoMAgQWVLzK8f/x+d6Xl+GgNibfscEJyK/2OQiTwZw
Iordwexg5oF2rlI1KTbSIE3xnZoYOy2zf0nsJWqkDilE9XpJ3ytmCtIdJrcf0xJB
aoKbrib3QHBeEqaVBEQkYDLwTXS46v4WrRFjvYdUbSdQED+aBSqHwstq8surtlu5
42Vf5FrKU8MOVT71/p96Li9lFv7B9s+nG1orAo+aDpqg7VNhtZZN7aQH8pNFgubq
80p73g1eFdcpMnarcNIDB5sf1nczslyb56AuvsIxaX7ikTFcKxvIAftpx8+8D/S7
yiXsnltTBHmbFhm8RIjkXuiM+EOFeCEwpgJrQHc/DdxShBVEzCFG5fdVzTvG9Ik3
bzjy1I5RA6IP87u35WdxQJz+qcm/oyi7QLTT5bGcqLP+a4Pune+3dRobf4lNMV7s
Q2Bto+x8gzr3ylxMwRK43teZ3fk52It1oiuiD8xwaRcehOZN1NMIA+Tm/vAdDzrG
94aJBqTbywEIAjS94CxVgt8HINH+CECpNcxzF9yN2DXCwLFFQnJMtfNqxoHGBwkR
YfHUQ754RAAPUM6WsYYXWD7zgUrCkW/k9qkFoa1rxokF9uU1BgTVxz4HjshkeDv7
M3fUQ0Jr2c7vy5juXHVgwjjk/3MQ4bXaoFAthpM1jLNPE9J8cng8vLvKG+yfyM4m
E/cTIU1XwhdR40Z4JvE1Mzfl33R8ATHSE8TBscGzxJkm4vFdGOjQWOXF9CBzJ9Nu
nm0irEItyvtL8sjn2+sQ6+X88GnWDg8SZ0SMZecYp+8Pm13jYjxplh+ymliOyDWu
sYfZTG5d7bkWVgzPG3aAwknsPJiJsZGEJ6bAiHJZp4T+bCeHIzhXkmj5WTe2lPyU
gKsVwSyVhhFxxzDd6e1ymkq6whAg4QpHEYXy41gmQ2m2eVtstyn16Hr/C4r10bSe
5Z8/WP/jmR2rifWDQAkMg0Pimp6WOZpc03SI2O7WUmDQxupWJIgHlONUxstni+02
NdaQpnGeKphV1KNRYOW/+vnx7nB6NbPikBre7flNiO7TWcF37id2wVItYjTrsyBE
Am9AIgyjfoL+ecG3x7BUrLbtPmAIoovLKtrzDgXigzacAuyOIzLmJXL8rOC/l6g0
tZUaCobU+ltUD2BSDaaLv9TgdxwLt6YnpgL66UMVrqXCGHEAH+61ZEyPsNmKWrRp
AUzSzuhaz1lkDn70OigPQ3YKireavVdxaqshhAiVncdo6dwC8KxlBTo3EFxMoq1o
3ldOqITZPPeRtgAThkHMsct02fDnKMWY0Nw9Pjw/9fyBRsxuwWPR5rI+GwY9Ds80
HnQ/iHgTeIJPtymV1iMEa6ePCoAOJ7NcmOS+hQL3X+KpblGGPD3dnOLf13F+yhcI
G/v6z1hubY6lfy1c30KUlM/wK6NRzhBiJyg4NPXh6sfQcmmKRYZXeuid1e00A+7e
vbnEZzvt2ALKMzYfiZisLd/rj4sWh66ZL6GtYIntzVAIGkyxwXHEpAjjm0pBx3Ry
JUHtH8jie+X3XYvH0Ne4HLzPcAjoC8OJ4f5FyP3G9pjccS8S20uF8UE//i+efKtK
jUCTGKf5Dbl5UnanByQpFYxoO7Gu38TefFSUG4mO0LQjHApL9gpFVHC8eJ+lwrI+
DAaDOiPMAvLoHURWQNoql6tAUYpiuaweLJf+GX8cdr5sjl0PD101zATARtuHi8Lk
yuqM2ziUr2pRm1ls1mnEHyC+Z/c9QgOZBkvuwIw52oDR7a5WuNNjRbWM0F6qCBl/
mZljJRSPqW7c+sTJkvBk4DjkZgrX6VLUGt/W4fITymSJ2o0SPedUs3CHf545guPA
FaBxxoliIB02BGXafVc8eRiz0Ys39/jdnTPeafsbW1XcLO0uXhwYb2h30pEd7hBg
L+TjyY6Wu8ZKuBogyp/1TUATqgsRj4tdD3juT3VmH7TsDQuW/lV7rNn3bHpW2pHR
bHHEdb4GNRRgHMF5IW2eSf0Pt0EofZiB4Hfz5cIdlBNxlCbfTQ36zTjnfjc1lge4
WLzSne9d7Xw22s7PG6FbfCNrHMjWHOL5syWAjYtODoiB7co+N3JzM/fBfrF/zz1H
dmCoH3RctZcTVKUxG2KhHMQ99DB2exrCProsQ7UYXdL4KKDPrqhKW7uMNzJGzeDl
p/5d4wkb68bHtfdu0RJFtx09MiH2VKx93U81Na8VB60j8WeKqc3WAQE+5jfju7bJ
OzfmKX5G9sNxKEqsC1nFjGm9GaQQmXGip6gIqWai/I6FhKHwUgNl0nV1W4QyLCKV
qRlG3onD0/0zqQrNq53yVB3pMgYdPUJgmziZLC8uNwegb+BbFjl/dA671GeerugS
EdgRICwn4jIK8wjAG6Egj8tUqPeJ5d3XthKy9Pwo/tkx/y56lNnMjPDARgYa/2ZG
t4KW4JngmDka2cDUtdr2m9OVN9wnbRjduzJ02y6tsH1O/AJaZCsT7ZO/lpmM9U6f
IdbO6c+AIqTvX4Bo++nCEOAIuVidyjYwBBghoF7ixJzH/9rzPuYb4htntDYrnRMg
dLjsKcbpHnmArWhOcvr5jWXfsQjgMgrKOX4BKUSJ2wxbUsEyytJ+6h1M0X9QnLUw
hX/kJPWWptUqsowBj+Np40TkFcWrHw0jI/lanh8Uw04Em6NAb2WJ2QnAEqlVVtK1
lRDtCp+lpttNAjiZUIhfRo0Sb6gLXA84mnYYxedYnConaV+Zg7b9/Js9VBsLjG8w
LgC4LVMT2GgIMZgRubduWlBD83CEgf0sQsT4K1hYkU+qqgT6eMDAgqlWaNKSFkXw
rWlF6GCRt10poDL+icyE8YVYXVRPsnINr4bdBr2KuGNRfUqldXafp9QUmQDvvFZQ
oPAKe9xmamQFmykNlT+vzsiskC22UnhFWh/P5uaNCuInXJO+W+3oU3e0WbkMlfhw
j0sELamSIL0bQF97KxLdcIxgpBd78sgubDyjD8+YlW0FOg9IiRljgT0Pow3EfSBi
ql11ZNDn0+8Kj1jaBmT+WjVIILHa5qX2Su++80CzFQUob6oKvffSfJlvfgpF2D2Z
1kG3RrFOe0FQxwruwNgs6gPnxewx4SOU0lkz9ZDzQoix2xeESr69+RsBTSBEec5W
i9BhnWuQ6fGanQbcUu2HaLC3g4kFh+wgFwoT1M6LtVftOMv6U2yDQSqFy5LrNzGU
3F+dcvCNJMOARje1s/qhFk3d+EqAVRWg59QifMJn5ZqouVUtVE1AIdGRYz6XKzfz
9SCB6sKRj5zDDlBpqoCmamRB7LPxbwDqRlY9T+/edcx6bz+gBo+qLMEsx4GPqkCm
wcWdv99so9W0TLuNQRRBIjd0BVHWY9CvOJlR5/dPtM8ebTEfr8ZRHYqOHodTIcGZ
z7Ip3myaKT8DTTyY/DsJ0qphhnEY9ksHUTpPvTe9uk6b1Ljq3qi4gg5hoET5ceYc
byoyP5IVg2fXxopkm80BUFM6sYa8HlXobkoFeqbXg1iEBkArlCz/k9yiAXyBmm3u
gHeHm4cbwwLj2B52Tgg7o6gxNvTRPnELeXCiBcslN+rE+W1H6ZpRyCFpv5/6N+LT
0fuUqyClRT1wmpxY+QQMpw3oqx1dcQwuN/xQOdMaYeSiUu/HZhs9RyoOIJY9lCUA
Pe+c4lra48NrfVjf7Lf5EAnUhVREMJWpiVfx3H+ajKo92Khfs8hlCYw3o44iTnWh
xkqKHySWx9/gotyCJNS37G4gs04l/tWaZRM3OKAwiu0tIw2LGqvlGwmB0yEiSvKu
TcGVp5wwLaPfKOpQt+BXS5hKQ5ph0ndAli3yMkl0VcVCpqP/LubGfq7kIrg+3WvF
tZXw8dLbKTmD8eCW2VNX9idKlnQiEQa7Rn36JoF8YZUKeX1vDTbIjgO6HwYQG9NP
APrA4KtAhdAIFX+HTg0nswqNSIeOL6+iCzKceGL3zNSWpKnHeKc5L1RUfg8K5c+g
bxkHEJfyw57WgxMcGCgzztuErKk3ozzppW9TzJJdZyp8i8phWoyErhFAffPEYWiH
lpyI/rhPfcnyspjvyfLbgxGD5iF06b8dXMyQThycX/6T0cQ0H36DWXsCU2bbPvh5
opWzej05kKm6OsiHP9FUYAxo6zd6hKElW5QGGD2hm+3nAbRBUx1HZMhSy2uDuuq/
7LgEKmU7o/yEuYwkExjBePCrPpmccN4Sc/cW/VdW2VR/bzbcj3kwq/Kvs8A55q0a
LaViGuFuoc9lK7NhLfWWP+mlQkWG4aFYnvhMX+SRm69hLs9bsCa5lAEK2CFeLS+S
7e2z9k3PJ9sghEQXSd9TKVfXp9J2uTh9W6BBLEW29rsggn8f9fRW9iOo18ByfvuT
U08ouckpEWe5Z54VaQ8k5cGbizxMIlhG56L8SvpVTORFAPYqLaKUDf2Zv27VanwS
mkAgiyj+AoXqaYC/fZlHyiVWqd/v9jXnK63OJiMzhTXmSLci51rP5DRqTznDK7pT
M9Qm7zjlJJBm6lGCLYhY6TtOud7mRS43azGUMxAAem6omq20OQE69XJlXd9/EWAp
cKTqci9pa1wjEjVgbtE4xeemkINVIqJvzAZY4cZ1NrnjKF68ujgJuvdYd6wCULAh
4bQOKtkpaCzHqlgKsdA4AV9TUXAdEMlKAMOKjGta3oAtukH2HcO5TwooJm9M/xQd
YhiE+rGFI9mlkZDCcCxoJOW2fm/sAriTnpYLM1CoSLqMJLffCH9Wval0kvyDyPEk
9Om4XHhA4PUUghn9sr53b6vYezVxcQMFQNHYqhSNgKTt6ARSYpgKHjWTlwE6/qQ6
TWEgAZL08x0avIkZ6RzXKTrTAMqpFfhEgcAol80/diT0UzBGlf3C6RFTVpYoLoUa
UVokIz5d3AOhMiu/7Xr9Dj4HzzECx+pDCif2PPRs7BxNKXhX8UqmfxL+nELF1aJ4
2SWE/Ze37Zwc32qurn7eUrVz6WHRv89zz7DPcMYkdVRp4res39MZOMMBaewE1N3o
sIBqJpn1xbBIB1l1PZ7bcWj+kho4HMMHDHPTgLIrrzNw8YYCAxW2/GXtU1nA7EuC
HRas+iXAZS2SdRNC6TclLWQhQYIVOxA9n86lomddI0/AK6UL5R/hu0pUbxSRKYoj
hrT7Ruzarz4oNw1YIozknsrfui7nmgbUCCIZn1zgphmNMK1cF2eeSd/BFvkotijn
Vghv8Yg1fqxAKq2MIuK6JsNNWD29xhXiOuLxUH2sReEPqMKCmunfJzUq88X7LF4v
M+CnI4kxEymRbvx2XYE/4AHq96o0ymXZW58WOpiYfXPysfrq5StYsFYH7z5L7QEs
M9GgLjG0d7lI55gHuTDexYVOadpYov1NwyMGmt237f9OZJ0DOGNLxqdzNpKgR1O1
Q0ywu8bJceqE+e0XayRTlqhp9+76G5wxUSpoRvmpPs8vYz0Em3r9oq43Naty/jyF
8LIRH0A3JbnogN6vzlFjrN8JgX/QH5sLfuFWuWMbbUs8nDt/ggVgKEYMqD3yVFmx
BpSrPfPBCaNlgiQnwQMb0qJvOd8e29nv4N0u9o2Gr/41OX7cG+a6LNsSuFIebMxX
tjMGD7fDzPw1nKTt+st00kbpB/vyt5QQvTniYIf/nbFHTrYYqbbglCfI13qyjDIJ
hbeGRYsjGiQXoZBGp7Tak5fR14Db/my1fO4eU3UZqD8dy3U1z49Zz3pH3duZoL2b
dMTRmkSM31Rd9L5lcuwfye4bpnIw8pmkdXO5X18aitxqEq0d9XE8MF/N5BVWcoSX
NwAGS9AK9OdRsoQwY7bPDwfUcfeeULzK5dKfCEzXS2al68oTvd19Z9PjhAd7hZiw
PVNekSWmF74B50dLu9DneTbsmnWcZB3QAK9Fjl0sP32f3+mp0UW0w6IDhcjpGE4h
8zgBrvapHOjgnjWBXX5stpat0WEioHEmSp8x9RrBvBhsfmRK1IchK6tKlFV9WohI
4WTIxC2V4XK20RtxxfDe8y0Y+vcGzuoIHeUDBjfjFhy6qIJ2dLhye1rEfOitR4ip
CwmY3NCwh2rfKg4Z1AYQvvHCFnf1CPR13A5SW4+cY/z7eFY9/xdXsPyTBNWzjzhW
wLAvwhwsuK8vFLptlqR2Uf8TmCNJdDAcTJRp3DKtCYcbxHDKbuyRXDr63umaB1hN
ZI2k3GnBHiqrEui9J4Ru62noxf5gKqwXBvIjp3CBwB6NPIv7SoyD851izYpQsFc2
u4zsSDxinoU17F9wh14rDeRI6zzs64ORsLrlzEfZQGtoLD978Q3SgW1Sv/qdy/lK
qtQ0MWRUdtRfYW8nPRNz0WnIlEOLQljOD2fdKdqevGvcIP9xJlyInlIS5K1xRTRb
OVDQr5C/EBvdasT7UTMaEZemKRHDp3awyyp/dt7woB8yixF7TkqePlPwc11lRnxP
vnZutzzK7Ad1UCffr8bxKnBNwHFCyLT7qfl2Ac1CJ0wYkb+NEdnKea7lCsR51JNi
LwPH1s/FdULFx/K5inRGkIpbj84YtWuN6tQWY09H3TgOwn8PL8yWX0j+eJMoqgWY
JqRVwtw3kg2GzRlyFxGcDyWuaTfw1+c8GyGrZPiw9ohUpSxkCHNd7D0iYtramS6C
A50vNTSDC8MayDFcxIarE4q/PjPFN+siK94cR1K0XiY2W2Mlhql7SrLbhOxGF4JQ
UCU02/pudMGUq5sUO828uJB9Jcq09g15/r5B+mPkKcpYyPurv8eHb80hfL6LyJn0
P7ct00PdgnFm86VoG5i/WE8DQpRK/UQzxsOln7FUEijimPwBw1qCJFzhN0U4mhhK
WKmu4edvPmJZAb2vf5c7CX7gpHMJ1gxrxFezhMcH15fg3l0a4zZqhpQs4Hk76faw
gMwWKQvrgXDdDc+nEaS2Lk+o38ULqLWMsb+MBTocK03Cb2+iSFLH2k7OXq0jEqIT
Je14JpVl63+Y2K2/xO8YVyEa7Zfiz792TeVJC4SPBkv7qdK6RIbwLN/0lUIHD0H7
oyD1wGaaXa3MfpWF56Zp7mcspzkeppYF4uAuFpOnFkgOkgDmdJktQfuMJa/K8VJF
dWzP7HndmplMuUfN703m47ShFXpelzyiRedbqtISNgq0EhUj3Bn5GwLB6LPrp4wZ
lr+rOil7RSz5IRZ9H4gUw2VeimRWv3Og7JoPbkGlaoic+UjQlQsXWktSLp95M44y
M7g1RJhDz55UClr2GaMIdfBxcIs2coZZJAkARJQs9C/sZp6PQ9DOobSBCemZqUhh
joPjP2vxqItngusLc74kCViauyWNLSSsjYZvcDItrMkmfE4X3USy5szyqiFjujUg
RWngGC83bdWmhq5pd08m9MDXxh/ueYdRcd2FxgBXItpZEjpdSa/uhxK5VrWODNSw
RJ3sDCbDUUhjyZWapghBoam0SYNG/33ffXb2RsBUZbFON1W8rof3RBPtLyIj8PhA
ZrIAyBNRDaiDCF6XOVxiFZD+8rIW4kS0agl6U8rLCBObNIA5M6BdxlrKlew5rhfT
v4/Y1OSbJ4uPlv2N66YUUfJYD+qVqoHBMYeDhuXlZVaRinnfgJeGczX0SP77xHPW
JXArdtZtEox3ct7e+9EjUXahRuu3IhByUZF5ZNpMX5JV/IfIjekFjebhqvO9cF2n
j3AkLrAJqLacQ8LSevz04Z1AxL7yryjgFfiHsQSgQ5z2DylMRT2MwIk2I7ADAvFq
BfhvEZX54hVyZ+7hUj+O0nxKWJYhyCVT1V1irHGUmAzr6d9H/0mwbEltV/XTx6r6
KdNkcCBeMe9IhfwSb3uBUNAnSuhr4Mczl16hL8yQp1IWpZ2OHHW0OVEYbY8BSOEB
k6ne4SDLd/jB4PlSzTomx4iTVNd/tLxmwDFuQcWc8S4NEOkPXLVfMg+ozUE/EMph
6Lp0W3b+E5oBEisnniKshBEP3SmV3EDIWkPRxlElXSH40TNMJonkHNw544pboL1l
J3JhDmiUBLFjoYCpZAfiflMdgv/bYLeXCsRtQnegp2E2U2uob3QZALyT9UQXtf00
5LXAQriYcU8UAdYena8hgEog2jn1x/BLqYeu6CU1HwKzsw70s9JUy6ZGezNCM1Jg
Nn254s2bf6o1cCqJvmIf9p+6c3k1gma5NuKorbtgCu5gWHppvCuXWO1kJZ5I4LGp
j+088xcKQCSl9oYiPJCmjbcuO00GcZhLXIR7MSzFn/1h6lNLYNfWevDV8yfanSpk
xSHS5YIyN/ji9+m+LUyF1aqVM/LqHl0XdKlZF76gW+2/9uU+gki4ckOe0kSKYfPr
GNdSjU5u4dwLLxQfJXVCKirEdKWPoSCxjw8KUxySjqGcFCa+mXfTFr1wPsxnG1Ip
WFCPg6hfIQ6Sy53PN2LUkM99GsBPpVwtIM8oHTmqcPCc8uZ4b3TS7C4k85ntKo1n
SWBqnbaJv3AnxfKOFLXOlPQZJidA+1CE3pGWwgcnjhxCAZGRNDKx/E2+bwkSMhek
0EkdtH52BREeTxVN3An9GNzrnqfoO7qhcW4/0iVg4J4a0ikq2pGNRxIEJ0x5vzr/
v1mO6x/c5kV5Jo3dDjFRRT/BJvonOfuP3AJyVVqly3c45iy+QtB8G2SD8FwOsfdP
ctg5fZhp4n7PChYamNIq4HhoE9jKYrbj7xGwGpiYE+Q+rwHvdtPgc9nb+w1HhEpD
1QAdYxS/gXJ9eATsQaXwXL50vZx9pCE8zY2THLrphTiT12DI1kFELOmIy3B9nq7O
aTO7douxdBicovPqny6AzCkec59OPt9ElogQFvkVouLMiC4DWBV9bKJtWXQfzjnS
gwdCdg0p32iIurTFGJP4oA9RrWLj84EeYGKbPfuLnQuAP8JUV3IiWrR4Ma/j5Est
NTl60Zkh01otJAe+JIxeGaKoHFXH66vbAuO+yMN73rhTO3uhtiBQ6h33kcDv/+DE
83JL2sCRvDFY0W0T4uU+16N1sNrVPTTSVBj6g+SxaGwjX7S/ncD2gWktRRaFRsHv
bx3LShUyIhRleP2WUq0cI8SDIt1eP4i/UEPOwpgs074xpGoupUBZzss+LWSj5H8n
boDfz0nF4Szj0uJ9dubk8ShdU9SqlfyMZH8hbYvBeWe6wG6F7L+IfvleC179K9Gw
p2JtMD0M1NDG2KJmo9zoOwfrRWuquG8zkdFPAtUArjp+M4INn5qrhDWJk45WHKhm
vkuVRivKX6kz0/AUanbT6Sv0ExImaz5EJcTvFCuYhyigfmlQ05V3iIrw7bs6028k
YJHDLNtSAlEZOoEbBeoo5eolSsa+xsJxOgDOXLgAqELVAoIsmnm9hiPNWNTvdzTv
3sUFkBrGSUR1LrbDqvFnQVTaTqTzL/u1xhnTRADti51zdHhwXpao/fH/oFZtpKlK
w2dsG9qmSLjl0AuSSn9bedzFO5w+nerb/icOzH3+OI/A1rpnDv7SzmNHotHCOcr3
69kPC6iL/AU8/q7uCi+tKueEKkZK+AtoymuCnLkE7MyEcSXgpjqyzM+UFeMOv2Cp
SavzaIs+3Kz49T4n4TODF5L/IDR4IwIdEl+ml+MC7yeoYLvNDLIXBuTngykJfS/6
f6Kqq22z0KyDSn2KG6ctIVhrCuISpWgEgiRNuh6T2F1ku2Jj8Qm2PG1uKwrsUi55
QqMMBxqkGCOb064a+cGxPxvGoSzMXRR+HPPpSMZDUvPULZ/aB6qy+mufb0fO0jLK
A8JYZfqOSrGCB5JG6hNa4Q8ub9oqtASCaIGoC5MY+ILddDT6+/M4FyPSM7Jfy98B
gLbJM3JRJzJVwrFjqtmKmSrslsJn3nmVIvji+npHrrycsRH5EZnlPoFTFfedGIwT
FMojGkAaMfJ9QEt/0fE8rCxJdxiBE5TwPI+K6kDpUci1KAJeToaooJhzeHqVLm2C
T6TSTliL1jjJS51MUWuS5Gtgc6khZzrWbUq/4XBDqw8c7iipBvUwM+PInIx+Dlip
jX8K9Qw5cOTRCJ23TTUiIvwN/ZBHDC4k8NjAykNXAOSpHLnRyAAzc9vL5p2evpDC
9WfrIXKH+DPY5CLEX7RAWopRT/+fVGPPuCclaEi1iUbpGWV3IkjInM1EJUbNj20w
3E0eLAQQ7Di/5GUOzmlLZajg0rIIq/gv7BHNoNMIKC36yDjDZl+s36ToGo+DFH4V
2vrL9CtFEREc8KClKq/TqCqOsqiO4kAQqHwOgnEVmKhvXRB5p006v0V8bX1+chNN
jH0hSRYp27Apv/oWTESXlsd8yZrwdH7CVTtHGv0qaOn9gDwQLsF2WsfqYX2+mr1J
WKvm1FhKJBV4jh7QKmUltOBFneCZ/6tmfh+C0ct0Uqy2P09SMJuvabACoDsITvsV
mNloUYDIZ0+HK3jMqmb6XDorq30jnv374qA0Pegp48f7UDdQsVrSRmlE+oDLhtbN
U/vlCnpp5w/FlzF2rq3vxLG7md3RTGooQBcy4elQddrUaLj4vb7ca0l8MuBBUDNM
0gH6BoQZ6GfZ2BsMIW0tN9ZjF8pMzXWJoTDQIeNsQn0sK2YMK8ypC/OqVHsAI1Nv
+qNZdDxbWOqp2/wavzfRtg6fQF8XqOXqGnub+uhSIejMpLAmZ1e1AkhxYsAEeGJR
eyMQjgZOvDDeoNQ4HndfSe01dBQr7eK1bCCryGdv2pScnMM+Yg8RuBkD777kZVFJ
gic7bzKu8Yi6objE40NQ1nJzjSGiKULYYwYvbmmb0KaUBvH/1r168qkDAu2C/N38
cQcfkZ5ppYLWmToy45nenxCw73FTDQBx8WSsLnXV3D1JKgh5BTyjBGDtmYpufyKi
C3cubmmFUusyKRyA0sdaHetfi8CR2T9rqZUq+bgIuS8oazN1XtvXBXBXaZXzuEBn
TmyvaSh4aHsybh+B4C8eZMsMIAc4Tti8231Uqhz6qQmDyOs50NHD1xnFXlgxpsk8
dG6Hm5HHF/ascsBP3ss1rTMb03CIZ6L4kDUn19wKiKeMMhY+ogFR13q0dtiY1wpu
1QjQxj+W1m6g/le/aif4JOsY7pelXgbmYhyTUw95seSkrN1d0CGb0ey5qL7OvwG/
ZkIuqEWip9tfi+PCV163xJt+cfqLSbNREzreb9GTFZnK278BW847ZplJlziYBJ+K
ejd+o/eqq42BJpMuCpb9RkQ1JtvKwTYcJYhO+FqJKE/tfzSpTiWB9JYahmFqoHR1
NnyOYOTCwZnnW7JL+j+haZM8ZWt47d0D03hdW0xOuHsiwW6sz4B/1T5lSFZn7RmW
0o8BEZnpicNIDoEQNYHfj7aOWtwF+citlEtrcwv+iFsRP3QRby8DFk7o8suXZpIo
hANcmEnId/KdilnbY+oHH8BAFeqkWZiH10jP+EeiMygINgVWBeYoAGD0vNS/7J5p
pm2OReSlHcXNRRPsLz1HGyLjSwXRO+teT99ZvA1dHM8XB/ggKro0Ye+LrL51SEaF
i8GU5WP1Ze5uMi94LNn/IjOsxcqkT9jdB6+3OE9W1CPBsXtqlElPtQNhhxcvgnvg
IIVnM+RgwCYw7g7Vml5R3KyLQp62hSGBPKhmrFmXUZA8KF0joaPj1f+GgijvEOUm
moYnwbbKumSLniPRkWvMIAAFqLl2icg7uauZxypfzGhZwpc9EvZqwKyTAWapLtQ2
gfXFRVwM6sjCWDEmWr5UDf/w6yIwk4d3ymC50dNugzn2FnjNB7ywPtdgEHvNtCdx
uy+EDA3D4uy6c6yxfNIS1wKJyxjvFC1eLsOLLKXgQWEBW4r/bmHcnmFPpVbkxRWU
EC2Lf7lHwguUuj2xlgzxDPgcB3AbgmKk2lftXUIfuTBFNMdYvddj5l5f/k2bj/QL
WM/uKJ+NlIWtGKlN45jRFeJpNWA7hlNp5dKKzyzMhp6OelLPChpOOhoXGX+D8/U+
3MRuCzNMsAGuqvsZf05ng7vsUPNIrK2HDXqvM1thZmp4tWs27+EUHpSIqHLQ/fh2
OU57X/CrUhPuuQUkRIDS2BZLdiro8v8A2CfjOTRZlZABg+Nrb7HcCa9JijVTW3J7
tqnKRWjSxfu2RjPWO0WZbFeK5VwngeNTSfZNt5dRq3V3jTEGrPQEcYSPaS5LSp+x
JJ8KuloAXD1+AkPCcxZ3rn9rdQr2hBOrjTfzWTF5zgRSX77G7KB5LJKreqxoLk/5
Jmjg1+3Z7JD5fySeWWUjuz7zvvyszOCuOvAjvrEyg8WIlilymO9gulI6vr5pYq/S
u9PWK2d6NuBtmQjIBaKYGPY5leHLvScz7pbOjsFFabo31bTVrCnIoK7+jV/WyNUH
x5vcGtdQGwjEGy3L+l4s2P3k/RY6/2QWQZdJO4pq4jT/KtGBBhgilSC+EJSQezzC
lOLP7naqyVRC6lWnftjOBKjHvPxZo9kNGRFqlzEKJzwvzOHXXJtCrPdikzT9QV6C
FNvlK0IqkbR6SfPc/RynPA1Zn0+pgcfxm1h+BbLdI5pDsk1OeYrzC6HfUsCabXpE
+BKISxerlsC5MuYUS2mrjpqOVEHSaRmKZReX9f6YyMIkYmlUQxi1dWLYtxJz/lZ8
gTYHaIygcO+5wos+XFsFfmmyVTY4xB1XHFPpkpQbhuBIpGZCuWfdXKWZ15m07qFM
Esm0sZNwcXLRs7Y4P//Uk4r+AbFH+0S1+BLYWnFroSYUXsKPkMjb2hl9G7Le7meh
Pb9X96+VV9LBaTqW1LlWtwpo2QQH8d17+JqTr67ydC9zx6Xq69K8w9JjI17tAK9j
5fQthS21VPGJNk1VcPZzmB1QHIZC1oWBLRWC4HcC3tz5Ppx4Yqrn6Y78pEUNgBTb
Lph11pzyJ9sbpC9bFSkJDiLXiUEWz39FgAzgNHCQjTmnfW7VeaQjq3U285c3d2V7
26iVlvYNqifOLefqqppAxcfRN6eaU1wyzFBhtxFgdf5aRYofVkW2PyFnUs7hltxs
sF+pPCtLIburt9M3+Cb+zjXFGKqfY4+KLRGbYwrBp77wXxXloZONhDRHNi51nERk
8Q7HqzLkLO6eLi8AFuVzcbuXCRdjAZqpZBrUvUp2we36hxrQJetI2lxWyF7Dl40M
ZO1rvkMRZ69kSZwlfwNLeMP4iSh/BYFG44pYMtmmH1l2A4xt/aRoLUq8df88ozpm
W8KmvECw9l8q6VvES4dvaQ4PSYAp6LG2DG3MMDTvUD4YLpc+My700r4FSZ9cBOZZ
OgVd5v9MZxjSUAmqU8ymJSTGz1TraW1vpxav8q9OsD64u5qCGkGWbJdZ7Sl0vwoR
J2lPjZeiZ8G8jgMd2Fk3ArjB/I4rDKPz7FshfvNNRbX6agTXRmvgu0kjrqi/mpIg
PqbeAgWBbQGk+DhytqnsMyPf2+3Knu+2omXXAYrhEKdns2RMUsr5hncE4eW4yC93
3ZQcFBZkyc+BiaJa/rTyjLJicf2CQjDymGc0oGKCLwRjlvsarHR3BI+d7mTfAPtM
zFLk2lJkHAhZkAevFHaAOMKhxqb5PfCVWKB+vmlmxZy3FnUItEE4BYRKmMHvor7X
R6PBWIwqiWJQaenVd9ndG5W7tPvcZAzjMw10VG935wCrVWy5Mvb7lUKpl/O+0vtR
I38/a+f0F8tB8OsHSIvGRlmPT6CSbV98B5xQavedFZNjF3b9ptGvsO2hndkk1VNd
cITqEIDJV0mkQ+idBl9Tw2JPfYSsfzljQvo9G2sH2nqcV0LcD160Uh2jjKvCgr+C
GrTMEztm5TBHsy8Bu1PplMTBaF5kU7AlGE1Bv/pMKDY5Amkd99ve4vjH6epQY5oI
6vdZdkWxfVHfUt3qUbeL5RcaFpTriVxNGfDJOD+oe2jUdoc5PL7/KPpMoZp9+Oeh
+eQST93hqqbaVZusbssSBc6gRZGTOskBKZMKeU8ZFNZJfeZZsvGrhIRMFsCc5MPE
epphYduYxgynI8l89v7ocCS+heGbRLVTpnVIYr8x3UAgbEgnF9Aj3OiBrHt+IniK
KtbLMsw0hyJWnmo+FQ2wZP5VOa52mBTXN4ei5s1xD63IR0Mq+hKgK99K34kM+XDE
5LiFB0kCSZ1i622PxxanDo01K2jGfnRt5D2rpAKTJqaPLU19K48v+VWgSWVNtfh2
Vxtbu3TJTfUyQM+PipYOu2ZiOi2dMD2rkQsYkNSL6Hz0NlUkO15ZD/0ykhSpQ40M
htsCe84KSXY0cD2tQzkRiqjDm2Ddvc2TlH9lXqmHYEu5F5ZRO+sGGai0655Lj4b9
o+aFxwkLxvmSmvF+B19YaA45fdyCoJ8srbb7jY9j8IjV7DhsHQL7Z/APIYzIBzBZ
SUpHTlrWBq/HMu2oNnh0lTgXZIvLMILEeoJEmwRJQ2TKhIWIu2SL996Zp+V0buZ/
Orhsv3ddVb7GZgLRTsLog/KJAgF0Q+ByxIek9T/Y3bIadlzSX4wSkRuSl9U1y2iI
+cM6AXCOq6R9xCI0JnwsXRHQS8z3z+znTjANe772aI6dMru/tr+R25kDkKDzwa3I
dYNLr+E+jGyd14i+nFvBiNMjggEsRgFD83OfcO9Fb6CpBbDvD4TtAkZq+oow58Oy
qwPoRd9z+2XqbrU/SbQFbi8zTsSgVEB1A/zOdTGle//73rOL1/V2xLJ5iv4accmi
gAO5oUSJnW2fwMW1n5XnhDmdAQjsdYW3Dc60KdlNt8VciihI8maAb9D2fEEB+K4W
Nz2KLonBERQqayWruq+2VlXnuoVC6TL3190YsCixH8XfcPtORt5iK0+803ger+/X
bFB8HTDEcvROmVwAhHs/MznoQ45EoANsmogPMebXLZ247SSQbZQV3+dOFKSaeDFs
jYWSjU/CuXVkilhrQgat5bo7uClyEnVHTlkl0Ss6mq7EcL7SH4NR9u3dix16PGaj
gdg6Rpbgi+aMnbTi4rm2EdMWli+hz3FKJQ9dMoti6hLKnFS394BI7JdOxEY1sbSe
rMpd4Ophm+bdj3XTuY/mrEyFCACerF9QmTEtOrUoSjQ/5VBzQJELHDdFI0sApaWY
aFpez3OoKheyZw1Q/9zNxzgLLx3znIqsjvPXCFG0hSFPg5q+Zk7lhYF0ACuaa37l
jwNGNfP4gSGRnSh4Js5Jj7UJRPijMEuyNJkPPJV/26ijVTmV0Yl5JNkakcqZiCin
vkt0wGIFnv6y2WMGQLSEeG6Vnm9Lm45Ti5FoV/SE2g4TjsoQPa3qJ7+DhGSZzYkN
bAzPrWZDKtDxGcWAGKPX3XV5TyIKu4+Ikar1KO3R4QvkGHrhoP+GndA5iwRc/d4Y
+RWjmk5rvB2IhyvIkT4mMaD2RuYHB+7eCzT5TRvc3z+F8Iq1VKFOdxChrzBTQwzP
RKqK/YOk4weuzqHDs1oDmFWm3A29TzmPT8ahn+g90AzHLVIjyuqg9uWVnCt4udIB
qmqzf5gXNaPHECwcAfLzZ4uTFF+e/07XqhEiN/4mTCS9UAkdFaDYlnkVsGfXWtkv
PcT4YQ8loWkPVWPQgWgOsxLZGE9SIEoQJnRNkVHGEIZ+00Qq+VSBwiluVOXPmXB+
dS8mrnZCxXOI4sXKkf5Kfqp2J1d4Eo6+BlbPhwV2yKftAKx1UK2DDEsPqxLPsBT/
VALQLl9e/9K0svDlOPtv9F0x2j2J7gJ7Qf5H/+wSloYdt0ucAYVkX4TJ9MBvX5Si
oug0nqSwf6xLoR2yFB1Lfg2AKLP2dEMaJW6QyerFvUr4HNUVKU9KhkjucudDN9/m
oY7BaCDYJXdRd/ei+XnfPQCnHO0Iq4aalJ1ctfONhWxqt8/3tG9pOf4bO9SZBFTi
6/G9sA3kI9n2TQ9wHipq6hTFVPX2QZSfshAxtjbVEoYMZ7Oi41Syk73Dars/A82o
EZNSxg198evfNo9KkwXOuwVzPqpWPoyIP++R5xL4SF5zI4YK4MPCpKWcVP2II7vb
LGam9t5Isv86nHOoeJqKOd6MSF0p7AgjnUkPz7pvHyEGfWyUBGFmiOe6Q2DXX+Ot
Sfe9AN51ePa1EuqGu61yepbvLJ294XdmweQdQ00K915FeoaBqLyXH/YXt5wUBDms
YMcwsVpoGrIP0TULuKh3eZ0qkYmUzIrsS9EAYpwL+0ECaIhR2tz4Owrxex58vQA6
b+BxfNDEY5mEM9LClz9FMwuFvliC/CnEkAGL6evRMKXYG6SgyFeJSB48nVOQ9a9N
wvwAD0PFHWROmqzGoTa4ekIfmsn96NQclu+YZxtbydvreGihdz9zp4FXFHUSLlOE
ibfoAcsLXfB+aQkIORlQKkpzuBx0Eu6SZtjRcxlinQXWRzjCmJ2N2TQjtt1YDQ+g
qDapAoldOsohir4xMDLn3WAuOeBcaGWWups8bBjJ+IT2wAvGlLZ7YBdqcVlZmGwX
NUhheQsFH3sJanAK8yxanopWhuxJHub7KFLzfpljFGqBKnG0f3p8WQD84Jebx/ih
hdXYvfRb+v/iFWK2cJb24exbV6ftKc4dAauTjJUVpEektY9s1gJcRYX8MnH5AopD
91CF2Ypqg4rqoEdoIfl5CsEMNULOo7xKCj9gCfGNf4AyPr0BvMRZY3QpWeSxDNjS
3b6ZWMd5vR6rddZ3UpdUU/FSfuiU/3qNY3yOAbCfafNKbKFbstcj8ENDoB4hRenr
f9Br4JNsL9AKUYqW4HVOq7rnLyR7IvGIqQxlIVMGKVdRNQtOK5mCFxjHbp4ro+V6
s07yRFYOb3fZszz2BTPy4hMRPm3rq/eoUGhjqYXWYykOKZiyNtg4gQpW44YVolme
I7MdOpMlRy1PzyhYTpXazTM2GFLZE5NO/iNW20+cSCtv3FWq1o9+pvqDX5E+Zajf
jrVoS694/bLAq1i+4BOaCNo1tYTI6p/lDE2cH2/HOelTYbBwaMswgmsRtJw1E1Ke
NeBaeM7eTy3czMepSC5Do4OpK6CFuNKj+NZTc5OTsFseyo8mgSUAitT9EJIamxCi
ZGAKgbq6T8GU5cJ9EdIZEXfYjNDAFsHOg4tmzSDWwB4UMTxnPs4d+RNbEKVhaFrd
thpBCCOk28wPOaUP52k75g953MRc/pGEhVSBh7hhv78oUC0C2iVxl9FPf9EqG7Q2
6BBtAJYBowofLv4KnwPR8A/VEm4a3f18MPUOxn4ygQAQsA3VPLEbBWAmxcEE7lDq
SRQpT+eRufnwdKiPylMY6w+Cb75lP/sTuP5ZafYaT037za5fQcyqpMdkanlQl9+Y
mlxfHJbROVBm+UAl+vEzN+JZT/fvWIkPhCuQL8cam437qhn5SL8PS/DvGZ+N4qNT
6izvzXiAb+OQppmlhdqCYY5W+2hn8ly3fO9uIbwIqd/E8KC+xF/AeATPeerujiIy
+vsx7l3hl18ThzpTpOafNofS5I0/ovdN0WTqFbD/uMRmY6l5AEXHkWRW+uloFW1B
eF7pD82PPoeI/iGZLT6JLZFMzCy3iFhfwP3MVVjO66vWP61ieppR5+PVZYRbJzhw
cS7Jn+0UPiK2bJYNzOB/Qu/IlULo7Pb+ZUv7Nyr1H7R+2404bceXCUUAROcZjiEf
eYbV3SzAhsoUWG+g4xY/R8uoPs4TPRq5aODa/Ra2P9olRRMBnq7SUF7y8NhglM6d
yfIkMgOQ1TC/J24oVKNXtvR9W9YeqNGQCmIPYn6lbeuVvzJjY9p2uzYEoBQ+Ixb4
qc/K8IuK8eN9Xbi/ZM4v3VQPvNLK3wZHb4b4WL6TN7w1fOUeL8IM0Gg2lIXtkIFm
K7PF1FHhdnb+kAvBSRDiAo9EuyKVGB2oaT9qAx+yjpYFRUytolbnkDxNIlUM0ps7
PXmYuqad+P9p8NFHXxaYdLFOjXG6NqI6O4tKJN+9/EyefU/vMvcUg3FxoeMn/jvf
bzFNsa0I4SujdhEpRmKm2zBAHfOh+Bl8R/RSw2BoHXcrAKx8ETjR14qk4eSYd4XR
Bv/G/BR5I7ujoLiC1BzQAkqyaebMZ3vcFW/hFH5+hyCATglUdiY69W62R48ffC+z
nHn9Ts4tn+0F0927n+tU/ZUQYumaOAOz2TX6RdKaBpQMtlkBvzBOs9ngrAogPB/g
PgpyfhlF4EpGEAhV76IoyRwBr8vZQIAELrr/AvfGO7KNznobwOcdzAhcbvWnJYeg
m8OnKFFvLKFKTfrlgQRGAKfP3jnjX7lTqFjoAVTGAAJiIQJ0drvA707KXFpJyq+O
nIimF4WhMnUkwDX9FJ6/k5XFXApjGTMUsyT/cXarIeLQvOB64rvyPGxESI0o2tvG
2aU+n9v/DKk6ybnnZmwMnEE6ETkXsnUin7tcVpu/5Uf2M1BWBZ8mTYSVoKz3vmjG
XihWY2qXH3FOqemvzuAksjN0hAwryzpC/Hb0n1O9Xp4kwtFMJk7LJ8ucrKbZJYoD
Fhkw4qgRpbLRpjtihBxJGGyhqwYUFqZXAGAU79RKsXyjZE27KppIJMWVsTU/5t/4
Gqm7pfp0F9VVLEvl1/WVlr5R+qt+4XZpFntXwEiAttAbyZcJ/Ay9WNzj9XCTaQRF
vJEEiu9t33Vz3R69i49gCgsCGXSiVRBl92RiPU6LJbzbjYHOBkadh+/fBgo/RU4I
FFx+MHYcAmR/lIIUSWHd8UOaxpBRLnSc9MEIM0MkUh3dWhR3MW0OlmmCe9CXKfkz
nTTiTs+cKGekt3MXQYjgSMj2AEVpR68rRcGscYcEi3qjDVM1/FhCkSzri9Xqxc3J
MaAo+79NimRSicYC8ol0rRUlzBtHldwkTuQnn282ArGAca8mFJETcZqxyRxJHO9B
PqfP3Ya5LuRSQ12YANWLeHrhOBHCS+hL5iGU/u0oFmHRXp1rSiBkG6MaJnPLwJy3
hDBhpLDwbzFveOsmvdSJcZxXYyOf/jmsvBlWq6lfrtbMC+EY4OJo+Xd2B1bPIL4g
yvj52xBh0ATGWdDhqK+7eJWckVHuPoS0tyTt01cVj6Eg3+qUrHYnU3eWJp5S45YY
eUiLiFY5nI94y4f++IoP60XcXHZBEzoaQ6RsjkvPP+3+V4Ez/zFFGwhRCPlEOW+d
98mBzqi/t6oy9vwN7v9gxIRUZF47UU/WToFZEikfVeLTJ3euNi7zYb+wKv9j01wB
Ge33yph5W4RO+jn7SD2Q70OpURNP8/K24OLy+QWrSx9xSOaYBSINWT3WgOJQKXLY
H1SI1dJFS7sdVQn9pGDlOO9Tk4Z7n+dPnw6pLDyixU3TyauVwqnOGHH9fY26IDqt
UKGf+v2gCdCqztQWzXU43DUircn4t8+BbxRxWCZMLqP3E/f+YRV9E7FSaCP9r7aG
bRb5KNgfzoWbCCNmJmDUAgduic3HVgzGMLrWkPB+L9pFW0LdbmlM9RAkse13Vnz+
MDmiZFlrygrcPDQSOk7vNMLFSDTxFg1xxvBlyT8zHU6JZ7ZM1xvHKaJYY/1jT1+q
tqWRVLBEnWJJSmsObRadWChicZFCsH3JZxttIvlWDyTpG7nNR7b88SFRmRbdGMPl
1mY7YkaVTwM65KrJSOmSmBwkEb9tjLFjw0/sYlIg0/NevVw/tcTXXiID8uqz5oQM
6zTdARpJ7K4cHEDrv3Zo6N1zR65cZMeWSdWxV8UsL9cuFtmmqL+p5PQFbr8ImSsP
TSQ4YFbauRgzqqAY0TMhyZYSS2iCq7Cxk1bNs6Czt1+dTub5CzkBGQv8zrW0a8VS
Hx6MyUUyv05irG7ZucDfquLmJVcD3ykr3uQS0g3pQXBpbwQaibN6U4DxIN63Q5f1
qRJbzQVPksWCZQ/vgIxBX+xrZD286aZC9dlCnGHuc+rUyucqtsxFEeiWOCCXZpCw
OoW7H1FDK5NYMGoX5mf1llKf29xOlWZdFvK46OMBhJmZiER5juyJW47EyyTkmjRH
aMzDKc5lAaqReNKdSG3+/8ppc0HW6CVKyabOHkhJeWg2QLDH1MKdhUGla05tuz7f
DMYIo3XzxRV6oO0j7rL9NwbEpLAahT6LzLBaY5EY4PRj4gsIH3idgw9DCRnZPeaN
kv1oGSn+remVPt5CzgAMxuIfwToNqe/Sc0tkpwZRIPl/xB2GKjequvhPofuKRYpr
mHrTcMfw6Pbn67o7L6ezEjIKi2fVWpG497IcSwZl/2rDaJgOxSV3Mqt1nBblih0l
A9NfwCbbN5kHc2/gNcx8YCRjtpemRkZb1q5To3GzDu08aVGN8kmkB/yowxL1CSGp
OVfbVhvWtceU1wXtZoerDWxylhk2b+paVZz02E0fULrgOoToKPrJ0YyNck6eB0lQ
uJPy9THM9RF+B8SP3PukcmuRc1qRCCpLarVcGPQZC7fGOu8zVlIvraomICX8fu8u
DMQn8G4OFx4XR9I9LCOg0zR6Gq1AnNp5vBckHWBe3tcV68O3G6RpfAgeSmy4Nyu4
XW/LpCGLNoDOeGczyBYCXaYnKw9cunHBnE+dscgayH2zgwznmnS0ePxXJhAHv+rK
630TlCEp/7E+UNf6i8/17hS5XuxO8ObQMYSxbHTKqLpZfmueMNIeTvzEpvpaIYLr
XNOwIyCNkdX0jGa2xbxOrl0Z7eHdHhPv5IQBE+UnJStq4JYrawVEX60n/ensuD7D
5OxciF5MlG7u4BdyJJGlYR2zCH+GNT5nRPbE5r46W1ecJDS/WT/aePpcyEKuMZuF
/7sFtYPgm5CKSRqJ8fsiZOrvssbuiA2PZ5is+LxY7wG9/MjoTRdLMsO+y9Njwxqn
yyOn+ddcRe7CP9GL3ELaCveMj2iNRefDDEYGKAknX1YpOor9M87HyBe8WKMbSo9K
4yLJfOdwx+nD2IzkbUVA29Ze4SnKc2saBsQcYE7VKta+0WIkWgnn6GMCHglVwLL4
elSe41FBXr6+bTmavF7cpkt86gL6SjGkHIW2O6LhwFtNxyPQW6PqxIRpxmvwuc9k
hEACMmGJgzb52zrDy1jNqGZBSJA9JwbdnJZ0HQuEor/ROH9YpbL9J4yyNDsCunfx
Jz+k8lZhqVg+B7A6qZRkcgWmd4xGOg2rL1Y/Axc64yhuBkvYksx8HDuJuj4kQ023
rSWP7Wzy6iC6LdJGYzrl9RkOep7RkqgDPaEW8eROgJBA17EsSqYFBdILLOHVbC+s
J6U28XqRX/M34rTtT7IQS3AXs7sUvkVYWONSIBz5ZKSt9eyPzsKdcOL42wGONqNx
H6gCtFXXniyK0yY7aJblyi7fqlcCjyAmM1381zaVQ4JTyisF7Y6tubnJ032hv6du
Y6JxL5LPYeK7OFHbf6vLCNrFSVn731d0sVZoJzQPGHEfQmK8LfItS+fsC7CDBjCS
6TNgm8MPZbjpkuK7nxVymM/8pFpoE+m91JfNPD3vfnkEuLDsC4BXHm5zO0ik8B5X
Gc1CNS13q69fHbt85EVmOqaB4z4XZlktJZB5ERdgi2ipMkOVh0cbZXg1P3r2AKEX
dp3ZZhgQ8Ha0yKlWj6rpjA==
`protect end_protected