`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
ddtXksX2+yylW5zu6QL2Lhnb2d1sD00763mmSITNX595NcHTEkwn0zB1Dry37fOW
FufOhVzEJp80NC5qZ/+F0Vk7Ik02dIR0elf3clrjeJRK85K4e3Hoo4xn7YbFUIms
l/8VZSb14+JVGURjfswrIyCUotIzlzVYZ6gzoZwDXIi5gQIBf/gI+KxNXPaKV+PQ
Ufys/12rjO6aI/pPlqSm0hCvftmBcnezN2hk1UeXgOIuKZnogjOsf0iJVX2aOOWE
6pD/psybjbnsNB6kH5uFTA5frkzIzkzl5d9+YDm9OyC+k84E83I/7/j+rk4L2dah
QJOvksSIzN867/4Qt8qYTQ==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="MvBXkzurAa5VTw+1JJ70nePUfoQXBvZOku/SMmg4TwQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
oRtzZL4VJ4iwysPsC8SXYCzXS8Fw2gtZTOskLcDV+1B9Nzn1zTyNtlo6lNICRmmK
ZRVu2BmCc2G+fmzynYlNTnSa7C0Cuel6FYpxCBlOuk3OF2tzAmLAuDyOH3Z1Yjzk
a0aHuoCdIRKv7BrZCdALt03JeUmXKPdOmIlkVGFl8yw=
`protect rights_digest_method = "sha256"
`protect end_toolblock="Jn9CQpRhJt4rnzZPRk+dOpzAubz7omckX1MrFd4p81o="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 3568 )
`protect data_block
gD6l00tciPUa6pDNTk/+t0OO0nC/UTtBwLB41d4inuAUA3i/ALrNyoJVcBnAmEQW
ptbcNp5fxEUJjnOxnedyZEuEBxWRieZFQnkRdF269oP3ss9Ge0d0UpCCrZ1w9x1i
zxWFI2bg3hUKbPMcwjhOuJQWWMjVIqf0to2ME1QU9hVYvVkt7sfpdjdI+FR6RRKI
hAxeIWnFrziF28oKoMR+qRUw4oGX31pBTd43LfjUZYtmd7NR/fBbg1+sH4mzHBCu
TQ2+LeG/Lx9A3v2FLxYQNa+jy+7eBipCOt+1ex0ZvVsDvL8Wb+JYNFM/PfWbtOh5
YKDLva1ErOnrFZZ1q6tgHpf4XfGHRWYkCq/Dh8FqKiWqLB8bcIZ5W7bzt1nqYzwK
Kgoo6S2KDzNpSTxS2LvdEMzhU3fJd7oS976u2Xz9QQYC1CMovJe8Za3fuNmO+2xs
ljYQXwwaSJd5FfBCnq8F4YWEpBZ6ycQx4szyEtINHhhTS3Kh/WZmTHhCNJ06HBYV
DpQBdSwBTBPpAykpKENB5LBIH1tfC8LfNV1TxSHlItcsfo2T8P+Wk29/XOxuKhLn
PVWGL2CJ7q9GRKN0fZc97YpBaKp2LjZg2wAc6RrQYZxM4m+0wksPYDYfKU/dJJTm
uUM+ore5j4Ds59gg24saIlBdd4LQ/qgNL05KVWOgA1pXafZVCGOV3tJsAr3GdxT+
HemlHfp38WX5kSM7bdkvp/lc1OAtLQFJuZQXI2VJO9scNbVv7ui3TINh2aReV97e
AMpOm9imQdQQlx1RzsFCzvVNDkLELmJB2LaZx9tNJYpW46l0JA8z8cDfhlQO6ScK
KlO9EHgWO5wNj+IoZOCIoqUzIGLa4IqGiyiQuG0QUdDlZBf6GiEl1I0BRIR97vSF
L0Vby92GACIW2RwhVyjX9dyscM0sJBtp9KO3J/6JA/4iLLeZ8K2ahKqjy/REC9Ig
rGizlCD+9eMJkkO5XkoHnv3s/rYapotsuTW9lZ05x3LtlbW5yBk/996b5JxURzlS
1E8vuM9gukGDB6DZ4cqkenmxDHN2HSCK6SP5ST1OKsFhYR8ycmy8h8dIJhQ7lBSi
zjrrMvzQlOSy+U2qpoVGwL9+kY0HZ72vtayM9NZfYZkA4siDiWGIBUYeIzCOuwfH
W+G/JlSqIkHakABbTqw4js13/b+zSCVEkMhGp4Majk0eQDvwPCaRjIwAzAcsZZlR
PFjnwS6+ZYMBWPTT/7anbhuTYoYRSkljpJDhwRSJxK15K3Lf3PD4cVIh0mlsyYyh
i4cd0oPVsLO0K0MvwLJgrOBCWfgwN92lL2Xuy4adNTJ7t7pyPALKqBiCp8bnkEAu
suA9TnoDrz0wyeZA7+oQlCSudJFtcsvEZLuIpaNWWVEfLrrPwgJWRec7r+REvu1w
mSyl9LvjxJGv/2z1ElRSjKdBAhrrTZxQJLkzgfopfv2okCiS29aNwPurAkZu1T/S
6TVEuSMLg/QY3DQTSeiSpFe4lDJxg8+6xFjunIsWvlvC6J9THWe8kfH8YpSCvcyO
EIvWFU9V0YH+mjumh6f0A8MVIwPNJnNhJiX69HLNSD7Rvu6HdrZ1XM/hsbZO9ySW
vR99nhCTbZw01PlTPQ+Kz3x3D4AHlzVz/tKs/qLrXVlWxtuAR/1hey6cWfgp/er5
EjaIuWF3SUSXAD4QMYBTwnFAMc9c1W9p/JPf08P2IawqaPttfCaGkhe+Ks3YXXyY
NeXnfj/7dTMBkslTykND5OPLDU0wvhAUo23WlBBmAkkgDZsg/8EbLiOfD6BM2W9Y
o4teDmlzaJ4+uxzPRa2IE8KAIT+Wg+nss4WQ41QKK60yAVnsG3QyaoDHj5mHhPPj
WvgXVH4L8BtnkFLStdf0WHO5D+OSLgBWq6iM5gsAEAseW5nMjfK/bSkfc2oZIM0L
0cro9+Y2uPnqBlBpeaJ/AJjsiJvEm97ETbsVc1Z4hn0Jw3F5TZwR1T6mc5BcTODQ
PNNMcuEzlWHDnUH5ADVnO24WRZmqgSEeqmPOCZ1/E6WoZyUADH7mXIRgid+8BTMg
iHISepd9oQ8wNuvEGHF8Y6mqitusalb17qpmM0NPshnQNyoTuRe2hFevCxVbL6RS
weff0bIUsapX7/IZa+ljgOUri6C+j9fHo+M4UFOhIDUoYHatwdGjWzBpiCrBM8CB
ru2jItYVJYw5alkc111iwkU7Xpu7Nr6BmYIi2aIb+DVM4WvqileXMHMHe+OVsxP5
clmMnXtbbVM4a9Pdb8blel3ZKp5CDp4LCJCoEFqWvPz9/hbTMniIgKFOeZk6yd3p
rj7pqWPi/fiL/oMShhGX9+Z++zTwrQzsnHClNyLhMmrxvZ9ys5qNJHbV7/X3KdnR
It5/dt4BsT56Im8a2BrFCP2HQo142A8mhA3UP0DYv0noIKaHbDRxjZ4AFZea5OeN
QTaFAKAIoPX64zK31OBdkxGm7C7juMA4Qy6X/vKZB9F0NfdTjhEF5ab3WCkdo1Km
MavDFyLXkrsUmNMXrbcqHdTkmwez/F3HAOTUwCJavatr54dWXShZ0+2NsOa4MM6r
RN1pKBenUxEF29sc9CWwir1Dc21Xjq5kCioV28KnVrTV1TFT0y5U+0z1Bkv7N3/m
YaQeQXMswyvU89j4n9xIit9mZHrcIqUzUUwHnN5SDbZHilDdCzKNVeRhPWtLcVgl
1dZBtTnyPpiFnjXDF2ZROhRbPLRPMsZgIQu2O1SijrRVtiCqTSs0TvDhMZIChsb0
OCbEHgSGr7JxTziQzFarCmnnRowMp3dXCXRw1zk3qik259+nFKiNFZafz2Oo9LRL
PvqWkiaXgoOcdtyeP8BhtTaXMI3bSn/CYTx0QuCJQ/vixtlBrLcvBUjHgp34Yid9
+TY0M985H82lmL91Y3QKgmozyFV5tXiuv71+iMg2YtikeVvyTTUu7+4UTHDm4oJl
rLypjQbKdDt4Fw4knX6hSH6aD/FX9cOIFArDsjTrxVyHEsLQZbeVdyPvAWTpP3km
gPKvO6unlElYQxZg4Ca+0tBvN+A1LHmlDekp1++lOVk1yj/jtqbMqpFW011IK8U1
jFeU+r8xjYVrMlfWhFR/je47biIsXXSCETtUhDq/oEleSCiErSMgh6c62Srxg5s6
b6MtTc8xeuP19OgyslDRJtwy4wgcAgtYWuGKZhq6tZX3hTP4iLmr/6N9lt1MaUiy
X49uxOPfjzeWGn2pZSCxS58jhqgg7a1A0SFCMdUZ7C6I9kSOpt76OE/NO7baxpUk
Q03uv0u7X4opjaw2xqCkDA2RFtStABMBiUUpREoM6RkG8wRj+vsJCqC+hSJS/os0
wnQLjLspDLOdSggLP1jL1Vmj+PZImppz3auj/UiE3taYL7Joi38MKPoulNbrjiHA
II+lI4aEMm4zWLeXmo4vZgdrr47fOjsRzZwSOBU4xJAFQXWqNX4U/5lndazpCxNl
I00OxFhn7KPF0SyTC9bJul2OQoiyrwjMUj57q9C2cFH9DvgrozQp7bKP3zuxWOBv
7RGXu+N0foFPQONWB73ztyYDYNnt7Gh5XE6os1w9gHLUQhq6RYppA8mH1dbndNIy
mrZjuPob/jThjjkMoQq2jnk5aX89XW7TUBmqCHsLfhpxOfjCwhnTNpozJjaRx+f7
I3FG4KM/bveRTrO7HjhUTFF9szW3d3ZwmxiWkqs5bIkoQEBcMmlgUu0Vpn4WTx8z
1GP5EUGOae/9tVU4SXnVGzKDQOdTzwmLlSWCgtlHRyLi1Ew2pvwiTmD1bME+uioy
PWjRP4ViECsR7+enbomGow+C8i6q9GsZRqxu+BBUxm3SmwfwYSQgMMEHx/HWJU8C
LZi/HVLHXXD1au68I/oRyOwBuHsjifanpGVUujDdnz7BHoN56CEpic8lFpg8EUOJ
ahRclsG8uu1XCz8KfX6ii+vVynEcc5geTtxYhIAtmVxMdo90XG9NAAgrCLQMbtwh
/tLS1a/47z3D5xcXhItD/N4JxXerrDMhUF8Cmn39YAApMV7eitEPzoaMfwv3sL2n
u0NK/VXUt8fsCcBKYzFU1jvHEuHfvbA1oOcLQElA3S7RMyNX6wbAfOh2UbG7CD2D
djoCKK/Z7fKEr/P+ZK63IuL6W0AIcEMqYPAig93bqAgh0MWpOMww5ias74EEGpre
PQGXvKYkAx+dMZsBIahJ3/wUawrGNmfcKCFgrfsw+P5j0nq0q5qED1oMx6M7BsxA
WSp+KSHR1tI6glbsAgQQ7V3cuNhXjO9yYna9mXhGrixbQnrGApCBkjr338TbV4tI
qT99tsFIa+2KiV+V9bWai8yRFkpxCxqVeqCa7psHIrEMuBsoIuPSgb1uRhvFxumS
XD6AaWLWX/51IHaQ6x0XzroHrQe/gItuZqO/JcQzpQS8WbHCQbVe3J4obx1wlmz8
ePoK4or94rAs/InSGS1YDZBEdsjJgkMi7l4oTJzmY9cQxs/OYbWWsWaV1agbkBKC
uLHkYi1cOfnqJ+5jAjKpmD7PnDrBy8m3d+mAPQWGwFIDWYxKzUTj25m3o+uQ0diy
e6SY8km51IQBpZtUpwb/5YJxxaVkiusdeyjEgPmwPdbgtLJ7E9NtBgnDe3lv2fz9
7RqsPC/o3CYpjXosYycmi2H7Nu+TqparO3+tAbTkNXs5xyOoovyXVyu9L2Jsl+Ow
OIfKaWs3bVq3QYp50fEwUoSDsVFaaxXld8lYzIbxhITGb8BkaigTAvJYGdxTpnkw
bcRPPgHTdQ4XzJGp33dkoA==
`protect end_protected