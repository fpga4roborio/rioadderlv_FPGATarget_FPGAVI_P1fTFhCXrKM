`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
ddtXksX2+yylW5zu6QL2Lhnb2d1sD00763mmSITNX595NcHTEkwn0zB1Dry37fOW
FufOhVzEJp80NC5qZ/+F0Vk7Ik02dIR0elf3clrjeJRK85K4e3Hoo4xn7YbFUIms
l/8VZSb14+JVGURjfswrIyCUotIzlzVYZ6gzoZwDXIi5gQIBf/gI+KxNXPaKV+PQ
Ufys/12rjO6aI/pPlqSm0hCvftmBcnezN2hk1UeXgOIuKZnogjOsf0iJVX2aOOWE
6pD/psybjbnsNB6kH5uFTA5frkzIzkzl5d9+YDm9OyC+k84E83I/7/j+rk4L2dah
QJOvksSIzN867/4Qt8qYTQ==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="MvBXkzurAa5VTw+1JJ70nePUfoQXBvZOku/SMmg4TwQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
oRtzZL4VJ4iwysPsC8SXYCzXS8Fw2gtZTOskLcDV+1B9Nzn1zTyNtlo6lNICRmmK
ZRVu2BmCc2G+fmzynYlNTnSa7C0Cuel6FYpxCBlOuk3OF2tzAmLAuDyOH3Z1Yjzk
a0aHuoCdIRKv7BrZCdALt03JeUmXKPdOmIlkVGFl8yw=
`protect rights_digest_method = "sha256"
`protect end_toolblock="Jn9CQpRhJt4rnzZPRk+dOpzAubz7omckX1MrFd4p81o="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 4848 )
`protect data_block
gD6l00tciPUa6pDNTk/+t0OO0nC/UTtBwLB41d4inuAUA3i/ALrNyoJVcBnAmEQW
ptbcNp5fxEUJjnOxnedyZEuEBxWRieZFQnkRdF269oMwTuGaF1FOkQhMxk9TrAQS
QJm3yoAcIWtPhmFpCDb1iZDcqooIPPA01rUtzQOhrA5Ztdq3VvEdmDd7IJaJQEXD
8fZSSqFH9Jf+KkwcaWJoNthPGRjol6pUUNx9MV8W0jF9m49Dr154Z+seVgrmtwAb
mS38xkpZF/Q6f0x/tCimrHKCWR4DKoVwxJLMXtw+V13mILudgo0u/eFGgUN3/Eyg
2BlAUCLLrcBLStNj7ZkuM+SUatbsZyxWH0T+XxOVJfRBAicpNp6wIFM3qzNKrOLK
yMWxVMTxTgjzpLbDmJlrJ2NY4Oil7gJg6s0+WJuVmrmC0x4RJGgNOAhjaLghxtdI
LTLcno9f7xZK7rWV0Ng7e8kwUUpBvkumjMU3uKyfKV6vCKtHr6NddfUo7Lxbh98t
RsFdkC3BtoFSUrGpH/+rIT4jW6wj4ORM4ardmmo2NnKnlSw+FSGlVC8RftxaKU4m
P+vlNP3yT7sMcY8/t1ksuDdGzTz6sbOEEJqR1hoqJThMYr6ep7aYRUgvBm+YlOho
AKWUZVmAHpPyyOeqZBSbegAOT7mqo8exX+sDIHSdV4/fGUiFEwhp3bvTo5q3yOTg
iBwbjrgNRBd+CUiZycdWpP1hbS1SlzBH13m9zcPsBBpYespu2hSbvQt3aQJLas9k
wR2zPuzKVGZRqpPh9JG/j3GvM+F8LsosuU5Lz8i/CsPMspCrClUsVgxm9k1cYxdH
3qSSXTnkgGgJlXRupv77DukXZBbRl7MOZwaPYg/MOPtmzN/FOVfGjrOjtVDlyNFO
nHvbGMAHsNMCy/G0W0CRcgNif+p1tTFq8gwwu1VNHqDQn6zLpozFcMD8i8xrQxP/
XJD0j//JhHcT0rkyrchzi7khzz0JpvE3I7TeFGcAipB5vV8mA4Y9YlyKHC39BdZ2
qVKrXrQHVNn6qQAS1Ek+qiH9aLqD62ImbBC/lo9tMZH7hIcChKMHRE1aEwUMC8oi
lzf/lNT/D6jJSZWL99Gl8XMWyqzvyHt5kNZ3R5uUQq2n5MpkCgMBwBhm4wZkeKD/
0CBIDBO0TjeX/mXCCKoTkVLhXgmuSS2FRHknGYy/cIQJeIHoJaXie0jMTSwjtxet
3nbxYHX3bn9v7FV1z2sH/9EP8AC6pRBEMUBDsScWu3nX55m1Dc4q+IOCXRBGjfmK
B2f0V93eB3wmk7iGcQx0eXntja/VS8CffrHNiU3kKaY8BzeE9Nn2E5KNKSbuvaaM
vyc5rYueHpkR5ay9YdsFUTB4uBxlLxe92QUwuqelwjP0qdsxQtTaHi4Vu7qQpxnR
7f3XapuearxnIAHDe3cCysOsgQsHVAMaGaSkr+tHbblKGJ2gc1XIpU1uArmXV06L
XdQzKUrLUBYQP/R25FIfrMrbmCXCKLsX/6iHsYxzfw6zlidpGJl7scfk8Vaoaqjx
p2Sni/Ddb23a5XiOCW94DIz9iJhiSpl1hRaYUPS0B2L7qxWYV1X32kBWwHYJM7tj
vNBho0znvcYSsd25VrsPUZcNiGM6w5NI75NkMOT74fi2E7Q98iJ6YVgpUWhuyHwf
EcUq4XSsIZ7bJ9Dj0zbGqGVMFG5Bfge5UVGABEvRTeBm5rkB1bi99ZApQ6tcnNuL
TvmcRo22JH0pjHoCCbNnevT0u0WasTdNmHwL7GlzMEzP9oyg7szvM56zlhMoUvd8
903l6aqtN0UOEF6+l32ilHX9hCpFmKwn0OMtB8N3OW2Nxv81+4YuuXnGwvMf3FBi
eiBD1YisvHNP3RtPOLQrzHK4vgHaJiU57IQcRn/mlQbnlFumIr1gLSdjt2W/4nm1
OCGHI3E7ykwd3oNgCA80oJlHbGil2R19c6+ydDxtQZ/6HUWcnILBXxvLa4Ldrflj
4sxTskRfPNyRyUnqj22S0EHeYtnTRZPZb+4UUxtPE46kIA348u9A9ERXUzN/lLNg
n/XLpg8cGRgsFFHWlOETbeNmZlvGuYapb0cXZAFRQO1td9Op6ERyZ9pzYpsSlfTf
l/hI8nOG4W0Cataf73d0hDd56ZWZULzKvzWzGtuVs7Jyw0/8prtNyprihiPNWsgq
aBkqUYZKOhAUovDKUKF7WBSEoNKHIQqvKUtl9bOyzkGRx+EnU6FOZGJ59N9a4f2m
zZdXnX06dWuBVH4oD6B50feNSlifsPAorihpwY2QcxwpgTfwp1SNJ/efpzELKjqD
JRvoSWZYthCXG/16epL/4GporCiqxl9yXQA8foAMzfglL10HHKoblyNGLgR6xyad
Y54jG0lEWvaHJc3+jk4dF/j0kEgZYrybHjEmqOGRmsiICu/A0bILoEONu5QvC3w2
yYgrQDga7YzTvTAekBrF1o66TxWYe5ZjWIScD/PRMfOTMgxKWOGG7gDO8bvxQ+b7
nMEUGpY05L4CGbVF8EDOl4M4NaZZ5SlRRtg/0ef8UM0Iw7PbgpxNpOntQma9X3tw
MFod9ZiFl3USO5XkZl274MoKm+cKUB+HjC1LTM8acllrMsVEHbr6ocELN3nksa+6
lBCqDGKlbndlFFBMlLU9b1HP7qcNIlG1Sw8yo0fHiOUnQ3Dn/2mAUC/rygVMvwPm
T1+F9tvra5vFW3g/RYLYHpW6z2hwsD4PeKek9yO+5sucGpxfwfPm73mMARB0d9Z7
ar1JoIuN/OU0xQHYkULcd9IQDwrxmJv6bvrH6pZX8bXZfVnNCIHOOuiesctR2IOj
vmfLUBH5iCygaqrJEi4AFGB+Gac6l1rndCV9qF6KAXxcqJIsBAtRJPxe08rI9Nmo
qR0h5pbb0l+kB74GvKxE7qutHeq3URSYISmfGT5d3hjBySFgdXrgYviaTLpYZoh5
diWFxgVyt7tSCFW3b+M3OfX5r2rQXB+7m65WDr8WRiG9HP2eISYFg1Qu4BQj3FNT
6uAMat4o+lBKCXXfZy2JecO6jv5ObhZt5YHcbJ5fJY5Hqxk4y9cmvWj+ZoOTfNL1
HvcWkQpRafCEMG/AOGtNbblVh2VG+yTjBwQpOXOq6sLdcxJVn6HVcnmE2wDmTwxE
ntxu/xc8BgpEL5g36rJM9BEClGrHeahCJ/QpkGR2jGaQFVXB+M5JBelcWfUnt1+o
Vm1NwT8Sqiuchh4JI0qjY9G2cTIOXnfJKUvOI+iWMOTxHs79rMgwOhEYau/vHnXO
jpsW7NmXPF6tGaYgOM8jtbu5xs5jmApAgy+a8oYqGSQ8NLbivOliHYfae50hxCg9
Wlxda5o9tp2SAzyojQljJMJGI8lxGv2GyjWMnd6wPTt6XdxpEvaakotE4FLbIkux
ud8ELQzJI534NiUbPAB3m9oeBg7nTBItxCXHx7agb3vy0EblO3siw4B+hZ2dTU/o
eqSX8wOc9luIac5kFt5VFPlsGYWIae+Yt4O9ASGr+rBkxdlkBK8zgS0HZX7++uqn
j9i6ipvAKhjEHt0vm6sx7GXiO2KxB+77avTKmZi5Yk2lzyTcE3GvutC8r2Px/UNU
T91mUk2fwfNJ3Ak0oX9HPqyokJypB8wsNQsIMn9G0gZljtdg88WxjblnzSyjbeu4
E7/m7NXo44KC4mfEeivuJtViileD7+6Ws3GWowPKN4vYAz/1J/KlPcQJ7iWCJxkq
fp/IEN+ipmqbNNgjoU3N28kK//we7JAONjdRu7zNX1OXMt6paz9NRjo8Xq62P3Av
LKrTzNJCfibwdBpODmCiXBBxdsecXAVEiQFfSr+4DTgZG/x1loMBhtKAjjBWr5kt
mzT03KbsiB84JRFSnHE2fqp+NM9pGQTCEUgyt/E4B88X2wYvzdfYE3imfa88hviU
HOYOTe8+lSqKS7LmwEmAC9ykmTvojPfDybI1qQFNCHQ4RORXtSHdTnBe2s/EUwSK
33M4FRnHhWNyTSFUyVGeib5V1PgSEH+q/SiEpDiX+sPuQDW17uJZavsl3r/7kWSR
FSFoA+2XH6/STmQM0dbqm5MM8fqffn2wZAEiyc9PCF+sAA8VYYy8K9pvLWzerKhM
vDnFSQ3x57tHNMr7VWhIXpNO+3FJ/vHcV7GiTQIFCsiSeE3UGsDyQ5citi4Zqb/O
93Z1RpLhPlsgAqfUyaHyDQo4xDvdP9RWWU2Z5BGfgYM8z+8gWHbaUsLmYHlFKAzm
gSu8/zHJaqub1anqGrbfsMdSFZlLdyV/7rJfO6qSvJ9v1uA4wemn7lBg+dQLe0Du
QPflO5G10KflfwnM7qkHSMl9BHx+lMTTzwN8/lX8cQLO5XtaGtArVbxn7nAYPUqf
87goy/6oFOUcOZxF6usBLUc4maws7XMIkxBpodBMdxp1w/fp0ByKglTrPkCLkYrD
HIu9SVVMyUj01poCf7Uny/khUxhMVpJtjtaoIN40VY/Xi+Blvbiz7wlp8mGjXk66
yRQWXIHS59LkKUiyVN9YJdhh3YPX7awFo/5EtTyE13EfKCGTq7ihgJpFrY1TD4yp
LBXNZ6E5l9f0Gll4KjSu+vuzzC6XbS8qLj4un/o5BkMt1asidE+HnDlGMY6dKhkH
srVnSwMTpU+036wGryOIyk6387GNkJlNjN7u0c2SbU+jWwMgJsQWRRyLpbMPEBbx
YgCFTHvlQcQetqEqZsHv5B1ZaNF5Z3rfxUENwte09JL4uq6hvolG6jzEEmyeya59
FrCwx3jSPxllVfhMwZ1GjgYoTqYVuL30nPfQxSgcXCwDedNFxJS8FaLr7bj9tYIS
MRtymyd+Qe+ZPAU+N1SZkSPke47Olx6Ko4sgH70elPCUrE6FvC/R7ThgJ6DBOTkX
Jb4s0BqjiW77w8ouKXXDZ+idXCa3i4gzOfNovX6cbhH99RjzUvKrhrLqgapW7YFU
bYytVhPInp1vQY6heu9PMP6w9V1W1Cz0WkK6cK93NeQZl9VytkTSH91Dafhosh6W
7synmGa1rZiycYbgSYEDNUL8Er/0tOLfHurLqo9HcDpvsBFd74JsmpkyHhZGMERu
ytmPj4QRtWQXilYMc2Rm95U4Ss22YJdqviFOzHPlA+HUnYJjUL6J/kDx3EqK3sRW
CoH5Cex11Ggr5t127Odx4l+NNWb5/F8fyurMk/mrL+TcQwTzEIeEY3VJoD92p760
ijJQwzndwQj11lp6Ll8kbwL2wDJNvzArFX3vKHi6b6lXHBlPGYpbMs84zkzbVoIh
3x3BsZE6vSSsw34/Sj4xly9CfXFyagMYZ/+1CB/C7M+zZ2p0Rfb9EdpNA2Mhdj33
xhVGVUH5zFaKpkvN6Iz2ZFLQoLlLC/V/7pNVt3t02Zj+rZRUd+2Q/ndJxhdAhX+X
tmoONQURw8T695KI97E3HwpVEmKho1KebJW5xMpQXwvLMq/0eOo2ieRyon/mjb0O
0CgOheU/bbKSYYxoixV09y5xKZZ7DmA/HlDzUagdC5WD09IW+dtkXszmlVOeV7qE
IhZa1QFTY7/qSEkgB2hec29AG4VVSX5mza6jWrpSLOKeHsTVdgsmsXRQbAlrybIa
2hh56JXB0CPd+aQ8qDZVm8jO4KjVOv4lOHGMKq7OfNgONv4jJiiF04/9G12s3OIB
XoHi9XSOpZlP3Q1pgfvmXY0ho5pJpmfbArs1igjpHQNekQv6sCOf17Qgyix0Q0fQ
Kbp20/Vazw2l0tKwMoEPVnnHnFX56CFxdsWK1EHGTZfyC4U/B4UmLTSqpt0x2zTa
ny+cY/TDPX8h3MB8iSyW/ITupXLRbRYzuVkn+SgsJoG/dz7N2jC1Ur4klMPuugZi
2aL1LRHUCDDv6YiQ6GhNhgU1hS3T47yZYCvtKRBuxb23rjm4tDbSLU14DfZpRUBq
h6ldFhE0m863IMCY9SikBT05Y8GdDo8HO/YWBIDyc1ROjpueuIm43lv6WK6mbr9z
VajAa2wN/xyM60II3d0pDFiX3ndUmwTk4Rr28RcKLOQzJob5kfgm3agSBC+Upw/e
HZr86IPtuXjQLVuPNgM7GXLoMZgSMNY+ClnK0AwWjxletxsuJmX1wJ064mhYC6VD
/YbcdFV4KSTKvc9QrxG4cD7WZZiaNNWr3DFLTDrDYBDniOkDGZngH3c86SV4+XiU
Ul5Haw8qi7ZCYXKWSjaZJX2j8Ji6i+dBmHqI066Y/wEGGhdQBskOD/+FWz/Csues
xlA9wsfCcHNcjIvM/avlR9Sbpag46qowLjWeyVVB9dWNvBp9SLSSLuv98RWxDQOo
Wn+I9giAxZzyjzAV5pvcEHZx43zMKEgb8VXdThqHlrZSFLdV9H1l1inivpzqAYbQ
NkE1Fi3cgB+4l35E2IZCQEqhzFLD/XdPKFgKivDRj4CSOp3cwxQX8THS27h0ex9C
SBBDbPgx3MJo99/3fDO7nqP/U3OZsDkfGfFx0Ir633fDDZ9FrHYQOaNhv60qKRg6
`protect end_protected