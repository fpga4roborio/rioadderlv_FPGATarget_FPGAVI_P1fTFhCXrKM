`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
ddtXksX2+yylW5zu6QL2Lhnb2d1sD00763mmSITNX595NcHTEkwn0zB1Dry37fOW
FufOhVzEJp80NC5qZ/+F0Vk7Ik02dIR0elf3clrjeJRK85K4e3Hoo4xn7YbFUIms
l/8VZSb14+JVGURjfswrIyCUotIzlzVYZ6gzoZwDXIi5gQIBf/gI+KxNXPaKV+PQ
Ufys/12rjO6aI/pPlqSm0hCvftmBcnezN2hk1UeXgOIuKZnogjOsf0iJVX2aOOWE
6pD/psybjbnsNB6kH5uFTA5frkzIzkzl5d9+YDm9OyC+k84E83I/7/j+rk4L2dah
QJOvksSIzN867/4Qt8qYTQ==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="MvBXkzurAa5VTw+1JJ70nePUfoQXBvZOku/SMmg4TwQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
oRtzZL4VJ4iwysPsC8SXYCzXS8Fw2gtZTOskLcDV+1B9Nzn1zTyNtlo6lNICRmmK
ZRVu2BmCc2G+fmzynYlNTnSa7C0Cuel6FYpxCBlOuk3OF2tzAmLAuDyOH3Z1Yjzk
a0aHuoCdIRKv7BrZCdALt03JeUmXKPdOmIlkVGFl8yw=
`protect rights_digest_method = "sha256"
`protect end_toolblock="Jn9CQpRhJt4rnzZPRk+dOpzAubz7omckX1MrFd4p81o="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 24368 )
`protect data_block
gD6l00tciPUa6pDNTk/+t0OO0nC/UTtBwLB41d4inuAUA3i/ALrNyoJVcBnAmEQW
ptbcNp5fxEUJjnOxnedyZEuEBxWRieZFQnkRdF269oNXCg5HRUd4JWF3ZKNjgvfH
kKCgbaWhxt6fewypYuyz32Q696quc25u0pEyslQvck+yrGb4fiM0ytFQarlXpbvq
NCutpz7II2T5zdUUCACbuaMSOtdMwS+fQcQp2ujca6CO9rYrchTKpWlPlWnAGrT5
nUiVnmKPPjMohgrq9TmPPBvCH/ToBUy/+sgSvcu5NQJJN+Yb0/0ns2mfE9uEhdaa
+4yM50r8Z7vOGGrAThXKdqWkHwrfneAj7uNIYhtlSNTgG7U7S+KYM6jjOHDTfI4g
llQ7WC9vzLPQ0IHqyEY9lDK5NbT12GdsKXOhOJYve98i6eQM6mAAbxw9DQwY8bgx
Z4dp6/GnMEW5pTRzIyEtB8tHRdUQPeRHlPmo/kzzkayFXOhpr+IDv+0eExDQt2CC
nYWNbjDsqYFNyPrPXmElb94DPZUTNSCDYmGog/8gXKyoWuLkbReYoci65f3hIaKW
TvCZGbxBY3p4Ozc4dRRBQtM1OmcRJdwYEPnKuURyP7EfLylxlOZ1/rxueJ9ZYto5
WnfsAO8JXnYiyZXqrtx2ENZveoW3wUI6yciPF37sMp1wDPsE0Dsmdy7ma34D34cW
dhqMKkq465e2Bn+DSa2+jfviSI78v3Dso9BPCaFCqL92qoRF0iQPwQWdgVJvlro+
zcrsd7dR1dzqBP2VfdISjbfoj/jxQS5c8vSZ3DYInlh/awyxbFik4uRadjJ8YeCT
B6N51ElxRzsiH405VUTe6NWPhokdPZaibCs+IZ008eYeadD5lkQIUsRz2+kuLIzf
R3Cf5GVlMd7uft63SJAx4Z9GjkqRf9P/ueE8JHNJzgL/tSW5/g2dqaRrgNYdaow/
WUmYD7O27zld0quQdx2IbPe1p8BWwZME1PLmfBpZT36Og9+N61Jf8MDJkrU/dXDA
9LykLSdnh6xelITuORHdmpmCNq2V86OsLa8Z12OjqxjIOQqRncgF5wWvi6PzE/eJ
L9AV3IvdMP8hKzISCl3060WEBTc1mG+TVpq5faNEEQqpKEeHe5amJcsKh/0aqI+i
0/xn0/bedh6zKy59OrXSzpPU5yXkahYlW+mm7tbVw0CGyqy3ouF1xhXai+eJR/Wf
Gaa2dbDobMhOmp9OfTBm71Fh6UhBJVt0NhpnBPM7YGw6ukYm9jY5/XlfZ7SNHI3/
zDERs1RebF6P5mi3bZyMmpemkTw8mWFpifURiWGldMI9xsYENaILJR45xaMx3shk
2Dp0IMgHKFKIM/Dhby41+A+ofOipLkhaIfVUNSz/MBHvsY2PiBVpty6YRHah39mi
TuBF2cTD5pXLj/GbtzFYb3rGMVA15I81w+mtCk1dGRBNtBCLoIf7shnOWkQmpk65
x3xQW/fukAlqCR8hz1+EVT+3I0k4EjM6hmANxolkmoE6YBYthIuwTljpyeq7u80i
a5C2TLzMIY6up0iQlLnkraVA8052EO49iuMGc4lkjhR02OcPPVejNNDZraQNIRAM
jTpOgfUpZnFhI84UTCBDgJkeEWtXUhoswBDY0KY8l7uXj5J4z6yZKVHN/ZoYvKg3
sNINKWpx8+pNdWcU94hpPJ6I368WRJ/BiCIwjkujEDmKnpUk5ptOXTxVoKKCyadt
nYQDomGqg0PTg/VGQKlJOR2jqMR0lgIOxmC9o1Mc2Pprmtu6abTaZshOo80pj5R5
v9jntMmKxoUvYZ1uoC2T4vp4eojTWj19dcmlSaTe6U69Oad8/Edv1bQPtZAHcjf/
OmkJ8wYdud0gL0YYS7f9BIedE0qxw3ETJwVIYNSyy1bOdMbue8rUd8b5UXI0I1UG
+VEjnTFzs83GOMreXMT73g7gH0RqWYhTZy7aknwE9R7HiE64lLS8RNMDqnZws/qc
KZ0UDY0fEkFLtIuf1MMxtYMq2NWEFLqvBGjQ7NIAmcwnQkQotnz+ab5b2pfm3kPS
VjpHHr1905MDxi+Q5Gi8oZeL3s6j75JB7NZT3lOYX9ApIDH+M/1XodJQbH3rkSLo
ETNz2pJwLOdwcPJbC0bWWDBnL2UYhTJMEzDdYUouLmE8tGotE4U7PRJE3PxN+Kp5
gRJ8x0yg0B4mMpm8OQJdMujcI6pN1GSjmztWQ215qVCHJMXNynn0sFck6VZRHV8E
WeV/5CyzZfHHQ3Nc33Owm1FGri40lm/+0MUkU6Y/2PTea3OfGjCpnqNOu+dbAQeW
/e4HHOBovaP5SXIdixGA84fXeT6volykeYhgHoQiHPgKq1rCRMGrRnRkCPilFQsQ
Qc8sNxihVi5TLSkgkEOrzO0Kz/qNH5xvc5tnW/JH4/MCHMm4syK82788d0ie3g9X
f4lBYN9kGS5EfxRmc253enJzEoKd9k8B8vcV5LoLrquR//OIDuSRAsSaBeVIJnZW
qPN6rJ3FJ60Kj5rHF6KvaMbPGP3KVe/g0Oz7igSTJTfIOtv13p/m+g7haLDuyid1
mSB38tH8zrhaR3DmgJ2iar+IG3C8gEOW/9KzMktW5Dfj4l6RC3uoY0D9C6dWucbf
Ydw3SlyBSrIOGnoWViv/xiUhK+nOEY+eUo3BGhNItqDglEswhmRpzXHiwSU8F6pq
zX3b/1BzdmU+aQoZujYo1RpFxJGxZvOy2MyYu/d1epoyec/BUPAGvSFN11SSpMkG
TLb5b0cZ2TYr70+/f74oPFv3qvNsOjmvDOPi0LxNFwxn7syR3wHoWZVQQQETXdcd
S9vv3u4BvU7ibVBjsiMwJp4GYonsRrAyGrQPRe7LzR+Y1NAYuT2kj2/gkA5jJtTS
kkdb89n1gwoG04lswn6GGpj0lStkpyk12L5NxbRg7k6hcO7SOdz9R9gNWcZ/u0iH
puI9UVN+Npmdzq36QnzIE/tojQKLMQgv0ckLaq5rGFVMTFw4U4H1q2wDGGvzjSLe
CIuLhfMQX0UO2vtiRn4sAwUWMRCSmXy4QBj0udxQZfVVD6fe8ifDdXtlhCa+kJnY
m10/FdnSEQzJDGLvuUpAe1Pms7Hc+ihy7NiSzrP1nLPCIFO/6bGv7H2pSGBdPS7e
2WEQeWsoaRDFZOEEmGKRNETR0SviQRrOEy1fopRPBmXZBJaeIldwjKNxKVuVkAgC
ljketTqiUAvTepFYgIL2pcKxkFD30Uq7Q14rryyfkTs3WsBtMbfdghik3CCOFuLp
LIffO5ODGoeB4SI4KRcoKf/Gc4ox4TF/47iQhUsO2JXQrx59GZDXah10/sceBUOY
yCGA6tJk6HNmKupObEKiX5AEyJRKC8tupVHax08GLgq2XniViog9Cq+Rc/0dY0Xw
Vr41BTkdG1z/Zt8qqPLbnetCKmH7N2D7V99nTsggIMyDguxeMY7pr7rENgQU/gIN
gGM7aD8j938XNKX4vDIUBeCY1BDZIQo46VQt/fn8ll5q6yrsxq3UiAGgp5SrGRZc
6esMhVjFXJzxsUsQIasBYvi2OoMUpk4H0gETosmJaZf6IubL8rtiT8TpLFzdVhUs
txm3bG0ox1LfIZFZkaX/p4AQJSgCVtgqw1pIaY3UOj1bz1cv0qMQEOi0oMICakkr
gv7FqZeGiRnhvz2ah2P2lR6hIAHSia5/XTBrinhwbVQcc+4N0gmJyZ1NpGJqUi31
5clH+AFHjVhhBP2UKXT/JM8CsfgNhxavNsYq8oIt5bMCBleNCJR6m8Sz4AVvQZmV
VeaJW3qhB/+RSB4lGLr6nbRqnXwnb1rJt4+lnJ16G6ZH2o6r454Uk/6PX3KzjRDm
HqLDggwVqUf8ApVLMmnzYwbKkON2DSetMGyttpBkj9IcS1k7/kCEUUwnrhKmGUn2
cwX3c9TCkLb78eGufXBPtJoVvlFpiyQ0sSCXbq/h1/Hf3AIAe3T3J52OAvixc3GP
YspirfbCVdaBNUBC6iTrCCEoacNbcK7N/IxYFdvDbmfhZke98mGydxQcd8LXXeRe
2IqTLF0D6K/KutiZ6aNhvkFekJfywmTuxsCuJSOoG4rrlfwXbmp2MJBI2CE3EqGq
GLdWLeDTrVpOxOLcAkIQ5S8SeLthkpXxEiTmpOWvp0A0Nbq0n6oLWL18jxWf33Yn
NWxpuTJsXJusiC3+RWlHauhB+Y7qB8GPRzv2Hzg5bRAlitHp9ePhShynI79za9gm
VjgTS/7OOyNiY9b/uhgp6msY16TnXjrZxiYpFGN8eN7lug72Lt//sqW0vxeoqomK
Dah0YD7nX478rqKN5AlA77UrthJZsLI7JGqgii0BUwD8xhW/bHC6LXiYr2OYQVL9
OyucxJp41OUPvmW3/yR6p5jStLOLESAVusUzqn5LtcWf0ZxkzZ0QuYoA09dDXMdh
J0ECDxdjjjbNLm/IMmeBO97EGRvFtG4adDx8/G3Mg+tqpPsX8hhWJ6BzsNvo+PUR
WtsPOfQieaxWGl0jydO+adYVV24EMjaR9ST550d89EFtatZkZg050vJ17//l8RI0
nlqwKA9cQlrK9rrojxHH0vWMHjB4X06Ysq9MkH4cweWt7miRmUS1srAKjmKK+WgE
0encS4Jplg1w5veM9dhC+dv+gaXD9Uwldx+AN7eBQR3mVBgwhKTc1O0oJjlrHnTw
Taz0B80fS/EBWqU64N57XELTtUJOn4yG1/fgF98wXluZGhD2pgbmaADvWEF7KVV+
sJin7dxATOpaDZYfdODcjcv27mOD9+5Fh2nYYQSDr9U1rRHUDCgF0WmMApxwXiu0
BQAACFytBvfNyQGvRpLCZ/CqLOyOcPKYPK874lwDlttTE9Cidzn1WItRggMuQkyg
9rrXqmG2urJuJSws7srrTR1t/DWQmJ6n1ZvRz7UAAa8lPD5fLs/cN8mB7Yl1qipD
ohHRlQFYG8gvi88t3dBZYB+4uYRgwhLb1dJAru+4Yndjov0+r3yW1PSG2ZRkl4tD
Ah4y6JZvdjrnbROE3jU9yVueDU3xARHlPd9uZ71rdy1xUWYj2Y+dYSCVD3IsvMRH
SKMTFMpf3DVJFqI5uLHOAciBlD6Z6r6oLxB2aczglNaD8bXJu0vO/6TdyA+HIi8W
DAo1ZNAbDQJYBqZnazE1E5pu2ZACRrVTRJ/KN0Pwjgzuc+QkIVRmiAy/j+FHbZFW
JSKe0jWT2QoNjcnlcvFYmT9IATOZEzN+aA7YVOxPTingE2EmZhaLTPs0+moJRfJZ
cIvjpuoCF8XrH1VEbicaDaq4leCqZydSC1hKhnulTU03QtA9RTcfBH003QnK2IMZ
wHnDxr0qY8qepRuW7osIB4oenpR7Y9bZY5XSFkjduBQEE2gncK1QLK8R5S4gaV4t
J4h7Xpp0RvAWMfvMm17HfLtNyIJhrEUcQ30w+UN2Gn8CxOCW9QELw2nvjsQj0vnT
2qqmc2zGZRdToiVLSws4Y6uCJ/eM8Al5GppVTf9fB3oPqDPdrTEtXZTX2GyIm4fl
CwA4M+AKUgZo8UZ1d2KZXdY2u2kZdwKPVjU3VnrQQWitt2Jasa65OyxD+MIMK+0h
RJDRvJCtunVzm8aTtz8K0EZ7nhvCE46IDKW4jsyh9IdcKqYITZWMPIjqLv+XzHRy
h0wKj8IinqBN35rXgbGsKz2RcS49PX5dPFl+zgzuI5Qaittfdj3jmsl1xdzVmJIa
KeHHrsLgmxiALuh5HMHSm81s8uO6e41wFsznBC3042VkXoXYjYVkwk9aIVQjr5Mq
DZJnxcO8VFEWgbJCz9ftgdFFWVX1tG3mfVQut0W+2YeYIE10Vla6qxL/IeQeXG6R
ntkApTQ7j/oJW6L71CXf9dBMzDYea35BG6hneUYSiWjJ6d+Tm19jCxLB/JLpWnY1
7ckcpoD4qXdBBZPYrKY6NpG4TpyZyuNGA4liFCCfNyORPC+10npFUwZPaxz3qbYI
SvQ+E1h1+ccyCvBC0p206k6Q7R1BYsrpCqPOk12Z2dmn/UX6RVfhq6vKOLZ1kEap
jFbYP/MwxuWIuXdH5qJODvuce0Rjyu30QI1QX2NWzsPzrINlo1SlVBql7xXWzdeP
0GG0WRGq1Yn6dlkFJMXyAJlcM7eTGlP7kK8JJgZC1FgEko3MXQkFyJKNl7Nmtrdb
GLj1higN4Oefcj27xQzubQ3qwaufnbA5ASqnhyL0Q1r0+LwAyAEkYaKK7DPYh45w
Fh96UR2sCzp00OIPTldQuH20Ynk457fZGHo8HowGBF1u/YIuQ3wevqAa1OzxQfE0
JVx9qL4X6Ko38skGG73jsRQ8DvLCiSgXIXd7l99HHLiT+QOxXVUl5wIo3+pyTCfg
KUanhaK1Xhf15Xc1tN1+PX+UCfKC3FL5d9H3ROj//OhmRoTwiOWt9saULew9gL/t
pA9APQSDPn3fleCQiFvc1MZVzJJtzqx7JuTNSCRcDd21fRuTKpVsBlgREHtUZAZ4
cY0wM/4om9KQCALJ3UiM7YRk6df/zYlJRyShM8nwDdA3j1SZh2ok9N7TeFzV3ddx
5bCPohDd91Mt5YSi+YnKo2a3vkgf52n0MNZVzl13TtpwR0T3yuYIzRV9bqhmLwi3
cpIoK4DOjJej6sfScMafjYrgivwm8YKjPNPxynFu9JO8bh8UEBmK6MQI+lAxw+OP
otYma0cusz3QcsdLQRGLkVTLedss2S/dN+bpQj+Wr/M89j+Jt49I+kEXYLJiixAk
UAyeSK8rFeqQBhLyPiZ7sDCxEHyMNKOm9RbzimDZI7Zr99fRQqWQwOhIeXWZ/9+Z
zkNugAES0HVhHs75FxlQv8X3AOBRS16IFR/8+JG/Sls+3y/x93CZt4d77tQ5G4be
fxv+8J8Lr0+6gF8Td1TLEJi4P7uPKIje2mWTpj2xLGJFV/tsLTc671ViajrIjycq
PJRDub+x1tvlMYbWkQXAvyMJ0Btx6Fjfp2zP3A6dE4hT26Ot6sHFvJEP5i6knWYr
UQhRxYcqDvU/tEIDYGGTc778ivohAIbIt7dvAnq8Ej63yeJSMwzQPJDPgQiyfCFF
4h1HlYPBc7YU6rFveRU+H/kDWfwkjwrk66RX87XSqK3p+rWKtpXfrmhuhoWLFh9Y
ESN3HjsRV4MyhVU4dfVXUD8gK850RI4FkUxy27uQI7rfljq/OFTQB0TSHBEV73oi
k1PvD9RSAIfbVWG2gNXw1ZjuC9rzxAlJjwlYgZp7KFUlBDJeCMMl6kOfKtD1+flM
2yT8ySpx3z9Md6+gWfSB1ZSC73o3Te1+I+MntaVyf6uZ+jhVHVB5CXF+2GDnCt4u
BoFJ64DMtnXNePVYsREGnqfQN9UTL3fzHgaScvqsRk4L9tyue0LsoRBOGi4z1X7U
rQJ3cXneFICulnXJKbPWzHpQpTRT7DsEvjzp31Es8i3Ts6VOCQcRHkaR8C5Cao47
x0EPp6HanEKYA3jx/TGO1ikohZtZK31C2q5z7fXIujvBtHR3Wd8MDDur45gA0lvb
BxiP47DduUfggw9hmxkZ9jP5En2hZr6yOo/kyQgC4ZJQXPTjkqMC5oki2kinCLKp
MA8EXN21/9ZFQ4AEUeMjjyS3C+8V6KVHZ46t1ilR+WbLrW5XzgsxdPemJooi9RFW
700NaQaWO++r7n2YG2LKfUY+KIxm6lbkL/MAWFMiZKS48m+8YVBj6OKiyfJkceQI
/LZatfLWjgGGfn6R5MRmHAXC3JlCmiGFPsIgMrNlOnEe4o1hn14DQRJFutZMEH2k
Pb7vBce+9vSkMo04EFgGdjQ6qImlXCwwJEeImHmbhyL7ULaxQcrRERmnJ49Sy6qK
O0GQrKxdC2exdTUcpqGdPxA6Y8FpOmXV8zKLAwaHDj8clJUa0aQ8/WvU4eHZsdK8
ryiQWNSHeGr+pvcr2D5Tbd2s26jtySdAr7Wyl25aAwgCkf4Cjfte/q4d8m++IHST
M6LYh64wBSzAWEr3BvEjkUl93V6THCQhOHBOs38b6pWE4l1qxNvBI2lvc2ncuYzG
+EJtkYVi4z2Utf6NWUCZRyb4AsGxL6RZXoi9hAZM85uxKonSdaqV0fkGp8k1yGK2
IutQMJOj/bHXRhjdcAzqX+zKQS8rhz6+HK7VARXZdXzT1qDVaQH13qeAwl8G2MgQ
Q5iPB5ZASrIm2UhxUlN88et6Pzxc4hgbl/+kbB/rrozcdDHPXabEeaoX9CS5Hyrg
eqPlPeZj2XIRiwEN6B2s6ty0ixphGM6nfKtFZPWXSEnZ3CaA8eUspCyamSWWd599
K646LKLREEoqO8d86vgTC+JTSxweYyiHbkYjzXwZiytRR9W5Hab9+JM3Lp3Ssczm
gXL64dSQpWVTmhY4LlOhEVZTvp8nbLk+3aoHZf5OJISYVn0GwNFZHaynHMAZ4BHW
vAYhngWyQrgHIm7lr4jPKiHjPNBEnVaieP3BcgJ8+HHagwgGo3pex8AOhHEQxR/t
Gg+bJOsdDA1YhA+6TRColqxA6Ax/G86Ryfrpcq13dQOhGbsInwK389bddzzqJ5Pq
EOL/LjGGs+w+kNT1gWJXfZnrdOoumk/mSevpJTk2SBmWfPweHVMNTOJKVpVt6hYR
Fe45naigLcXLXslmK8SlnOwjMpc0Rt5er52K3VDiR5CHMZ3o7aL5QPnWW+DvjxDN
zQi0G4V2EFer+ZSIp3aPv/CWHF1V6zyCdhpuE8sVoKMuunIfgMgoMNPQwWMkW35v
nzoxZIkKRMhaALOuuizCnr2rOOZnhdMm+tdJXSOZD03ba68/Q6dKBDbTL4oABGVx
zxXu8CEOIZQXATtwGUeUaGwoyspxwA++wblyF3zUi9TdNpeQSabm896Xzke6GBD5
8Osfw+69UyOdcFqobSN2ASUoq3xP73kGa2Cv7AsKMLR9+/Pd2EfIbhRrX3TmcQZH
KyE9nml3Bre6K7D82VHWr7JKAc7Y02Gy0rGHBm03SPi+QD39CnQL+R7hb7Rhsw3r
kG4zbf8vC+v2uJhH7Skul/bkzcYhyuOU0hdd+mjAUbwZ5Yj5UjkGro744J6txJ0T
ZQc4Uj/OFCs06V8rVERXSicm/cAzE+4XQcTrdMR0hcqLSCzZzxyvP19utKX2ZJ47
i3tMCCu6YEKcfYIQZckxwfFLbmMsNKn9aTCT9+DUVy2y3oL0ZE9dnfxoj9Vm+ypJ
IUINoZC3ieLErZuYrMpuOOORDULq2943sK17SJMgrGN+2ZIAnV5AjKFdwv/h75TM
eC1fMj7GAJ4x23e6UO4Wjin9xlfaQ5wbgfosjvQfIuKx58RZgiYbaklaSAdWaFYC
IS6a4WjATHuJ52aSDU4/q2MEUiUgx44nTnr2C8I2LUxiQN5RPLmLJy3QV7CfF+8Z
ZfgPkubb6fes1VOM6ybWUmPJQlEzl9h0M41b5MRHBUCtawNHnVLxEY5AAXoB3Za2
LyPpWTTcexpDL3GElHTs6wgDlMDGjVkg1+oYn9PHEeqFAYxtHjLN8wnBimY5NEKT
VPKoyWlc/E01Q9dr6dOlYyBDftsF4rWBfifxRMomgmFl0ap2JBMkA14kouxXlxn0
Yth9m+WSRcpDAKkQqy6IYmX+cHW7oYQqAgag33EDRN8NC2FCEV1IgFrXGFm0K53j
qdo4VBvbdoHmKBBUGWDkbcfv4WU6u3nf7ogDHc9Cp/RydPxYbSzi7UMK+vUUSW1+
RUgCAlHx51dplm3pYBi8g8HX8wf44WzmrL0Ex4ATrVOOn2N25qz/vLU4XziADVlz
n/CueK6d4GWtjOm16jm2SgTffyJk2A6w5vskJBOwAYLHYBB2iCorHjn5CZNAi0ao
onadGoiAMOLcocTQUIGATvayZrsBpYFHjGf162/Ije6nHJxomluOqHciP5d5bWxn
acRhjabdlB8NkXRDrMhBWjKVV2M8Afnua77N9HYoUjqy3fPRqoA9fYlq8DovXml3
iwLXvkAR3x/DZPGTp8icAvwSaezgfW0s0xJ2ny1r0IfoADMNtxAAj/979dU3ypJ7
ViRgS5uD6wgHJ1yxTlIWFutM+qeF9gv4pT8nZE5mutoCa50kEzOuPFjpK2oAvwEI
JU3X/18fjJWd8AuKp+1lxZnjV5Bzms3mFIbYb39yPf6i/sBpBEFzV1oLlbESp5ZE
R3wEpeGFOj0Ooiw53wAep4JRsbspFOnOS965Vrf/ADRml5AUysntgCoHDpbGIMX4
1SX5zRd8HgutNwlCNZyBgxFrPh8VepsiaSxOo+RbP+3/AzYYViqdTVENlRHwEP2K
40wlMm+Yf4UYrMIbgUBwfj/PYS5ITniHQCM4EozaqLtbLeNc5AENgv3Nij3Mg38m
PpbA6DAGExE8P9U5uKO3Gssd1bgoXfY2A4hk953uKwXpQiq3vbaGR0ah6haoUYe8
64dnJIWgp1j3VLTC9LHUW9V/IVpYXw31YZLSInQ1GpdTXsP8YZlFj0zDTC9bLVar
79Qs+ia6o57JjFDVMoweA+f4xzCzu9xIwvwYgJVoZ8pWBrqE+wlBwMna1G5V/Wus
Gi4rgRY4wzIu1xPEChcwjpELp3wNv3P4Ly9A1X7U3r3kz4yfZ4jQAQRkktKevagL
3pWzUIiuYmwAB9+utHdF6IzybcxZSkAS5W5g9w/xKVLSkMQi9qumgg/9so8FdKip
t7u8dL39WG99XOj9qOLRNIpShWIl57fHMUj9GyINwc6T10Y8qn+3L+2zgqRC5kJF
LF/R9jss/y9gQSODZCYBv+Ms30MVIgosMJ0/Tobs7OAAlH4v4VHhtUaI3sN6ET2/
OixbqKlZwke4cY/YWYXSXwGzYq7U6ADQwgGl5GSiNI7MRmJ0dXGkcol1tKBbsqLd
77rYJx1AApTyS+qNJkL8ID3Pd9SteIb3p3PTB2m86dxoSeAHYIwKHW6VAn1fW2II
2d9Y56BSYlksZ5rqIUV/Xm/yLWUQrClEXSxsLA0Pm9HAHA/rni0vDm/Bwd4UbOYY
HeG6mGI43Zsf4NYgAIdvuCxC2YsUDEVxYEHFNX5ZuotM6LXKD9BEUA32QjjXb/za
nOf96j/8uXr13n63E9bHWjsdJl28f9Gls07v5eqEmCX3FgIRpoj3SISiiC5gILd9
XUvP9eJio8Z+s1ylJdyTKXFWJSMZs47u7r2RwZr8CwbKn5CKAIkAk4GbqakOfEee
tr8929ushNNX1Z53GarMMR/o+e69D8VPk12itbowktcb6YPRvs9726EqWs3rrcx4
ZbZrlCvoIMQML08OTj2ul1RQrilrO2XcMkxoG08+lWe3kGohP7NwDPMQ7naH1RYI
cETA5VM5j2VFJMDaNBUZSH3V4z9ODktjKVOJ0YjR82/xOKXInfIOd2lm4QYG9qzm
7U9aQcXVD7S/o3G+/xu710NQVywV2WNuA2xaKSZd8p/19iOgryLvZNC72y36m6Wh
7fMCrD6IRjqMexsZxn/qv+FmAz4F3VM7pAmZokY2islwNM44Ibfk8b5QkMvlrkeH
TO2Umv1lCgURqvaZUPhUcQg55e9TUoTyAzzHMRlvdPaCGxur7RKwBJpQGYsrYgQw
fCCSOlosd5aedK89GqzTZ+7bcKoUEMxSMXTWK7L7IACb7RUuCGvcS/sYY6580Xa0
Mt8neMA5Gpb83U6p5AaBsUnTCG7PRQ1hf3NBVcleYEKtxaCXnPPotv+1pNFdg3DO
d35T/QOlza3ez1lFx4bBN/3fTddR0jqjUMlN0Nd2m3VDgCexg9IGNKG2nciRtCf+
WHvhZuDmB56sKtQ1sfguy+3ZnOio5LTFR+9heew8OOhymYDyYW6Mff3YVPKmGi/Z
gLbwEISrm9IffoKrqu8EhgLQ9g0dioDdXD710350vHfb7s9P9PFL6pLBVIdRv56I
DLYYto4AgE0MqnlAkQAtNOjsTIDBV0ElZhQkFufm2HRNp5xPbw13g2Io5Ab7ZNzG
uFFBztpz71YotCbD7wo8lZx1mxZHt762FCbhYs4O9WCR0yb7dnf+lqY4wSGcuSgw
zOoUzkca+wyzoxWaF+Cu2l1WoFQxn5amARHOlVQ3vWqgNywbIQ+i1in//Ge3GJ8h
nL9obZyZBwBgxRDCCGuLWSKu+SDftOWBpUAN6LaFp4bXbBomDxIj3nVFpfRmQniY
eeVuXp+6zTTEo9IWaq0A7ecjVs2VNCabattw4EfLVl3Rg5aiwzb9ArTPjxj8W6Lu
uPeihD6xv3vSBjEFceXXGNoOsQe9VNWBlFdErMgASOajO/CDabVizoe+nHhPtVa0
/Vi2bMv9AtgbKj8PezqouoEYdcd0GKKpZKAQEXzZxhyjVmNUS4V+zUGgwufY0Xpo
JTX2/5JFYIYSyZH+Iwhnk0yWGECbP3lIKv8FmejlWlhYKQJEzNJEBo/0fTWG1eNf
tMFrSVuhqvZ5+FuAsy22accFJ4FwRsUwLFRuRo0YkC6b6VfcroxLLv9k2sT/c5qc
ooidpICIkHv9MspA9hGia92UiPEzpMSgQssWFEtlEsdkff4E5kQ6SF3D3Xhk+1m2
0rSwh8/SLyZAxmTen7cc5CNGx7Dvco+ZQfTcGNZMRWZiUaau/AlH5QO6gCioILwx
fveI02qeVbmuN1XEz+xpQ7Ik3k6h7hmeTjn/Xvkju9DZAtOn6k3wLTDZAxBp4Wiy
sS4iKadd/V+A9AYRMdm6asj/2yChJs7lxMrWMM1M6BsYG9pV75oyyprAgqbt6PoG
nhCTqV+ic8Hz1Z6LU2VeJaT8RTRZUlByNpZU+m8hp68cQrOcwBkGkTxG+hIyW6/3
BS/h81OfksD4oZPePIXtg7L5h2/AN6F2SMIgMFSJTWdh3d3+Q9XKKH6eM4Pc7oK/
e0vXitizFjxN3bD9BPU2kKLBl48Veqrsc+9cj9g9TsI78J1p0TewmxgoMtg6NK5j
Rvmx8WtkA2Frr2tQLCeQsu6zTiFxaHAQhKl5W+4PA6x8hsamyDhCk4J6YoBrS9OM
rKC0c9cwrS/99IgfuS07AJluwZ+G8K+pISD2lciWMbETSHGECjvc4Xd+/trovLsb
C48GCKduG9fSL+CVOyoG2FEd73Ck2rqVyDc7AtEaADkmwuRq1XHUjERVmEoI5Isx
Yg2k/qrEd+gLtWKBFsoovux8xrv1BGEf73i6Rht9nNNAOZslh3mYq7JgzMb2982o
14qwKUkkQOPfE8yRKLcEMcZbjW9sfEw+pRHUdq9ZtPLWms53sv1Pc0E2eln/MXQ0
K7Y3/H9wOoow5OdGYrUMh9ePQHVUT1sbbHbjsl1hO7uxHELF/xSxcwBs/wd2mN3B
YExJsIr9Et+G3+teTqR5klXSF76i9kB+Wm2WiVrQiUNwRBnHcmdSWBtNJyQ8qUSK
zYDen5MnUjG6wRkPhSRGNWfHrOu/V6f5ElHrOrBX5AIitifM3mdkFTa3jKpJnp3W
/skMVB52oLafqIN3UODRe6DdH9lKIwawkpblmW9igohdkv/gj3ajOf8+3fFuYF3t
pjj07Wr8m7LPkiJ/uTPK/llvOfTUTUJp7BW0RMlnedC3blR/qUp3hyBtTJv0XD+r
IfZgccT5WnjyKpZu0PWpEQaOwfQfgd0VgB8+VKJ6y6uwrI003DBgh4SVqg6N+5y6
0GGaSidVWMGwJ6S6PEBSezcKcEfP7JnahrPwTAn1o0uzuiacZtZbw+PDTvfxFdlV
+zlVAYN0WWygG01P0Zf4FlQyFuTEsbU1qI7H4SrQ58zkQZ3EAfZJXqLFTADMVwov
hl9+OFN5Na08nRZPnUojns/Cqyp8F4V7Mybrv9irq7xz/42cqqcEpwlF2L5DsHyC
WTJPmYClFflerVg0Kj1ZsLcpLlLMGm+su6pULcjJOfI9e+4x5AxoQ7mF0z4gOo1D
DRyicxPifVFaEQY4kRvk+smS1TAOWBGsNxRMO4VymomVXBI246ceCjIEIww0jlj6
Z0SV/6g9UlAcrd9F0q0yBE0vK9G5bx3FJjs0G15rs/Dex/ucudzwe+oS9H7FyF05
ar+7rhb+K1LnslPh3rvsK+w3pDcJ2sG6iYT4wy0awQmyK4L2twaf0C5uQ/glLtv6
mrIXcGoGAcfrQ2WqrZ93vWANWVvNxQr8/PkniMhwwq7vDg9IcAbzyUzFIwWC0t3w
Zsqixy+RsmTt/h2USk8srzml6GElIioxWQi4qsZuT6Si5LcJ3TJhXfw8mYUQ7RwP
EdLoEFf5bljUea7fsOTO3ZeqB43Q/6x2fEm91+rz66Oa5GP+UTJ4gRnk8dOYlwvK
Y2mQ6baxpbyljq7eILQAJLfrWYnBGTi7TTsnyvngjlIkfaj+aTYQcO/2FmpjfpmX
YCj1zi/+5KXreEw9ZCwuUCsDJfC5AUsNVXqcCI3JV7TslDYNTVzAKRAbTdcNjmGG
MLUFkKNPbQGr8D7jRFQOH3YI5PU3fzDhfAVbHHVD2budaN1y8OrsI/pn+4gL+Nvr
Z5RDYDLx757HarluA+Ken/m1S5royBKFUZPCUvdtjpQvoxhOgSxQ33+ioToJaiyC
pjYIsyVwVngMNmCMkbm5W1bmQdb5zO/EEnkpSMfYOStBNI1d+4RVF37w6lHLAeCf
UZkz9ztEwjrSX2CHk5Sl6nUaoT1G6nR6eF5Z+q94ZsxolhoN6NBexj0T2KsEmHdh
n6EUd5NFon2P3wdYFTFKAmrZyQqmcmaXZqZuE34lzzNRaV8/aJya+HJcdGiSeyOG
hEewIkDCJ5DCkXqn+gdLd9gJ8JkaPpH4kST5TVD/ULR8fzSgHAo6p/WV/x+xPYvm
oytXyJWRirHn1sNnk6Ib88IJulf/arIW5OFOroDhP22auyT2gGULQWAyx3YLagpd
7axMSP4aDCwJf54LtX0c4AjowU+B9emKeMoxXhLGmR5d4VvgrAtvI/S31LPPZ+rV
9QFozPFVkOsPKCPokSBwRflzqKpVv312BRCu8i9PdKAmXaYoZyIAnm0XCZagc1WR
3+cia36IgjDqZdeyzrGs/BbqJOikAQP2rE1K0Y05xaRHM2nZqaruxhtA/YCjsFuz
GZtdKxCT/kKvgiXS51ezlzquxL/traGESbsg9bI2buF1N/2BSD+EoW5l7vqlqClg
hLSW7fD6gc3MihB1W8fyBxMnPWZWgxOai9kiG7cZoznkRvJLS+N1Bq4RaIfroTe+
kNaO4YHEJLNo3ZtZmsLliN579bCqChjeppwoaYwRGr9r3ib6HFgdVUu82grGBtAX
ZLzHoFn6nsykumg7diAuzlJE+3eKABOKQBF8ebO779QIk70/3foJ7X9DJsn3caKc
qvGHoKszD8d3shkNOSSwNleCIsprm3N+3Oy12gpnWH6UbtEdZUeAeNuxAmzq7Igv
REtcwzroMWMWGts94eZAhZk1Td/A+vbI7wEF3O/Yv+dF3cUDa3XCaGicHbioIzzb
ouegs3v0Xp0SeCAmkpyclBl+B3hdwuRG6+mXhfv6ssgtF+wBXU5hrWTLWSKjKZ+g
TgYdnf373+PhsFkautpIJSBrD3n4YvahMK7MYt5f45QQ+zysYZNmsKWg2fnWJFFP
vOY598cTSKlHf0tMlpNaGsjRSo/dPPt45EDImiA8NzWSmUWjU/U2zMB4tE3N4l1u
WiG9JhQg4N+PTjgc6aizthhPZui2lDGTzV9AjcNUJ1f0CZkNDJIOZY/rDKjelZXb
SfyOzlLyq++No59uFUkoIGAokXBc2aWw3MXXCEktDp3WdfpmVhi3WHhUpfPm5HhB
RVepvUt5H0NlvPbMWu09WlNUo8tQ7g38MegqWpPP/gdbusln/alMf5tWp7hs9+BE
xRImqT5gnEnwWY0lfQJ2kxVN7mbQ+ardJNR7VsQlbOsO3jBTWK9mqNLxtC5DHk23
B2mEVyttQXPyf0P/1c4a9MvqOaYOOn9Of9z3z8NxQhim6VXZ1hhNo4AqdfSHNE3a
NkaVikkZK6YP/8r2thR62xoy1zdfv+DRjTlVN3WEtbTZli8jC9/1JTcPvVRlvlRF
LgU+4cWvPRic4arcHlGCrjqMNWzp+x1aBIqK0glpjf9rXjoZVNuqO24FfNQGfQby
M6/u0lIPEdURmi1zr8bt9jC8e5a6AnDz/nfNd3xu++9diWJ0kX2duqGeWKqUBqL7
B8JHYHeTG1XsQOJ60hllPo4O99151pcgXarOIDSGCMSufJtEmzYWOputbIsgbM44
6tOu65uDdbOjeEin2eMLHDhsTpV7M0P8NvVviCYtGWHSGMjfiHYbQYpmqmQf+IEs
8UEJRKfZvBt+dFwbiEyVVsRyuEFAeWnkNOPgXW9cLaIDgVjkKgdgbIhtMmFFRA8s
KLh4mCUDKMQjzbVECOflgMxuQPg34PZzxBXtZ9BBMrt0oLyjX+SqFfX30K5Q48sB
lG/sviSlCaWnyoJNEPYwNvLbT1PMOIoLoh8UL/Gq+bmdLRmo997IwaNZw6bMY9Qn
yvZKbSq0IaoawQaTq1CegSu2dXubJIcurXD67nxQEVaIQ1n2Ry+vXB47X6itpsrP
d2fZzx9uZm6tz2N3ZIBGQk5xXsdG0dz7Ua+zFl3fHBgpI0ewvoAYDS4qByyw6Uww
CAX8+Kk5Bz+OMerDO9pB1gyw7mEf3VI2qzgNcJv9drw88vv6cGYqnhXP6v8wQ+Qx
5kSgzsGjfdckU3BddpE2KREkE53gVTvUi8HOtPpLNS4iSY6KxlnR/dp4Ikj+iBXy
15tSrRl92B502pBXY7QpbpsK7BCvJeIcVYsibri9esGmkFdBbmMD4mpgif38x4Cw
v1NoVkVkclAvbd6XzDS/Aa4Anp/9bw3i0aOzLLNjoJPXfH/yWW0bazo+cZT4y0Mw
TT+emkP/HU6qe+gPV7TFhABghOsyYnJ0nmh2/PwPOuijj7S6llJtpe0ugL8H26vy
O4EBioYo/wJBwi36tm93qNzvrbees/G7rNMYYu1ynRaiFvGhqAANY/bZT0DCxin9
YdHBjN4L+dDuYBQaTLgsdqF6p5ErP9hz2deWoB0LpTGJjxKHpfgKF5nOLCZEDaUq
mmWNEBgzQ429M0SoeKq5pBBYAFuHcKd90v0xb5Z/W2N1/Ya7elazirCOavPoYQCD
6XFgN373XwpJktdarxLe5FhwKRI38zPhlfh/IFelhXuWJHmMqGBQ/7kmUNUibIKb
UfIeSRUpItmXMjf3HMcsj4Faiuvso9DxYK6udnhnMrG0ZuajiJdr8bQg7fdmEjzc
xd3it42p26Vq6n+8ewNOFEx7XtLGP855myBmTGVMliz1V03VXP9y0AE49Z4eKMCz
lL3CJK0KngxhiXD2OoeUDAOa17qhexC/uqHla2oiBlWathTU0Z2ymkC9DV9/1TSs
rN3E1kuUfp9mipun9ULd0rC9f9NGwd4kfaqbaZmEiCMDPYP+9IllZKaAvo0c9Jrj
ocK8ipZl7KqUMf7VzQjajSLtd/NjngSVaEISHfjpXjAmbsHcgDh0iSEmUiR7AetB
dMqVro7u0Y0Hkb7SHx+F5D045EKAluqVliuGXpZ19A3ciMu5gVG9yQ4k2vbqqhMJ
3I5VZFyC9ulSCH3ecT5HmdU4ZLEr1IVSeLVPgI2CwJWQLfb5PUFxDR+VFMOAudJN
razAxBoBDh4Dzodkig+G0/rptjZnB0msLnr0f3hmW/lWMLOJ6xXBMwG6ty2YEaXJ
vcUUexHLOZT5+feOM3WooNmbF7qbBUaWglkxJoq5p4JvqF2EPAULaPOSICVTG7rR
ivHqVohEigz1Gjj4NrGBAzzQS4M7hBJzepQOR+p6E+UIKszAkFNd9+QT2e5E+iVW
9I+6L8hXU6bFkrnejHwtwrd6CRe4nyzhhKIrWyYey/bIf28kVMkLJ32utBcoMLWA
tFqwE714jXrUh0z40NKu3xy9muqoZJkCskSpLkL7WBoJtYQn0X3mOj1k8IeGAG/O
8BN+7RgMAHJtlfhK26nww0tm9j/fFsb/4MTAsPOkyZDh/2scbwr5WxUs0vG6nSqd
IA3bAH6Jn78w5Yi6RVoKqICWe4eNqAprvnf5xbIrfch+OCv9bwGKIuQWLySPgTeF
xV9nso19l4ZCW70wUAFlq77BdTLlTRkZQdlE/rJKAPjDI4UuaDq3J4DeZARobPD4
82YwFvfT33QwtYD2gL0MOmvZwVn3HsJ92XqGU3MKXdwAKKeYWxZnTKXFmPAIsg3f
Qf7ZhX6uaxjMMbZSM0xNymWGj4R9OdX5S5o7hplIwT7BGVl8DCMjU8hp7xNKpnHW
PAqw0SCiXRLv7GaQu2aZVtTYT76aFlh8mRbDBg5Yf1vDoIXwB3XSCiwvnkMSHYgy
4dR9gYyhXHG1NneEHnxa2WXPU0H8XvQ5fVjkVVjw+AuZ+yckM2P6jB6djhPqIgXy
yR1AM0rL+2AXRwDkiZs3kYzZEfgoWxEoDr31JbbZpAZzp+snZTns587yuri7w6Nv
kbxgpsarc8Pfq4EunPMH4vKVSzWztmGFEkwfLzytVPoX3+1Nl26DyNfeR+gP/peK
a5PXuwo83bgvKHCExU9aUkoY0ACfFsfWTN+PoF9KjXYKmaR73ZcckAd+wQxfGEtH
rHuPcKIQNZMD1MPgc/VfEk8baQEu19Dabd7hogsQCTwKtitg/bNkQghG4QQeVLhG
WDZ2btOmD+JjSDjBLcjWkJIkflvYcCP3zT4eCwZ70EElC7XRCXStZiW87x40GK3o
3s1z9y9zPvvrOX+7yUUKsaIi/mpx3V9lw5rVr1JmDehQ6y/eqEvNfySiPtKXtP7G
9ROpWJ4OzNOCgZUCmwY11o0uZcrM3+KTpcoXRi+/YJYMmM9JY/6c1iSMgFjPw2qN
wM20wAbxb13O+4b+sQqp3gDOvgPeNaqUm/qa6q13cfjboILwAFohvKX4Dd2H7F9t
kHTP36fO4oEcHXKDW9/OsQMLmxAvc0eZTkZS/a7KbxJU9lpsny9X/T2cU/ifYfTu
Fr/alrgChntm9oAwvsALvII6iQwKK+0EHPhr90D6+gFDX+9GiBL4Oo/U8HInPbDM
u5up5/xNVDi8xLQCO9tCQ8kvzvNcXOB6UgR7uXddzAvpH5LlgBGWZ0+daRYjB54M
B0mmPzb6Vp82faYUZjgopzNNiO6yamorxAxy8ozVe57xjoZgNX8Tkuz3x4/UAtG6
2kYxRzgjfCsoigQ+/oFotEbCVAL6Dy9xYSI2ypBZmW0SyI6Q+tejY1wA34iwkWMX
HQN4VZL1QMsE7qXXpkea1v8phamuWq6H8BYQwqS6LmoQTRXyZqhnnGp1KXJd+kSN
5+oAZNLHmSRj4i0GBpeWhYMI4Tfr/nfcT1wh3nDsFTZwYLPZJXfbB4CyWXUJyuDF
PxAd7A5bB+SHH2FaJ1+1CzgOlO8KiFlv+poAerivvrR7x2bdS3dL61camstV3S/Y
xb90mpeAmViZCnBjH5E3gGyIaRvA6vYSeyCGjWHUqxIaBcKnOTKAp7st+zc4aBi+
mDhMkZwfL+MDABj9I6pFvqQ4Mc2dZzunWe3HUvZavwFCSQSmenz/XqJpfh2zpytO
qjI6Ze3dm/Ai3shT1q3vDxshnc80eBM4jX2Wf9pLEVajmHNTnPuwj/hJEVyCmDUG
wnYNSIHqzycqwlM+Mn56evQ1rhl56/qMawKJU8uXTemJdhnGnIhPyPTV39kd1V36
q+qm9vVWvG16wPaqUFaoo7Xq0l5aWl3qzuxPUJcUYmTVv89nZvH4QzAGs5OQ4jAE
fyAdW49i69lOmT6yujzukaQWrMj4dzitkk+SCD6k9HBXy0HrQJr3fwaAiRFyuPBT
DmyaPNjIBE7rCebjh4xfkOyLUUG9yIv0wZvJfLg+wERESRjdIRWXOZdTe0hXdeYP
WfOkvFe3CTvC+NJneDJ5f88x6sBGg1PqygiZdPUdZg8zSRPERz5HZIFDuyioRWoO
b9O7uV/F66hGppPPMSsGTdTy/IMls/7TRVasQpnQrbsBkR13fq59hAIcYmqguVtx
UymCw+4jXYZ9VXxP8nFJYPzgmpZOA9B9Bsbrcf/8z4jFIJ95KwhOqObzwv2xKYkQ
gDi4SFnvYA1+wLGIP/iloYupOVX2b0stiVerN9q+KI8JtcgOoGKFkWeg0edQXJ0E
bJ8UBiphWBGdoinhCKlNPc7YWfyd3AykSUimTjeMDmumWWv3iSgOZpxlWS2/WCrY
tlmyV0foDoWYSLYSe+vkyrFTcFeEOB5YwMFw5x0DIMrshdsnYyFjBdgMBzC4Gp05
roeK96+bXAZm7APe8V7229xCm/eVdpuJbd96vXqtlICt1oUpUEOGlkXSh0NKGntv
17snvbn8Z9848aS6uey3d7NZ7LKLzZnJ60ICeEmgka0s07Mk5hs7TwZVJcVaB1qm
/bF9lGn92wyzMBJjnrqVDU0VApY00tlVqurW4iZ4u/8WszSaXmMYsFdVrxY1mBpu
KAjkWhf8Qy0Qy8kwwCUvqik/D/t1TNOqAj2JITsHo1GJ/VCxYJEBrC74phpKcj9k
sBPUcVZt36Gtcz0LV0cQQ5mA9JxHse3UNCqLinHRJunmoQM1nK3pKb/JHt7K2OID
Zd3I0a9XoC9whkpcDs2WqF9NkJeR8h8TUaihlkxXOXHvZ8NJ5Raf2Pu+G91Zlqog
uviaFQVOZegtJnkdECqfq+HHfcf4AAIUQqcx82LZCiY7pO7pf1GhXxPqznneHVuY
K2WTMQDJzjmdUAbFgmvJkwTIu3LQTpSumDIMyPYbeMcJkiafIQ42zjSHSqt6BbFH
uyjSNsFQq1Ucdrzftl/gEkHzVr7CR0Z1g6Sovt6LLjKfPaywRbL2osfZuPLm3e8r
7XXWdMhjX7MNmt5HFrzGgX48TSwzUamYW4gRJp12pc9Z5fVgIXP3d3wptEZvw9O2
15LK//9teJliPadEF05rtemw0jsFLFRbcC5ho6Nyn+ZvJHRL51RKiH9F/b202nUI
eOsYpPE+hgUl2uvAaabah8HcWzdqwdYKmeSIzmjeak273WNdxLSd9u2DTxAEiJpl
UDHdFrlQSTkeUhdYl2p7PvIAmVWlhPdi5u4mvgffG0oXduwxiRZ5ClxY8t7kYZqM
eXiIBmtsfXKTpcbDCzWS4cBI0l9FEAv9y7bO/zt43Fo7ceOMHPJ1f7EldnM7iCxt
BHINnmubw20+AsWdzbj0neN9CxreGqX7UgCwFedVoN2IGtGrS5EfagRr62m8PZdY
/Cm/PwPb1fs3QY1OqRCLae8iXsz4i3o/Wnc0k+lPW+KWseB7kbMlpCBf7acX0uHL
W4i2GWdDF9W9wEeI/ctuyPV0u+c5rft4FQkZ6D00y5i+ZSNFoRwCFveHJNpVwHR7
+92bc6eMENeOf5I1AzaMLsv83TtL2KzLokEwaM5v3/Luv3KlBZ69N2H6SfUHQRMH
mzNxaKMkUDTY+K8hKBoknRF4Ov6UEwCz8FJ0BbjfN4bx9WVfBCcJGsRbuYvDjoXZ
h0rpVZ9A+mwy7vrZewmUwsbeBjDelXlYwMQJob3iH7bxOw/eD4LYGQQ9UMtXUChZ
AXbk0M8HLvQh7v7L2XtMLqbGz+gBswhtTPQcjdBUUitXuFFpTqs4tch6+3sVN1hY
0McXpZbSy2tJm0u+DVl5r/Txfd+zT60BMQSCd1WgcjmEzKdp2PRcYlk6RI82Ckf1
aaYEpBWI1SOSYgCzgtutZhOYd5OB5kS+/6EUd+O6jfSPADKm+5BlLb7zBhZ+6qRH
gOETjiYzjihfA8FpeVBlXU9JNZlwaEQQk0HIkmXbTa253StBZLKD084V3kT9HYny
bIlzRlWAtQ8czLPsPWkEi4yh3rVgj6bEC2C6+Crr5H1VEFeS18ADmy+TduMFyuaH
sgWIf7Hx7zqbi+xk9LBb3crCQl1t7VfHreCmTx6YsOpGFzvKSpLTrbjncRhgCjBg
ULq/lbJCAuzWZ8x9JdBcXmRHHzC2yENmcP5KuqOhe6MZw6tuHvXorxOVxITJCL8h
Pd2VTiISdftxX/hnMCZDHW3p/FrwAMi3U/jsAXoxSSCdYQ0bkiOxQUklc8MPwEMJ
d26P3r9W9arN3NuRqORdprJzeR2PXfG5SjcxMi+jb2dLXs8IhonEGshfgPg491yb
dw2Kd+p+BSbkmeMQqqBe/TOQDUnnDxx+RsAznnMkLgxjqEhtnL9LvSrMe1kRvSWz
U2Yc4uVqe/6F8m0Pg9MUICxTJueXqk/4OUt9Rg0gM+f44bBDdDi1dOXSqojJuNyj
WPn0U0iySPzrR9sG9DQMRGU/xjRFhMo7fbSsHy6Bth/69PRm/hXaZWFxBu8KPy+6
Ee9B+7KQLvvydhn2EWfxu1kYYnk0A56aJFbzAz2JsBpJmHn2U61HpsdKCBHaTOJ+
j/jRHj7HbVcggqeiRTWc23jlGfhZ+l5XyqSR5e+a009x2tzRw1rsitHwEOSmVO57
jHVa9Bd8stJj75KKBX9CxRS3AlJR/BUiwBYgf8fwYwtLPKxwqbF4aMp7FlAOXafR
5a9BMebk+HVTD9b+99vSIoZ1RvDEzk8JgM8z89LFpBycqVmZnnvgHsh57NzNb6wI
1PftUFGxCg1X4/SzxQ901IePj2NYTWDIyPXNgwx8vZ3eu/XSJHDPZSktuXq9bB3r
akMQsxKaNDDX24ZTFZL+9KnYzukfbpVCfjiwiNYAyILm4889C/mgWPmsJaTChI+C
IPUSZNF8RKf877RYP/0rFdOP/TZBKGG7fEhwEjfkAF9b7AdtvrgGwccNUDpz0XFg
i1TQAogj+SVEEVY/nnIoswwKxZb2++aOy65VQFj860TlzKEwNiLT1msPP7MWnlVC
7dFQNqt6q3MNjmNPj+PRgLCYwqfelSzj84dkah2rbA/obyz4k8TGj0gOPOwV+/o2
TsSWclrgV/Vi4N/006uSVlzSh5B5Fmapa0IVlACDBVjcr+Jy5FI2S9K0W0cS+slj
LWhYDjwHeOuoAE4JvdOs7ZeAok0u442SDcwA1V9Y4DMngdK+kY9PTyjN/OSZzhlp
GRR4zYqz1xzMfOT+/EyNLUYsLOJmJ6P4lOLk4G4tngVYp4WMOuIuSNP3V2OIL4jw
S7Qy3DOURLhIKTt6hIhoCh6MwgBDHJ4wvA3FIcgdeUKSmfff5iTvrSrjqB/baxOY
ysI1lzFc6s4skc6q2MnC6Yc18CE0KQw3tXwkstTwUvaB2PW2nF7a44dK2f1DYeCo
GdLcWEH5/1jaUyAPiBm41PYrUy7W6mJSYHBSSlSTwJIHRlC4S8Q+MtldxXku6Q78
xTEoWZ8BrWWk47ET4JAU/vSZH9bDsCd1bHyMYIqLcs0jcOX0chK2yGAa8sP9Mgho
meCQ4Sg1hBzodXbnoDao6yXmymXOkSU9TYH4kDL/fTVHhGqVbeujOAEKAoyKpRX0
jIkxGO+cAnovMHIsOyBZEEzTqvif7vHC/SbEirFr8ztF7Xajye2wdGs9txq4I5PG
QDHgZx15XCttm7E0knmsG9TQNrjAkEJHpcHcmPqhJEOdKmF+q/vwrnrE+G4GUlZR
CeRRWErLttFoo6znrAo07fn+HlTJqQ6RDMgj/DgyZB5louX1nAj8KcOfQKI4vDWX
90E33EOaRPecui1t7LJY5FbjgHBd4hkXofMBqPDczsmXiR2jkpdgdZYAM5XM1a4g
+gNIhUNLG3R9oJ4x6K2wgnLmJdn2oz8j2GP1hCjYMe0QUvumE8slBMmoo+6OMVdf
SXsxxbfR/7/eVSs4eM989AvZzaATlOuQXJmrKWOSTnHFVtruCNjjQ7wdzcs9LQ+l
vQgY2gFVbFOfC/T7C/UKsoHji26K2TxmGrWWG1soopE9zKyEe7f7ced/NXzaBX8C
3qjRdNvO2rnKa5IOODmRjSuVT+60zxIhzTyH74gg/yUe4xlr/U/XssIwkGw6cWoS
28v8eRRVSfcuWi7xesHHg9lXU2S45gegxqvh3/gYYsYUKOxXLslQKCBvXFnrQ1Se
pMg5mWx3H7G9Q1C7YR8QYd/XzDDBORGZ9VHED5sMAewJi0zYbp4o2n65uyKQdnzd
BJ0nmJY6iC0/A1XibLZtzs/Kf3NK1lJvj5mw5xIrCbWG5NysRn8LU/votf8Lr4se
LvK4RuufbI3oWejigYFVpZ0TWhaBsvXw807RFmdbrcC+r90OnZ6RuxNjGNgL+Cel
yhW+gz6dybm4kKM/8v6u/KU0JKElq0CWJx8tFQ4uKiClUzTY7hs4Jsc230KfVzsd
6ylWOoU1WiDmfx/5cHXFdxE3lGozYx+XK23rXN6X1rKa93VAahXMTpoQcDbZ33mU
9pe6mo8O4r5jdHCKJzlp2BqkkiyEWTetAKe9U0k6BocK8dLAmBnWU02iy9K8KTKt
yTKX8/v6skUVvT0b+5ydZlXszhWNQRFjV+edziRfUppDt5KVAE0URs9ntmQgcCyy
t0GH97XR+pnDFpJr3bnYjhYbhI6xep2T9cB2ACs+TsKqODwgbaKAxceLJy2qqYA5
5eYa1wFwLQHDGNFUy+kMWvqLHoxeQ7N6RSu9rjfqTjPX8FSD4X8mUVzDed4ADOqI
0AMPpjbDtN+U5tDG8WqWRsnl2fbWFlggappWYK4eWqPYVEHpTOsmaiIvgCFViMCm
HZIiKqOWI9ERa6H+T1o7Anb+md4bu9xjp9UggFyCwK8uYBqiUvLJwZlze74eRzJh
BNetHdcejVz9W+RQH2YLdgijv9NmK0zNrYrsNRw9H3IqKmRW5oxliRN74SP7E28L
HaMaw1J/Wc6vRZQaL6JPuTVd5XFdoHZ4aB0CC5z3QKszKClIkh7NeFf7uZhq9imB
ndwQbsLdm3hg+M7m2mx1244MmqFpcaXYt+UlOSJBqGv4QV1+tsphL+a62zX3pGWh
pZAQnh32ta676iIH0NxBC++wkaYBRC8yqKMkD/nJjnm3wPCPXNTsApi+9nuRwUD/
nHcNQmH94+ytDUjczM/8e+Ty5OR+hjmTKwLQfY5bNXhITof9vlKVRJ1gbt+aVlbd
9qiVKkhtXdBWUUQurgC3wFJ+pVMY+J2r6M7Vtco4yiPAEOyFbSLSkYhDHbLyE6S1
3F0Ny/OKNI170kSAuOjIcNf/CKGwlDRMshr7GruDf4SGlgHi0Zf4waE+3Yu+tdq5
bqIont8GVpK7gCFnRUIyHj9lh1qUfsZEHJfv4AEKaiJABa9MqFo2OYMIIpxWGAnF
GkvHqWNkfJ2oGDj2pNDYpdspLfFF1fvhTgTawo7Of3DqKRM3KoJo/jjx3y6hlfay
0K/k+g6ac0YNIwtHE7KBvDXLBs5VYA1KO8Ly11LTH4FmPprhCuJOLpri2zXADncZ
wwDEKU5vwH9o3t66D2HAZzQYIaFI+ofQVOmbUvSOFxTj3RmC+QuYEMS+oOTMul4t
jBCQAaxQExf1C8A8VExJHSeKTzX8YHxY+sxnRaIVy7W5yp2TlTgyCKXv7a1PZ4ur
GB7JvTY3MKbB1EAkPKUX9Dp+kvVfjyc3aNutwZ2kikyTXoo9HaCGpcvyadZ8L0f8
4tklccrkEvLmLy5A5q+qiwPyLH05ZYe+XCwU3f9drNamEakSq+DPHc19x9Fh9XTl
i6SS62pmKnSR00U1tqEFTD0WgCrkSxqglUTLC5thJXMG1XJByKObX3DKBE5HruUO
9mD2cQ6hSizpSIN0VEF94AS1MkUwTmMsz06K2C0TDUe2DEgzcWTpZR7Tq0Urbt8r
sMwMrgBGxFNe+U3Vw8sgMDwIvAWInf52EFYeS6T3XTcYTFphaJE0JO9nfJ+srEPS
nzz3zKPBICQuto/HS7tu7IEicRMiJwfDZZ3o3IEMkc9gQEXFLC6ag92JmTt6A5mU
RPMU0ZuiCOpjPMDCeaDXP8k8tF6FaKjNJD5m1Oi12uMH3TQg7e4gF9Rr9ncn5ZEZ
u9k6YO+ESZvnr1e807nUthbo1yF7IGp/esBjM2XgfoNS/BFKMchUe0igpZKAlFse
AWuLiUWxtQD8KuV0dr8BfMzxaHkjzE4U0yyrgV9c1XFpVesxkCtdXuPjd23pQCdz
WJuLXCGxfRoLuhyezVKt+v+hxtN9kpBWXP1ubRtR89CXF/5/j2W8qWzmt/S+LVvQ
ROaINPROhHTjXAuoaQ4jCP9lxdwEPJtu4qhffW6TPgnqLn0pjCT9voBBgJe+XChA
L55NNwT5d6eSV2zyYilXc0cK2TYNWLZEfKyhTWSsWKuOjwU7IrUXM7MSMfdJ7Vzm
pIYk1kcCElIVGaFP2nrW+ipWfDNNBTFAY5gKk3klAY0Q2DA1xpgx7XQRdVGgvX1G
A1eDwEHddknfDji59PUBVzzxVO8mgoBKhEe82kbNJsq1b2/r5b0k3JbQIrZC6mav
P+vLPStn+Rh22dT3Vte9LbzttqNRoww12Pqdm/lILbl+S7UfvxSZ4ByUXn81TJYT
lkq9/c8gASirbqQBSQvcSL4kk71D1qTrxGM+j3B/KSUzHpF3KO3v5EhtSe5VJE8l
0cYj6Z6dfLj1ROM4igfIdU7FyejAopXDm7dJv7TNpiAh/dB0TXoa9Hf0ByG9csKw
yfYt0MK6kfkZnxz2J7NXWT2JNEkqZlj7ieabG84XOkoJJ4mPUPmL/LDqF6itMv35
gkToNBoIpmDRxhOZIGLmyFpYQoFTVcv7oz/+VhLzME5ybPXA+ZdPdtByLPpvc6j/
TNT3TISm07kfZiqhQxZpMij8VQqfnTDmgCkZB95wUBmOagAOes1hgJbYjqZbzBqs
37uoiK8cQjTBq0q8iX6/IcjAj1WxXSpcH/JcXGLd+77WyVXXHhlQ5I9pioIYvUOM
uCvQNpgLojqPSdESeANeFZyj+r9Ale2FaLP0ivbmZxsLnbh6pHwbLTkpjNrlODFk
3K/0zw8gbqBbkw5MIjLzBbzGAFQ0/R+dFSq3FZsTOGhaFs6BbT9as7+S8gXHKRTN
NxA6M26ylgt3Atd1qOejzXgQsaNBZTo+8C4ukgotSnQ2+1DKtjitZL2eCtR9I2+2
L1usHenc0Oxbh5C4DFujyt4lQlwM2wFCvP2ABBrvVieSpW1zPwkBpgs3OD4JbxC0
aTyAfUJtR+ViygcFKbjCuDHmNcxB+WmsAFTQI1R4W7DEjsHrGkkUVkF8xv4e8qZ2
ExSM1Ix+9SzBmzRDl/NtO91RrpK8tx5hNNxa3VLU7cynNB+c7IaN3VhmXPgbsVba
7NGDtVvrt+9OAmywmcUQ1m53yZeCq2f5gKGC05bKXvwPSCVDLm1QSyzNJg3kOwkN
kqjit24gfokrtGZH+ec3I170/IyWZ8ig75ZM1M9zDBdOVlU+Yw8GB2ej/NLZedJD
GVUqkMIL4H3NVaQqtiqhOVfNBR9agaHa46FHJpR5ru9px3L05NfYfJweGgR7nN8J
T6/ep6PVG1G9E/qSZ2BkQctp8lOJybhyhu7m+KLeYq8D28eeiB9idAlcpsuaJibw
Yp5Tt3sNN3G3+m5DHJsI++QXMYUNWFPCTcQmX8RK5rKJrN1J6vVNDKv2EwSB6QcI
3gwzsy0s48xgfhfRpI7OqjmhvASqvO5WDp/yXBVDLRzSrvfpalj0UHKFz7rYaym2
N7oxYmy4QumUJqkATbjp2IxII25EVorhGoN3uN+wEkVHsADfQRP6pC/1QbB5fb0O
zu+pRdud14vtKpcPdO8SGMRIOFjAJdpLTO6RNJdbyB8cA9H73TSo/S0lfNf1LKbU
upOgMV4Wt4ayhh/yafdTsheoxZYTMwyhZzuUHLSAEMVsPDr7jUzz0hlOy90XdNiS
klsmoI8CyDZByS6zzWRYTs1lTfRgra5Plea0MGHTmqAJ/qTeqgh4AUmEB4TD4s4W
jeS/S6qwgBQfUZAa4CUjxfBnLWAFGGJEV8qBFOX9sy++JMImxVr8SQ3ezbqw2ogZ
xZN5S2Bs0pyHewZ9cCfEe/t6Ql4zakZzF1jkDsl9vVy+Bto3vku7zhZg6X0BgMJj
k1c7KHEjp7MTnRWF4nWCY+oywNgbwVNI8H7zEJfFc0XMaZhB6xPpN71E1HjcKGLx
Khhspj92/oJEjrxxxX35GBosc0PvFFEHDRJvPfy0M70pzJYCr4NpDHSHgIHh/N0v
ZgIxLNz1FMVU0k/zo3yigLX+TiqnT2PFIbWd1P3L7pJePsr+ogf4Al6KJApeifWG
gBvB63oacwMxzyJ50ZB1J6AMcBipptL0U8Bw60i+NLgcIzag7+6fcqNBQJpsLJyP
/5p0mW//tPiCMeMVF0nJ2ypscQuweztYOmIXolD22CrUCZkRbPWXepLgVpPSr/Ux
SGYOO5usri9pBx4jF1T8D1UbHn9B88sc01QmvYR81WA4mcEqmVITnzaHt7CdBTkl
bjkS20aIAXZK2/1MaH6ab5xumjljUQ/KHgcamQfcN+Xf3ewE8UloI1k0SlFXSoj1
RyCgVYBc25XXiELPtt+5gKSiLleutRq51Bg2R9QFIBaIj3yPOKADg3VaCsYmEfqq
HHqoF2hNj6AVf1k4C9Y+kDs32TDAgFB5S5a+6s503ocxJusCi0HnBlt8LmBhZ+et
lAUIy2sK3Lp/pKTiD9k+RgOxPNrCCv+nMtH6pMEEif1rz5AMWdrObA+bR9YRGCXL
0gQZrvOEj3xjR0P1ONZvQtlXWWiRjEFxUr3qi7i1ja1w14WEiHlbnYUIhwyXAEMX
UcmOYsnXrKJksx83+s7ITs+ZOEoaCxLZmbfm+b1eeTlUScmhaMANeZ8cGdu2P3DS
ztFmRFKBMLaO6a+YD7i1/r94Ow0EM6UjzwD3eQoM4HfabZm5azW7EtJLNpvUnzbg
G5DY6OWgrtcCnATQUciG9j1wDpkAWLUKRJJeHGa0rWstlbCiKb41D4IPNiz1ELU5
gLZG2aeiHg1yqQFRsoAJ3ZsiCoGwRtmIteX4mUcSQQNTLFL/2etiBgsfn7qYnF/K
zDDUw/bfi6G2L24lfPMSuWicOEQRVJxno8rWZAPt0qm7S1lnkSq1p+TN9jJ8YAAZ
n4As6ldP6pHDgdcFQIiyN2mRVZWgkKogtqJ61t+G113zqntz5w5FqoJUpvgSMQzs
YY6/5QpaclMf5DIFlv/RPG78fUklWSJZOiJ4fiEMYn/PNGBeIJDgpiCoW9iWoiU1
hPRNuBMtHWP9ardX9q2YndpkLs1D+D1Tp2QQJ9zavAmYKz0vNhnjt6VxtoBNq2iD
EDaYgkoaoG6UXDRFDiG7UHf40LfGVW5XeGu5MBjJFDlL+5ACwZ4gj88Wmu5bI9oO
6H2YKbmv27v25u3thPWbTon7MzXnvM80r2wsq7pBlDD3DtI1YzZbJDbTr4yoNe5w
2619CXikmnY89hlSrh+2W9vGRa1UE6WWTOneJrwsA78LfTvAW3jnUgcTyygT1/CO
GHQyk7D7vHA9uFEJO0PRVtfVDolKySQ3AfFms1cpRezwjFEWegqZXbkcJ0FBsY/S
vu9gs7Zb2cNY7y2ggo7zw6FDXct0aguKIgL0MTWLt56GkEIHYu2XQHmTxABEGWzV
6w1mfgpoKj/KetbAvx3+DrX3O58jKZZydV2rolyJNJn+tO3jQUAyWSb8sNPtVbK9
DCsb97WMZpOVclM4VDMiAUtpEW8WUy4rf2NxXncqPWvf9z3s8h9H6+PmV2X63gAx
tbmfH+cgjpuNUvt9U+Vp7gSQ5EVJYukwqjenMawWQWyAnaQ9gfugDiPFZdZNdhP4
Ef7uQ09SZwUTRFCiqPFSJdsW7pn8Q3b6Aas8xtZYCb5yLBHB+if6epmX7DvhLtST
p41fn9HNBxUWaRV7TiZyrBEW+YImqEVGUzimqa2qa5+Js3YUQ0tQoThYAnyn7pno
k/lSqLsQu5shb8dNTL61roHXvGam+GWa1Bw9PmR3yi65YJhuOGsk0H/YGdFlnto7
BySdxJv58V9WGFiOEbrtqQpE8Clz9xnt9K1PtJitaYQsGwXpUsBmPA/uDxHAFhnA
ScGjwuumUXEc1LEbqBMBLRo3Qozscrk0zMaEKE6jLB0xZQniKxgdiO2hNyHl4bpo
bra7slxQRzhtdwyXGb7K252+8WeY7ZCxK3rfo6ccjtWBecY/JsxI9RX/OOe5jkDD
KIQaoy4hMV0mjt5ofye2Yc2AWBwglSkSYdbHxr2i0VmtdQvOyf0gNEFKm65+w5Od
KHMl4gG8987pdyuipCiUxYz8GTa6/HUcQt3dBkEQN/xUXrLq/t2M3YMC7obyUeNp
SJWQMeE3DIsNy3EKg9c57F7l1aJrgsW7xENWfqJKW58SSH19vopKbHvu3I3tEXAX
QeAryZTcTcG1sFY0tZtFGiI5HCwQhEQnBaR0KCLm0UwZ/wcPprbvhPArBhnKM6+w
RdgdQwdD7xCpRyJA6b0V4v9gT7G4PEIeLqfWW2uq6sIWE0WAJHL7f1+Pcibo8aCv
0wSl3TjGlPjslXc8WOjVnkqYcqt4SBvBtiOxCMFSVf+9eoF0kXWDJ8C+eIC3ettB
DjD0plETulW/RXIXE1JURJkmxSriNG+O918FZHcJCEqXqoHDN5VxOhRR8SRICref
VtAUDBkdSs4AccvmKir+Lt0TtlHTRJrxhPlR0iKg5zhY79pWwqm3FMqdHHeJp/y8
HzyomLDeslZlX82w5qrFkBVQ0JyL5eXKpitJaNHZjjRtM6Fl1iE0MKfXy1/j8mtP
gofgc3BI/T15dHhNKuWbSgj38uqoRwPNt1alcYlc+vXTN2S8jX+PZk9m9hMyML27
CUGmwKKGoI3enDx7TqHrCWenEpiuRbwm3JS3VcYhyaP+zeFdgOptg3WvJyDAAArL
IAemxiB/eTxTb5pJRATh61L5K6584CMrXU4nwqHe5787oaRA4oMQa8noV6mh15VK
Kn1FR28dzVO7xPHylLj1BgV5ripOUBiOYDkIdnQyRA+hEMmPav5zDIZkuIQi2RUP
xHYLq2hqiz0Wzs3rDHjvIScxXjE/X8AODnZPFP8ED5d4ZIKlJNVVYP7N1/khH/ed
pn35Yi7a06vWfIoTVK3eNdzN/RChecyDOXQMlobrs7ChZ0pLWEmVHwIxn75dJrmL
KySl4CsH6MNw0oZKdHl1jc0jmPWDBuCj0q8QyTpgUmdWJxAFTTcnimhbdtKjLCnh
Dezt+6NshwGafPfD6GWpyBdqHN+s7wyAsWOyiKj9JoeqxPrUq0QPyuU1Sr/0XsnL
TBo+WQrvu5BbVLf+tCdw8LXGZRNHKnqWcDL3I051eibPh0sKlUbGlfvF0bloClzr
aHjKrMIsNpzxgr/TbBqIm1AbQ/KKtMzpHe5bpQv1xa6MpgzLoV4lZ4PB2zkftVaW
8gi6SaH7rGwEmM7FkvA6kSLE4HsNR7vEIby2lCJ/1lGWDPkWAXj0fBbtDBrUkg3a
fArIc/cqTs+jJ1g6mr3l3NqNFVGZLh1NZZJNe44XdRVlQC7cXr3aJEWtxhTD3SdM
oyjJgXrATyqV3uUY1Ix4LdU7zu58zt3vmjY5gk3JI1qUsiqjzNnTWV04R5Vai9Xn
dsQE898/S6hwPiX0PnVn1teQvGmjSlrqhvge2WH84lZUq16pkZ0zc8SRH/+BrQKF
dAOK4c8gM+u+ktBBpv00JhQfsVbdJYHLI3qsb1AC+VJDatMQ0KA7+T0EzbjtI1SF
dnV+nUGbdFe6IDmyMUlg9v13n5oNVfi+VKQjBFIblQ9HfD40AN0ne6kOmXaW99jj
ljCxnocolh5+z74ljGmeR6Fqyit9BWMObdc1NT+P5hMmU2llseB8PTys480BAfMH
lc9QyucGxlNbqITPVw1jGviBdGgn7dn1PObbNRCbjQN5LXZxmCgJKl2/OXZEa5r1
oWZMew9KLr1DT0AGjlasI4t2xvmVQ2l6GgoFLDNYtm5zLQZXaiK9TqjeokQrDT9h
6YraJIMlWeK5qY/IdiaOSIL7mvXoeTXvGi9FtEKxzZUP4T1Gnyd1RVJJfIgUyJ9l
g6C8NrEjImCNBBwFE5qhLw1y/fyEtESJ+0Ksc+y5LojFx5jSasWC0SDeVZwp1sYq
J21QViGBND/bfvt/RDXABFcmEK1groTs4UJCUStguu4dc65183uCMJGnuEEpFXYV
bH6E8xeb0nhsV7S+vIXOWUAldDMX3ZF/zPklZAbKUpZcj5lGv7pXlFJk90359DGl
6n15gwKGXBZFRPp+rC9R9vzXcWH22e5e5agqHW6q6IIp/l1dwaYkp1zfQrAxk+kC
9vxAl6VrTMp2d42mNCSAS1jKyY3ITs/f8AsupjZLeHmsLSr4v31RtmZz9hrhkF+9
nzyQ7X5AeVesWm2qzbEhjs17DyVJnMJBzzVr9EZU5K5c4SQS3+hbWK8nrRgZG2ol
ZHPPHiUEU1PiARMW6Jmlb9/VDBtJl8bz01DoPewZYMv5IcO9PS3nezy/2LvUjoAj
l70AqoHbYe1/G/lyChO7rY54G/jb4Ai7jZ7i5mJ7+qy3tOxX5rLn8PNYrsT4HJzv
nYy/9tsbAYkL8LT/PtaV39kpZo6hReICM6QufEMUS9+rcgAAwKKWyx6Mz0igOgzs
ojpuHsO8Q7rSQQlp5iaR+wbgR/B8CTnoOIUPgNV5V2CFC2EPp2vUxCZbEnFki/Hw
d1RIR8rdx3xjhslGB5sk+PbEBMDOHqMRkFXdunsbJvs=
`protect end_protected