`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
ddtXksX2+yylW5zu6QL2Lhnb2d1sD00763mmSITNX595NcHTEkwn0zB1Dry37fOW
FufOhVzEJp80NC5qZ/+F0Vk7Ik02dIR0elf3clrjeJRK85K4e3Hoo4xn7YbFUIms
l/8VZSb14+JVGURjfswrIyCUotIzlzVYZ6gzoZwDXIi5gQIBf/gI+KxNXPaKV+PQ
Ufys/12rjO6aI/pPlqSm0hCvftmBcnezN2hk1UeXgOIuKZnogjOsf0iJVX2aOOWE
6pD/psybjbnsNB6kH5uFTA5frkzIzkzl5d9+YDm9OyC+k84E83I/7/j+rk4L2dah
QJOvksSIzN867/4Qt8qYTQ==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="MvBXkzurAa5VTw+1JJ70nePUfoQXBvZOku/SMmg4TwQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
oRtzZL4VJ4iwysPsC8SXYCzXS8Fw2gtZTOskLcDV+1B9Nzn1zTyNtlo6lNICRmmK
ZRVu2BmCc2G+fmzynYlNTnSa7C0Cuel6FYpxCBlOuk3OF2tzAmLAuDyOH3Z1Yjzk
a0aHuoCdIRKv7BrZCdALt03JeUmXKPdOmIlkVGFl8yw=
`protect rights_digest_method = "sha256"
`protect end_toolblock="Jn9CQpRhJt4rnzZPRk+dOpzAubz7omckX1MrFd4p81o="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 3184 )
`protect data_block
gD6l00tciPUa6pDNTk/+t0OO0nC/UTtBwLB41d4inuAUA3i/ALrNyoJVcBnAmEQW
ptbcNp5fxEUJjnOxnedyZEuEBxWRieZFQnkRdF269oPC32l3y7dGQrG5H8/MtKBM
3ZqcaC020GN1Dv5vr5CTCTslpVJG/ZHpYK3Xyy2RYaSz4wnUHdLti/Ama8bFCqA3
vwdC744sHTVAxLlbz6Bzjy/RdJY23lQ2WZVjAOldiAEYMHvW07oKkmK4nLRJVFio
El8HwOuPG+sYzEzF9lGZdp49Isb2umlxRs8vmljjbpgUugEoanq5YZdOdnqnxlSL
IqjRvnKUMo3en2W4FMai6sK2PULn3WFFI76bjb30McCYiRYeKZvLJZ39fxeuRLNE
1M5mjBfFqGEqDmBz50OvR5F1IfsPoDdeL+PEp07Q3Gb7k2SmCsrFJZjnDwnsYwTl
OOceL5uTYZe5sPNBa6fjSdSQ+xpUOgrrdADZc6RcBv+sIIXUJj7SB6L3pvqbjbBS
kWN+8e3pi0Dr7WWT1+jTGckcLUGnq51nh0R1PguUegP/L6cstS7MuWSHGqnGkDiq
KFT3ch/iXsweflVhrFAAwju4D7rx+xcmSv3T6hnhPh/wampMQdk/Az86FaMBY/8B
LDie3Ye/Qxr6q6n6AIFeX0aAmR35iSWhQETJQr3988oEzBG5tOhvfVscclAElnX6
UpHvd4WicASJUmGepx/VTbjqMacnzV3RNGlfdlqDpaj+NgMyjqvOHXNdRTTJitVI
HrC0X9nG1JcVRKF+mdnfmLk0nlj638Yg0oIR+kAK9ejM1PMnK5HY9JAN9VucSf8G
bcS+9VaNdhGK0lq1FJZGQG4B5EDT0+/VgtZwomA2nKyKSyV8oCLhKnrzwSfK0i4b
xhB7vqlXmD9giwMtkLpdvXsUCG1TVzCAiMdQR3pbKQK0iQKhfxT6WhBhK2gVyTmx
m1Av42Vc/yh+Dnu/K2YJbDqCOIQBlSAHBtpg0OOme3+w23K/6kmTzFaUlvuSVFdR
lfX4lZwNlHECcFNHzMfeXIoJkbVETk9KJU2nfKBtMZAnCro14fkKj4XZ3AWjM090
d8SuhHIbkUvIEmYcv91uzD3frknSX+toYqjOxnFGi2a0cR5/oiTHlWwljaJ8kqMZ
pTAQPwdoSMyVTD7NPElohA7JJPJ1mp0T06pXNaykucsGmf1QKSYV4qLAmgbs5Mtm
HkyUIxt3YHieKaPyU6Ali3JpAv3dqXG5614nv9IIkcbQFDWCnRyq1gW6RoBmZuLR
3OvRxnRDFnQWZWnYyJvYoRpbGvlr74iNtIWyXq8n8w1cMjSIWFwfN8B76Pd4TRIb
ywB6XSZSVdPSHxJPFewTF1UsrYYuZrHBY4S6LlwwVsXod7X4TZiSKcmtIn/OnjJl
68u/CYvx0v+MuKv8pjh973DLkTJaPJEZgBsz3PlFAiAKSdaYEpS4bXgYr496vEWS
prVQ+LJ5GxUKHNRqnpfnrpxo0FRd+D3J4T6snOX5ypFkL6WqXPEQC73z3aGNgfxR
N8rwn3u6LX33tqtPyp5Tbl6lPkbiwPmbcF5fapnTIAW8vmPhjFCGztBYT26zNCmF
65fzqvodpOr6lQAzKL66x628cKvv4PIdajn+Fjm7NU48z/CFwjBePYdPOPZzAWJH
iLUmRw6GNBdjbeWi9mz1l90tbepDgY7rG6NpNg3T5BLAJD8txZYvugRVGOeoahsM
0i6B6U5uOOr2RuTkVRMa2dt+7o/gEG7RCdeth1DfS/yA0ozn9csXipW9W57R2bdZ
AWdev9ecqxYKD0PiJxpdqJHQXmUAdXXR3652lcbYteok+h7O733i7qrpbfzKUsum
14Hn/WQqrIr9W1J/NaeaCcTQV4iSjNwqmo7iroHX2kRhc+QT3WNqgNq+TD8Zl1yI
KvRspZrVQydOkE2zUwtdkVPmHNQnjmVXoAY2F7Y+xld+Egf9Mg0gzO3UP+bz0ZNg
1wcCV68gq/WF/5w0v4P9UIBNAV9789BAeXTWeNbf/9DilTdCkW0O3clZ3oVlDHkP
G2z0Pi9TEhYiMB9H/iaQPIyIIzJPhdaWnMsU0VPNM9msmXBeWPUeO85ZhKCihgQa
N8Qhcxo5TYXYYDP9mate+lsKGCKdPRP4Djce2ZtFmoya3lo6DV7XFetZExflRUVw
jZFXy4p+x7NoN2DzVHTs9iZ0+cYtTpcXxgNyqUO50H8fhN+mk+8i2sV4YPaNT8aa
yOuf/UxNTXmSgyoKxQg+y/jhAr5kJGSRHzss34mtvR9b36oCgpcwZXcc2JjmVTrO
vYj2ud630njbS/rCpwK6Jhfs1kfU9s7fzLkGCbZxQ15p89FcH8gixgDpKHnoU44E
ManSMNSmm1BbOSk1EN1kcxP/ku25wK+m1KwZvCyrGL9+cfgEEdRnJmIUx1wHdIqd
Vsi10zv8L4VDUJrqo+nKzpsAnIu8jfaFZEmwI3IeWIzpI3I7ODAFNhQ0NUCDpVVR
d3MWZFepuskGvdMNM8OWlOb7Y0GfXXtKWpugI0yR+cmncYgH4Oqw1H0QtaqRtoEP
B2z6cJj6+pExetZ17iFeU9YJK90lEaOb3wDWUWMFck7JD11OsDTjJdOExaqSQx7K
zCdozGvhQ1H644A/OqR9dSJgFyq2k/d7T/7NXt19GKCOaooQO+H+gbms/vZtMG4E
scAjDXBXre+RcX+KLAIG4GxsAt36GJPDUFtXevsGtxxczfdE76daVxQ6zp8ik094
IU7hDC3I+g+sr2TS7nwVWZqukQ3sFfSC+F2LFJYYJkJjD06qpuYgRNPvpsRVMuMh
xZQdFrsJfuLi3vFeAfQvU/teVrEWrz+ykHteypa9kOtFcGd3pn3M6n/BV4B8y8AE
RpvyTUxWT6cb4PuZ7OeuSVdofvbe7ZLzKgqRxKDFxxPEydsv30pcJOZ88ERAyZWT
czfctRKBMpi4bInVBmwZYOqR7Z5joz6+Nmf/IhiAyToXZ99SHHQ8SYicXzg1I1ak
0lfJilSao/pGOeJ+PsrWe1I7xzsZ7c43PCSY/rJ8aW57djfXvFrqY09q2ZnhKdZs
Jj3u6mkSYuNaUEkGjE+fA1/6ZDpOZK8N92Yds4l2MR0is6DmE/+0Xin1Rt+6EE/O
xgWWeUlKY5cT2HsV7DyIFpc6FY65go5yjUyCSZL0qAVdymZ9xFyYem8L2+1LNmMo
qFewpF1vbwT8Kv7vlRgYX8Tiap5a0uZmxk+RnMx40RZ4LqskJA7SdPemfJsvNtgp
wmuMNO7eVMmZxS76J0J1TuB1/1J+lNPUKA/WWbzpWU3wvOElk1YKRgudzquFFEBO
YgF2znlY8y0ZQ97B5d2/WR24GGeNi1PCYfiuYv27FCxryT/Oq95YlcsfmiP1DU4k
bZ7cqxbBYqVqQgfKwvgCkZO26yXw0kSYXoPHGYg0i40+V3Kr+uhZ5wZKrJiSqcN2
PTegostGVVLoHT2rnorqVHcrXaYIExDOPBVQz0nIGDs7Ja6RhjhlzWp+9db9Jjvz
dDxvI15SwCoYnX9lG60wP+9OZSz4ARjdFvurQdZZaB4qq5fJqh5eVud33CrXpU+V
M0/3gWqeRPERmbD9d0cw+uumTeQnlUE+5ro1wrSEoC4FAqWu02LsRLVx56wNJPBr
WBqfBpYClHSPD77JoE7J0QB9Km8C0b9RDUvGMPULHGz66U3xysfTEZyqv4Y5+U/1
qJ656qqVCOWzC3Cc/ku1faXvHcS025/fiEN0yfHNWCpL8DJaMJirgLyjFANY0J/8
g2jy8scqSm5UFpKXpLXFIJkizCnBJ5kgwfEXkMAOGOrsodBh9JeSMWB+cloC693L
4u8jy/Kvt5u3VUJ3FSYvjutPG++QeiG7lcgpQxXRxYcc5vOEXGdaiAvAyR/T4xmN
ZdmZcDGuKxp158A4KUtp1veNmxFuXq2QkY0i+T1Cnb4B0wAGZCNp8yo11DBtF66E
XF2EXPrISLPJ4vSvbVphDsuar6/dB5duIeunnw6x0qSe2OpCQ5IGekgxx2KITxge
8Ld/pPw91hC8NQTktmTV+nqLEBUw5ZJUjcQzfeJS+26l8ILnJa47c1mtW3LXyhXh
bL9HyPY1wZ8DmqIGbYU3k2m2JuUoTplxPf3JuPj4LE3N17WuM+HqEPy/zJqd5Ur0
a+jla8Suoh5LZva628Td1XvtVCH5v6j/OPLK5BVPZssUmLhIlks/O3GJR6oKiPLP
9yL9YtLd+zUrHPKCK5+eZw==
`protect end_protected