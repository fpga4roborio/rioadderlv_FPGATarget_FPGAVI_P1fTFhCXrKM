`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
ddtXksX2+yylW5zu6QL2Lhnb2d1sD00763mmSITNX595NcHTEkwn0zB1Dry37fOW
FufOhVzEJp80NC5qZ/+F0Vk7Ik02dIR0elf3clrjeJRK85K4e3Hoo4xn7YbFUIms
l/8VZSb14+JVGURjfswrIyCUotIzlzVYZ6gzoZwDXIi5gQIBf/gI+KxNXPaKV+PQ
Ufys/12rjO6aI/pPlqSm0hCvftmBcnezN2hk1UeXgOIuKZnogjOsf0iJVX2aOOWE
6pD/psybjbnsNB6kH5uFTA5frkzIzkzl5d9+YDm9OyC+k84E83I/7/j+rk4L2dah
QJOvksSIzN867/4Qt8qYTQ==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="MvBXkzurAa5VTw+1JJ70nePUfoQXBvZOku/SMmg4TwQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
oRtzZL4VJ4iwysPsC8SXYCzXS8Fw2gtZTOskLcDV+1B9Nzn1zTyNtlo6lNICRmmK
ZRVu2BmCc2G+fmzynYlNTnSa7C0Cuel6FYpxCBlOuk3OF2tzAmLAuDyOH3Z1Yjzk
a0aHuoCdIRKv7BrZCdALt03JeUmXKPdOmIlkVGFl8yw=
`protect rights_digest_method = "sha256"
`protect end_toolblock="Jn9CQpRhJt4rnzZPRk+dOpzAubz7omckX1MrFd4p81o="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 7152 )
`protect data_block
gD6l00tciPUa6pDNTk/+t0OO0nC/UTtBwLB41d4inuAUA3i/ALrNyoJVcBnAmEQW
ptbcNp5fxEUJjnOxnedyZEuEBxWRieZFQnkRdF269oPKuKAsu3igWd1+dKtSxJ7R
AwCTdf+3PkcJMYJPRX3VlgnXWP4lovGSB/4EFeyOLZ1A8rP7nqeh61u52GXFCSA4
GqJsyKTWtihvhoRb1cCIZ6Mhj83AhcOCAE+5hI0DZJiRiS/pVE+yr7ruePZvY3kC
VJaEXofULLoI8Fnui3qfD91cLSgg5CCqFzCRb09B+CxuRXH8SqClnKEWFWrsyZm5
vw7f/1h1K9I9TDlyp9qe9dYSEhAtvVTSa0sMk08QnfatWI0gK0Ol/WUdMdxsuTYI
+A71KsGyT2ra65ggeJTvxtD3SJX8wbUOqWhufhWHf0K1HpAxxSFb5nmVnkbc3jIC
lSzM+4hSZ4fHmQwSr/Z1KDHt6qVQICqUjOQq/vZP8NmwXohnz1svwUAAcBR9iC2Y
eP4zdBKghcZWC6TRncs0jzIUN7tZ//CBJqwKnkpY2/4+v4iTOwgtpwpSTjlnl4Nk
wPKemvGx9QzAr65DED8ySWBJeei2efrvlhe1aemt2P01Rm4XNI8XVpNxKCyZ3zNL
JeF8MWgLXQAd7p1aCAQ4Ll4lBO/YKOL/kik8x6GF8gFugH2v6bmwHk66o3XQNLSk
qJy2A02LcoL+ijbDtDZl3Paxqqt+k7ZhkvkiIzw3yLUWvlye9SX8hjxJZNFLGvAR
4XxGC4dGDfJQAEQ5eS+bjeSX24VMkj/1Z29w1xQt3uxR/Pr1pp6frsEZT4Fp473t
eUne38pC/owNxC5QwqlUUVOe4P1e9g4/unkq1Sad57qIVi5u3Sn56iVGdFfpXyW/
rZLY5u8ibGZUMNYm+3AvF6p0ZsvRL3Jsf3NnXI6HR3FX8otBBQa8mf1Qnd8gIvjF
7HxVWCrYl5hifyn7GycrrBdbxa7o5WBfR9+cIBGA9tb2gUP1h9izg9xU2Ah/rgif
h7iDFoIAx/dHdvln3mplmx3D1M7lmQ6+HC37C5QYMnhUM+SdZYRQSI5wblmwJ8pg
GYmH0QZl5SSekW9DkKn13rZFG+WuGaoTuK3hlGeySTImiGE95PiWE5gtNRThnVWf
+YDwFgY/3Sal/DqQOdCQxMcMtU9l5wCEYuVIyZjD0anmS4dYTgvQ5jQ04njXcRz7
RAFWor7IzxY9Fl8Z/tI1IEIh3JmkavyAdiNS90GbCEfAtcFs4Fv1k1+CYg1fH6lR
1TCpG2jFUMQpnCESlzx0Z4KQ/+28YuwsYofsV9IAb0K6BQYf5d0DENdYZuSmje8T
a+webxjJUs0WEJi24jOhwlxoOENDtyhuiLGq/8fDRxrQfiC4g8RZRQgkg2Kyb1DZ
2h0tRWWz6lKVw/gAtCgJVton8IZ1wVcNWtWwu9cYUvxSGZH8f0mEcriw285e012l
FP1+lIIIkt0f1hb3oqj19ohHFtKGyzlKUAFk2moPX/os+xTuD/eRAChDaS78JO/F
YVtTMqG/8zC1QbFCHwB5hA4lMccX821Cds+kNTQ8nJWIWxAV34gx6VyLo1ljhDX4
7bRWB+RqqDkfDDHfEqjxzJ7TahzJr7xftXcUKTqJTRePvfR0bC58lcjTPjDqlsp1
NzGTJfzRecEi/uL2j9drf6pnO8orO9vi2fOu3xgLoLXh/6/nslXDXONBLqxWOy8w
Lp7W5SqDITN9Ug70U23IkQdxTYzkw6J0ZHi8ePs/2rbeNIvt1G9fdFudOiFC0FUs
VcOVwqKpgjDNWpd+35VLN+spacQI8y2xGyX4Yi7HCRYc7Xmn+8SM/wVp9Ur57zSC
e80805OZ/CzLfytxmDum2AUd0ZMuFs1f6oZfZ4AzQX5wygsha6u0Rrz9iwRM/XmJ
A1uwln3ZU0Jh2shaYFrkFsAeoiCwRCk4sH6kIQpLikLcWxuPoecTT7k7cXCNiB4L
HbvoJJo4AAYJFFHjiGsv7ONLYqf8UoZtUSXsTfG7/fNCA+OQMdq8Akmzr+FOZPYi
uETeZxeUK9E+cLeq6GUtPesfUn69uBfAJ9xYfXHw77OSMjfgnEsyPWule/HvJQgy
N4F2Lk4GVcVVVs7LY6yK3tLLwJmpgyBfXKdXlpffy3KgrKoRc3UGaTn2MFX+Z4wK
lUfBF5Ot/AOWXVDC3QC8kBJNJJbgtlA7tttbVIAsluQcIBhEWWrTmZLqzweWcIGn
Rm0Pw/y6na6R05huxoaeORMrf5ubbfFvwkvnAyxAX/zNrOPzWcII1sY+ElUYMErs
SrkQ8FuA8wcgYSJgosk8RDde/lWivyDHmhcb55vdbRvvLezbbcNAC1HyhqGfNUn2
GOgoTb5i1zSv1EJMCyyN7m8NvSkY91GjmycESP+9msfdvshM9dFltkKqVIgmOrDL
JNCmxhiLn/abm0a4NuRY1Xvrd30/AY/WMARUgYe/soeSVqxDR1fgqu7l9qFdZh0N
L+la0BW8uUnxO+Tv5ddSQz2iGEK9sCE1tdd4kFvFToQtQ9BT1POQFl5TL3oS1NgN
es56gxZNMN2uXDFRj6YtGucI3CSFfat0BFrBVCBjB7aVux5CQ2Z42tAU0uk8ECUe
Mpn47xaWYSCgDMVrnoXzNJUqfc4nIhjd5dCHnhYGsp1bDg4/4q+tAQHS9UZwpwNP
Fxmy6pVKngJbeoHMm7LVIwzdxym1+qQaBl2aVcYd1m6O/9aZp8q42OLrJ0s65iLF
nw2shcBNJ3j/LkcrsB3/d2LrtlpDhGqeeqZIXID705iX1De15DCVbM4RTe9xim5v
XTnALsMUa/nvMokSoSrxzKfqgxiIXsJNUAZfTrt8hZK1iRmijthBEGorqBfvLtyR
9go+d+p0VNVIloAONjMLIjMXpQGffi9QFY6LS9dngcK/Zi0+S3a2AYgkRnnRcYjV
C60DAOl6sS4DHGsUvfX5g188MsN2yZ2T6N8slMcGOCYDws7jgx6nfcyC+/tW3wl4
K1jmFkxRsFD2HDihWZgIY0QHlb/6yhq634BZcUWosXwZ3B5U51IWi2tdNWqkpY+T
33Z6UmbrxXCeGvjW7UN00nQVDjSIDSwDkxTD/Z/loz4eVLeL1b6uL4eN6qFnR0G1
enPC9mU5m1P4SRiY1UMMoTr7Cwz784jK53MzkDjF8HqnR4e4CRVnl6jb1U7ZEIw1
eFZsqQ/xvhKvD0gx9JDQk2hVqxIFkR+EgLJUj9PPPOBtcSzc3X+kiKOVLHQRLgDo
avOEPjmbhj8MpTCDrJdpvw78gGH4T3BVtG9fFuMf2u1ZwXcjSBRatg1jXn59oYBF
m9Ny2UHjtWvBJPSuLwSP6ayBkO9zdzZXjhXj2I241z7EFzcAYVdsT9uyH3T2tR2x
DC8NdZ/UwGQGXUsjYwgsYhxgb/uJbucasCTNRiaTWGVqK08v+nnT5sDm7bh+TXdD
lvmE6c4qS8KsuWzo216IXnx4VOIAfbCTGImBqrxj8O7PhfnfEHgpa1XVXKYE+vb3
d+ImuZxsbDzX01XlRCpklBRiAw606JVbj71i8vl9f6pyGp3DVWSD0pTCIEHZt2eM
xbboa2nQrUBXNzvg1nB9Baah9q/bTz+F2rc8NLKKap03YFSWPxDSV4aBWraJxtle
+FoQOnSZu/AoRnsk/+gjqCWd31zzpH0GFCBRTF0DMXKMh7+viHJSqO1q32OgJ3vU
g/SdXRfQpBnPi2IX//io+HAJmeffqeSaJb7M5vCIrdyldBuiTuwybRu4QVPF/9+I
8fUwAW2mmqRjmkf7mkWSitwuNsHad5XC+vmHsZz368i1j2VVWV+7z1PElbqT4Ho0
vgrmO1L6VvYkmUH5FkO0okc8RwA+vRaSpN3Zs/OXxdqWjn3XBuW95b6mcPOQ1wsp
uipMXQWBU6O1qPobel9OmAkv89JWpEn5EqqaFiynKFxrtZUWywHS5IRKrG+DkHjC
sMC5bEB4lJxDredEaED3LM5offskqVoHTkgNlv2lircg8T1re51OG/RN7mDg1shg
EN0cPvu0C8rNbWUqL9COJa6mAd+4pPstFavcOoAG/JjTFa/udBSuv0B73ZgCYoot
X7QXFGAeatU/joCHmnCTwzzIGUJMJJ2KwzDmkVJVlDgxUGJ3IJpRF0upI7s7cS4P
4uwHv8L+TX0UtFrS1Tru9iHLqPW8TmMK2J++xMBwaUh/ANvY2SMUpHXoQ9q+vCSO
t4coo6yMpfnOzjffRJqzEXHKdL2Q61zpBvV66bBacSNuxnjGgLk3BWKRjHZchQSm
OHPX7swze2G8LUXNjhgByCs5qk3pBPzPNLIJFhyTao5ZNVn8IyeXL1uBMIpCeu5X
ULZlb2d9JofUywdkuYa57jYwGU6qBu2Ue3Hs4MtqUY6T9cfZlKjIdEG6Xq3TdCHt
/s5NHXWpimdEDR6D/yqK+pa4yoXzxuGFIssKy3TWhZs4uSKjKIhVCr5cpQtUa1i8
JHgB6WbUe2c8wKiL3OHaZlVo4NbFLxTZyEpT3BHeAGlXplSiIMSczAIzm9J0R7ho
twOgY7LmY6nKBTS/nzDPU5zf/FJnT+WnbIvmXDMXKPtH0/ZdElZzVYu2//1mmzOd
zS2n9ri2hU8uNNdjqVKJlApRkyOuI1eQSIGg7Ifkwziw50qJUh4IQG1gzL6s5kW1
Nex50V/S3oNCXGyRvmGf0HnuZcmHpuMYbboCX/5tZFqhVahmlww6XKk2q1TE0QwA
GS85jrMeXWaB2k11VBwGYS4x3ElGPifsdGxvDtmNwZIy8DkOHv95LB+2nGGhcDMp
JiLOWRWqYq0viDQL2IsoQEdvPqA/oNst6yn50L3IKfEU/vf5S3tJfd6ADtgvS5JC
uisn7ykuYuRLXrXZ7GNsRpIpjPI1PvWLnOE925fuZCDAEuHbJyYX0Hwydr1p9GYc
1bBpmbQsZN6yMNsPzjvddLX7HTY6qBvyFufZKYp3yFDXgHV2leZCq4Zxp+WHyaRh
7IJXeNZ9H3Az8zk8Yhl6G6fMYq/uy47PEJBvNeNmkCdlo5AILLchx33FrIy1ZkQl
kl+EN7GLbvQAsrEdsHIpV/6GA2JOzLM+6lWMGJwXhzve16I5WJG8JQRuGmDM2UsU
3CA6G9aPNUyiz6bma25LS4NDUKzTG5z9XAmAXJiKwyRJusf9s6gOzpojGbpgBO9J
x6D71bmoYVgdsa2gN/OgC/Hunubz97DIpxF82vnFfl0tLp2W5hvGAefPlprVvA6R
owocYSIspqZA4Lmfqy/CrfMK4EFYquz8x9fxsTd6xfSacXEIvd2DxHVML8r0lXSn
sLIhmrBExg8RfBQiKr1nEYhdqaVCF+b6/GZamWkzX6hAdGfJNE9O2rXKRT9sF6yO
zv8+EBBxy+VihsaDB4/K1uMKdujW95KKT483bXhSRR4w8dVHB+w30+SyGeUc4VVU
h4nWKsycuFiOWq1hOq0HWhqzbthUPyip44hPWSgEZ2DGjns5AXIX4qs0iaDV0fuF
JOm+5/r/uCQhd5F65QCUrSoHBkbI95NgpUi5r06dTXhADG8A3miqk/nRTLQyaqiZ
IGsGkFRCus0t/YfbBlno0/0+9MLgACndYIkoq8UjC46piREHPU7+p8YuklwHuFmk
7j/1raLJGNCf+kg8G2YHi+aq2kz1hEJiIxmvJcMTVDk6jzjl/MIcb4zFW2Ci7FCU
7wnRx+UmW2YpUyRtE9wZDEGB2Cc1YHdPpvC+VqH72jCoumLxLT2sJm587aLc/ppe
6b0tLkR3O0pa/wKGvcc2spa9WA/0kQMcIRUuvxJRAat9EyqbmEI03ZCgHdAhbSUO
3tPLxbuELQN5kx9wnKqyCRJpomI1QNxZVUJryiqkLR5M01tnFhyx7QoOAMu9cRtj
RccC09QGoy5gD+DsUrsOa0W8F5pc1u5zmJH6Iyd3EpU2D9LXq+r2QMySbst8Pb4k
q4TUp2Wo+JioiRlgHvHBWQmuYCp0V2IMf+mztPixBJCNU4IPHBgztQKzy7EDUVAk
TQ9uTwQKlxW00eL/md12ViSw+76s5DOPwecp9GLSgpjcGlQzBvN2siLwte0AHMzd
AcetVIYorlYnZ2vuoO3E9pn/rDqsMQ/IdN3JulnAm9xmxvT3RA8vuocZmYe8YiAg
taaJk7OlpJQ3B5wPWLrXepPImr5uFHKEhxWlfpSKkI/cPJABXXPpmCblbtgqz/sT
IQYP6uUK6F+0Wx4tagnyabZ+OeCmwdY2GgIfi9O42p6h59WCosaIxzcbaXbvtmEs
hThAMnF6jUDXqMLT3P2IaCM7VRmIMZxxgoXyAJG29gRVebhBk+3Y3ZV4+a0ZTWr2
MgcMV+p39Miq64cbLDiPabcu+Zyb9bz0ovpyQGVSeGaUb/n9bL77QJO3i9BBAwES
8dpoIotCXc/+h9foY/mTMhx0gqofjuuTW8wxr1ZySuipaXVNP4UIHhCKN/ItPi83
FVlzrYWqVZ2oSWf0dLpuB+FzF843hgZkw9zkSDOFKJN1uTOWzh4oMDVjZh81hmTh
qRw5I7drT5vpv6o7W9l9s5qNByNHraGv57TauS67pmIdjmr5FbQHrKJAG3cUmByE
/Ml2mryRkpycTc8EOM6ikZmrNcjKHAj/qfge7C7Y2P+bHFZVv2kB5rzbQiwfchz1
kiTyJic9GupWWr083GSL6yYs+PUDo/k4zSGx5j/USb1hLDrxdaT4edee1Bm3bh94
Pt1cSXD1PDVyaUHkIGlvV0mBcpWtmM1PxCAEHRVJY009c/s7ia59QLbUk1Mt84sh
wy7Q5lRgXWky4FUmP4/C6hAMkG6hFHlz3G4IJr+iVBBXwf1r8jnPtWuCSmE8dSgr
4fNLta64560iKCte4u/6QuPX8AEGsUS72WQK2zyMWSIsZOiDkWJDYSRb0o7i50Wh
nHZ/aYSGGagEpGCuuOkYVEj5dqT2o0TJdGaN+rq0psVO688mj7Oeg8lFW6WzRphx
0JVo/Wyw00sPCoYhCTkXEDyyzUjF/aI765Y9ih+jPGVaMEiYWWva+maxBalwsD2s
Zb/wLDcOJvKlO34ITs7zV2r7gdf1NNTbapxeaXf565AcYcLxE300eTdAxglqoXaF
HIewhqBQ29Ue2hlIjlxEkcYEvD9KE3EonaBU7faEuo90Oma/MQu6jVoqJVJqPy4P
zG1++JnjoyT4MAwn7Ljl2HYhSmJnnqNETMi1fwBZnhwdrjCf/7Q7QWxO6rwn+e1q
sUgQfuHqfPQn6lOIfaCpib7JgR3b6W1W9prqR2qzcBXPmEpchhIf3+uwCdT0yUYq
tfUHvGgjGbX2bvrfHHQoeICOi2qGbzWvF+LdJz/rpIIOVeVSOI6n7Nj6FFOqxX4N
Ygx6TC76tcHEGmuxAHBa8Azx1jdqKTGH1LmRffJDxd/OHJFm4MDAt4sSVJD7JXeG
Jmz7Pb3PQGUBpLF0FKxGirBQ5Z+uOyi7du5bmS2Y4S+8HAG9QAzwTqUo2HgVd62l
NRZlHqnYIYaKtVq5/pN+CvxnOQEevHGm66Zf+WuGXKZAyTLSmDoTRNSKGXEil1LB
p/92TzxqdP4Id0afTVk/lw9b8o26ggH0yR0l00eNnMseBPPAJnZvDrVIOxBCv8Ts
/3R0+u4VQhLlUtCSwmwI8hMdFL9i1kSkNEcLQF3RmgTBf09NhPVGGGCSsNlFpo7n
sCEbTd6u+EJT0YMfwTXVC+RshSRgoLS8ZNVSbT+Y22lWAiVArp37ZRAjF2fqZW6y
MZNerh2baOyAjiYI2VajxL9O1BO+h+2HGtsASXNlVysPQRvAiwOOiuSnPw3FHDWP
l752IJHdKJPMZLrqLF/NFVKiWokoxlu8ydmvtcidaR+4GfhwbLsvRiy/OcJ4DpDS
nDNba/rjqP8I7F+2F0Q1DRQgA6D4BooEICqnBS835TataIDLnMxC52EoX5P70u5Q
0RU5pZlk3qYMz1hLACWDhger6ny0R8zZTrAE3hYSVhfqw9Co9k7wQI1djCNz1Fbt
TcELk4HarErCEt7pdUm6s3bF/vgzxlNInZ1IIWJmOrtB8vbbGQfXCbUMIwu16/Dq
y8ZzwiFUCwBzxIE5MjGfPd071Ii1YWX13MUNcXM7RMeh+b8EfSLPxNym+qfZyb+M
JY6pBOumCL35REYti94iCaW2f1Ni+mp2XD/6p848jIYvFNo39RlXKs1cjNB3znyh
mMfIAcnzlb9qd1IgcTYxxcteZ0rnEMV6oLB4dou/T4KBq4NASAdeHg0kGw0WL2wN
Jhb5cctPEP/Ncgr2LbDz4BpKnbvDMAGs7ospZdcvYKF/xFMU1RG2natTxa5RlPVf
q3w5T9miI1hpdumP/9J7poRmRqHADEC98ztE5qfnCJYxaf+XuFw0OZ1M4iw23xI4
08hAjeHyiHH302iX+yaQK6gMjp+wQ5URnh5G8ozHqqBLDY30OqhbybyQVIIwnoF8
ia1LnBFRmxTHic0qTNiOjr21OZ0pG+8elw7PI6THO9VRjKJVmuqAIxVXQiQ1uunY
rK7wS0j9KfzAcmGyVpXzrcPOhTbRISm3ADT6wjIecm5VTwYJKULVKyYxD4M5cW0z
NwACz87WHPzInX80/t540azP21GZy94oh5F4I7MJ/YGu0M9rxjJNs8VQ0Fxy6nI1
242h0i2h7Kjkqk0/AsW1Uw8yrTdvuwYf2PwBS6QFJMPgipZCfNEmfXCH91Q86m2j
SPMVuy4d9b2PQ7FbABT8gV5xIDKR0Fq10QC+df4vrPNxoJcLgFxNNWkMf5o1UOc3
V8zeTPS7j56JP3ZIR8ESoYs8aZTCzqrxFWLZ2ORcERF50f1i7NX0LWdlSXvIX8jB
NWEBYu5ofToVxL6vjaiqWFmsixEPn1fgL+AOmBjVWl2xv3a5yiwHdZ+tTujCtWfy
qd3gbl6qHNCrESSEbYLapUel2txjukDvONFhY1ywL/0iTrDfYaAdE4rSs6M86FW8
xzgZE9emAntW06NE0FIL7k8AzYQdrVLZfQMZ+y2B0xID3hAfgm5jWiTN8cX8YPcY
QQcdN6PjWR6ATFmC5ZEeHCMcQVMCwvfvdv0QeRuvKmnPXh4RsogdA/8+IK0o4NLd
PedFFy5Opjj9awBlXMhdijY+M39a/BxXKO4JS9LYAI86/oSS4p5xZvoHyc3PRcZ0
+OieYRb5xFZxVea28GHt/sD5FULqRgfcvvaXm9OH9zG+qA8WaPsuPymINPRmHy3E
pPcX5EHgDtHPurcf/kiMlSH1YpufdXrDiBvo9sB2jxdtPPrXN2Fh3g+UFP4eD8iJ
Ow3RunI9sGcOmYltYJq0PJTDRDuAxYPRmkmD4g4VYpf/27nvf4Swr11q9S3l8zyQ
7nDfnkQQXLlcI37mP+BDFLo59igmEO494tpK8TDMRyfcMBakrSQWSKJdRpJYk0a3
xbbL50RY7kqoLY5rrOGNFaFf04WWKBBc6AjpW4VRS9fYzr7ujjwJFtBK1Nc8YFIp
3zgr/9XmgfhRwNZK6VlwnFf+0W5Ep2G8RGi6pE3FbDgj/b8uPuiq6hdnulGUEEGf
`protect end_protected