`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
ddtXksX2+yylW5zu6QL2Lhnb2d1sD00763mmSITNX595NcHTEkwn0zB1Dry37fOW
FufOhVzEJp80NC5qZ/+F0Vk7Ik02dIR0elf3clrjeJRK85K4e3Hoo4xn7YbFUIms
l/8VZSb14+JVGURjfswrIyCUotIzlzVYZ6gzoZwDXIi5gQIBf/gI+KxNXPaKV+PQ
Ufys/12rjO6aI/pPlqSm0hCvftmBcnezN2hk1UeXgOIuKZnogjOsf0iJVX2aOOWE
6pD/psybjbnsNB6kH5uFTA5frkzIzkzl5d9+YDm9OyC+k84E83I/7/j+rk4L2dah
QJOvksSIzN867/4Qt8qYTQ==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="MvBXkzurAa5VTw+1JJ70nePUfoQXBvZOku/SMmg4TwQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
oRtzZL4VJ4iwysPsC8SXYCzXS8Fw2gtZTOskLcDV+1B9Nzn1zTyNtlo6lNICRmmK
ZRVu2BmCc2G+fmzynYlNTnSa7C0Cuel6FYpxCBlOuk3OF2tzAmLAuDyOH3Z1Yjzk
a0aHuoCdIRKv7BrZCdALt03JeUmXKPdOmIlkVGFl8yw=
`protect rights_digest_method = "sha256"
`protect end_toolblock="Jn9CQpRhJt4rnzZPRk+dOpzAubz7omckX1MrFd4p81o="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 29952 )
`protect data_block
gD6l00tciPUa6pDNTk/+t0OO0nC/UTtBwLB41d4inuAUA3i/ALrNyoJVcBnAmEQW
ptbcNp5fxEUJjnOxnedyZEuEBxWRieZFQnkRdF269oMAcFp4NYn0/p/Or3KFPexP
XbRymFxTtx7yCbn6iUHno2ElrwJ+OIU2dTk+T0ajpHl1LB4DTjd+3Cp5vsI1I0H1
zC+hhj23EvFG9qk4eFBiWrqA52nkBRGrXeneBJbLCazJoVWi6QeIOoxawJaU1ZCG
1ptenFuiRTnkrREEDd996HVL6QCYfcwchCm2/4OWKrtfVDhuTK6mQZGKE5rGf921
sozWw3kEnJLBNVAeRq50Ccavrx8sBPKRRfeVsc1CG7R2VJEj3tX0+NClIcBzXSWD
0Hdt6+txOWG7SATEb/AMJxedN8cxCg5twbl/KLllkxFBJ0Knmf+WvZ4iz9ETTgvU
2ntKlpHYc4YUx0p0KIEFBjFi0/c95Yt4lIo014LFygYOZqGK+6gG9UdF4yqAYz8B
UcH590cIdt93d8VahM3Qerxw7dnUiVzgek7cMqWt2hBit779ehxFoNvfO9G1BYCE
EJ1tq/X1E//bD7F37tqO8SxRJgmytGdXnkESrSbKYt9x8w5ZbizYM5ryb6EgM7L+
m3XkCZsVH9fpEFZQWLGa+xrz18pqeVzrle4IrkffsQo79T55SdAC2yR27aGX8QIG
6usjSha6MbB5kQSlxLMHDyOAiV+ZcRVRSdRpZUzYIOwF0YzwMfP1PatXGBJTbzyT
10Bb0+Rkn9jw7kjgxer2CkddpWdRedycOx7MAHzzjACP3ylbWf6q9XMFjBOmZkPw
k1WwoIcNcQgL/YEmCj6LjkBNjHRCylf1QR3VTM5aq9wYM7gsGONYgB4pwpDDhl9W
o6jbJtUPfV1Bn3rNxQNrT8olV/Q/9UBpqEQKL8ke+JpqsdosgiSLEp9iBxjgbtXY
l2yOeAxqO5d9fgSTjvVJhFXxeWWvDtGrSBsg/UKmvJpt2m8BHACo2Cy6eMM1TYJx
R6Y5G7UUAv5+eo9JPWsvIOY1+0j5KcWTln1+OL/7JyaufxOIeOevbidK/ooDKd2y
Z8RNG2ocB6MS9CNsp183QhoFLc61fS18P7Eed1868uxKJktZ4xciPrp7gGa5g/cK
TMsNNyIArCJRTjIFb7OR8U2M3iFHEumM+VP7zyhbV23n70dmCz1qUPL5NEqDXTsl
w69AliEkVdcimxnQyKGZEIo1jw7aO6xgFQf8U8eHGqciBkUQCH2ULgf4if5WsA/p
D2uxWW1yn6XYDVPz/1TZwHIEwqd9Kk30ZcNUDaFYeQ2OG6hqH387HrdIRBi7YFC1
XTXLUS6x+cUFUGjZjhIM4xhM/kurzTpk58tMfb2TN2UudlkWHgXDGF6XdTt7E74m
xtHnfnLTVDKzqnfXOWhyvSyGuY5RQAnT9umtXqaStidLATCjvINn0MM5FGJDHDh8
V94DBAytqBqGKhXChmj1/XJTlzyfy+RBMoMcOeDdgR/Ye5A5pfiZP7ki7xBtQaO6
+zudUpBJYTqYEEUs5+CcrC2uyQLS+BUxJ98rlE90uhuK6Z8dpAN0PKadiQVRsXTQ
W9vTH6AihSERb8IRo7kGCaSVjkYdhHXvamTd1QLObkNni8Z8KFvOcWhqI+jlUr6Q
d26pCijq5Noi6kyziEUtfdl50/Exa0IYvFoyurQlgfviZbLznTdXKncxkdPUv2VS
jmSRBJuw/CnK+2AXMZsE+Mb6lDAxAvjYOEkpPgN830CP/ZMLzyMNl2menEL+QfuJ
aO3ehvB9r6DuH4WaIxeS9n0JIhdAOunZjtktrS6RQE8YIeH2QCR+++9WfOkkkpwA
xnXoRwM5zmLjlDSphbrZchWpQIN0vgUY8TpNtYjTT7S7/E04IxtIGKBK6ueySe1D
9Fm7lP0v2So8Tpm2WIchIm82fKVoQZHFnrLLGIGgwv6zDCjN8mSWKZ+pCgyeFQRZ
OBHy6dqbfxlgoLG5soY/+9v2NfFmGuOL/tOfWJCI46fChKK65wnxi+TRl36lLBNJ
fmp6xypz9RjfJK3FlRodlK9bv/Rob89g9Z4Eu2iynKPxm4nAn8RHMalbNWkn5TLa
6iTq65Fmy66bz/Z/31NdxLqWuaqCuRybPeLOKWxo9zzHo7/enpq92yiWeaa0MRwW
Suuv6HTsqvPHIIjggo69cTKwzdODKwhBq24ZLo0skg0TZtheeW++FU5E3weXfR1s
XGpyfMn2k5sHHfYi76ZjXAnHMsQjF0oBvGvTScONj2qGwB58dPiokHDQfsSrWGdk
UpJ8uWDqUhQd5EAg5ujyHaQpknDgHpEaxHx71HDa0LSE6/8HPurtjHshwc1OMAFn
hRnZUw65ymWrkakMWdlhEjvViIabpomOLTfdSaNXfUUXXMkc63ppmACN78ZD9Pos
m9ez5kcM9EIA5yyWJjQCFuuZbmGk8leMZaIVG0P4CvDUMiXGRyi61tNz5H8dVVAA
Du1gWTobPDdA646rLeETGLm2v4IUceTVFn/+ZFC6V/I3dxRhSkT9gXjvtdAcb9ZA
3wcWuGHRCXPVp8vNR8hVI7opGPtsaXPMA7iam/u1h5cbxFpHUyuzrb6h7FGYFQ1d
6zQAxYtiBSnKxP4j89JHz6/hbUenb2vHQjVBbcZRb15FiPB8aCu0lP+/utiayQ4q
fQiz2zeP0vLTqM/05uBPjGx/9Md7ZZat7Aw76sUvL4LiNwNZpYz2ae71wWQOY0Ix
sS6JzQSVnOox4ph3DSEFBVuNCXt4/OKLPrH1OxJoBVkcWKyDJ+o0HnoM4P4h//Iz
ap59ktT3WWloRKtVwvfKT/XlmS++1stcOzKRD8TwbUF793jTRH6b9V830VnkFaYc
zUWEZ2vDE7E0B0DTaz1SV0nrXGaIWn1gfCbm6W7AgpcsL7ISh8E5HtFd6y2Fdjpz
MnZQ61lnKWog6UNbKuap2/X0KQtteTez3FU7rZWG/mdUIDEY8jKKEpDkFoMb3rPv
CsKdGIxzs+G/NPlYord7fj825Kq6gX2arhplprzvgR+o6mbeEpSBXnG88Q7AAVrZ
8WY4BvljjDLW4FNSw+eYZgYWgCJsxTiJ7RvBgxmiJL+eCrLC2aKx8/3+cOVVQBNL
BSv2rzIh/m4Qq1MNrKyT2lrxIjoCBXgRoqvJO+sB1LXKJ/y04W/bxZ25Pc7vBDdP
BXiLah/xc2fuPl3mF6TwF6MmWLlo+bJbsAWTrBryGbF0Z7iGFhgUYTp+gJhI0T9r
DybjRpeZkZKT1Bo315lpb/WEIsrA1drrki2ADmQZYb2yv3Y3iyn+4O86SJPdE5IE
pEL4E8DV9nuxyLE+NVP8WZVR1eU4bftXALAi4mY9nCKP3ps8amLVs+ZSN8Ibkx5f
uhAoUBvRHYiCs6e24gbDGzmnuGnTXxoxXSTRSH6vFrzDCfsAGd6FGzDjowBwLrFS
moT/UOLP2kgQ2/q7SML3l6eH98vY8TgZ7klqtPMZZQ/DcxzjX+UVGJsxc0lcVWfM
Utv2x0NmH6lAUZv2TQilBaSTAMAlbx9b2tDw78GP02Kl3t3fcsBq1O/CqNJxQD6K
1Gf61z5ktrKio6UHxNtCDX13pGwmoCxMrXS98duGOdSyo5dSTGyuLBRdMrfAGIqH
eKStqgrvIgKgR0FuPLmMrwifKcvSpS/lWMorDHV4vXS2VLdTFTDPpgKGZh56sGq4
CcOtfJY8IfPN2EkBlojVliQfS7cHBDjRYOhYk3Ta3ujZ2R2cJ8RhPV1nBVcGS2p5
tWAPwR1NpCHCN+yd8esObQMvzc2WCgIElxqtPGSdccQHPvi5h+JH3ZgDsSfQDDDy
Q9K1cwSrAF/P0TxtM5aE9f4hJguvn8AbfVFyH5FeAm7DrxbufRi/UGugzkyRlSfM
y6gC/dWWAqVWMgSHUZmuJ6zcH7SKBACfS8D2SSV8TLwRTBbmBvkE/zqzkwIxEviv
nrxnGfbjrwhw7Ki4Mq0jcbYoa+WBc2Ii2KltMFCqM/C2jGW4BZztcIfz3PgVrANg
7O7ISAWEc56E46i04LjfaWcb4uRFmvSj6cqCSkU7v5ZEl7u33QbL5FZlRy5oDtZ9
CWKzxNabX2EcX6bm6pYGRhqsdtV3J8E1+XbMUnRuNSgY2E8x3PH+FSDFczMcrGs4
rEFmivS7Aus5Yp1mNukO2x/xlrQ1rl0qBs2aMD3f+AUqxi3ZeocRqW2F6A9eIadh
SeA7DM0VmM6dibMjynftYcYxzHV4BbM9HML/mf6QF+XuE5POANVEriuqM4uyni2h
Qbv3l4l5u8Mble6lGS3gKITMuzvu6bwJe81nOeQdtZ7uYpkTpKG7MpLbBqY/eFsN
B4jHspeuI4sT3WWfY37KLNc25vrJbY9jMY/Lgk3pbjlRK1PsO3psmn4uoqa8I9cR
tLIZoHO9sdkh44ZFH+XArqnPQwuQZJh9AMJAeLNuaC/azVwJNbpDvU4dOGP+GLfM
hcqqeO5gJ5VrKReq9ArMIP/VG9HMC/8fegJVIxDRdjdQa0upxpPtQUAT1XegzUuZ
/uOcNSQhN8QwEU+TruQqB0k6PZDnSpD7m/0CA+FDm/AQCaWcf5Rx8SmQI0BQJt2l
z93e4pKV0lVVFD/tBZfAbQ1eQDCcXpur2gRvFcIC9WqAaaw8Y03kUlznTCBLuYZf
PGyBKYzJXbIt+BAqy/LANr34OAETlyzwh7W/DHzxSza+v3RbmO1mk758+jdRJ36T
WFAoBz68BFdTu5U3sG7mMzBNoygX/9wJ90I2O3IzKC5HQwEBO4PpjpPnd9EAnobh
3Atz6ZR2hvGMAfgYm5ruBMB1HaoShULUOm/2u9jQMkdhUbzJkjaOmO+6JMlm1RT/
gPX4mjTLfQieN8lc0YmYyqHguOsP0nNyAKHQW0Hv3FJ6hBdtoLWOT33wNNe/OZs1
8OHBTA5EkSvPTbBFBPMTX7z6G9PIQyXd694bcNjtlREHEqzIyHf5QFbx42u1eluT
3lcwRyE0g9DjI4BcFrNw32azUPlqbkhdiXs1sfF2BCw20aOyDa+x1xGafCm25zDb
XPiyjfH9sGV83d/J0U9jVdf44kopH4gX1Jc+C+Rf300iFKQLqOoGkA7pWFjmVLAX
K26Ab7ld+ju0y1xNjNEbh7tV7rWzsrLuEwfMIaoFe1Cz4VJfQSVvv3RJGWsSItPg
aO9qypd3nD0xIDFGqrvUXhiFszT0zyPmOOfkG/hB4GD2NP1EsOsPCClIP+owjt0N
ffSUBsoAPI2ybA+5Vcrikf2rpylzf3e025foDqCENiTeiGjQbyfG8zTqXVd9x4Z6
Q0VoygZZATLMEc6A88PUvDuo2iYi5rCkWj9wmTBs9Q7a8hxqX5/i8FzxGOK4H7tw
ypiWiFPoQjLfOgepetlP3Jc+qPjJfH90tXjDxxxcqle8PpGmdwVjFoRon5KGrgXA
vxhnqgDxh71+M0hu8Pz38PWjZRY0UUA545aQFau84AM+N4kpUrTURf6gZaXuqMnV
5FScOH8TA/30rftkVgM5zMMHF3QjvquyJmxWskROo4YrYajdiGHXhh+17nEluOnz
tVUUujXXC+tB7UxLSKA+36rEpkGl/ybgYQMEVzod7IiOep7+ppd94ZPjXAfT2J34
3snMp2RDjHbb1hXUkHrPxfXrzn6Rd+54lMLxu/Cioj8zGOfXOJVb2I6JwARA8ugR
z1zKI0RYv9DBezFOx/ln+/HwDRRc5qo31V7NjN5bbtlJVEZkfkke1WQAnJV3L9iV
iM0R/i2v0ln/T+tJiFGCNqnTwdVzo94wAIlkuQf+6QG2fSoq8RkH3pZ4lMWT060b
NMTTNDoUXaV8aGZdFnwY/quy8yPIcbUOeyHmM6ndjxNO66xNMjjbjBGwOgkZrHEO
rO/naNB5COLTaBKLS7ybhrWrWZMXiLI6GJEwJQQFczS386B2seWzgLA2jFyPORuk
UifkdIVeIrLKH10gdR3D71thB3gSFCh30a+TXDnmLTVP3R5Iwg5xH1JhE4oWnKzF
76lE7JBqNY1Tvl3XZxUYc8kS4HESKiPgDkLzBDUKajefClNO8LGWSLIxjcSq4qKv
nMXuPokCW1IlUZ1vbl3HOsgYLA6sCJpIMtfcch3NvqsVtJqhwXc3gULjZWOIRvyw
oWMfOpy33cOdt0dlvoiu2cs3IaDw+l11qmqgKQahwOS3cbc37QZv7s9Ztarx00wt
QwusjyB26c3czDhCw2WmtxVMQEf1zMCmWXIH4LpcqJpDd6MRW/ZsqQdGRr4VoTzM
ZK7oCY5zC5rmvYwrZmxb3gxpmslG7baKbjFgOyAU89HZp+6YrK9J8/u4AFlpfh1a
+5cmOuAZhmuND6RE34y6D7upJ+mhzouxPpzcNdmhDb2jql20rEuCs6rv1OKGeMpK
N59OL/sPdLLJ/MOy/rJl022FAMqOSlr7MEZ8U/IyJHen3k69eXSFmZB12XReMVkG
H5QP5ZxEYLrxjtmwjkL7XTM/8mk4SeH7HlU62XDQXI56Z5mV6lLZ2BU8ttVOEC9u
UGml4FO535kWNdoSsr8pYDcGQrwRiHh7QqHjDLRnFFpNAxM/54ObDj6lTmdHS95T
LAshsIe0YJBPNZBPtjcYiuBcDExckfdCURIS7UDspMhB7nwwc2A9iN7h1xyoYVUQ
CYwnlr815ZNBrbKneS9sm0jKsQi1bm9Jq5uXZnit+r7RA6nN9o8fy76mWHM4qeq4
DXdXLlyLcz2eZ9aNt9jCwgcKlVmnoLQZ8kh0TSWiNrGe1/5KZhSSUXKISSVQHRcO
0yJqH1W8zh/UIHYVEVkHBE4yE6aUfbMb4g1Tdou5dpN7BFs7YqwGc3D9DK//h9MH
OlOVmWPbF3Mzco2huFosTk5dM/ylIzdO8q5TBgI7L5JyLkPSV768HtchgYiyD8me
LEUw9rDizjtHp/DZzblmwRkRdvnmwV91UWZGV9jwp4qOkbf+6uAFu5grdYB51hhV
H8JQZLYUIeWpxaoYhiX8PwuSMwZFu8i1Qt63W54/zqZNK/7whx9yMYoYeYrx7J+0
U8qWhKUrPujJcGOMGbpWt0x1y2yTz68H1ra6rMb2TybT+6j0II2SD4x6CWH2iuwn
jHtssulZGxiNKIw6F7KruhxRxRvQtS5Di4bEmy8qmnx6E+1uLoih9fVJvI9R4qcg
n7FnYV7MlZy8cye4QFRLKbkISeOKZL4ugQ2Git5va5o3MFmSkJEDJS1h/pQLX84T
Mb9bCNfRyXZpoEpstb9yOpXkJYNDA4sVC9HF5F/ryCuF9oAdv0fvmecbfhWKxGLz
S7b2Fv4K2feCIdKHN/mVybqhT7lqo9QCgAYwSsA9oN+A8PYqIzTDWz4/KV2duR/y
gK5M2T7mcRUUV0C9v685xmkic4T6mVYX8R5WS3RroJ6Bw5GiPvtkdLgJZOrO0ELo
Dq57cwyKb8iAQgtI/bjYd/aeTS5qrPRGV9CSt/1El3zn7UaEGyU8oouhCHk/qnmZ
5YRzVejMrqeH/0db/BBRUqGQzbaJs/rdVeIFhyhkgjidVzSHg9KBO8qlx9exOKAh
WlqDBvEeXb9zvcn4yjP8eAl7q4+pmjMYvIZyGW2fY5RfsczoKH1TLh0S/7mn8/aL
6bHHNM0kM75McfdT2q01KOydPNJVWA7VqdLfeFHdazugq/FC6wF3y3yGYwO2KfSB
pPTmBEVBkyxhEx47x77PoyISS/sUb6vdsK+dR0Z438ZnkboXglJYOwBpDBEugYAB
+aGjLdlTX76EN2t4AgyDoz7eEud9FgMbwb0xSrsoRdwPmL1jt+B7gPs5TL226h6l
SSspHKOu05fTooUNy8S9V7Vfd2VkVUwQOpsVsppPxb0aj+L5CnNC4158/J4dLRFZ
RccSXjTUYIneCCBU2OyHvcUfiTID7IJqSj1Nevp7MWratqMmQs8qadGG/iSvqnfm
E5PF6lZE+BcjpJS6/4toAmU/MUpNbrq/43w3xqiSbknFCndj82qCAg4efF+isXzC
THc5NweokiJXtoQHy8v2novpdk8tBthGDTXKgWZAgQbvm0LyRKN1PHBV1ZbIWzYr
tbhsANTx8P/OorX2a5HXP8N1tWRRhK6q7dx5JkEFntBiOoY+Ffg9NhXDaY3XscD5
ym1iBzYbtOv3IdODeZh3gbpWS/rUtHE+Mx0Mc/3/KMXtfZY+MkFLMbu9cxR3lV5e
ArqvpOi8hybIizbDFGJ/iKm9PUrGeeJJBc4rI1VTbENaGI1qaI11RugAB8YCGlGp
z1l3Fboo84N+1tsqTDFhDXaUnQIsSXlNeYI7NKo2dqE3c0GEarB0N2+0DnH11klV
7pKEgcJxyLE4jwG4ZwHdEh4s89o33/FqkkFQ9/yofQntveuGi88+U4+rojWfGe0K
gsu0zXuBevTWFiM1jCivQotMAi1ejIEbi6g9SIZmknYFLS/ns/ap4l4aacBx8ETW
vjpnefPEAR0tzIchQdjCMR5pfn4rjsLqk6AkiJhq8fwczB2rjT7zZQXfMRgiii+0
5b2CiD8GuAXrNpO+5A1zpeOmjr7d3pPeXUXreD9ePqm6tW/Fv58K2cmAqAlXpcpO
lz9g5MZxBMa3gthnrXTcd7mrkF7Qc1nibQzk6kAxZNIOM7khQhXUGtmBMvNAZ7WU
ceSLxn0DR8cqNc2NDQdhsjhjsOX6NnUcSOLsmPdBnUUgmPU9jBxCaento8p/pOiL
VvQIDh0a3ym34uxiDOcleja8uMcZPqm/PNoPYaksZfqJkOzk/1TKTv4/tCuaseqK
aztJiPRFgPQc3BpOIdyNY86E46gKgXUdqsBopJC3Zcmp+YQSeeEy5S0cco+VC4VF
sA2C28NZv/LTDqEanBuzfjHZmOF2hyq0AeacFLnzAA2UeGZ9fz+ZUA7CMtyPrwsv
h2Qk8+d39ixLleUIO8FIfb7QmUoGpgD2xGAW6NpVT620zRmZkOh4He9RtP62HMSx
lsEQ1ezy9SDUz6fifkkBYmznHNbO7V5M9z5sS6JKWDfkIBghU5uVBUM20j3LVzTS
a+a8MgvL2aCv64GAQytlj9T52ylP6EYMsfpS9sWYISa08JP94XempAbHepFpt4S1
PCyip4Itl9QZ4rqv6JxmXNmD9SDbSDhlmDu1G7JNTCukZUn3g5D+50v2z6O5JZIL
lvbwd5KkMcmf+iSkFoP+jUnzojZBJxOzRRa1AihJNRDe2mknUSkoZGHK14zjLQ+w
rwXGUiBkaZibSlw49VnIV0gKbCO8JwLmkGtYge1ErYpr7n8vZE3wfM+cWWYY6eyE
fosk3JzkKwyzmGIMxdQgj97JgnouM6cui5Zvx1ky9ee7TMbBX5kA0zENlFhnwqBC
2BZGwrr9934vCvJ+mtJJbx/zUzLjevsyo8mSs2MQxnn0/GY0iNWgIabT7gGozUQD
lBt3kXo1HN111vSNZLetmpUffG88vG88KBzMKi31ZXsjDfYuHOcwNJ/4gE7jLFRy
sW2WhSjKXBe2FDnTe+XDMzvuyuuwPUstr7YFxOrOlDEer7Lp4cSpp+q3LvGiiK0F
pjziZEd4fjE0YK1VU/nmqWzklbRmkgDWh63ph/7Sw3+lyLfDdXjdPQeTRoBETi3s
tk43nT7XWPxv9vlAXKnhGNCW/ihoaiQkrdm6r2fEosk94KZj+fxoTSq16xGKH2ec
3WHV9VpI8234+IwCX1coZz0yoeb1R9Nbhnb7lRsfJilFa2OB9m9zYaBv1sLhKOLG
km8+h5P/+yN496tVx1SFyJAVqrGPV44Xlpjg+AqVchbhYpMPI8cLXgEXUJeQSWfV
fySmzByT9YN1e5JnaVhfEv9p0vJQRR+iAfGNcKX9JAKb/NcPEQeuS4FoBEpsRwjr
pyHZMBrf8OXtgBs5QDVKCatN/ovtoVEPx/86m5G6FPOc/t1Dzv1VkYjpsOiSSrsw
PNaykeuv8DIzmonLiKearFJBpUiUHnu5Cmhocdyy73GSmsdpCkVEO5pqhIJ2nyhF
qmzOUtcX1wx2oXRGqpuux/boxjER3as2j1LcxoRVQUHuXq/LZEGtu26Zmtr7oFWT
c12vgnKwiiIbxpRTVVCD/FCc1/OPN8yoh432cYSvvMsrzNi5UZWq7cjgYqv6S5+l
vvEbBymd9pAa/a1w7PJjrvJF0uSW4JRif2hH+t8le2/z6Ct6gJ9MGYOq83dn9/IH
kLhUaq4c03+t+tJ0YWaRIfhfYD7YI9Sq6M7to9zmG816ABPEym9dTqu5QJWomfMW
KKNErqlB3NjBBd9TLqqZ4ZSTtuxUOhLtPqr8REVhy87KeGc6ihsjzbzfoYQXD9pB
jnSI3wD1pFmzdHARfOJKzmTOQOBLd6uEbrR/ifqkxAXNt5imeyCdBCDHOK5IL6Dw
1HdueF/I7BPzqYxUAaOKLs+TB+EzskjgkrZ56ERxt35eqVXA7srOJdNAM/yhNqSZ
WiTFAzjirQ2mgQKnSx/Psxj0S1wUvQY+cC8qmBBbijnky9tHOpw8amwARzQTAXnZ
y4by/ms722nG8zm6LTtunErskm36KQKhCaVoopFlj5CGDQsEGssNEcZCqGZq/Ro0
UZyubjShF//gEJDTXxjlvCgAt+2+Rh1fSA/n5fHy3fRVDBilB2/geMjVe9pUPnvd
7oIQyyUF8Hh2IMv1BOeeNLgPy89AdtcC/DFxYtJMo+E2BUV1J9JCKNENSGva73q8
dzHUO3pOA/b1tz4+NHZc/6VHDfRtMbkcuxVKUDlgnmY2ocZCVTXUsaoJs3kTVdl+
iB86Cm26R1491vy3rl14kIUy5pQJ+hNe0wlNCTaARKsdpbjqUEQwCwLLx+Gj3SGo
GR5tFS0s4mHzrztj820v4xNBNI3SEeUDiZPDfyq/Rsss1lXJZ9CE3XVI09HyGb0u
CyR+QmzHQK2BxhZWwCfXQn2V+deqv81yhbQxKy57vxFVBw9kYRGHO32RMUHnuw+I
99tWH65rSIjDcuwAd3GNydxkCf/PDtBbB8wWPsn6uscw9e7dBs5V46Dpnvch4vLp
YP545hSsFc2fj/KWkXXgy4C7cC/k1AujX0gj4Rl4E8PsID/23FvUpSxEgF116VdU
wHzNNYVDMG6CvCOs55XLmUsJ1wKUNgnA/4IydyeD3ESYz7hM2c+k5tV3buYfrNiL
8QGv2ms1bHqzAxA6znPZtVmd0/l03aPodEwXhu53YDwUhEThMRV4ZSGqzR6OIoA3
I1g54lYDPnYP8sa6Kll4jOgxXbVB8RV9vlOR9XRP/y0mW5NOtklBLpR/omyjJNUg
7My5OqIwo5BHme3zgYJlMSpTY03FDPy55p5tBDeEcpscModb1a/9jmAoVj/241uK
pGlaR9Y+wb8U8CK9nFuw0dRfubrS9Ap+sUaQjb5hLnXwBwCMihu0A3sfVkuAW7dK
P8jyfalwkO77S979jhGocztTixIk37RI7NXho/Jgoo/B0sg9eEbGQsVP3zZjtAQt
zPL+A/WNdajAgVXnAiwM96EWxjB0fTAiuBRTxxllrONYdg4psHnXKJbVmH8YKPu9
oCjRYuhJo78L+Wu8TBCnwRmHzF1VGmqM2+KxpswgwpV42Rlx8R8BKgZxH5Qc7xNH
9nOUnsmZBHvki/KdNQZeXeaJsxpCRNe9HzYH5Wcr1oWM418koxbQ2Lr5/CjOn1zV
8LtJh+4EGmG/Vs4Ae0zsjllPxY7AHoIToGVhNriq2BQT+q+3+M9ip/R9/MEp7OnV
m2NZ/WbbCMTkDmc7+aNgmn/10rNAJef9XcMEaanNN0AzleKDuiV1Nx2JjNYagdQw
ZSgk13CgrhsjMEe9nBFhfrpPSQzeDVK8a4XOyex5aWdj6+l/j0Zf1RH+ZK/Bsek/
KgC2dL8hcr5umkOvyegcdzkhwF3+SDynDqVgeQ7xQA0XC6Lnu4vEi38hgDRykV7y
u/bRHcoqm6anXjhjMoMGLqRIN7qR2afyYUdTjEnvtTHObNty/GFhyOOPpISJk0Mj
v9kxgN0ajhmIugtdw39olLhrNdvgE+OxE9gu8Th56XaJmwwkEpdRdVHnqAHoG7Ni
KfSG2IS0p9SUL09LRoc/ArJ5UddZ64rjbTuwNW3Hi89NObr9UX8jetPYVLLdolob
unAEB0FeZscmRoaQMJbBDlN2+fSfu6sHRgsrZ8Uj081bQdT7oF0zB+3zo5AUCpDS
gcgKhb1GKKFoamGc3H81EtEb/6nyUwKl4pgauHqZKLbaRG2bUGZJpZ48PoZPlgAT
EL/qNPAeCkuw9freMMz8zd+GDpG15KBGuiQjLYa5Emq8EaM4I3J9KfYAryQdRh7U
KHxkotgJlr2DEis1gwsftEz4Nksf/gu5OW/XEri6I5QkzXMadPwJ/GqYo9noKnFW
AjBQgZdhXA3V6E+AJpi9VzItKaq0fFaaHUKUjkO35pdT5ncN543Ner0yxiYo8AaF
uj7s7iYGriSHOLzzw+ItROoAR+zdzCXkSbnpB1ItBs/If1ArOSqaMgJL70jCf5Lp
fmVEmLGfpmuTsVjGlVM2XjClpHGSvpfs/QkyjYiXmwCfru9DygIYpqkwv5ENaoiB
ydw8QAHxpSla7Uw1a+q5is4B6lTxCKfWy/w6lKciWfV24LE6N1JAOisiIwCuJsKU
va45PirUYzWG+fcZ+3HEZcenKLJQqyWy320cdctLCYyjoEQpXHSHt61avqZutwhr
bzq/UiKixBiTKkQ8C6sr/XTZDkMUNSm4LuIypkttspuLOnt4XuggGIqoP/KOymm7
rU0I6bL+Z/WCSTDagXJaJbm+1KuKbI7y2exwEa7tl125GH6fIZ62gFUvaktl6Urc
K2MsLaVOkASIzoNOwPaOTkONemoBgo+3k4R1VUHk9eHDnFOwjeIykI+K+Cs9YQJY
ZUUihABCXj1/xQYXR29aZJxDLws2oSXW8b6Ws8Jhv7fRxHMzMvrYBlnW56OpDYP2
MvEA2txZGxCMk12JUTNyoQlwZ3aw7XRv7xO9d8DmxXKFP4ce/j/vIPbMjCxNkktE
AOmkq4WeJj+6xbjlOOMyHgASsbs+2W80cdzSl16lZ/dWJCTbZSSzaH9IQGaO6ZRe
60w0loj4nyh3Ps44sDDfdVpfAiox9lt4lq5ZEUyNmZ+jVz46NAsKtsTb31GCK5QB
7qDmVM2S9QQlNAX4XfUSdG1VtISWGoXBWkHUK/EQx9lq/SCEenFaxq/ry+fLBqBv
TClAsSK5mCibCjdGQq/jo1uLuS347DaXsh2xTYccz9sRj+i4U0ER2YPhSVfz5oWg
0ktUS2SJohHDshQM89oXvW1nvRlaoEFrQUn2J7QgJF78SRiXWbG2gvom5kKPzg3s
5iWWu5DWBf383f5D7WyIDl5D3Ft6XRE33X9DPufie3hmkOX1lm/RnIoejRjit22d
6qRl6DQhzi737nAPGYBwtXYY7+ohcQcYr+1/LYQRyoJa4CfTVjYbp/aLHV+/pDx2
GEYKJKu3yXF3agW7CmZ/AN/AzN6iwdVz5YrC9ydggh4jteVZ1oAmzzHp+hTAwBqy
8YL3GdFTVEW2/RKKOHp2uoU3INLofntV/uYkgKgSb3pavYA3H7VtjqvAgl7XF7PB
GtZHuI9rDAFpbw0HFh/VllaKgHCSgKT7LC7TaoUsmzsjjJrOLXcM/o0v/x4EC9zd
mSy34O45vgl80ce2Ndd+K/3+K8j3xbEQDerv0QG+SeIW1WORANnxE3hSVobAIc3a
ud+W5tvJxfQWVjZRxEyBSRzsViZNbfh6O0Q/l3sm+MA8j6uXn01GM/4wTDv9zQ4N
oGVKAl+pyEpKWHhH0bS27gaZxxKypsrA77yxcNV2+WLFnk/bgfpUDxpXHWWrmEFa
YUIhIY2z93Br9J4V8ao/lOzTZ3OK5pyrR+nIZUcrgu257WQlLGj/rJn+PtWQ6IrK
+LXVcsAG1Xy2DzpTgQWAWSdAhHu0zqpy+n7yZMBiSiC+xY9uqMZIz6NSYWMMyals
xDeWU1VbBF/3txN35EipmLPsXdh7gz51td9jLwJiKt6/7OPX7x4hyBpFuUKrk9xA
yn2aGnKPAqmgbwF2zBwWB35TxaoYfWUZxUrC4hw+G8NLLAF3PrQosDJX+hW3sgqW
3SiZCZkhWvj3M+fNsJnFFSxHso6csQKY0dUY8LYHRppGA/S7fFuwAYAX3HYCp49s
DLmqInN7XcZqx2O9zwIdhsFvUDi8S0qfHppFzGvzXbqOw4XQOy6/wDB5lmjB/fPX
cpMCDMWL8zuElTHHobyQm2+Z26oDxKIcRo7v/6abI78H1PDsYB2lANKaDA4KRhMc
YsTnJUdzbc+nCKoSsIdVkM3o2+QktwO3pG7gtVamAKBgFvqDWvCC/lKk6yks/rYT
wDlyAfeAg3B0jggAvQzNaYHqDk8cvKGObBh8zITIiFnkx3XGH5yyrTyDeWiBcfK0
PllGr0EqOu6bT3aEwri4rIBY6aCHDEUEHuMooz37bKEo5G7Gi49+8rcNZnumGqrw
L7PBCkCTcIv1pfGVNmtQijZECgUk6eyt1C/80ejZ7mGUwb3z+VPeYL3jlmOHZHpc
LjumVkjYBOCYgGoK7hlwLNhzJtgiIhpZ86l/OG11BzurSaV5lD6A8JMLM7O6ILVJ
HsxYTpD1gZpmgAtzM0gVig6jgC/qpKWF9Udq6P9CS9fR1d+JB0fjX+7fwMJTum+q
6J7MvF/MGY0JyWfk4JDrli1/krAzGTWgWJ0YHcZES8tsLIhw5iEEZ0uYZUqhoXEU
sB5wnLxENoJmvRzBTslQYI5XPbcFwPWmsTNKLmRc+tZansSpBc8bXVqNY8CpQdNS
Wif6dn64RW+PI6Bwm1+WKZ9134NEzKH9sjUJsMdiXsVFLxw0EX5veU2H1o5c88uS
VeEm4bOB4X7wApkpcGNIMBCyA3V7SW0tllxpIe5IWEeckmD2y4HVER374ycvHXrk
sQ2C+87tLQwEay620VElZwOFWGknKlX24CMXXxTdv+qh5GEsjGA5oSlqViaFtCTy
K3+NDSUdZBwVaZVJqwy+se924QxySa4+QLTbYW6JV9nTul0+T/niar14nRynvtwx
XHVJ9/bHG66QEe/hpJQjBd3lpV6c+yeMhEISdWTI+d7t3joU0o44c5sPnlH+2MKe
yaiciI8oC993cjeMlELqlJwov2p/XX+jCyYQJqAv123S7/14RalWJXKJLGJqHq8v
h43zZ/Bc3FXdU2Lf8grQ1VGvrsU8HXA2rW0QfgWDU+vHUf/2Pxe810P76QWASa2D
XD002oaFb/SNDxryw37MiB2AdkEGbfwfXA76ueMSnN+gYyQpLDrLr0gIThKws9h2
5hpn7ukoSiE60zKu6N2ajUGUJDJ5bxzZGejvZkX5neqnYQiXJVl2xk3/5N3rnOnr
yMKjk6hHa0DVdcWdtD+G0cop/ugy224l3Rq4lTsRdgwm0mK1CBUYnMoEtralw/Mb
dnKS9xdXyhlRhPXyTxicePC7LQO6v9Cvw6TfB/vLHyPnMX8qRT7mKe7xD2CwtPTd
uC7q9ZTXvL2XfF5JPaPGVHw95GnqEmIwmkcqN5xAZmK/kDYsRwkm9HoIQLORgM9Z
5zE+fHqjCqYRDocAxs/ErgG59GDVZtVdMkZTFuq7Zj6SfJFmtKPi6o+6vNqtNvGY
o2YTSrPBlSTHJXO7c7C5bp47N/NmNug5auyws0aA+QwDa4a7NRl8i6NMsNKA8omM
Y7CXbByQ8Dz+GDdfHAMCG5vxGCANisHCbpAm08Ywa/0FwrXgrVl4OZQuD8ED5ObL
ENooOamPyGbCVCmOjFeCtwoHl9ow986tdHrm4IrtPteIE5zkidZk6NUJv/19G8l3
fveLkTWrZ5AcSLTTKyz6g41WBURjYEEdSM9MCj4EjIXbntJZG0gmDAD1m4cdE3YY
VBAlT+w80OaMeCQNvxo2GGGZzbNri8+QDbParWI4vO6k4pQelC64Z81yPruecd7H
rUWFdw+KE98OiiyIPusQGuQjUyvnzjCeNzDT8/p0iQ2frnduyXwzY5/durj+p78c
nsSYOlKrBrXIzIWIzu4AEss5yhU4ucejDXmcgIkU/cA6elvPph3PyiuIasQ2YvOx
JdtvWQ6BTEMXgpquJlowbMHHdbOipChCF4J8qf8sSYEdJIyag7yTT4MJIOWP2pdI
sEvvSHjh9C2YcMV5lBuFkiD+5uYam99neFFTtrJcfilFbiaWZdBuwWlZoXf5d+5v
VjBoMI8K3piVusCIM3+wZarvNieRMFL57wJJBgxb6Nux7i3Sj7pGtuwNRp5KJi25
FGCUBFIvBJsRKURQjJTKdnmvcNhRiUrTSA2jl+z99sqM/QBGCPgZDSU667ALXdSb
S90BFB3IEfTDLnhu/mTjB4TnmyBMAAitksDIjRCRvzwOQ2qXY0KBIVsUkt/dQ9U/
OP8/ogWS7+H89VSnEvfr59EXSGXpMKIR2JLVlCXRd30zGzY59O0J7flRuqm9VGN1
hU4MVzI/i+xHu4BeACML0Y4M0tQGQ9aWtS6mL9uGIb0rcrS6ovkc63VKkQE/BMfz
fac33lLnXIDxC0ak7YikcQgvf+EOBwFOWG2qZSjEUnWZWtC5KAAubp/GBPD1GLgr
lI8bXoU80xRFHGWDbMYW/47XXMDoKUlgKEUzP68yMooIXYgPgChl4CYZp/q7cOrZ
iplWpD7RedwWUSdwytq9gV7kQHiiMmdojNlqSldGyKE75NkeqlAkGbyX5K42AzRp
aa0hmoxT7DlsCW9fC/P2R661pwZgVEkLLUekAlxpKxdx5mROo+HYuu/RHKP+yAm9
de9IXMppvusPVDJ+LKn+alYezZcRcThnM9lSBon8XOoFV8jiidU7RpwLgEmSWd+1
kI64heMVqWN4o590cFih70x1xw5TDSOjou7ujkzlV2jNp6PzqaiY+6gaI88jin+4
yIBhRPyNLscziJDhCbuWuSG4IL5LMiS0PR5IqGm6LDfTR0w4lj1lYNH6z8OBI6wX
zN3o21CpRyBJvzBJ/fvt1WCR4iZ2e5ZfPLFOcCI2U5HLHhIcz4D5bEMpoyzfjpR2
GP/VwekSxyEW/ZKaQAk+ASA8Flk2Et0lqflqlWPIe/jvMJqzrChS28OkTgNq/rLD
wvG5ayv2vRGqaWGE2dCi19kUZaqz8TuDWJUFO1buwxuU12c/xfSi9qdSPU2IWpJa
8tmvh2NKqDQa7Y0ojOj9j9qOBhht82Dw/j+HQ9Vo/Epo7PGTNc3mNubTOH/ZiNNC
ofGxTifFQXC7vdmY5ULh650Mrn97TOm0pSnb3+H7/6AT3VKZP17SCsr2jSbhGLrz
IcuFlRf+1lm95/xs4JFb3DPiCJBtZ4br0k8i9vHcPjiSqqoOaejP0y2X3vr6zDN3
Sw49fflLT4sNlw35wTrae3zNp9+OA23I3bn6aZPaOn5cptXmehDYe6gJpcy3aXSC
HM1cOLHr83W/1nhxuHyUOjcnWRxymJFbePET+anqNfoJ2wipB276bpuKHenMDyuG
gLUgScxWqSgqyKMKO5dNF+0UqsW08cP/zomaque/COgnRWGwMF6Z0y4RWGW66hDW
xfaxbT9VjBrSylw0qOJbJPNRsQl0bYWUVHAcWF0EM1gwtk5hzKlICaJFhZioxX9G
MPBk392T3UYL16rfm/YuNZwqwvEXyMJnWkESihO76cJbeKxyg1yg02ED3gRbO1m7
YUKodbRRefRkWRVZ+CrpRGzOGk43n0p9ZmoCNEZ4lc2fwnwV5hLax1Tg7ETxa3Ob
73f1MvuuEPGCcEZb0Mnv2yaNK6XBy/DIjCoVYKH4xB2rZoUHTROZYt7OVwJCWd6d
1MoTf/UnLU92lRUQWAKmYeQWeJ30pPGKWhI1MD9ZdgkT9+TZ5ePvYN5bOK6eESab
vJHm9Z/rUxyntJ1KfY9qIJusd/91cItYXYApZhRqG7RYIkRPESIQt7hslHEY8VHz
kpcguvhKMMOqmS3udBYiH7kGRyXY2kfn+T0pPkLPfyK9vZIMyWkTjmsk9urGsCiB
FtbfHoyVa7qH5R14TaXx7kyrlQWeONgh1l1VYiaitTxaKwmBwmJE2JVAJR4s0RI1
ewWBxN7XPnOX6wWX3IMvzEYcb8s/Mh0nGKajwIVv0cstyp8RPAdA2K/eGbVRgPsI
t+Km40U6AjTHDGzRvHjILgMP+jD4O/D5mK6vPP8FQEDyMoSQ6zm3UwydakLQgmnZ
8x/H8DpXrB0ClA3LGRhQ7Z77os1lXa1ifYPXyl3uPYEAu8rkqLe7UR2eAg9aA7kH
LPip8wkQxirQpIuAIwff484pLLVhumxL1zdpZsydcFPW0Y3vEGUiuPU7xk1SnKR6
YdGbIGdmWXFj3Cg6fUKMKDECDeVwjP3ULx7jv+IAIxf9R5jVW5nP5G/Ov/drvFrx
2QTm+JXI3qpyDlZ5FG3Hp9o7DQbbkGLsVBiKPdDOA0AGDeX9jqYBu3XvPg84cRp9
R6bUY+05gQJ7PgnFSqCIrsUMmCzzTD+zBQexIw8+dqWNcd71rdrx1WdHRt5u+px0
JLvG3xY3WoTi2gQ9YZtUXHTrp9fmSc+Pcg83GPMszdBjTUQ7cyE5GydP/XXMeKsy
/DFq9Eky4nEi/V3PnmNYhad1SXjNLPX/Tm9BTLc9g1SXaBaNcYHJy5Zn1maxvIca
/h4zKDPm86XA2q9D6QjdXNNANWcHjRcNcOSGa8n6ChuwQKBROj/SgPNpviMhunYo
U9nyPvq4awT90y0wv+52zDOa3A6LLbIdXXegDvwZD679F8dw44Gq+vfpJ627STXD
THYsBlL1UpdpNYBVedkfcl0S0tzlV3xGuUIVG6iqoA6HUlvXfM43zpbPZTOZPHql
Z2/7g+58yzgoI9k4lhrKreVpGQvUjDL0r/9NbteORps/FPFjOGDexx9S6r1JsEaH
8WmXpVXoeAwQhFu6gkQS04LnBhHf2w7ZQyIqaRmU35gojwk5XjaqZLIIgAT7Kfg0
Xgk3jkJsagHy+UXlhLckenLHVXRrx0sbt7xwO4b5la3oJIrs05nBvypW+7FPig9K
IvDx8cB78NYTPbRCzTZaIwiWeMZk1HTxgCQRzLvCy7x3x0LzNvZeAv9lFRxcy/Cm
jTbj+0Cy02Fk1JkxRHwrWwFrBPl5/ZS59g/sWP7qeGV7lQZbq0H428T2Q5oYS5XH
EwrcIq2CAEFOxkBav8eGPptCuO1A0+RCnH2In6vdgaysjStBiNSsxwhaFoJXtSH1
2kHb8sMJA4z05wtmVXWSmzPszeDDbqsJMAQdG57OocKAA2E91Ts3pjr29STDQISq
fgLGBN+/5U7pC37vHTPUrK35u84p+rAYlWXvt8+zGobl7A9hGEa/pzSg/kgdZF7G
qwOKsD5qnHIZ+R/oX/aIZzctqp3Qh/MyEJpTDM8budZb6XklWuXepGHu17T34GLk
yrR6SBBWEkEAgZ2vPZU1BcfEu80Umg0baE590wwuUuLn7eaascGdNUl4kh7a7zR7
TQK9senFso/BgkZZ7cD1S+d7SzVYqsPKLR+Y4bnDJT0WKzZWkxffIbUnCE3kKEpC
uHsrJD/ZTZeR8SzDXkEJZiIw5KrtvBk/D7P20B2LRWnEBfWuncPzn2FwLF7+qTJm
thvUj34dWPpB+LSu+ZoP/9HpEE0IZYWtsneZ81eQMpXZbr8RQ6w3PjfkDIyn44nP
usSt9mPq8mZjJkmJ29krqeuffRfIKhTSgSz+NYEuFl1mQjXiEB/3E8BwND+PWyxq
RbH2Z+avbDtKl01OXA6HnIR2L07VGM+iRPK5rfVTEoFqHCKzEdMQchP9AwPIjG7l
OdiwQK5CWVAWkV5WTTs9z/vOAyzCrvwGD2zPB4SBfShIYR94hSv3ify28e4ftWUF
5tdkHqZ0B+DaFq00Nlc0eWVIbfBorquRo59mSaJVA5jOmtit+3G0UfYi3ypn3FN3
wMQ/GgdeP9JaPs2s0GDSnpJm9rkBJZ7MboNWIkHUYaoz4URk7kCI3rXwtDxGQ/p8
Pqtqi3uWl38BF4kQFW5o/z2dETPBQRiRj7VJdkT9kbBg7SpleOJlD3E1JAb9vk3t
YVjk7Z431q4NmbJ4wQIEJy2FH4qVFc3XaQsFsaxlylavqfrEXesOJvW1oNK2sjtX
2UQ691afnLizW+8QeN/hILLOGYBYgNxruhzYTa0VU8VgYLmtOPsA8U90XCUd9TQQ
4Ji7ooKgUOqTTzJK1w/8p643RF+blViC4xYPC+Bolkk3r7WHGfW2SWxhbXqkVHfE
RCd0Ox/h3jgr3Goi3q4e/btTdTYQpDjwnHXB/VLoAmTp0XsgWOzAx3ayPKno+PxJ
uSP/XlLb+9q7cQhsneEyBja6uZ1MeTvb8VOGJW0HFZ6L9XOW8/EfRjxOJRiNJr6f
1s5fqSyZPt5UxCc6JLAzaEw1SATyEUta0dcYkXQ+6nYsmV+Z556NWZ/7g7eqZt2C
4a+Q3yFCIlz7qX5FugaMWBQGdGLw0pTHrBWPWCibjrqRfHs2ah+zUQOfacotZN2N
/pqidDcE/+Ql+Vz7G/TQfMnrgarzEVo8qrpJ44ncZZVo3mSxxPz2Q2KBPVBjzMtO
R1Jfqim2pqyPsBiLlpNgy/nRJW6TgEHo6KXL5GYv0YC+GGut9COoPnoZwS5Orqfd
OH48jOpN/+6DZqjvMawMWvVNUUjqYM5UcZ6MxrtLO/0bKaR3vo0+Wbc1ErGhNrDx
kCazF/q8iTgBmdEifiynJpB+QkPLKtLSQsEXc/Ay3HJbrMYQ2IxdxK2+NQrBAE6K
1PAHAXERyhOXoJzbe20DXBTbcGrKdJE15f0OjOto43X3LvzI2hL9ggKO9is4P441
xrJBKyGnUF56107uJfPtnThkNQIooLNdsF+sbSsP7Ra7my56Bk5pG5t60iKGlfbj
PafcnNq2qO0g15Ih3lZSRr9jynctEy2w7tKkIrYmRzvnQUldeBjiaTG0bgK8cdlK
F5z5I3aqYcba0+ueFU6o30D6GfmhhKXpKxdnj5Qu2S+Vy4CUmEG+FGi+xWDnaMBn
CH1t5GB2Rth2qnGyp0Bfj5LiReuUwUFWs7fujwQcvyC2NKnFbnx/Yz3kExZCNDis
+Gl9id2uP6fLj8Vo1e76Iphv7JgMDoY9K1dWzXvB8dyY7leFRLzbLZnZueT1tIct
8zfXad8CNVS9V/0/iFFeS5MNYZg27MOyBb2Z0mRMxSDYLRAiKVa8hqSKiXe8akWL
QKSqDHILu7SDohEXUJ5JX8MOLNd+Ef5MSINk8E1B6EuCD4Mvcwa7c2CoRYgamXzo
nX9tzj15g+rJd2OGc5m5g5bNcOaGF1sOc34BM+mg9XVe8zG5WlWpgybcPM/4w9lm
dk1hxGTTq2q5yGABDQEy5EYiMtePbSvJWM8+9iLkfz2mfml7WTCXYR6kzeRXeqxl
uy7ovtGRQHzrXhyDY72OEDtHT0GM+NMU7zKQvNEVbDXINihHYvXyw9F0iUZPgdNw
CX8SHRfXEgMP/Wi+A9HBWx/U9P0lS/Z49z6quNLm+ZZ5E7Mg4VqbLY49kklf1dN5
rXhPGe0ZwY+bxsA+Njjo+A0pNJTKonGqUTJBHHbwURpFbola45OXI/iC7oBvwDXv
69YCDr1WWI0ZjflGtKufDWQLV2G3llCgnZiZk6yg4Ff9WnvPWgG5Ym0QheqBACxM
4drtGdTv318wAgLuRH4ugf3JFLSl1r5T3qUWNJD/JxNdl7wSN0tQiSneMiQo8WTg
ihCYz+WTISUqHeoMDid5ycqBNwGitX2rBywd8uVdEXPeYakhzxfhceuFrfMz2a/C
AViif9Lpgpn0XYOe+wbzChGYd/Btp8DzYKuEPTSNBXZzvh6l3cv/KjoYBug6sxjR
9b+iyzqYNJ+jXYFldF6bGJzPQ4t71jZdePF/AyZf4ugRotagf5rTSB1mERUHfrfa
85QoSG5yxF9h+XKw9TEascZthGwdFZMzauS4ZobG3F3qW9gCQRjF92cl4Frre+c4
D5C7XlvWdA+aEyTQbTYvbWeSrSSVYH0dN/Wgt3hotExsx70J18fmNxYK5dXs67On
8JS8F7iU3Nqr5cDvX6hoZ11mVeSHczf1SvRa72sGN5/cCaEJjMd6V9VGwV9ezCWG
3l4dE/jiIIjH1u3ZWQfWi5kxPoMDbswyqHRn0Zfe7UPl7EvtVCp0K+H5KTqBRW8U
b3ech+aOQWD4fDAvXq1RsSU/0YsITxmwLdPRjjc1NeYHIBN4z+6ui2PJDKAmHHmq
diaWiCU8jKL3bPXk6+PBnS47GDH9SFbNsRHAA7moc2TYLteaJSdPlT+AhDH6bxPm
Dd9dQGe32iLpXCvO8mVGRuWgCvlqz4KL6SZZaZw/BJYxQzkroow12gv2M7DHWIO3
F6pROea/5ixHoxZBmKAZzBL2OgAlLbZ93gsXuMwKHtiPc7Ps6A8uay/uVFupr0OZ
54p/qP5hTVR8YDFkAcd2TkcQHl1+Yt5bVZCViiILESvMg7fVW6KaDKtcvAXcPJyu
KJF1DeOaXDVkiE915N3X2b9uQJYbb/REFTPKlfHM4mUgBwMxVeGEvQMx8rGu/tll
frqtGZNcH+zhl/crQWHcS6QpcWt4TFZpvBnL2vFcvQQTmMttqzhhM1hq93mS0e8+
KwXiCq6JKklyLks2HA49xmgcCZRJfHzS++cGedVo8bNk+tjnlxDpV2bG9pYwW1J0
2kEw6+NDxDMwSSDRCzJmEj3NqwKNVXJiDwiC5gcSzy3zxa1OaSlBCFiWrdyLJaqx
dOhux3/oFrSvtnAFuEwP9+w2fkvhIbnLX0KiCiISUsiXiFWIs0ShiqL4N+fCWPzm
Xs5St4rgEByy2lq+Ay+EsPTluEmrhQSq/keXKk6XcMZKlzo6q9eVVVwTtKWkgXHh
4O+HFwHWPgdhSTC+i5qikQ1v0aNOfb2vWRJefdnYU6aOMmtw3PnTppsc2RK/7xBX
T/rcPx2jUCpVLJPTQcJy3AatnBehLPtTtXjCAyqNmGDzq47ztaclHfgECDzt0Ybc
bTns0ZCXvZQch4yvpbUbjAzvSIldNVK+LiLSMgVhMQ4FoOc8It1H/ttQbX5eoxgt
IxmA+ZuBf1RgF7zSMI0m20nRXyuSbz+id64WD5YCxXA9YX9Vcz2o8tJGxwxRHJpy
kfsDwe4wefrsDLm8qhqhR6KsNLP9CbfsPKgc55botrHZ1ht2WzLyBBSnOLRtYyjs
sshDUOXHtCvMeW5bL4HN615rHjAZn/i6Yhe4IPkPYT6M0YuEcL3ePZip2AxC2w1h
pXgNyAKKk1XTIo9by992zpla3JPnRYS9HQdWU3S2JxSpNfguABx22Opb1vHlHa6I
Z44VIoJzrFZFTYewy75KxWYC2L0j/Ur23kWRii+ZyqEtEdzvgKAVhqwRI0dTWnA0
NKxlu3Xck/6kZinLxvQCZjC0dA33zWCTQ3b4vDfggD0chaHJ3LyuyhatUPex9of4
sU3xgmO0Mk5JpHCTdi/7ps04kBIIIzX6ljsxCwpAFb6SsyXWAPRADhonKoNexjqP
cQPZUZf9JoJwIbnrFIgVqN5dktGwE88lOGuh6Ct2aBvP5Kkii9lDKvVg5bWKAXCI
hMCBvN2t1UJ2odHSy7+nMnUR01ZlfjkA3zg/zP56j9Oz+hX3sK8bghuM+GzavV/8
eSXgPq5agBz5bfBoDDSX5MqfJupBMAtCnzMdH9AJjgcZcmwi5hKI+Sp04qWyrU60
UWB8B3G82YhUd0ccnJDhZ1+NG0P9KC1DipoZNiQkX8URz03TZSiWJl3mAPvOc95K
cla6/BEXlVN7jLAvqLTtAW7BS5imypPV1NGQjca9xaKUo51eZ9yRWMbaVTaIBwG9
BI0F0BybBdcn2ZDp51A31uNL7n1pjyw4m9rqDv5hGaQGQiRFI+7pjaAImewVC8zb
s1VtqiyQjuYRdfj2KBTUeNLsA4KAGSuCKVJwgEqZm7IpL/c+tQdusgiNPReHrTA1
qail9AoRtQa+WpZGNVVVsv3SXS2afB37Bl+L7JvRNTKYU9wGzXg3qv4b5+4oFU2l
5kEW6D8knXFFDjW4jBYI7sFwQLXwHn8yikdp2M+LUO4rFgKgCuXRlIBi03/P38Pq
0MykMipo9zgQFqG8kvF5d9XBjKNhJt5z0r5am+6FA6JhfV8BMtKjb+uBEs0hRiPQ
EV11Cbq96R4Iuqaw1FCLqLogJgBGMYyjzYR86mgCmYw9IAS309oQaYZ9oQTxNxQu
4u3L8FiHksLWkW7AEd+pg6Gi4t5v63IUyKehiW49zUP+39l91w0IP9CI3hzxnL+p
9Z/NYRSLIjY3WhiWJykOYfktnYbSVXtfyj5hdVJttbhVVYoDKWK/60WGSz8J2Ooz
3hsx9EXd0kVjWNkxgKwIBrDFa+APYloRmvMQWCP5YrzQ1nqiKJcWqtDh5CwwEThS
wB93pjMEvFRQp1ncfQh4dNNy1tJ7PcK0IpWfr9IiFRXY/p4XjpZAMy0aNdOrQVRx
en7vLvrXO8FUn9JKWCedl3hFubCaB/NaZ3xqVB+cc5cfT+U3kkjPjEAfzDNFTvsO
9//nWnUNK4f1PS4GNTa8y1xHkQehB6gF7r8Le22/AQH8j9EfnxmYsO3wqMpoBv4m
6p+0QDRt7J+CeJQ3f8CnOyD8zQZ9EHc3IJYSQkJXd6rWOfXvIotURJk/u0FAdouI
wKV0nqpdInUTf9E47tp+y2IwB116/Z3pYY1+yIpI242gWNSAYH+YkMothObK1pdK
yYYCwbHuSTTnUSPj1gL4Ddtx+kPFsM3seyfww74vKP54kkIz9tzVIlNECQXTa7Yo
51U9CQ+7+wmjGJFILM1QSm24EslpVD6llRH7FwIeMkuw7Kv33yHV9G9denZFvqAE
tQTK3hQBI+bdksFJYhj7pTuAhWfcXC65/ATbvF1cDOw6HN6ZNrufJZeEh31RKPx4
IfAGFi7l1ZSqYnh247XIvFVujCL4ELiDDakGnqXIyJQNkHf/8Gv3PvrgXaYLRdxA
ChdWdGAiX4i+SkHQ1VrRzrct6gloTw3JyAnI3k9dnGqVYHRphmDUeYOffYkNsjIU
lNtYWCsGXjLJoqKWr6bhcM9NkOaCLXQVBtXxoYVnnavW1zit3PRdCqnpP9kkGiq2
iAQMn2lksQLpvAq0R8CNN29/l4i7+/v3OTbJsINv9QT1qamI9G4DU5Hq06f17X6R
Av7TyZIBdp8pjmM1UzT+IcKkXWVbZLdQRo7agMr60cnusmRiOGzh5NATRs7HS09Z
fFk8N5tFEePBQzW6oLC8CTphfp5L/PN+wwLmDJ76u3WDjoOCpf60N8HBwXhzDzxz
DIn3RPB2EEJWrgpsKAiSDFmHNV8NTBl+spofPiZGDPIEN3MjwuXpfueehfkdFk/h
w107xAumb7uR6zHUKIelQFcebNb0QZflvN6CZCtrPHjkSywwe3FcpUzLSp8OtCob
ORAlEZHtVndlFtWVJ+xtjJpJW6AJZ2+nQMn5MIJTXNyexd6cliR2XLaLWcAoIzVe
txfiGVbzRqEXQ+Rd+hOBDhh0ply8vxO0ae/ZIUQuBWVo4T7Haoq3I43QN3k9EJkH
tIa1trmLvLZqkEVkshrVEM0isY+h1xOK/OTubw+N68j5jFpS5eo+auWOriqaseV/
kosYKyFqtCCrvJEZ0PYQkgHEsC4HGXdgiJXYJLpYNFuJ8I27ebWgBoDY/ZfnWvnU
k6Xc42Yp+F04hfBg4HWdkEPzYHgcRWS1yk6MplY53C9LXoG8IPZ+d1FJRcTTJqcX
fP2ur2+QefkH+XE213lhKz992Gr2dVWXZePUcskF0Wku1w0GWLfknOxuV8V8Ef3F
jlK0oawZj+9GlOOAZ3pRCHInqBaDegfVmcd8AGqf0Zax2vmdJrX8RudLzfd2qIkM
q08fuTHWRw09lMNtsSkGb35+1ERegljDLOf0/HWHjARdh5aHWMeKwyYVYirFCRHX
twivA40gmVOzRZmYuOXID8pWdJjtBiXAiZNo/hVaBRicNeHaWShR+V48m0QHvUQe
RISfKhXDTNL8fzPkWzMrTX+NTDMqvMj/P6pmFVwzAAlu59aWT+dNDRMv8N8C4816
Qd5ymZlwOtg1u7GTE8r6xTYVquP5mZiYnHVyHBoArXIKW9NEBhkWLk/xZlwkS+l+
VVwyj7VDjNC+SdilAMqK7bwDV12koVmBjbf3WzJCDVojA61cIK/uYIoNog8WtxXM
jgEc771Co0FuM/c5hgsWvY7je9nKl/S2ZW3+RJbmPGEOqraXUT2nEALfsM5JWel+
WzXWivQcbvRLcG0jYO/y2lpNbENfAmRV3P4k1oc/yhpUqFxn1r1BFWCWPtxpe+ZD
HSQGad/Oh7guHfAdVXidYBzx/PoxyYOmEPeGn0cy2nfoedv6uRTZBqplO1Q80a12
4xFkYPKxFDGnt3ITZO4OvjCySfrAIQAS6JcB9HkKdVWKfaI4D2Fa8RzoBwOaK5P4
B6OTRIOyJLaVJGll7PsSj+15ja8J/rr5U0vbs2kTlENpzNGB6PJq/Ko919st98G6
mq3lw226AmQfFL2ElB1Lj24vzxNwWUeTom9+ul2Vn1U+jmcJMk9wZhwpEVd2/x/I
yongSTmMVVZNatbqJoWbeqk8vrXdw0yMl8U/SqGSq5m7Vk2/s2SwmthWlKZnZNFL
WOQqE4sl3lbFJz4bKKo0UYDbZJHZnYH7J9FsICcBwMt5qlp/ENhxLbFYVnDN3vNm
IA+jAdXp8PW+TVcIKdm8juhofSGgkYLRXmhpY1CxQuASszmho6jJCjnebXEThFZD
+3mHzs3qgIL/BQfmg7tZ7KwpZOFAbWpA33jcnN6+5VafpEN1LofmQRXBy+NecD+1
eKAPw3R9NdZeB+9UBsbnmUz+UVFlWBTP8f8CFKg1xdOAG+LwJ8ZS3nZ73MzrxL5T
0+FUzXXKUIBOWJGRdhjYBOGEU+FvCHWNnyYIgZ+Qx3oJ22eeY18GSlG/6ruiHPPe
uehenaxgwmpgFltEQHedzN6/SqCaSIohFo2MVWo4M9RhxHXNg4rBGQbP+VLJYPp5
0vpYKX6MoUyi7GrI2O83366yT18eogg4uF/knjrWJoQfVNIczUxmTgvNdkAhhCaW
CXDwRMO1jAhYDzOscatAOG7Eq6WyPq4plGLwb34As0XW9Iz5Cg2Z1gWwav1NwrXI
hv9wfnoyG4UtXy1DJrzuDMIlN4MGwXW88/2XDx/dLrNYj/XZhlihhOITaX9zuldB
S3TOAnXTZN3XyyWfhy9MEXVIUDjm0tP2hezCYr/LgwIgIaQfVeT7IUEH/XbZVIeh
kY69nUt3ZR93gM65CFMoy/LJ2M1I5VNeF6t5dtM3vK97vhce06xRc6j0u/oxI/k4
gH73Sg9zzCcjLDrAmd2cNpsYSISE0yxGYG0bAeP3e7Z47D/OnjwAT7tLmbQrU02L
cFbhy0HSL5woEp3O8UNy3fis7HbzNld7Ralfr/dulC8tbj2gRblqwOxF2KDIiME+
EbxyKKOZtgxyyM+8vsz7jAEuRiTtvL96qReLS4m8IO3cjFRqz9VU6VbGcJYAQlbU
lr7w9+Vg5fBWLMDZBT9QtQGMMGWBYA58w6LxT9iEDUd6H5QyHZDaSHp5RgHsuWmq
OMtyqkEz6h1yi6aJZ9hFFD8FbTUGW0qWyEHSkN2j5OQnZHY7WaFtaczsnq8Kfd8H
3X7CxCbx1F0W82LO5AbegQxMBwfSOLRkbEd1UwjEtIpQKNMJGno1YWUkF09Ku/c7
T6Loag8TgxpGmJZZLiPM5qA66KEof1H52xDoVpzFEg1OcN8d5SWWKXAV5Ur0LtTL
zoD+4YZPXKK7E6MGXIxYFp1DzoFTePNtu7VQTd8P3AfBNry/NG7GBBblCihBqReq
JYTJA9ozarmKhx813C7lOWXbJnWz3hiIeZj3W7MRpZsdbwjy4swSHbm+YMKuBLq4
mjGLi59fEP+LjVgahHXO1BiV+N2PggdEp3zadJMiyXRKA3MbTkLYsvy2syZ2DINA
vUdsr850FBs90FzvSfqqzW5QwAyLvSHRbNpRkTHnvof6Cp+BCs1tjqweJYsbNVx+
TqUmBA2XYtMh6e9N3LgBsLNgG5YY9sf1Q0m6wde1DiYtDq8G0PBfdzsazLhoBwFh
C9lMIHy2FSD3iyE+Lg7nsICEuKWwuURQh/yx3KpDX0g16CiCR//im2+5x5POsUIX
f0nIwKc3sjMHAFGCcI64ihN/0YaeL6G1+RIWw6GphZwELVRGsZMZS6u+BvloeFCo
GbAXp5hfTGYEo2EKiPtQFkYjOCHrNxm4cL0N+rPT7V8IJW6/ea8xF4XQopcZITp4
rKbdoXyqTOiYNe9FgQzZvqJSREzS7s+uOS8opOkyPIug6S96PiOxxALgKUdOTZSb
AQSy6v2fsZYsfCx5PiFtY+FyLf9TLXJtKdfMaa+FIsdI54OTjYuPBC9k/XGGl4l/
nDOGTtFnJ3laTvB1jGYt44nqXwkXbpA+pMCsqMbQMYJKpM183pX/7VFoA+ZrvlBD
zy16J38+F7IV6eSXj9Gwo6zg+418RhKHn+HHuNz9Uk8uPSJoVGf6m2pDbalk4ZBc
gSaBRU6In5J4906GCTmZOYJVlNuOXxTgyAp/HP6u004ojJuhSsxxz1IcVxdUij1o
iUnu9RjU+I0Lj3g5Qz+AC7U540zXEutVCYLBbspdcxLs3SedhwJBwrJRowSKltQp
a7xBBjsj73Lfo0kQn2unI2tINasYFKRGQ/MANUIMObi0EdKAwVZBGOhdtNpgH2ia
BOeK3wzQljJWy4F4Fa/zijEmJ2CaofXkoJnk5YWSvKWuN87VRKpfdwQeDbtT/leX
78+OZaxxyfRj5AreaQ2cfhuFKxU2HZlPV6mbxuNVkSUIS6hqdwQc5i1DYm29nI/4
PtsXXZdKGmzmL5aoLY9hSXJ5pAcEMsJhJ8LKuCu7ndXUquaJOIF7asSKTIudpDp9
FCoJXpSfmvK0U10m7NZ3dIYIXsXbjeNHLjja4SFmFN+aSnJ15OtwUUE2od8THMIP
FwOLKhivr1zto1XNjtwsEBUvOobv+pRSfq/uF6+S8001kesqUGT7XsrZCi5xC3wo
QqESzKs57EdWLyl57SbvVdc4X9YbDzIpyGb3ikpfvidlBWb+vlUcDQUKTPYU/BSY
pEWzU8Juue6juuquDz2K65XSijQMhXhsvq2msX8XvhK5YrckIL9YEd7zMfSBXOc4
I8+mPbfuZ9QYtNhluYFpS1XTsLyo31cjIpc5wAUoA9Tnug0spl5fc9qo8D2jkRQS
fOac5fYenE8QRPXHH1Yxs4mANcRuCFp2mqGZZWFjz2dGha7/gjzrSFk3FW5aJqqC
ddOScDypJmSotCnQmkuhoApSPQkLjmMcK2HjtFd+ELgEtwDXlwKgaApltyQKBADr
rGljIvryzYXrbR0FlnhLyedR7KXBTJKB9oM/HSkV8YTyZ1vn7/Hha0tI6LOpTJOm
X7NngZ0ab4EOyu7BL65/wzHoLprvHFjH2FNZfCB8dZq4JGVtsdRRuT5Fn2qLt8wT
m5Cx+0H6tFEw6JSoJJntNJyPBg6Yjtbc9zNEO6VsUmdu4c2a/uWpEmd2zPRBq+Du
XizLqAu+Gyi+FhHXXnhGAh8lugroO1s/6Wte17zsD5ryaDBo3ejC/BogM/0ESYjU
dVy3zRVSTSBemPJgg8+35MmRT3ZbdQpI8FsInD4P5L/CCNFdd7YoRDqqgOKfYXr2
HugQLKpvEFuwVNKVHuhEFrTFb/sv9PeDk/chK8HoX36zQToRkSD91nGf5SAkTy1H
rFSzmTnsUF41BI60r6fQUibreNmyfOMZ9ToAB/0dLMcPsojNQ60TK/kqnLPlvuPx
QH0ga6K7WaChiVhJSfWrf3CJwHx2pRXabTHvs3TdRe/B5XeKsavg5VZpxHlF8sJr
sjP8KCBqwLb3+S6SQ/yWDgwMNtvZot9Px5L44oBHeesVnyvBJl2EiEynfo8h7AQH
slFKpqi3Mr+Q9vJSMdhovSJvc63yeXCTrfmShg1WYkAkmvx5WRCKQrzC2MhlknI9
IGFgOiY3NKQye8heZtiotGedAOnFMPfh+POjrBnTCbAgPn0yEgL0uj8qSCPF2hpt
qpatqnI/hdk8xCm+7u0Da0XVcK0+BMmi8BlOq6wHxc1oN+QEqm48yfF1mv6YB6T8
LYRfeTHEBQ4a1pv90ee9nkCHr/uT4yV8W+wlNK5cHce3r/dM+Xc36tblFi3QITMT
XwEyOvXpHIsRBZd0oKDEApfyZXRYy0pnc+ocfSLfJkdCu8O8svsw/tONiE2yXn0B
LiVj5J7RI3/iPEcPY86dEphW7LuK3zQY8RfB0panvKZDYUzfQnF86c0LqWfu6IeT
49lM0XOOrz8bveDtCUZQ6+nskrm9mXi2D2dcw/X+rsFz/iAs/gifGOr6qNm9CU9U
xAq0Zk3bkJCtdSauegTioG56EZp8FfWvwK9471tMiwFWZC0wMZQtKEtmC7Rj5snu
n8d0oP/GeEthZKKRsI5eDZ0h84Dq/sJ3KX+2jxvRSa3DBZuFow+9gfgND9LrR/fw
dWFPqMZri6VPnLR4L8ErZZKsQKn1g5NAJHXn8dNGjSeyaRi7zjo5i5Rc75ajgIxh
TCtLIPFXfuN0+iXRzgKJOAYCsQtPlNsQbeQ3xREvjuB4EqRDDxWJax8mQtJLI2JT
VGLh5ZMyvu4he8x0CJOWtqZ/um7udQQ8uBFhly6chKbgdcRyw+jvQTbF2nVNH61G
QnK6whPc0xFMUy+xhzYn3nuy3O/VHcrrsJhHf2sQJQmnDTDPBa/Oc6nxGa4QmSXl
iwndlDlaeey7x0+UVNg3IAeP0vxZ5AxvQHfn6p+t5nRghGc3G4WGXjdynhU44+rt
v1XNJTNhNigoeqL7V5DzsRG0rlSEbZVua/3UjA7MmuP+khZJsITY5IhIHoZ2U8dw
E4ARh+DyQ1gSUet3UueMNKJs/MEhrGedB0T6NL+bsJ8Uynd7tqa7wxyM1/sOIA/4
5yiN7XFn/NmFvQeM2J1BtbUFM+5lJpjr/4J/jdsqfczhjhtw84u5ADtaGcxfTWS8
9LNOap8XjLpe2xjevg0/L+KTxHN9rLLLhWQRlb9kmlBAvA/5bteokGB7ZlSJFlEF
68Q5wUr4a5kI3fickR757N6TKPAghUfXQmOIfoRZUXFP0aa0nxMvbDZp2tADQcXF
qnGfndl0L11PTNiCec3DS/5trskGmLTZOM/4LckYCDO1ceYow4qhakSqgGSmvqZd
0lbbcSDvIuKKXZHieS7zdmGP5QFmylF3M2ozG9cGdvtrRcsHU7l1MHyj2+ZRJNLT
dJTE0iaQaP6afbFMNBtV7bXlNVRWKvSuRG8fnatBTbo2Vrgg6f15MXVrpFoqtZLV
9uzeEUpbVnjpYQv/OsAYhugibb++V6ZM/p1VeOLrU4Qfs7qehllz250P0/HJq/rK
QKGM85suOElnZzNL9elH68eW4GAjFuVksiNCn4OKjsMlu1YQX5QPITYMD5i0dgXQ
niXbjbLRD7UsYmJ63nWlGWt07D/JBRlFCGuzfyx+DnFC1Q9B20GPjWEwHFlze0PS
xyWhgZ2RF/ueyttD2RK/fDHgnHXUghcKFmuhMR7qTvo73GQ3xRGl6m0FaKYUf0td
uPjk1u3w5uMGzJjUO8fMA88Lh8hZJVMVZJ90wiQjRbN4LXjcTQ6OgccrG5fjRb+f
F/5nCaFfsYc/PppXt+rQZO0YN+C6BrX5iYPWocF886HaKM974+R5hEVX9nTUa0Hh
J24HCDPseGkpuT3/OsExF4uzwXQngQHHHwr330CDFSVjjD7BAMXfwjCw6PM/Bi85
9n09YbrkHqpn7n3na+xPk6Gs0vAdX5ex72Ddj/3OVJ64eEiI2wHJDvVLalrw2UlG
OcQpyeXBf0PNUNUQP0tVv2l14C3zQZA7/SA09W6YfV5l7h61/p+wl8X1VNs5Ceot
LWULATMeY8MNI9pq6PZ844Ge84b+FN1ArRp1yUWTxaPgN3UFYqnZdjuarFWCy+oo
8BD9h8SAtxlb9z4beTwbUxBylGFUxN6MBlw4BU+sx8U3xTWZQ0ilXjyk9SbzoLsh
lT/b6nd2vGTvccVFGwoH0tpMTDoEraNk6aFMxFyECWw6viANSnio2syRmXalBUx1
Nuo4QBdHJkO0vKQRIv/zcCsv/z1C9BLDIoRjzvOF9xEzGR19zxGm6sz/gTJn7x9T
oBZ9WMZAB12D08tWw4YZNqrDcu5TDTGxl3ZATfoBPpY/23XU5nY/Gg+A4AyF/j9v
LIn0xRA3HPPZNPMBDrxu8Ph1lqNBkg6MN4M8KZn0Qw99RBEp3angkEpzRErEvpa9
G6NaaYb42NLfcPjyLUVK2lvOaYsG+Zg2N58NiYmcMHZaZ3oTJ1lvi797a+hGeXks
7SAt22+13VH/Kyu3Z+9oKBs2+e9D3LUZRNlY6q6UTJWbETOeA6W+w59FlyAqaRV7
nsQm6YX5174KYIysRsPy2oN8XVEx3mo+rDTO8/BeNO9ZnTWeMnQjX5JDCPKf4YeH
sVkzGf6se57MrCcmC7Lfu4hEifigsUhAecLYWvb/gbobfIWhrAjoI6qs9ByZJLUT
9z0oRdW1AngVovlQQ0t59TfP/cwvGQrumR0dT0HmZ1BctKUZup+o5xHMXw8ptpWk
GzBObnjKGXlMjHbNbl3NIXEgk3eK2WliM1FIXXrn5Eq1KGUMa/wXS9+aGiF+Bxhb
Fv5PKHVqe3i+Tp8JFQTbC5+IS41F7eJH1OFnH49NlGGiB0e3BPA54UENEj9CX5U2
x7eP3YFULrA9/u9MRWD5thmnx+4BE2+JCBkWYvIxbzaqcYchSX7hpLAOe2RJldiR
EbcyyoLWjw8jeaCtDwH63FiXyxnJP1rUqhX2Vw/7j5qilzVyFsbtyhIdJfPe5uv4
DwIAuRouwqBlFY+5+WLZvjZAqh/W7LprQC4YhKEbvbeWBmW+IoezfHywpcyNc2wY
pOkhCJikWXHZ45fphsPeMnzxZF4KmGiUuhwLSIqEdFVpoFie1oi4cA4i9+UuD8y5
Ol76GWG486GBFctRiNQTnKz08Y95GRuX5owf1/Z0sf2dl4t2YEpaP//iRvd/lfib
tewL1gRZQ5nrbKJSpVBLViZCWXmVTILsASXlH4IK4sygV/xuktKZOc3uhhXa9nzC
9yYeMjsCvzCiMMobjvodPfjm/ddxLJEclhQdlKeD0mp/zVazbyvE/FdmHkqkQBgY
8jW58Bq8r5sc08iROo2klNufr/Cphx9HTDHRf/yrQPUDp1TeCTsfNZpGgZfs8DY+
yWkrmDJt789WMeN70aEkXGC2hTNNBlqOAhaT3jNUis4EiGDw6MC0W7XQlm/c19p2
ZiV6lQs1vKxzTUtMJW9lPFLQEwDKL82Gf7iEE9SCqQABmJhXh/n7AgSQDpAl7Ahx
Qr2f3zkdspw0+cHe4NwClkfFCma4FuYHBe2l59rFn5+JMwY4YX7ApLiJIAhfp7dD
Klw9TreayfYsCmBWrk8O50bH0l0NgWaX+yQ6onQGiSxQbKpjyzdA3H2/h7YQk9sp
v/8svypRPtAtO/KftSjFjeHIKwwD905Be8YV4+f7eXrKv/SozbeSI0MI3wjnmePV
k3XTgDUtAbG1+m+ZYiTV+ih/czWxo7KS7c+WMIuU+aL4ZgHLqdxcNa5iCLvNBNVV
+L2TJSmOwC9tAEU8edOp5C0TH/OMMLFy2Vhy2/+icFvQu7FX2W7pFnD/XPAjLa+i
AGyGvT1hIEzB0Fvx1lm+BaltQcc3TUNprrggFnZoYgzGY6AWZ2wQoZUStkxdpc3D
FQBJep2lulMgT8hlOH4akGFyg0Zw1PjNQdBdzwWH4Fgn9Akf5lH0YcqAigLATnuk
YNRFfPphb68eeSwE5TcbwWTCsGmJww9iXf+dVKzptP4ymwy8+x0S5eLxaFuR3q1j
7Rd9uCBe/mqQPuvyTAV0UNt+IVY+SHywNqNWIRlMEEMh8Bu/zVJUuTzEjZdj+hm2
IwCEXJB+248fD/IRbnnUoi+tXCVQj5nfuPxnCDV6bTzso9pW7mAUCDMb+TggusRJ
qznIr/5ltIQBT0KHsQApZIkR9UN+rg/BnYuPYDRD1Tb4CxHoB0pHmsnPGcl5eH4p
/CLTl9dkG/txUIHX490NIv9/oAJDPNEHp4P6TjZ+eXJNmrn9IbbbTrc7T7tOJygV
OlnAoY26rcrVcI243t2QLgN2yyerNOoVSa7EbH1T2qSeAihjngN1z9D9lScrcBJX
v9aSNh3uXLoq32zosmu9udXRST7JP1Th1F9ugN5wITQQzxteLu2+z+mv5CtJ8LGy
ByZCXd27cT2p9e5SjmJRqo+qMABwBKqAWH0ko4ZCqf9/GWSdCvVNBUVRldA/tXeT
gbCEyDbRVzQMkTI5GphRxZqeb9ZhK3LhYjYkkgVtfVYJFO+Zb1O1hTmWLY/kAmxL
JIi3a9/ojdSPepElo3PlpC/WU8HTi33jm70gcx9JPe+dE6KfiWOPkn6g6tkMGMAE
MqCBywOrp8OYdO2mHENTeyCVChb0wGA+Nf1GazT/9g/xL0YjYWaGYWWZL5xKUQjn
VvDKuRQirlQP4x0RTd8jRgcsC97FL4c+9NjDuy/JzTFvrdz1diJFt9E25LzpZTBI
TO1+aWpo3MZGFOL4Gyv0mO5nio5d+sRICX+DZQhK1lPugRVI799POlQMUW8F0H17
UN1IJ+NFO7+Uy+w642UNYPDLUVb+8qG0oOmcvorMA8xZK3Qwc3fXRw/I3KSF1T8n
k7OE+7FBo+zHIR3Bk5axvKdA3qg01be1QfFVaHDSyQyv2YQDTyE2ADs9xwAxGULi
N2BrZFHuzfqNRMgwCTHfbvWdfvFK00upnf9WiGtpv6o3PhcuUmqBst5XQRxLUZU2
tHeQCEjIq+yY3pVBrfD+GMNxmDCoau+6cSV4NwXoE1qjGTjGnh4r+VJe/5p20oiS
5/VAj21b++kAskay0UYvjI1yIVZuaW7uaH+SKp3zcT2/P3M7kC6Zj8N9L5KqbyDg
DtkW6r0L0r0+yA4XOqPXsK5s2RHkGqTr8QD8t4XsBqyh2eZsiUkVmzR0sJFjxgAM
tJoz5BYDDK0viBko2porFdZczh9bDuW99zCb3LzIVpKH/UOtQeBdM7+nxCj8Slji
ibRZLy/UT8J8ticzeGagAJ03quUtvMpobrfqMcfvod2fW2pd2XBR6MvHHxfdCFb/
VTUWhi/qIsy+OHZOp4mfuUbZu/4gEO/sxYuazC/vF1iqg+gZU2x+BrbysYb8x5bR
nr255Jr1GpeCp4P7wjJJUVZBtIozLTEevCnDz6i0508vg4lfX9Q0nRpAJsnDicTX
xTrzczY9715hHpinn3OY49ma4+R1J7rWwKrxkyYaRUkGlaTIyYk75j+MMlNimYnC
cycl4awHLV/oidmcMDYaZDkQtLDXBYi9Y5PGB1XbUhnqmASgJmQZgeA79L5U/Mlb
WKORxJnTwpSuQeMqE7WUiMBmxE8GrUIPHpgXIgPP3dBZ/HJlniyj3e4rCM0NPwvz
ibQQ0RwohWawPUk8U5zfYC55FkG14kli42Z69/QBnKJPYgwMgLarEjwpVxc89Zsy
f6KTZmomJjCknd6QiN3u1XcjWBmvY+QL82TMW0Xtghja8ZzU9SFOqmVY60UcbTqP
bRdO9vCiL6bJ5NiZ+/0UVRrxxxNCJpaDikztu92iy97SvQiFv2LxilOOHp8aKBhn
ItneEZhXh8Fp0WZ28PZRQjssFFWnGLwCEEtmZ3A2tFxKQyycXPa265XfSHWnMI5Q
agSEirw3wz9a8TCcs39SFEbu4EI0ft9dmZb4BZ+wS/qEVtG5sx3KuX+qHl5lyOWH
AjVSsePyxXZ3o+Y1fYb9GXVuJFG0GP2oKnbAkMcPqNWwcQkyDz5TIvUHkYxLyREA
Wnk+kDXL+AdeswhAKeribZWB7LcNZfUf5X20Hp6V8upu9UnSJE7n07Xcp8DUYY8y
YKXiPTkfL2RlsvUNCw7WMxPvxo5ShnBRbssmweORDKOAHirLJ+PnviuG0q1aoOEy
O3+BXjxqiFFpfMWNNIOt6d3xcfMSsxBBhUU7Qo4svhOGW34BK6e/NNi7+1kbRX4F
jsm92buKV1jQseZGZWs9NPuq6Gum55OAWP38lnauU3Mstl8+s6H8JoD3CYYiZdiG
6EReuj8KrSnYXZYx6sFEXA+UydyG6lMCB5l7ERGdwuKolteyVbdZXzDr/tBBN0Cw
WKaTkdHwwdL0AasQpXiZqSawEploMO4vD9MCv5Tznj5CKPcS0VwEFBoKevhcXerd
yqSVSlJ+5C5hnP67achajlxT+ZRUUqbXPbx7co4J6j7+Eu/DqueS//QY1MvF78qi
Gv5A7McNKG+Emwj5JtlIbr+aB6xKra1MNFucZHDpm3tFJBPVdOhxrXEox93vGXUh
xKSLqNyXh47s1ZQpI1wdryRYe/+yzSsmf/E/UP9V/UJqLhUSKpKLkhKjbV0pkKEE
Wzc45iyq0b/u12DPGUVhCmaB6XZYL9aDjq57dMe5OjyDIyFjeXwANMsJcSQEy1F9
0e4d0m8Ux7makHTpHr/WQR7Qsz+Odl1gT+1J6WNZK9u53AxVN9mArse9diUI7HkK
Pi2+2lFdmnIU/1DsXRGIo3KbDnrG2gEaNtZSI78hfaABjwdkaPWxwrLPnAsbfLGe
4ortesjP2R2yq10sCitWplN0PgMd060XKu+xnbR7g/6axD20qzsjk+ntJySnaTJE
FH/rQOOXX/vjY2K6eRBxdqvWd2v+HUtbwBooh14fl0JGLEPSSdfbc3/maAHEwhdN
xqNdy+5fBGshzoKmOzGKCYvB/DGlrGFQ5/7ka39brRi+/CUTcLQvFCMT0XR8WxYe
wTvisxDhvygcyv7InKUnEKdRuvBIFxtJiRRKXttHjozncymO/Er900+VjjQlfgBP
1QJ/PG/Lkpg32At1ul4G9wEzO/Q1huPfsw89V/aT4h4FYjGJBg8atcU4WT5Dn+ST
NO6SBl1+9CDtP47jZYkW7k+1F3n7Hl+n9a0zEhwO6s0anXIA1SOuox8dPGKK3FDz
agYys6y599jH8uWVaGAEti4+sf3DEnvlAt8x3ZziR+PNIkShfAqUqY89dyEHO/YT
lz1h0RRW4fB3eZKKSbIsSw1jh6KStMtsKuEfnI5OjPNLsz3nCAPff/u8JtIQHD5o
H9Vhol3QS62Bp+6TVGmjMsUADOdZMHCkwRThU3nOOxRbW44Aca+K4czbf84IytW2
DC17TXdjO324VZkXs1Yio6ZiJsXfzYXud5hUhMeSjWdOgaxy4nQmj1dUIX73cg/1
zfOvYJe8ClgVF0ybbXizGfyF90HIe9iliBuTr1nYrHF46HeGhfW1rkLlmhfar5wR
NWku4JpxI98fBugERyijGH7mmh4VdaJjAAiXFKjVasPq/WNuOY69yhxXCP3OkwUH
9c+r3z/mEHK1renQlbbZzhHz7+3Rs48DPKmQya4zAUYLNCOCSLVZmiaXXzFZJCkN
x3/N94gYsjgklhUE9e9JmQzGks1wEJVEd54jP6IThNOwVz089ygyLZD2UCSIHeyd
6uHyMWO7Ma4GzFKsyL0hhrIjTncJFHMgaR1mldapZIkmlG+r9ic5DOnvPwXpHT6E
SdaBLGQwcX86f5UPQiD8IIzIl95mQFziKc0a5yuMqpwBhUbHU3Q34YsP0LsBHq9k
eJ2U7PMm5MrJN6QRxwuofPJ5C0NYrcmvWemesAlLMfDJnoqXOXDl3UM+CDI38mL/
cfYWvO88je1MSrhFaRREbEdc8FTZlAwNEzLQJHwga2GSybCY6293bg8hGRmqDgoR
IwyFa4rfN1yFDFeALXHgjgYjP/N39mB4yeWR7PwiZCVMfX+NOeaMIp8ewYzW7aGJ
mdvigHTt+f4eco3hC/aguyKcx4Bz9bO1OntNoZS8wDCQt3nHC3xlhw+g8Ww5BmCt
3dO5olYrvrhJJzgaonw9LEKOW5Jvn857HMopd6vM6oVdL/l6OFO/fEHcCMBgPj11
Or10yab45Xj4R4GRzPOKAA+9ZD+LZXGlQSduBFD1jROYwTGQjHfGYYP41DxX6vsz
0amRpS7Y6Ir9ueDyulUesiVqjc9vEJ6nFRP488dxzDZnal0sjn4EZd47Ov2TAi9V
FFbQQw6+20DOWvTjew/HeCqSXRfzH6ocgz280xxtP/5LrRvUvvUR+ozw+dmmrR5e
h1cFZuZC1dxrhOoYbVuZQckA0vhd5uylUG2RtJO1jwR0AAHmehL/k6Lz5WXaBnnc
mxMe/tUTG99Wt3/PbYUQuBwnHYOZva6ofcBpjTYULjOPajxCWm5OLz7UHZueT27t
ubjK4L79/AjY6ytci/v99sKDZ8dxz6OXaHavCFJmkLGurKYx2oWfM9z6IA8+iRrC
5MjzIUx/aoayIK4owH78joBY1J1iY8EOpYAdZDs9NLUTK+dJnbkwBzNlFG8TyXkp
s3A8SDhTa/CORyczlp71obSMbK4eL2v0rakFa4xhOMTjb4snBL/77tDi2BXlLyIL
3tOAJxnvOU48HzP0mdfWRnukrQR9ITf4bukdig1oGhCFIV9Y2EV90A5f9+QMuTjf
YTj0WdKSi59AXImQjMRyEoxzPE+PP3YTwSw3bsJkNRP+hBEo4GLi1ZWRISz/a1hJ
UTl+aL4lj5g+TPz6f/5UQk1kuQ5B7a1Uuq5rBqUBrXECYu+cGLp/lZ/nvO1/lUWJ
LeOEd/lkzSXx2+qShvIo1Keff03On+e0hg2LeyeDDmQg8zQJxTzPpqqYq+Ouwh9D
EIRfOjQ3PjmUhNTr55OlFb/JgXJcurEv58KEuNjZwMbE107zei6E6qRcCC17sd/d
TYAhhM0prsJtyGYxPGXqYIWdNNfC3MBXs6Kq620MMpf69MxhwT6bo1ligRMu6Sjr
bg72YDHxMR0uiuiz1NH4z9SNwEUxSjHEHZVfENA0Kx/Y2lI7ur8JpACfQ5OCPpMe
2IyM/goHeLF+jYWmfG5nFfR8mYaHxHKRullG5Tb7MavSmDFZmLYbUrJ1g57ixihw
WzQ14Q5GzJ/P6yEGncySULPP3QSu28RlX3qaRMKhHxAq+mdNTAHlx5PZ9fzAr9Za
Y4LPyxbF3g7I0K/N6tqoWV45HLm2j2A83RiSmZNr1m9ADWx+t4PEKNGotbrRfBit
jkV3czU+2JJZzhgbcnpIXPuqfn4bGxfdOWytSDteJsLsFJJpXfyjOqiXjXIw+QWb
u4W5NrxR4NOuNM/+xq9sv/JECLkMC4DTKHbT+oJqJLhlf8cej0Zw1Zse5xqTrqhB
CN7n2YGSk7Hzf6pXrQR5695skd3FPUnJX9fbasyoPtUJnUBIBrUT1z3SeCij5Vo8
C8A5pDc/p7USdEYJS7awHSYNBnD0SQEfc9c7IwgiBi4iDQEq21qMrtT4JnALP3Hc
hOYWYMDsTZiNWg23UlQ2pGvOVkQ9FtD5+5UPyRtKf7J6K+l3GnrvZC3gyaMFZvE+
t4iT7S2KnLh2rcKv1p7THCoolvZEq0q4PgZmu4jWgd7DPQ6fIRzJz2eWAqsq3Rew
FyfRY0WwCkUllYDt6QMziMmCRGClMmyBDXL+0EgJXeIYPNRaPZnxW+3jjA423vT1
5RjCcPpNjL+TfuAASj6/6IUiIuO7CxcSXMeLbzrmsswv9471dfDBS+W++6qBv0DE
/W8+UpU/Sz9VhDxy0QeImoLlQSewugBQDLtiEapSRjnckpvqMznKebgS8s6qhoYN
L3S0omuRUkyMaOpjOlL6qe0OZH5romXY9Q3iUhIKaKECurpepDcianpG2athdLJD
+PA4rVPVVcqKcGK6T8cyW7c6i5PSsKbaEp37QP1YvEzQflx+pRRvmN6VcC7zXsyS
WHbzpFSiTEevitdyvTpWXVeHbjJd4VkARI+Zn+vC00F09IfkK3wlWWAyWWLLFKB8
`protect end_protected