`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
ddtXksX2+yylW5zu6QL2Lhnb2d1sD00763mmSITNX595NcHTEkwn0zB1Dry37fOW
FufOhVzEJp80NC5qZ/+F0Vk7Ik02dIR0elf3clrjeJRK85K4e3Hoo4xn7YbFUIms
l/8VZSb14+JVGURjfswrIyCUotIzlzVYZ6gzoZwDXIi5gQIBf/gI+KxNXPaKV+PQ
Ufys/12rjO6aI/pPlqSm0hCvftmBcnezN2hk1UeXgOIuKZnogjOsf0iJVX2aOOWE
6pD/psybjbnsNB6kH5uFTA5frkzIzkzl5d9+YDm9OyC+k84E83I/7/j+rk4L2dah
QJOvksSIzN867/4Qt8qYTQ==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="MvBXkzurAa5VTw+1JJ70nePUfoQXBvZOku/SMmg4TwQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
oRtzZL4VJ4iwysPsC8SXYCzXS8Fw2gtZTOskLcDV+1B9Nzn1zTyNtlo6lNICRmmK
ZRVu2BmCc2G+fmzynYlNTnSa7C0Cuel6FYpxCBlOuk3OF2tzAmLAuDyOH3Z1Yjzk
a0aHuoCdIRKv7BrZCdALt03JeUmXKPdOmIlkVGFl8yw=
`protect rights_digest_method = "sha256"
`protect end_toolblock="Jn9CQpRhJt4rnzZPRk+dOpzAubz7omckX1MrFd4p81o="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 1312 )
`protect data_block
gD6l00tciPUa6pDNTk/+tzLxvdHE2s3DQL3/JqqujQBC/Ei+vcAB8wM3doqg5vTg
mdfn9XB1bLOis2CVSfu295W2DNwHfMSTc/8BhCDRnTlLIX0UCJs9Za0+LoM0rMrV
T7EjVWppbP+Em6PkVKCwlmIQ7JKaifJ+Y+kjw9HCGboYo5074hY+K/CBbfsBQY86
6WN0Tz12WdSSpD1yvN1Cmmgljq8RK3d8Ri3D45vaom+QRLUnZUGFtxSt3CBNkALY
bhmWnXeWbLdOu9ZVKvlKPrgKkFq9009GXIKsKNs0ShRYhoHCsrfbmUlHyWrMCzTj
lHitxvfl7wm6JgBBTMdMZ89I2Z5RS2D3I+rzpD85YUbMPXFpkuMohZTSdxSe89br
qdC0LyxXwMAEyBVVeH/1IOfx0SDkNG2oVTZy/wyRKJ6/73pbcamWYomr2yyG68dq
gTvT2bxuyFvE6YEjdx+lSrI1vEB+opQYJqYaZ1IH3H2C8IrjFYiBCMc18zXkaO1/
qmftOf835XJkT2fJXQgLR2kHjrr2ux6AuL2a8gkuVKzfQoP9DgD0pcxE+SMX1sDW
8J3Jtu3be/8xMvGZWdbye3aECYf62CgehsLxsz4JjXNTroNf+QXdQvxJikn959zB
RCqOvfWyt64B+coB+wE+/Gnx03J9x0kskR8Q9qSO3PqO9kOEFuvQM67w/zOkqXcl
UwY3fvO/NHKodgsPXJQt86voALanAAgf6rsDqzPDVDap28piz4Y86PmZTU5GJmHF
xnpKwg/o8XTo7tsCdxOu91CvZue9NxHSfrjkvUT2vmi3jWOOfEAAR0da7jHYMwnj
fE09YFWQRLoslQaQvupkswOJnkIVnRiQxZcKWv1YdF9v8BPuY09h9t6GYrEz8iI+
xwWGH3ZZy69USahKh3HH62pC+L+3R1pUzSWhKUnoTpd5HUzCHWib2HCcjZPzk3F2
NFbjC/KmLGJdpIO+18lpyEEQO2G8Br0B9KCrRu/00f4DtS5gKSweMMmkrEPvLHOZ
0NI4CLeiCvVxRK2v7XzW89DctxT18wib+UvsDvQQBHEMlMaSDSmHE4tPSdfXIgzH
J4BDJ0vmXWEsSrofq66muqzUZ6PmGkwIbB6FDFrgIkkYj5ry/Tlsz03TJ4p+7zAs
6RC/mqPIsHksnAAE8tq0ReoU3lbW9XFzkdhJtm72t442PU+/uZJlqnuVY0Dx38xQ
i4Yonwryznsf0eqeswj4IJyogDXF7UEUFx1xYova4+k/bB/BqKXQaZEciJE3vQA3
wdjuCXmVyktPtJ9Tr7G8tQeEWKZ8pXld+6IGjYvE3kJIlnkIK0PIU+FFsWy5vyWS
GkyyBJUb+gwDVEukF6ZXfhZH686PumT2778FuUWkOobL8dgJz0IPFohBlYZwvVSk
r6J6eYWxZTe+Ovz/5LKQEfx7gsoHz5ERCVFJwldypsx+UR50gYrCewymCrLA0c5a
pKG1LRLfn658Cg5LjaxEcSzY7PbXp0RqZWl9S70coSv26A07G5FM2Sn77ehuA+a+
gbOfIa+hpJ/SU12eztW3c0m0uIUnt7XicLEhrrIS4Na0PrNnMnjnDBFLlVFLnDZq
KdiioDWI09wShVFaZ2GRfwS+i6YG26EjG5HvjUoqPLxdK0Rk3L9EwBdSqO1je31g
uOF2s6/1h6DYi0zD7ynNu/xzJcZogpHMDmPzeRVLM7MNehY4y/tti7aVZ6ItGcW3
5eLx6qCPiq7ECgpWpz44vQ==
`protect end_protected