`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
ddtXksX2+yylW5zu6QL2Lhnb2d1sD00763mmSITNX595NcHTEkwn0zB1Dry37fOW
FufOhVzEJp80NC5qZ/+F0Vk7Ik02dIR0elf3clrjeJRK85K4e3Hoo4xn7YbFUIms
l/8VZSb14+JVGURjfswrIyCUotIzlzVYZ6gzoZwDXIi5gQIBf/gI+KxNXPaKV+PQ
Ufys/12rjO6aI/pPlqSm0hCvftmBcnezN2hk1UeXgOIuKZnogjOsf0iJVX2aOOWE
6pD/psybjbnsNB6kH5uFTA5frkzIzkzl5d9+YDm9OyC+k84E83I/7/j+rk4L2dah
QJOvksSIzN867/4Qt8qYTQ==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="MvBXkzurAa5VTw+1JJ70nePUfoQXBvZOku/SMmg4TwQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
oRtzZL4VJ4iwysPsC8SXYCzXS8Fw2gtZTOskLcDV+1B9Nzn1zTyNtlo6lNICRmmK
ZRVu2BmCc2G+fmzynYlNTnSa7C0Cuel6FYpxCBlOuk3OF2tzAmLAuDyOH3Z1Yjzk
a0aHuoCdIRKv7BrZCdALt03JeUmXKPdOmIlkVGFl8yw=
`protect rights_digest_method = "sha256"
`protect end_toolblock="Jn9CQpRhJt4rnzZPRk+dOpzAubz7omckX1MrFd4p81o="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 14352 )
`protect data_block
gD6l00tciPUa6pDNTk/+t0OO0nC/UTtBwLB41d4inuAUA3i/ALrNyoJVcBnAmEQW
ptbcNp5fxEUJjnOxnedyZEuEBxWRieZFQnkRdF269oObX4kH1FtdcAImnMiXJyOk
jpyOH1kwFsBT8n6c1FCUx5bYv81O4iY6aTTz7p8Vc0Rp/g/lQGbHuhBGhEhNQbq3
bj8TALSjwsnpfdw4QX7WE0n+Px3/yt1YhsXJyCf1dDXQUxoO1iRpZq5IL/CTcLo9
Xjc/wZY0Ce+FHcbwaY6MJyQE5b3dbTiCRGwx7th8Fmcf/DEYLKl6AUjHYO1PfkWb
SLyuA6eRhyR8FPYMzUu/6MBXrB2MMT43ygrkp4afktCmY1cKvHoVQ2N4mnj7TzTZ
vmtn9Lv5OpJqO+OBzrWbvfPQQKBzyBN9Qmv414QLabkuLTPAlgT14MixIOEM8CD0
LfonSYucpIzRzA1s7LsUprsFg5jTvIRVKNYdW/lIEq7Jw2mslIff1G+810VdbfmV
eRTqtbOgyyUJIK/2kVKJB8OIH3CT9UXpvSACNm1dlJmXXpz2E/Q3V2GQVHasN6TL
R25gv30lq7JBiInQgp4hhL8Q90lc9MLX9pS0uuHjTIUWeTuaYc+O0QcdFGTNBtzh
WDciUsZJs3s3Y+dcDUC7FDyiIecMbbtIb8WVd8hu5cTS0K3gy0qrpk5TdZbOuzlJ
0bGZqHwPY07YcxN6TOw+OckDrhiqQ/KuUu2X45gNTmKBJ4UQT1mYk/gEqmeSZOPm
0fOPpngqssnyvqQDhhO3nAb5IflK0ThIJp/7XGyNdOItAWSIFc0v4Gnl4m/6Z1MN
D3jGfJccGeVtWfC+oim//R0J9EAxWWw3IozmCRlN1s6csf/ma/UvxWqNDnRIID6X
02rn2pd8BqLybt4j8pH3hdhXoqJ2vffsN3LEEl66i2d/JMt3E//rDPVfBgog2umc
KV7yGoAvEIvr2r/i0F3uC5wGt8JqQxyQBF4Z2Me3f3hNNn1jvyRjIaThjWgHWaEf
Bi7DinDgYaiQuTDnSGTGgodIR9QTlorQCZtS6cFxsUa2PLseW/n/MQkvlndiW2Rd
5Xq3rmYPPPUXrKA5XhE6T0xphlB2R9olTWw9DFJZW0DckMyjcSKNW5KJnIoeJTmq
Dsq/NvHAG8W9OwvD+yZMH734WObIweZownmloJzULJ759LG9W2etvHxe2OOqtUUB
PbC5Rx3pwzIr0OGx8p20yRenPBfXMGsyBzXhVkrzPPUIqnn4sLyWZtpjHDPy5TAr
OcOEIKkURWSIm/VIjYuNKPVocuzhtdAJxZtj4fT36Q7d7qTxiuJ0+fCekxfild1f
yLD5VcqIDKQQYFhvFdJeH+wqkRxWJBqLW+VPp48riV9CI9v+YQ+pBhA1SG364pBH
v0Ae9AwtJsEMMr0WNJ38ZQ72XDxXOCGmUoOQq6L8TFFZBEMMnEFwguukUlLedM4+
FMKseE/u1TODWxGJkA1eFpgn2HfHECowXbxNRETCaKwtakmLtiY55dS/zcbKLxgF
RkIWhQh1ol9TUOmsJav3yv23PWanYpuLLZ0e6nZpGLfxWRkW3bPzRNgDqv0qeRgI
jAjOrqJ/kN4jHIjVP4Etaubjhu2PsCGdWXwvGQr/rpGqv4GRE8ne8bylPJYMC6V4
mAwU5uzW3Rm0wpgdZLuh1T4N3MBySor/k+/5i4arF9+8Zfvmdbeov3mIfvdYOah6
fO64p+HbCK2yG1vvEvZ11HgPHWR2zNkBPMzd4D1aIXMgljST8qUwnGd9juQrQhg/
DoJ9M5WrrImFf9IJjlAsDzHIvT/I/RHopRmkNcnyWzv21apsblW2tSMW39j+W0xd
j0/sJ71et/Lif5dOfOtEXGY4fwUxYIwVZU9OblUmK3IB3jAqp2B+W9o3rNh+6Lb2
Wv4zp3F6x3neqnBoZS0yZUb1B9f0KidDvsgEHjGz030vYO9bjxQfbPHAShRYsuNn
L32YHTKFW4scbeikN68HvF9zNIqvnWcMOIdWBfsmAYqHwzIee90HvDUTfkr/50tr
taiSQHMEXjB10D2bE3KJafHgKZ9gctzXkkQV3nKrL7G5hmJCG0EpIB5lstg6qCSf
EFuEZ525ku+dzN+AvjtY8zLntlxRK5o/pg157We+aIIQ1Ur3L/a9ryYX1V5Xhstp
eoVZOV1m9DaUvotI13rwW8fKigfDFEFDk4UhXUeE7/21uwxcamu83ExWPRfVajr8
il4N9GYa/BigPpRdfMTZpglPEUH2ogHZ29Wq2X4s2CaBwTPJX49GdXCsSxsHgdjK
JyBkphSOJxMFFb3ZKMjoJopvb32rezG/UA2QnGNO/pLlu4oN9l+22Du9RMX6ZL0I
keWyie1oCVDHbVnlQpPDt97UParTg9SkOp3uokmxRRf0d+6R1GxEzP/6yCnpfeTu
LxDY34w1BEX1mzvZ8re1xS0JrJC1/vIJr27S3OjS3slFioYOzNATf6+0yVe2xIui
63nNAYRnWM168z806+6FIV+osom+RFky7d9vJbk7R70b05rvfrMOmybIIE+/QTW4
QfWFh1uQgxrR7BUO/bGkHlfyeTKhorgMA6w24bTWubS3f3Pt2KPNWOjas13TyWyO
eTGDd80eTqiPYblskNCzdNGDto/pHFIk9+TkQZkgJodFfIGUmZ20P0zJ3gV1vnF4
dzPlBZ9Gd+NoaAFKrycgFlpz2NmYNg7AL3++af6Oh7FUOrpiJnnlfCg0fYtNsFLt
pUyO2KefYwK2XcPA9yebZzYvE+6FWBnEMsJ8dtY/nItTP6OUEFFSSIJCj/igXbX/
q2z821Gkqag3P0BnhgfqnTHJiaxMp+hpmtW7DnyWorA3PdQGtA0111Nn9n4pUDSS
2YtyaSS/r5G4xvtfXxeNRiUDyu8HrChK5QX1MBKD7cI6g24ywgxkxZ8Gt9Hl6ZDX
ZM0Z/bVPcbMkpaI7O7o61G/Dt9Gg3X44BDcZaHhU4SJxkQhTDqGKmHLnC+ptZhtg
rxEEMIiW1qttACRic1nM5yO43tk43KSgsp+cnaMnp0CgZInZQWvMlkzyzias9bMl
kYQU58pQG3IBYZ7eukdSu0+c9j+AX5K3GwI1ipGLUEQLeutyCPFs3y9J9+CbagBM
vk47z0axuO6PxVRFTOn5Lxp8NjyFEWV5QVPQZMys0gVC2y2Lrz2ifHf9VFGMK3hl
Z0oaPV72RkQdb5EAUc1NIoYqfmoqzJfTnOvgq2VjGFkYtkWua/FaG+xCUivj6mmA
2SLLWwwLDgxhVuOy7civ3At9xDYPGLjrG0TA2A0FagNgjacB14gtUoiFBSMYSWY+
sa+CD5b84ce2oz1jRIw+B4/InbTc4c+DDoNYkN3JDD+7IdmfKmzAb46efrw1dgyO
VGZmoLPJamViERomaPVf27pgVfiwPz06Q5blbrwrqLeD/P1lbji9ElGgin1clPlq
5jx/k5673XgEs45cnq1ETfaJpxc1fn3OY6RuWCcRYM2Je8w8qbvb3wwLdwdLtRMl
dtdWkZ9gv6NrBNSoaLMqulctUs4+rH7T+2pvWNFTn86Nb4a3jLqOYTev6xhstxjx
h60X1xLI0SW2dsZUiKVCxvXMs1QpsNHaNUXryeS/4R+icWRdiQFfdEYMGOl2Yi2n
Lg3y/X7iZS45dTxiwtteCcqFF6JBP1hPghV1Ghgvy5aHjOKobGlFCZFOFGQMaYlm
nSIp2OBm4K3LAU+PYR45h30ASG3zBqn/Xf8SRGEgIPYLYLOvjarH+cHndGYzQzEg
4nd/F66+O99uwrrEHAZHuXHitNiBIXY++sF2AZ1kUJljLYUBferoz/xvUt8+c9u+
71FRSpTgdYPMzJdqydb3I28+koh4MZKdGFGq7Tm0RPraNAMoB+1Rh32RMTBp7mNL
JLFFyEwW4zK9q0VhUNXrDuuOQp67Uifz3wRoO+Wk+Yx8ztmVpHcIQD+dYXylcNIT
YTffA8+7TAbWt/rauM37h3pcojRShqEjdXhIVm2yDxHv6mYMBVpYvbZB3tlMsH8J
+uhkMmwrbLS+hx3XPwnwdg4BeZGKhTShyDG0320FqRdUQxMwYIcV98ZcaIEAGUGu
Fopn1yVWH+qy4ej6lb10UWdJKwM8lAEAYdyNC65v5jrTXyap9O/Zb1/RnAhtXpK0
3nH6UTK2bD4O0Sn44SKBacdLctjebTiGJCH1L0BlQJwpN2660zXFfbXrWKVgzo0A
HMf0+Hd6xWdc40zFkmiNiT5A/qN7JWBLbTjQIR+VtwC83ffb1WnaN0p2G8bHAT+p
a97yhKPB7B/cvzQp8XDmfcY5HXNSc2ANDSU76wsVVVvdaGhqFRlgy8QN8mTSOXov
woI/Pa5GkUp0IY3TCEfVP29N0FKE3T+pw/7zu/kgb2ACDvs1jCSqBqtAxuA3CCzc
0BurNeptZ2ooL2UiPMUE83fRTeDPxarKyEuwa5U+drzySqEHS+Jp/ijN3KGf0qAW
wnuIyVWuq0CLKOFAEgGNLxnVESQZG9XpybMNBlI7/iR/wVbJ2XZ/P65eCJQYc7C7
Miql4XfqunkWf3HiN3gal2WWVOlwdeT0SU/LcaMrzx4x+qQnHvJQCHkNPzcFQ9zq
/EQ/kIOszZVNnwlAzj+AQYDoZBBajg7UAjZ4SMHidm8OzKNPfaXU3FH8yVMe5wgU
Ym3gsv/xVg3/TQ0wGs4KK3NhC7inNeF4xrbaYtE611orWyJe6Q0ybaOQStnJDMDD
0QebY235sja6rKpbRQtWKoT15zqLhMNHvPVNQ+qdKtTdc5VZZCPOMrs/nuKMOWST
Aml+pw5ggpz3vd9P+YiUxlDsTOXTLlRiviZFILe38y2RgrKEbWdsAIiv8M3Vj2/k
a3L6ywtdJBxYLOcOn8c58y4KP9XR8bFBjb6y/B021QxsE+KzQHX/SZvli205DyA+
hzxUk1sFIfFasLbsBAZmsdyJdy7crqjNyXX1A92sMfM5A8l2nNOgh45zC0BsmSKX
cja/8G+xO5rf0LvroXcBDilxt0KRZyoqx38iaQQ4COVSI8D1OMi3hwlyxKMUs//4
r8vthNQsDIytcumVEOGNNFdG6dojzKmtgqyJ1sDJChErDr+DFFkbWETwu5BIGQ64
J9TvUBBm1H1dukXyfZlKCawONFRkSG0nXRprDSEC1NincZVp4RK8hacRElCFe3qu
MKLjeBWsjM3dnBevpP8NdA/wtP8O0xFCf/WaHmmaiyNfSRS3csI8xmTTetU6scxu
zgwgwg2z8INh4Hf/fILd0FBf+LdF7bLveAXP0N4Dn5TTU/04W07Q1+gztk1/UVTz
OPrvzABnbpkO+NQLnIL6Hj649p2Vni8F5XmTY0VWlPvGhQ9uZkX4gxipZ+9WWISP
ZPs1EeN4O31onwIniVZcJvZIXTmBwpmFQmnfqONO08hrExEX8CQzHCeiStgO69be
k0mMlPQcyiS3tkP6PwiQyvTedlUUNln58WE53+l9bJM9EqYLykwThfuoOCZ3FxVx
DwyDy3qQSdBYlVHHlcbPMWotGDalauQiLhzKxLyQlKusXks/aKkP22acIAE2s731
1u7w1IP27okIAXXMyhVlMYDTTW87fsKA32S0j6TlQUkHAN7S7wNjDQJeUEb/JpSm
GJq7aKWfZzUfHe/slgJXpgpFCt5/Ea9FOdH+TOzaaBnkOhUaOjHrbkwVKI9vs3cH
097ZkOb9C+hywRA0ncDev7xdWJvNYrIqT3Gbs/aa8iQ3nP/wOiyQ1BIoavoecktS
mcywyUap/TbPjDVTbDwHvC96kg0Kg1gzzdQsDu+4oLf4k7b0xPgcEUtm/qH+DuWv
1JY5mon2B2d8Gyq7H7+S5gi1v+i5ndZBc3XoE2cH2JAcyTf29HTMjdAMfKnpHsJu
6BWGqH+ZRFRS7m+D9xZK86MEqwQBWyobGI6w0S6G/fdZmhMcPFA926g9SBEagekQ
LLSjR9i2dh6OeORxbujEgKbSMREUmcwrzJmuiQNL2fE2VyzRXtABEiDcOdFNgzk1
w693Jl/OkcziOZcKDDFFt+qYA3TspLl+ll8n6xvRDL5XRS9DEmWXTvsGeLPaROxz
4a4DXtW2bh35bF6azx6Dlv2wXNN6t7IRB3aWmRJ4Ln8Zb60z1y1wbvEVY1TEKeBQ
/0SngcMntKUooytf3juMJXpewYZolWSK7GW5iWkMuYBv98XZkEAlMVUakH7LRv8i
mGu3Sy0X2fGipgoLJIybr94VBFNuRiA3xkQC8u5/XsXiQt2OYoAJEwz1bFcDkd4c
EeliQ559th5N2q/VbBlMRErwXX+ap3I4tX2Ih2exYzEgGC5XaIf12l40Gp1btzur
MPjN4aIJRYIxB6/dhdraZKpxkWGqsTECm5MD5iF+rUHqvorRbLKEW13rlayq11NH
rHppv2+qwuVHH8fa80QXqsdsCGm4PR+OYRICuVmRsQ8gn7xFLUcd2KP81r/Lxqf8
5XZRbRPNW3exJLiFTV4ps39EoiRbMWUrlvTtfrVBGDogrS+WN/9egjG9Ltp8awby
WQMuZKgyzIaGPC/yR2NHGQfmlOZYxXncPAzz0TyJEbPIsjumgW1/umxCh+jXpkwU
Tiu8Eaqpr8yR6Wibh0SqELR+9ksYr48J0WjGr11LtNrEup0IGKaMX0DhQifQHk4c
NEWjjeDvE3qPMggRuYKppVoCxfrGoyi+6l2xS2I8IHq1PbLFeixYDrKre/S6i836
8Zq8D7m9xzVsXiLr9H3TRu1xwRvzOuuGvmYhzkHkm6YkHl+iGtfzeIG1sBIpskxR
QmYw+1NmFWft+gOBqfwM5xQDjQE9djRUCQRN25Iu+viDj5VMuwj29tvp8pwBDEFa
wDE02ax2c8f9G2gBGvaqLflUYOzPkXpjeeOIhJktZd0BUyVi40EiMTOPB5sYo7Su
1f8koubCxso65ATDjH7xpLc1vGGo6msVMM8K3AL46btvpHNcntw+xUqFRNB13I5a
zg/hqTDpAtqlzfN8qtAs722bB8aHXj0e+whMcXtL9tVrc1OzHUX1jZwn3vi9VV6T
896xOdaKMyf66W6hvAHjUHo6hDIZ4zSMb9BL4/cPwfJI9c4c/BK3Kq61tCMIgKBp
RUswq95qmiDT7WIUeyqkdl4oHWz2g9MNpcj6oJ6F4mdun7t6Sp4ZcrAGtwbecRqw
XGcilpAKxNEKznq2naqpCXgfGQsLU5iIODtphKELNeCyzkIoaXlol/tTxy6tKTQQ
xXoDbCOnLUwjCGIyfmef/Z2GIqoKPjhfB2O1stG0UGGYSXdbDDPQhQmPW2khO5ho
wdGIWspJ59GgrI7xgHKPF6dYLIfXadVOs4V/gajnmMCBhgN39e7J+u65nZPAThZz
3H01trgv8xLzaXTQywoAY1tdmXBkqtULizapwxCMpBh48t8+NencSc9aLC3mcTN2
c64CyDW2jFokgNZL0FNmq0V/hlHYUG26/d9qEqawzWQG1/jPhXaPqf/2joKguSPP
lyMCIepgU2KRsVeM6XPQKvtjiirFTMatr5bGp3ehCpR2rlPflCog/Ax67oNpIory
rmDeK1QYKq8uYTg6JIMWucfRzvjg+sZzjN+SM7yuvbw590PkXx7IufyW07dCgjUv
yhelwDJSGvyU0rB5o7BooSF/WZ9qusRBUo9KJEyPoUPlvBiXmk407g2PQ7Clvxs1
n994jTc7QqB1DJx/dh3bhLHhfwrmxBxpqvABnnUc9QvnAMpnyxides+sYY007LEk
Rml3Q3mGU4dXdYF2sWCYKDsDHYmKiwPw0wSrqJy0AR37z7LYn9kDmnIfl09lm7hz
+xj1jGVXyT5MyWECvuQ9XAAq6m2exe0lUnEF8WOMVyT9wqvxG+v528WjnBEJSF+E
vIWPtRPCluQBXHv/fe88c1wTtxZDVOhuywzIC/+iJxrcmTdZcLuP7x0iwqXl3/UN
49ii7GOBSVj6dOnlzevWmrEZX4LYfj1hwHyvkYuuhidorCOKDff5Hmiy8J7yaPJJ
0qWJV4++T5OuYPqWTkQNZQLB7jYe21bD/n4DiEtUT9NFjxtD+BxdAOl7vr31w2dB
lwAq/de5drpkdIhNwD9cu1Nmjh2Lwb0l0O8TLmWBTg+0/OXX5+y0oMu0cjyO/Rs0
kcUK1ujVe+3DrQd2AWvktXnjk1UZhaDWO13GUilXC6h/lLJcKlGW35vJXZQHjNLW
Hopkdk4qmQ9ICZ0LuprhgmLCoPVGbn2wZgV7lDqf/Vk4o60q+EFHC762oZnDCnLl
tzwcoWCP+2TA0Vha5IF59huNfnm2V78pthJY3wED4Qk2R81p96tCmBeQRhxMUnoU
OX18ssc2OP/ZxfEt69ucYo8eZUJT8LXQJ04kLW3yzhGHVT3ssFdBbsh5FwjwPaBr
q8AcW/oWfpLhB0MqYNNuwLrx698z1dFIJsCabM73Jd/tBvNuMteK06Yz33aD9uvd
QLRcT7ZfHmitDGbDSTrntBr45ywJFrWwX9Zu7iqmd83EtGyrGp3YgommbJAzSHq0
svAr+0qpeEmM7HFRe4uthKlpS8nudTThyaVfP6iwbRjbQV9s9+0Tnm+tnM6JbIML
x8Ui13X0EQvfvfWKThkiKvw81BQOc2zHKO54dJJTCWl9uVkVmjXm5gn5F8Z6DvDi
qywOyLKi6nTkepUJELljy4HQ08o2EWoMwnhI7RBgzyyQThJ7ukY5/3qebOycker4
+pk4qVlcMBgu5KCErB8blltRDxTA2M+P94GChld+t8Jy3IXv8R+PxrCoL+focnGw
GHnIwfxlEOqqD/7Gm2DL7n2EFiqLBbuAzoAYfMAP/W0wIjJWJcsuUlBnmTp/CX6L
uNey1gK5g3VlNdv0qBSJ1oDU4ZLDJ7FM3r4R6AfXkxnVm24EIPjgI5Gq+uWZVpyR
ZuEx6BGJDLyPIMYyfdkAuBmAir2+XFlBYuFWaR+9xhGWRw8GNpvIhGAzTwDAmhcE
68JFZppcNXDu4Pcc7miDbGM1eKH5mdCJLK2cQov/sc4miO7aEg15hoqGu0XjAiEY
LyMY/hiGD0AJTuwfb1QC3Ne3lTZjfZlQy8iDZeNbh8IUHXDziBBydaxaD4I01Mnq
3mf209qWKfN3i+GzvtEpDyU9D5iNrAHoUAOL9tps3zB+huY9N9ErmAMbbL9HPxPe
nEv0mAmgRjblu2uFugJodrClBbG7nfp0C7j1JAGQXHZqiNMQ8y/gqMu1QZmL4nov
UTaO0pHPb6O2nvuWr/4O7MbCSV9N/fdkac7FnedbsXzIm+v4l5VdRbGlMEnR/pdg
XwVk5q/z5hChJSDQ7QZgnBnXHFEag0NDXog7Y3HhGATXadnOz+BxK4UO9A8LaM39
UW5zwGgvM5FwtX1nEnCzUuunM67fbVDYF+iOr4GO+jJXphYNNxd2Kq2X36oa4mEu
so3qivxwjQaK8pGHvbWOTC7qyUGHX9NZ3YlkQCLAz0Z2s5ZcU0OuNEr7yvUhMtp7
scnfiJH/Rb2ztLIzMj+gFo0+YT9S2PLs04BvLHLkFN+EB8zdGh4gpNmjlXQI5q8q
M/NSV7n0GMyjxOeTXbb2PDOeCR+dycgKESQJyY1o3UTr6qtqTXRaMOkP0LQ12lDr
DeRA/e0+9OwzI+enVobRZYPhzQoaGWAxEtOV9Rqf251MMeETSOYipou5vg8Fg8VM
nlSB+nBjP7OwQ1HWWvN1MGyBW97qQplNX62yq8TpG6OGjrjoHcWKanta+AaP0C/I
LSH+qBTL5UrWHCQiLpD2ApbRhrQ2FSQbuzNdbi2NgDGslihFcQOBtEi4ixWkqKDT
8Nzu9HHPnSrCquJWrz8+QY7ByGvFmGzzFwYEwXjrusWxsdYginlkQHhzG/Gne1tT
EQHejuNw4z/mqHOjphoLMQaCWCCyOAY/Box18TWx8n2wxvRa/KqdMNPeolctd6fz
AwmPj92AaWTD0CXCT/GbSPXLCOeU68rPbOlxyGk33REMtXtDPO/iprY5Jnas0sVC
8jSbC1zLFi4tq5/qc4JBxdZSce8UmQF8Ol9FxoQxLFGL+ZGKD/rfIT7LH2X+dVXU
LarSDqbBx849yx5ezSbhtIb5U9l9y9WY+3gmekd+gVjLpYdTWqdshSxj2FTYhej+
a7KJ8OIRHHk8r47nanzEAw7fNqKhKKyjsbUZ2liPllIRWkuBh1jKZfRQjKkfMVAv
KNW47eJM2PmMg9HBFJB5TvBV+FnUEZ59auXaKf+rIJvGb4NRF0Vh6gNCnvqjYE/w
KAaEnBnrNPjyx/sj0jBGivzodpVpEzqcK3is+j9gQVfjj6ErHLIpXzttviUkvG7X
bqDaq2U7E36d65QA4QkiWHAZKMRuyjeg3WEkAvQQ02hUNf31Oa8+g12atqok2Q0I
JJPcYseJCiaYGpZ+yiQDNDGa7WpjhFcpUJIhqz4tdPNoblqdI6hPj0fO4e78xhTP
pkpETDabN/9NdpaiYNV1L+VqxPk9i9pXXhhPt+Cv+LGAJBzQlc7jwwUWkUgacvLm
ars1USoAIvGVx/la4o4DBHcujXXlMnb4KCp/EGQqGoGRzs2qSFruE9E+fspi6Kaz
JpfDngCKQtCzov+xui3oAsVXJqRAJZQXlcufOD155h8lu6DZkK7uGP6KYooWqZ9k
2TvPQeJ0CbAaa/yNPXvl4yVhaRewEeiUlBwnNMpKGRfmM7j9anG2fUOtuWtPKRjO
7wdhFUb8ar1OZrCLd015hCCGq+tE3g1EZJOkjsEkqxBEGIMHACQ7kF7cMZO3rhxM
E3OQXxS0W3POLUfpGhKJp4XUI/G5nz06cLaqfDruXxXSAsp9truUKUoJBIJkgp+v
SqFDrc+XjkySBYngLKOQhIwyZ9+cRizpbLCX72AoqXI1RgbMDvfOeEmTisofNFSQ
eYAfRDA+8IyFcQww5NgpuZ9sjJpugYrjCWRe34PqbXmlovDudSqAtTxQIPWJ3Eb4
0aGmlHaFe+jLF+owktyqDdDpK1Md5sz7XNS46slOIrmchG4Jpp/Lk9Luu4Agp4lR
8fmwMjubZxgMsNc9vo14L3pDNBp8LIwCE6B9J8S+LoPQC6mKTLeOY5MKQnvOQasK
mEFl8caUGdYZjwNe64N3ARrrOBpx/OFA2Qvd4ACxntjZcXbcDUP56WezFIY6JUpZ
FV93KhQG9So7uWGcy//YQR+oYjif0oMkavJpJOWvJlKjeX+puaRUCVmqJiNI6ed5
LJNO1OvCDmjnSZ4ETmSo05u7d8nV8skwSahv2QP5O1K2/OsIaryMRWYDEzPobm2D
ff4FJm+Mzyi6yjl2ue8VGRJ+PuVbNuRmU9AXWdwyOSn2V+ufsHCvLRHJPlISZbST
3E21TEz4+DysYrs0KfC1PvRgcSoy8GBeNCizWkD0zUiVOv4Mz3SYDu9Neb1+6+Ny
qaq4MSBQW07u4ObIeMtGNopLnI374WGXQGfu/lD2DFATLKUukpbZsk7EyVMuFEVD
wHO69ICTAZxcgasjgaeIe3ILpCLjE88iE6altOK9dZr9K19L+E4vG7I+w5DjVBZG
hyzATD28Z/kpAodEFR78jhAJ8udtTxaiGE3fgFqpwmcPMqSvullQ5dxGneM5IS/7
My1+yS8gk/x/DQnzr5C9shYlSkrmvjwrrk4jiMb9aLIMAEeQB/Mb3X0HP/Axq586
KE095gZeuz7GzCIl0ZhOymXVh3OGT8uz04z27jtzQe9Mwu+IMPHTDgy62aHmdkvW
p9M1v0SytDQSjTsBj7Z4la6EZXA8lICjF2Dmgt1EpOxqWPvmu7/IA3YkAV43DQg9
g5AarOKgi97txILO6Ub4nsdKOqw87tNK0YnFnu42wJuPvoekinZ4KB4Q5ZTjgUa7
lZs4atprh0vfsVEnH36TwSnf19X6TKMe9dcsxdOBIhsuLjMeAhC2Eya6FRRujHNq
O1WJotl55eVrgIixc+JxjB037HqC8a/wp7PzmwnbCc2wpWSVpowP4P6kQRcLkYiA
mfZ6BuTChDnsN48PKMR5Eb1HfvhdBL1Z/+QTaFLi9Hb7eFg37HUAOAvxuPa2oRRj
4wj7wakyFEJNon5aHLTne8t+0/SRtBdbJtU5wd3dSjmAkeQQCmZFhcEHWWitHbov
v50IAzSvvMMQyV1iXXHWonnVMNRtc2Vw7pG6xVV40YggHdzyOlESvgyXLOUuH2Q5
v+SiXugKIbg+UXa5PGHwnrziZSl/Ay5TFUoISnvcPwvivS0Nyy6hAmw6wvCyVH5A
DW/OgE7+JdTftXCz+yNhKXQK5KweYk6CoqZPFSUQz/LLRMamEO64XldOmPvzYsFH
4oyqgUoETMzyXz6bXfL4zz20q31Op6v005hFc3sFbCDhz8qlfOnlNdH/R2qlb1SX
PbiHjnoe9pHWYk06Voqo0oQTbtPsQo/9Zc+dgsTuAxyMh25GSfNdbd/2DCStHEzD
3RXlLkrEC9ldLOVMnjEfrfshiTmWHdSGC00f9dDk2UOTt5V8LNo/ZXwC59MTveev
5w17rkoVlGOebKJHj/JccVg+JhDNq2Ei/mTDG7RGy5nuFBeu9xRaM6S80FJAg3c0
nvv7JRt/xfDxObidFDaoqlfjO3qQN7KXR+TJxmfSGpWONnABNqAFkt5kaI9BVIhq
1Qrv4lRacaYCypgYigriJu2vySSksyMtlH//RRAjcKSz9brfaKtO0F7+JRhqs9RH
TYUvIckMlYE1gpLC2lhcQDL0eU7t6GY7L7VDBdHhXN91bHL38imn5fuFMhmop/dW
ecfUD+DQhw3sSPYkpf2lcPart+Th/wTGMKT8gyRZajnvAtd3V4lOjp/gLXn1q7Z1
DUOOmriepWjvzDOj82RfQHhPh5KnO1Cx/y7vP4NYOTWfT3yuLjp+vsYZ0DfybRw2
SscKLD4m8IvGyyzCZNUmkLvsVR6u31lmWk+95zbUeL+YYHOy6FeMbBbFQM5W6RLX
lBMAy5MtRufbjPlG9bs4Oz/wV+1Qfeu1ViaO8fxEqcY8kxJLv5OtIMLNiWxELYuK
rikpIoX9tpB+CmcpJ0c3RCft5NLR/74il55mbYfDnSKDnSgh8pNydSIRvlclbbj6
VJtQUQ7OR8lSzjdAVlwG+Qrswv3yBpIG/3sRuVrv3s1HXOv92XTke3lT072UWgAP
oaNQHjW6XYZjXQdTZFaHTDvlZoKzM7wn2wTAxTl2AH3dlq00UmOCBzz/QC7eyluV
rcRHdwYHnQ6dxihWdFuyGirf/lZsZ3dEpM/usEd001S0Q/OY3iNUgxMur9s3z6Gs
nWQdeSJclissEYJZlVShZbowA/5DI7tQYSB0QjjIBdInRxNE+ZbzKJ7g2VlhAz++
gY12Y547JhdMZ7KSXjZ1D8zjYFnEmcJf9cEh8n9X7XZzoE1br9dkrXe4jCbC4JMD
e5KeE7P2Jj6EWSVcw62P9XbkfJIrYScoWKuN9uXDUkrHC4s+rNvH/O2CPcEIw6zZ
TngRttJW8i/4Qx0ZDrOXOkHWBnRyXvnIlrv85AHixzw/sHQPLMHTsl7KAPcl+veJ
h396tza9Tg5cTwynh51B9aPXuRDAOrgZAYLOgON8wttkvYTvklyvKPAlUlWn8JUA
8ojSQ2TjYdhcWwNypooXG7Am8ISQYq+dtNRgxhvIhMXoq7jd2Xt2R+GkbhaWuKt+
dQO1Nj5WO106WUbZdpK05qSrG1YLD8Ftqau0FH5aj6Hnokt5kUtxdwxNLlMk/bR4
1vMvpmZCztXFo4+Xtcn45wOybu6j4ahjbjibr/4fetCfpQlsdLtVecAZCZliTuS/
kyLFV3d1asiTFS4dsj9z+rRJ1peR/b0VbajDgW4jheAcc28UW/GKzc1HD8q+EPru
WsLwZubG4uGh2fHQtWcEASdlTf0nwSwlExtiNAi7o1xcf2T4itQFH3457S2MZFbf
Y2FoKIfCBHDuUbhbuIWLZCf85YqLVj1JwPVTjG2h/+3L+6hrlvuEnXyMPBHg2h7p
//X8+4kQJEtB9pqdyulE3mm+11KWMvpfJ5y8apGI64SMK7ox84YXEA00EiRzMttf
xONmLpSkufZSdujeBH0IiBAeXCtzpeeu58DbE4iLvF201giEk0tzjub1nwXjSrPO
KdZCE29UP63ZmZ0o/bW/2EVWnDVOlvV/woRggX8Vao3Sb6DoWQ2hJh0PZ6aEVTPs
zpeLHYLhZ1asvfkAObQb+9QA38v/lmjLcaw5laPAor4vGm2VnrKgb2rNG1xIDyqk
eL206CNAjMj9HHH55KeBf7kv1DcsD4JzQNF0lpl4ED5IBt/FYTDYOA2Tdznw/mDO
5h4Bt2oHnJuaz4m2l00a8x4MGlIPEUTPwv78X0rqksWDAuLYoOYxAY74S3ze1sG/
c6XWb6Z/xH9CEvWMri9HJ/zwBMJc715ZlyYzrYZ6DkMNPOuoIRfy/B74bOEW5zF9
lkpEYv1IqtfDVUqmj+xcKFxxdtbeFDAlR1jn+u1wmUin7aucJb7HJa6DdRCDO6kE
1tlS2DMo5+nU1iQUfIF0D0sfab4laRFPkgPsBRAO9WKQnJ7DXNtZ/nnzlHvpih4X
8ykBAYkC+rhEEzdchHcTJQXekuIhVP3uY1SNhklFQh0PpVZzBeqFQVRpiyxIOJmw
fa9yKKR19mik83HA3FfjYw0fzWmlz+2lyQiVMXXZkRc1DL9IJSxlFOmK5EBSKkzF
S6mOehSHv4ZPWciBjOq3cO0bi/VB9CGBKnj8IxpN1VKUdWVYlwkr7pCAm599EtRV
y1TvdqjA3gFwVRSTO8Sp6ReYksV/yaEKBgK02hHmD3jEN9tWtu3hojKPNyoWk1dl
xuE5wgW37U/nrdiUXJZRAjTX/8BsWQ7uUXtfseXFADYO7TrTT6bI6uUpLAjzmyzq
Qj+87XrVpvCtqsbopClYhnpwoleaenVRe6pa9Qp1SmaQPtlD1bg00wPhzeunqqPQ
B+ZiA/dinr81rzvI2AESykGvctKc9gGVcH0ndOuCU2l7jfd+HjAX+bV0Jgm2v910
q0kVm7dJTJeoHckgixsrRP2H3v71qighb6GLzF/t0MZSTRSYqgD9KwcBpapU6cqf
C6g1gitgL75lhLnzC9qFKoMlGuryJpW7ySm1vKBTcc3+rv1YkcsMxYsNzd8bSdyU
7eo0rlZvJF4NVM6eEoCeTArvbi+bx9rly5JAWbRPVm/rCpbiqQW/y9N8KD2cYYVN
AsIf+osvl6M7jAS9bT2Jo0idwCN5ffiDaglYgRMvSGiovr2rEQEvkEql4KRyriav
3HI+knQoYMpZY57DQplqj6U2M84J2cmo+I4QRKvQZGRxYSVpbnoQudMX+of9iTOS
+sH9purjxBQ9DSrGAlbJ+ELOvs+ZyDPMqrh6VYp9DWvILtvV19W4Z+aKpsXllsL/
7UzYBFfe83B5Z5+pIjlAL3RKMu88DQlPp5OAkmWnBG9eOhdvpm+MVwrXCBLTkLVy
Fc4TT6h0N/HehQ4BsBSFxI2TTGiQloZuL/6xxBPcFgaMQCeFYEeeb1CabnN0MVtV
HNqXCwz5E8xhN5iZfBssCUWl3URP1NDKvCRw16p83fd3BZY8XryILEZzHb2kBHvn
7oALmEVHHej6Yqk6uQ+LUHh0Dx2iwyNPrPxQRef020gPxJvvinLQR3XwbxcyBIS5
UPDoyM2aCqo5TQFu4svWAe/Sj7LWgBFW6cchR10f92qKMO2hL5GqJTkHY/R1dFLg
a8trdH60WsYnA14WHOAEpoSfP4NI7QiBm+39KjKTwxt7dOpQnecQf65NdNDHGev+
U31FXYAeVKbFkSgQEngjV0mXFtrjEOf+kXdqm4m7i4RUlCMYH5pYW7VIiOsGvHCe
oghISKERKHsnPPycMd8xdAOIdDvrab6bt6rFZIR12c/2O6PcZOfMiDLfP5wlJH21
2zqB9VOe3pMG0zaxR8jo1eSOiSotAl0qciuSCuqRN+tSNDkZxgVtpE9paOMSJhYN
mHKt1wtF0qV73Mjj4ikQIMLpVO2eSOFhQqwcwIsaqqGuuwjt9anP0BrjAL/lrKXz
HycgWV8NfG0ENng9fhpfB9ZuWHGQNuJkfVJJdsYDow0zmXbVrQDTIgo6ttfcu1MD
mMk2QPdJp/fMnxSzBItI1Amvm8/tohHghYcR9MKbBkreXaM5VJGFkA+tQa2RGZU4
vrevwwy2KfHcWBRwWXoGW3NT4cHkd9PNTqYq3PpQEOi/gL2PF+VeRq5nm6Xv31C3
HPELSh8RYMqN1zxXg8Rri9gHz0BQA6MMs9BTAqoXUr7p8I2WJnaadZpwYeeoAzcU
EaZcQZrn90kJ0Eet686Dyx6l1ReAajzVIAho5AheJbWb3dzqouUL6Hewp9Xe2B/5
DPfLmq58EgsNQzRzlRJTxA0N69QPSTl24xULtYv6Mg9xgb7RbaPydt3NZpwM7t0s
s4VCnHr1vcZULsL/en3e7RdeXxqJ63f6Ly7rSFza8dlzYBXUqsmM4WHF7EuDIqir
R4F+o5/G/H+7iEHGXZpD1ucylgb/vHG1lIrCLnWd7CJZD2VtjVlHxgdSvOG/tYR0
MIM2g5s3keXZQ3fY6HDyL/V6X9oy1NKzRtNn6nqVXvStpwEL6SNyqKH73rRlewvG
gd/Ldk6EwdbJKdLI3MbNLxnH5jQyDEUbDkwmSpwBEFMwMoTLVoZxqqyndvsBwORa
ERxBIR5uMH9tYLTgnvgh9Lj0o059Tw0i3YIU0tcozGw2+mS8EJatCnON5D14ZNn1
BBjLGXGhNxGF8w1Gar6uNDYOuEHEn4VF7O8LyEZrk9nGUf6r9y5pwA8es3O3n7e8
8RfjlKEbTUeK+fixgd4aYyXqZyeeR5cq7flx5BcUS1eDvipd1D5wC10MBALwBhRD
6XVroFJQKJFAmuUDYy1CJv/N0DkmSHtSEeBGg+7miAuEkncEL1J1z/8Wvmmvd2QF
yfxincLifRNjslIgzpbFvlyyvDKfFReFJUBqB9l3RiY9htSH+l8jcBbBzoENcm47
nXMwa276uvzT3CDfeQKjCwavuxI4poCvte6BDm1AU3cVb6IubNsMpeoAIFPtAAJf
QZ2stWPWPGLdkQLcjSNl9o8NK6U1TtjGt9LeadSNb3qWZmENpZIEOl0+hgb9NkbV
8pgUsOEtALHc4grUKpdHp+fgayu/Gxy6zuxM0coHkpVzj0qQiSmNb1EvJCVrL9tF
TLGC4hW8x3gGAt2Kg3iSnPB3WZkDipUXztK31Koyi1Pj+cfws0qgvNsaztiaxMhX
jQPLtnurIPAIdOXN2DZScfB+gj/iI7CvdqKZofsAPthz0K4V8x81nZrOMkzKPB83
3MoYGQjYeizpvwY0JaCUpkiGbXo5ZFuUb7sRchyQ43GLjL20t2zutGqK1JofcWKK
tNK5QNLOe9GKEniBS+TPR53DgAkNsMrRPLJ4aReAomsXZfklJaxn7Vdq0BlMBiHW
7W32Fe7p8HIIU5rpl6dNLP04GH+j3Y7qYzth627liUi2oxbyqZkNdhESjBL1Tmnb
gj9DqOecVQCZLsWyb1UC2lS+ywTQyJ7FTyo2qzwIetD+wBNOptVJL0o3A120U8F1
vcO81zE2oM4WcYzbA8X0lJUTiJTvwub2jep9iCqgZhcQN6/43FEW11rhPyN8zBjB
xq20M7BVFonZze26Jx0/ruEiHYo8LrQBlK+gHZKf5eqQayPjRGDPQDKHV1EK5LzT
BrYzXFaTLYQVTcBntbnNDRIUcxo/M0VWZSsPyRpGBj6RTMwjsYVwb0bqnCUK4WmH
cWBOxOF1a/ad+YM6T1MTLrphZ49CbLh2ioYSJjZqKMFFzTtE0sCXBhl63X85EQ3f
kCDKN+Fy6XV3UidHxAyjmsnEgHOsyAm7l/Er0t5uPgw2uIc1WNXghSJGL7LSHg8+
bvevpkMxK1M59/SZYYG+nQJNYAT96hxoqmwUSPDAlD+zgU+Ne9k1QEMGW2uoWkwR
lOvVv67suV97Vq6uE+YvLAhmaSqioQBrMIwKf2+7umGQxEnpN35GGKYF2eLPPVnc
Y+WDJJZ+THULcZWDq2MxvJFh3ZODFH0zMis1FHYNt/n23hWoOTS1dJN1PgvOUB2J
2PUbhRCc5qhQpn+voF1Ds0RtydOqZcbzQDsbe3u9H+Yf4AJ53Kb1GUdTX1NBpclI
fWD37lhPCsE8J2pR2uzmvJMuU6U4yeuLchqXd8D0YzjeSrPM8hxJiDSX9y4Zv1cL
bXAFFuF2amsD744h/WYO9MstvgCjRhFFoPpJLNNTwuMvcex1ZnXgBrRVIRP5TIUk
4I/bHzpOyT1AeEKk+uNrEeoCF7sGnzYF2yJvztZQXeqk9OG35I1ukISCS1/CfldX
+fygN2B4yF0MEBYlkDyqyI+SC/HqXJIMNXrzI5WvKb8xCTfeofmM7IwW2OqwuRD+
vjIQKcElQeZ8bdX86ce1+jWZ3us6CbL2ABAG7XjlK9YPGQj0Y8eZa+bCBA1bPz9g
HGSOnJ3Rqm6uyfGGolcDOw0aW6+h5Vc5l2FmND8bmTtIgXo9jTeg9tCvsDS1ve50
cuWAlkjsgeIHlmqDYYuhDib2nxv2ujkcw6udfAGpqSydyd93NW/9rFq5xcvZqMM+
5YY+l3+y/vz+EChr/CMOy40VHhf6UEoEeVrAwWgQBeqDhvRVe2RkFfXGCsVe3ABq
/JZG3miRoAuf7G6RtnbGi5Z9V12AHIxr2DOSl3a+u8i/ysIUYfksIgoHhHapukQ6
HNcyzSk5NW0IDdrrpxvBzcPoKt5VnHN0/A+/4rRj1Zt8NU9wmr3y/2GZzh2iWiSZ
TnpOVGUHtKkiXo5gKEmEGOqYAPkF2RrJdTAd8iGxmbzCMXs9trf8My0spPJ5HshY
qcm7nqJw7PAhO+8pwzFzIUCcIlwrKzl415Y71s5pC2W/0eGESG1tAlV7YEVLT+xE
N+thrIplr4abzDocjWh3T8rZQaNLjlQVqQqtcS5COpRKN/ePAVA4UfWSd0MDboZL
IUzNX9QcE+4MDQ0Zb+lm4g44EaQnQOGeMd+1v7KGFeJsCwAwok0Zc10iGV9en2Bh
+xjsiZC1lHKM3xMmqsI+QUWMwN4ISam+KVmmkDFQ7M9ivTFPoQcnx/aR3tpOmGr9
e01oC8w3fGqEIjYnGdEGvcpPB6gnXoSD5qf9LOrSMENUFNgGss8UjO5Aa7wPxC5J
`protect end_protected