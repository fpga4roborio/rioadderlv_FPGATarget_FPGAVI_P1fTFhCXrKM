`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
ddtXksX2+yylW5zu6QL2Lhnb2d1sD00763mmSITNX595NcHTEkwn0zB1Dry37fOW
FufOhVzEJp80NC5qZ/+F0Vk7Ik02dIR0elf3clrjeJRK85K4e3Hoo4xn7YbFUIms
l/8VZSb14+JVGURjfswrIyCUotIzlzVYZ6gzoZwDXIi5gQIBf/gI+KxNXPaKV+PQ
Ufys/12rjO6aI/pPlqSm0hCvftmBcnezN2hk1UeXgOIuKZnogjOsf0iJVX2aOOWE
6pD/psybjbnsNB6kH5uFTA5frkzIzkzl5d9+YDm9OyC+k84E83I/7/j+rk4L2dah
QJOvksSIzN867/4Qt8qYTQ==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="MvBXkzurAa5VTw+1JJ70nePUfoQXBvZOku/SMmg4TwQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
oRtzZL4VJ4iwysPsC8SXYCzXS8Fw2gtZTOskLcDV+1B9Nzn1zTyNtlo6lNICRmmK
ZRVu2BmCc2G+fmzynYlNTnSa7C0Cuel6FYpxCBlOuk3OF2tzAmLAuDyOH3Z1Yjzk
a0aHuoCdIRKv7BrZCdALt03JeUmXKPdOmIlkVGFl8yw=
`protect rights_digest_method = "sha256"
`protect end_toolblock="Jn9CQpRhJt4rnzZPRk+dOpzAubz7omckX1MrFd4p81o="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 11488 )
`protect data_block
gD6l00tciPUa6pDNTk/+t0OO0nC/UTtBwLB41d4inuAUA3i/ALrNyoJVcBnAmEQW
ptbcNp5fxEUJjnOxnedyZEuEBxWRieZFQnkRdF269oO0t6rUBNO1Yf2Xd0kpTzZC
FKqce3uNDlZyDuAQ86z/zk/BG8aGOjCLS3ox9yEPkbOu56TY2/sLzJEFuAoOkkBf
tMOv32qSXXM9hJT7rSglQIOKIBbGfRgKXGpPqCjY2q1xWkuwxT1UuCPPAb97tcYE
HXLkMhiPl7dqtUozyrJzzYjtUi2m3FkB5A0i/Mdi+cQKus5f65LxUTcGRvhMv39S
krlgV0N7afdEVzt1vHPOqYKqjOz347CwWlbgp4VjnvxRvqD2QP5P2kyCPI8B9c7Y
vEZYk58hf0KU3tiD65HRyaGVG+HP4pEudVdwrvVguBH2hSe7gwasCZHKomShS7Lg
1/n/deBtp80Vun66zWAzNA979CZszG3zD1Ar0ZjhJj7uSK5lb9NkUg81UaJgJV47
k+sav/a25Zv26jv111rblCVw/mJH5tIm3Xg45VEDUWXX8sVhLzNUa/fK//c4Kbpe
VAUPkoXAF+tIXoD6wYm/aaAqqHPh2irf2MdRyDo7pTKK9CtoQpDhyH5MdVX6Bia1
CkZhEyghgnryjdfuSZqT/n/vCiIJi2ki+3VIWeOOUa3ACS/V6XkjCPppOO3ST0ET
Dft76IvLBfUgZGk0gGGJxJdQEg4OXe06qIvNsTPeuC3kCMmEORrALiWhuW5EsMKE
Kw5VjO72ZjoWBPIJx/R/7DRzHw5Efj/cNFOUZYCCQfZaGCKayrin31azW3Ac7VTh
YmcWZHJe+PyMtDJANBzAz/z7LMLfCs4DC26ALqHpVAw8WlRONBk+yEhs76O6l4l2
0RvOCSGPq5sm+/1rx9pwd2XHXZZs7FMWnMn9kIpwxucWS59jKoQQVVZ/rPXGGkV/
b4BcH7ms2743obRpe4ytXw5vR9TyZKHPZNeDUthbVVXgF6KM9NvEMEVkMdlqDchK
jRD6eX5fJx5Z8ptQsWk/DhpmciyEmDTeAdjkp4t7/qMfBr7wQubBDmL4ZL0Zsyen
RMJeeruiNpb6R6e7ras5yH4pCdmr9jG07OsmBzLvXc/BQIGOQyBz4DZ2gHunisQb
tqdh5MU/kADuC/QlPDbOS+e17+6F2rd5C2Frzk8X+3Ib3aaFTz1Nnpi6anaXPtvU
8N8Ag84QMsNSym2bj1CUhx3eIBngW+ADWeXIAAo9ODOOajLhi+EJ8/BNmSDzied/
ORdyx6IC4CchZ8FqHOAuWE76+4aDcIBxKUG3kx7NxtDHwT2PlI8e80MpOZbL8bAr
J5V69DNU0knJwMJ3cc5RhNn3bLylEgjFbj7R4TxKuareKdZ8GQgbxwOpqvgmZ1vb
/VqrXM2OvssuaK20WydHGTz1bD+GWv0YlP1vWWR5pIObKCQLLMrkA/HXDmhPniFj
F0KYW/bBxgWFx6WMJAiLlvcOYlbRMeHjsQXpjrH6GNXgg6yZ8k4KHHSUINNDAmbe
0QNjfHN2pLOqpwmjaOdWpVtxuuM9VXSZY8mJzkizUP29VlkgJtSs6GVe+hHXE2lf
NT/ul2kixor2Me3/8jEaDetCyueyGCFB80RZybNj+8CRaw610D9uj7peaFt126y0
DvFvCtS3Cl4Znzy/fy1sZXcMPe6g5xHpTDcXtkHe1NuhZM8Ag6vRf3Rwo4KCy8rL
hms+LpYqN3hnQK4EEtqTzP6e5W9GrMI0E3wM6AxmnArOflFuC10yMdzulbdLKN5e
s305+WOHbak1WdjixtLySLgb9FBfW2SZHtYBfLdiexbkeIpaU3yY0lZYCm2x2KSM
lRJ1MuNzzHfKA4AWTWS7NGrGICPgmaSX9nPOOZuezYgzRycNTnoJ23+OHSh60c/M
8HyuvemEi9gE+lJp3S4oa/L+4zE6NJXhlypAt8t5Z8vJGzZ54ELThi2RhSEv8ioi
E0BnaohqDrJVJuJbnojROBWg31p7Q7SHJaRsK0F5KxbIhg4QhZXzhKrOpy7FkoDj
8xNJVja9vfwdYVSDWG0N4YQrRF3vmBGiQtLX9s7aO6cZF5BIYDo9k2fhzEELyZ7P
M0JbaSZgJYSBCEz3FZkNVb1tQ4B32v8ajBhRpbhV7QXW3ieG3GqdMltoZN3ROPwU
7drL42hqn9gRoPR8DPAt2S62gJBKjT/UJV4Re/BO8U9fACBz7v1+7j68Td+NtL+A
EKKgHWTPUu/MVsna3rz+MEOziJJh06davAB6XftMwQYp9/MN0st7LUTNbvJrs6ff
jFIWd57ok5QAq2HeUHl/NejAqEUBjy/GfEro47h2GJsSghiU7f2ZdDScItpkaaMD
wZOWDm8Sj7uuWNp/WPdoj0tGhigEt9fAADljTzuKWa+LtOxslxpJHOswpUrvYHcz
AgEZYwzTnd4IWg/vDiDU4L7cHQ7BAMrEty80eBUBA0NQD0aJQSrLwmDuLEJIPms2
qn0edDhrcI20q+GPL/ZSlgYw0n40s+CEHbO6v9BwPNZdmoPpPXgP5lsyO/ER3g+p
KROTIM4E5UiGmRFqauemlzmg1atq0BttWbyZ957iMB5yLX3bePrGFtPnZOJ5iA76
+RiH4AUCyDQZRWwAEf5kON8YcOfBmjlaSZd8xW3+ygY1FRO6jn4hrGKSZy6BudIx
plvyR3DFn3pfKSGXH5uqbcyRfCbhIe8YpFlep7vWRXEvZ0K9/hUc01fiQMmBGhlK
CtlmKT2Ig3XwJAYRrhGSF9s3qMXS+vX30ETnoqVC6gW49tag69PaynoKRkzpBlYq
rK1zmkw5OnQ0tkC6yWbihF4IT+PytNAR6y8I4aITUsvdKVDuM18HuJEzAII0nk5u
lOwWfaAMe0Hl5EJF8MjmFMYcM/imlJnShzq+xNggUWWzkPGJgxLK1Y67ZV0s3tU7
7l2t3bJJKouxHRswb7snQ7A+KKMq9RVcXlEXzteWIK7uRmh68NGXLbOCEYq+Ve3i
NrGet/J1S5lL8PIWky4WqB/EzB7204zpHKV+Dxj2d/AD7P2e5zBfDLibQoK6W0ig
NgIGLEpRko7M0f9ocBwP0iYRLZJJk+8K9Sd6kPu18EG/xwPWZJFTlCh4d6XEex/F
X4vZM1cCs0nhExHLhkgpAogNEULSrV3VT0XbWTr5rM+nJb6AQGtP9EbkDydHfqDB
VJMkWShTG9NTJfAMchauzvBJQw353l/u85Pv4+8nZqtYCNy3QLCMGlKDPvMXQk5x
qkMPLhideFIUUEDoLTMPnozOC02msjI/u9ideAtVdrL0q85pFUXonE/IE/r+OF/b
uMbrJlybmvKWExVOXeL1eIC9rg8lynRtKLtsUMH03hEKOEiP8xIyeDNGNi2ewmvs
nSw96hWx1fHskIrNLGWW5eYsNYYWbNiXKSRgmsPHiFrarkz0OGAeCcKgiUByJmA4
1ZQN4pqjW7iHvzSfpk5e5vlZpHsHVIJICPNWVou6hxxaxctKTzaaFErK/8xf5lgP
X6X+uqDI4WKoeBb9eHGxKlzRiCFm1xQ5CYjrnjVd5DP2J7GXso1IH4vTHVznqsZX
FTpCop7EXOyoXDEZN4eSUtyei6ypi22aW5oRqkEsMzTJPLxVoNbHVhXzscRhrNL1
nObt/x1s4Br9SC9d3sWzgTShYTUw90QJToA0mZ/jiYEvJkfeED5gRebnLdcvU7Os
0y3Ur2WvDLC5RVHvg50NO4cLphouBi7DvIoaPIa9XV2uM2jrvdsMVbvTBQnkD1fC
3oBuXESJxCcm2tcL9vcEFqrwz0SLbW92u96r2KMLApF9OKzd0HeVyieIhvCGngme
5SgRxQzfePxOS5AdmjJIM4/1jQE610zstqZQzsa3Jg+eTcI1ds/0D7ksTv/IGTTm
dZVX5Zl72k+thvua+RLKJCwWSt0aKHm9+2MwIgHHKOjUThZ3eaunXsGvRs/kVJnk
BgcWsOIf1hB6d32GVhhBMpBV6sQIJFvAWe0O8aQ8xIi8wF93v1kFP0u5PYDL1zCr
iudetJ9hiypJXanRjYffJzKbDEqWY26UcPlqnWTMqLkSiZ8pGYk5F5nDIP1yN7QP
bHWtfPzloWJkccm8UzMuSuvV1TUbLClPjHa5xZgq/2LL/iJw0mvIYyRyi471l3WL
w/8f4t++jGaUuQfvL5nVvTkoLtsyELwKcFwDhyC0FUZF34DY54jQtWAied+a0Vko
kI5SRcOv8vNrNjMtlJO71MS2Enatms/TIqUaYS6iPzq0+MQEJr5ixVkLdd9GU6KM
Zsd91reNK5AJitVFVYEWie0Z20csoHEAJ3leCzGQnTeFYdECRXbley+YF4F38ETm
1ftifr07PUvMm2NN5WUnPdm8ad7E4h03VlrwrjSEoUWE3XMMGdfD3SQH8dt4NSky
LV4UWKkfhrmc3m3LPuy0v3cO8sWbKNeAH+wwTeKQBNIMouzpJ96dJ1/2buCau0Al
REu7tQyXi5lu18LopltBtfbLBaAzhK5sgBEtLjb1xSZnNv8DD4Deg7pQ/I9aTowx
9Aj29qEai0dfDbEV81X9noSp4OQRTXd0ZNxOWQafEcei2RWWda3cDbZseP17oCIB
3iQ/HLWw+oJ3H5020VBUyb+bmEBY4bkMVA+6GFUVgXwUiUaqMx3A3VR/UBE7yS5l
DI9Kh8xBDCUW2c26zEAoCPrWHQjkLbq0CZ9fb+YecscUjBqalhZqdUHNe1vO3SUu
q8Cy3ij6BtnbvAcYzEA1MzPdCgG3OVMbKfiOMiVoaOFoH4hXSbJyfv298ZPr7Pq/
f+yGJDLNC/G5HhkOJgsqhrDMWWWJA4ExC20EN7LC8prsuBEPIvRr29a2kcQQGUn9
84c0wDCwk2NmjPveeb6hzGmuqm03hpKqLIZL2vXroLKgKOKO57WJ4HKImmegVp9m
cB3bVtumuosbqnwNQmIMpSjiAgB905C5Ya5BYw6CXApg5jm24Pnq5u222mDz3KOb
gl2DBHKKbMzoZnjUdnF4gRlpoifrawGe/s/Y0Cb61nva9Gj6ezssjySlUCT3fxha
tfgztRknv6JE1V5SxMUUrymefxpuks3Y08jm/Kpd96u5n+7XTs+BrdyLEAKphUho
jB8WzytBd+wKgJeyLeITeLwAzPY09lYt8Cyi2tQq8cAK+a1S6heG+BI1QzK6hL2/
MY/TdIhlODL0obJdRVHxx/+YTeCHGcH/jmR5hqP5jhs7zV8ydf/IDnNxlhgAYyFT
B4FayiZshieHBWr9VpnopNNV0OPH9bnRNx7i7CQ7QmzLzvHfuxaaqfhQSaLZRtn5
Bf9s0z3/SqwdtoItxcMu/1nBhhxr89T1qkzS+TfA6Zlxy+4eHjM1KqhLBP8TS9XL
ToYf8Zdn4yAUAw9eV8oebkcvbuJVwz+aWzpOE3krGY82ppsQgaoEbh/K/fBvkxhg
gdvEWUx4JDJoRYgnFZLVzSRl36zrOlLmUtwfYjcJB/vKVZgL4KKbKLnq76KN+0R3
maWAdcSQTxOdIRgKOra8MyASzI7x7LDUuYb2KlX/U7McBIzsoTwD1tVeY+EXEn5N
FoB21A6/vxWqR8I+WD3uTtn1y2h/vN5Z7x7igbsBQn59IBhEdj6UkE9EuGmovEBR
m6vYqxseKW96PLPTTAscFjxzCBltixwY6Er48klZ6z/L8Br6Q66n+MPUPI5r2kG1
zJ7dAUuUEsA1E0Z9SLDCTzan8Jey3ukTw1NOByF+4XwZKSW9MZRPJKfCskeHv+Ae
zBLXI3JNlpfL+VB4GxJF4BNvY8F1Ap31qvk9d8uWwhO/TCzRW5//6Isft7+jdJN4
N92Ncmj1MigCNfJI3xCnrsohEY8WYenT18/ir+Z2iCt5lDEdH7DLB7N68eKfWRbp
mngIjXsRa41z2eQ0wQJZWfJB2Zu9jL1VzuYV9h4DmXwbGxN+ttJ1eYviFTEqdVJi
KykB2CGMK7xAeevPv4TwzlgfS9llVi4dArxVPup2Y6NaMcQWLFVchOOyxXRHixvw
L8V7eJUsxiVCZJ9QPlqxmL9/uFK9A81ozquGgFGavdkq137531i/1rhXGVQS+TPb
IvtcOF8hEfk4zR+I+dq5uvxTo7QRfv8E8WOkvEU6K+IiwTdZFiUBUEInQQg0p3YI
7wRugJZEpHWJr+RH0WRMY4227VG8nQHxduF/EjGTHOHoJYb2p2Hr4vrlsOpPdTG+
lCZQs1ve1YK1N+AdOUWVK6BY2YzNNZEZEH3Yh15RARnldQrNNah38k9UNlDyD+37
crNwVZDg0Nhm0WcUTNm8v6G4Z/mm21SNepRvZMAyy3blVrkefufzTS2o3XzahwBb
AY7wfp97DJJ9jEB1ikxaROyebfVgVNuT/1t8TQvGWlx5ewSs56TP+yX0u5VdMiw0
vNiMGhpltTbuDTf7iGYDPYsrsSK5thyl3GNKzLssz1RB/IkEOKYkOJSGqIh5HkCe
QeH//u2DU1y9E2F6exnwpHDTTmxHban98jku6/t0Or1SeWckI5iWkTCAyFVOLHLs
oGn0WYfdv3vmzDUjGk7KpLUDGmhkU5JpEIOZCVQ3jl//XlHcUaD+j4cnDv0fsXD4
4HDtq9HBhUO7XOXRvwp5HKhuJJ7/yywrBOX+s9SNyQe4TkHem8ZygCVfQyl5St2X
se4Ska4sYwUFY38UQgBpkGZhKp3KPC7jxMkLILpLiWJe8y42bmFLKJQ9H1NJIXWL
sUQRr1/qnVEJiPTocHcOoklIg/hn1PNB1bKusp02yXyyzoQ7tCAhzqIBjmnz5RRu
EdFPJTzfQRrJN2thydynBPOzCr21sW8PScnQocQhEHbs7YHqJOWGyTND504a5IkJ
q3KFQTz5gi7xwerhgDbCXJb84005+Jcb0hhY6dt6uwayyDJlMASgKVUmJLU5Qgf7
KXmiQvwD4wOjnoR9L4WdDxBes1QsxIgrHeq6EUp6cMCuhgdTEMO3VBD2R64tiKm3
Pt5gWEcnjTmhZXB+6g0hoy1rdm+yx7YHN8QFbTMCP4NXwKQG1nOk2MebIDAck+at
R9ln4C261F8cPBKyfUSI1rVtaHp9bcJPpCpeFE/cjz0Gry8b4LB9foKk6VoFlXA1
WC/gUhtcwPF7/oi+PmTNx/IjKJQuK5+m0W5Vs267t5G5YYSMvRLb93ccbapUUYLr
eDlWPoBoSlsnIkvN+xPx1BlZZnKklyhOSZmcptzTzRIPfpsFTJg8gP0rDmUzr43/
hk6MtQPpviujIgM/I6+zxc3UKEnexhbf4+T1dFgAakcU3El/GV6lokalHYZVVip/
Vaqa+UWErTDVJ2N8ltUDJI8xK2/1DMCgybUwCzmQoePF/34UGAUSMPTWZ3NiyrP/
2tgJDIucVByjzG0ZP1/JKOpt8xEOzVMNpP1pzRDrBCSqovvjOHmoTRmawbzyAKHO
3CAFp+FCsbp/CBaiBH6T/jk6uyWZlRCmT61PrWSBxDxFpMAlFGyDV4HIuCVmF57O
HmBkMriRNVV69Xnq6V8Zkgh8jl1hOfS9Zcm8lvZIg6fYxHjbd5Kzqy5B8j8P9SQR
bGplNAPP8qk5EkY1yL5gT2tSQ/jo4/XSjOqBUqYwRc0W0aW/xbRcUzW/AHoXZCd9
YT0vQGu7TrKZX9qnsO+eBUPUhDETqJbblSck5IIAYpMUlLrrTyhbQkW4aM+dtUNK
aQPKXoNBOBLr+b8v7Z2tu8QdQAtUsnTV3+79p3p9MQpKDX9boW6J4mom4eg2LkNs
9qvJPJpSTZiy925X3DGgFUC8VoWstrrJrDLTCA4B/cvAy0Pjf3H9NY8K9c/YAsJ8
YIZQ6UF/FsfcYp4j0vqzzAB95WHo0xs3Jq52m/Q+u5FXtnPg9f85MiQnULr2fdgD
s1okjuDdGqfHvW1sUPdjOuAlSQyJmJq1BCPJSPtAdLfZFs9eK48g2FpnseofGrZA
aFOcxVWx8Yw/M3RnEHaQHRnqNZlzN4+9Upx0GlR0VGDx1G0QfkEELVvsIWUC+f/h
I5PCrM9VyZ+NamaSWVArEL7Pg+RGRwDeV2KEsxgTTnZweHknaGRGDIKYxgA+FMBZ
wfuWlAVwuLlDO2/Rv9STEUkDXOe4nEjPDt38ynzJN+O4YpSaG4akqdNMXnTdfPbq
rqKfPjBOh60ANfhQEmhyuvvgm5WmmVDlJoB+Xx91hDOKsnuejEyC7YXDWXfWBlV0
kOG342us25b1CD04V2jo6rzHfwN2a9eaZiAZEx7WT7AwOZZFCyIncGnwvieNPg/z
UYm1fOPv0AahTsJpOPaqUUvyBNuTVS6cJMNO+JclIfZF3dNHRILqaEzqi2DKqyQt
frDNp5si7/ev3rDfESo/M+EhNpGk2I0WyYVjCkVtQPNsB7sV0Z/tB+HYPNgD7GkO
LpDHzKDyjjxHCYHzFwiEeSCoWPhfNUWcJNgDQ7cjBsr9rsYKYobLN+Iuypq5roMV
XyeazxG7jtpnM3EmP8aCMw8dWB8l/U0PI1ny6XBHXKcQdk433zRTYCD/O87IChrG
IeKCOAUUJ5+mg/JlgYZQe3+ezCFq7kH1kkvcWTpz21R9sojND8DJ67zV5K0oWsfX
fsYRnJbTula2c1s18gLCpXINN25+FjQVY2/xln1KkMTzfyhWflhO3sgAc79Pcjc0
K0aSuZMl4Eoe4IcWZsu7VN27KzfOpZO9YQwXfx9GuVslF+DOrvt4I7tqghcIh6Jl
qYPm9K1kEfTVAWKcFnEnWAPUlJEOJ4rzmhVEGb+RM6YNCerKnvG7bjeOTmrX5CGE
2M/Si+7ZJcSgurZtf5Sv3/CsNCUziHxnnP79t4gI2RSelGSIuyluJoQShkNRM+on
O7z9JV/zSZh52Lb3/5ieonX0kqutkpX/9epDvOub9+xFQkjDsa5H3GBcj22J69Ku
PXox+FsMGX1Hdn1SEScXb7w483I2EjhwZknzKKiIIsSbEPr4f1cNoWkvibXl/ICb
ig7Z9PNEb0tXYVDzTyjbjQXCmo25zUERUd88HGIJkoiIMQnjdL+O8JCpngkOI7o5
KN5dQBV+KG7QRY0afwAfV1GVopsziCBaeU4XVt56LJ4UkYaZm77cAaIltRn+rb8i
OfnLActd1IvC2ioBjWoswjNcP9E3OeLMXeL6JYjyU0OnnUw9Wcq6MkdMBo6fzRUl
YkOlJO6XFxrg29O/QDDDiTMFz4Wz5rjrW79HiPqAGit+GUwxdvjtKC2JH4F/zHgI
5/PWU6z928TlncNfGCXDokSLCAML0CuBmN2dOwRF3Sfj4YqoowQ81Y2OVgcpftXT
AoEZ8zM98EHsb8t7sa+5EVPeyNgRGY5HnqSvNaNm+70pRBBAyyMeXsb533n3B5ow
0CY9rKcNGDr7hmTb9UbHWLWEYN228UExHDWCiPW2fiz63mieHZlNZJqd6m1+3CtW
nROA/U5H3tGuvoyWDocVedWhBH628Fwl2coWnpsiu0phCQ644DQUrU153Otv9+g6
Zt841M1KbyAEV+zUnnf9fMU1PA9zVfM6a06HgQeXezC4xwV/440SF4GoEkWVPWSR
bQFSirXASwVgo8ZC2e/0K9jAIiNjyQ+34VvpaMVlgqWAS3W2Zfn4GHcBSiRmEous
sEk/2cq05fz1stHgdHcuhPBRSeHqX6p/H0P9LHeLb7+c2lcDYdDdN9+t9Wt5u6z1
KEZ86DVNanu78knRK5sXBItS/rOKcO0hJtMMfBnVtxznOHxjseW4Zek5linTVQOG
JAyAQFVs+gRJ7vsqUA7OTlne8YnNOW9C+d3Wj9kdVUY0iikCHvBOu4Rj/O8Y6/ef
H5qZInSj6lPCr50T9txw0OUzo6LfpXhxgZtSOmXh8t7EsKf/aM2jYCoZpIeOykvx
g4HMzfgdnaZptvdyDhxxDYcup1voqbCXRn91rJ6bq/RF0grco6+g7m5orEqi1Jkn
sYaVvZUgZ836juLfZsWafcMPUQ6H852GBe7+bWfFeHFRqdhD2HgMcwnpFt+LUhL/
NCNTVAJMVunE2AqD2tuCUMAJaReu1QFQEcla2s6NroeZ/ydpC+tQP0wp4YiF07n2
61fdsrTZm5MHmQQSo1dAeuvZNFChaQbZdCYRjj/I/UvHsuOs596GpuHR2XywtvDt
5SwU4KkPnjLipLfBO1kTJ7msD7GdS7wSnK9u25f9Szl+oyDFRkrjPSt2zJxzavFS
RnAHUFzecjC6C5CXLyVTCMO4UwvrqNaI2J5srfQUTd6SnaZowldV479vTT2MC8ZP
5b5Rg3iTK98BJm7EVszWkJCNia2wScfyXKi9wq8wQvf2tIk0r0m3LmqgaWY/gHxV
9XixsCsnfzZTkBqT2hVMahBcuCDWiHVlKaOXR1aq5/feuHLiFvgJ58p1MsTuia/X
tab3ylusp2mQoajSC29JX0L36MZDKAmzvb2bGY7+u+oxV570/nOhYRdXNgqUi8gF
sAkk0r6aZfHyQk7BVFD4EJdMtUzKWB5FPshfQIjtoldnTXmjGv51kMYaBu1TBwIH
VbzrhOO0cjjmxEIR6kf1Q70OkNDeC2SEKEKQ4+19BtzLcp6MxQqxYeFCug4APPpL
OzrCsmoNM2k/uyDFDGyGBgbJ+WhQ/LDLSd/BBZvGeqzrBqnKv0u6VR2Bji4d7wJX
pj6SqTyLpce3JQ36wkVxvgj/B0Yg9ZoPKjGiOo8zTagNoHPbsNJ+nIZmTgOHmhvt
yruawXPmuOIX7qcXSxd9CnDsk2RWWsJH7ZZySBpgiDXjwA21dA899AwYXGeGFZ0i
2hr/Y5mie+qBRnAl78116y6Sv3t155WZzSvvmS2UQqznMzVnyGhptsQTRodwSgA7
n2ZSAI+GKaTCVyQE+fyPVy3Zp38N8mrRaVwX2oyPczG1QhiWxvaK2oNB+XO5Cry4
GB5EbTQ8EAlZEdc27FC3wiH+yAiUeZ/7xDBXmfzaPxZbe1zVicD5CwBhzuzZImdv
yZGAezahdWrHWQHK3VfQz0kO3xnyuyGBgHf9AVkE1VJA5IU1z20oI4XZlkTN0zF4
v81OrhJ0+kFPiaaUuKhEkxueTdyFOXRssTLruLJSfUhPzHgd+r+N87DqA3VeoUIS
5idfZDy0ngWE7ncmrfv5LkD8HyVh1wxBHZQUnYH+8tLYyDc96iuap/SzZ39kvPlc
5BJytKvWceRmeiCuhy21dhRK1SSICUlUuDUm8egub07WmJOutSgQZW82mH5PA5Sx
69V0M5gH9yyTeue9+qcPugEnFM1rBjHD3wtBeo4MGstJLUzg2ari/XQzpvrs1RG0
crbHN4ooeNipJsww3SG1WbPXEYZXaS2aEziD5mU5y7ckLlsv/H3C9aOUKfviOct8
2asQ/lJI8zvxEIS45xLtXDOO/iO3YMLgrsKGcSuumjnfrJJAUR2qaavB/6tTNNto
p2sx5QLopoKmLIS66og8sRTZNjHt6hTmrL2YLh65nWUpuvMHd+482gNNdvsvSPpL
Y/pB5bS3y3WbESGJN1mgB1qy3mv/7cZYVZRflopnqcPD37GII5NYH+hHFnPEV/fP
FHcL513uPbEp1/rUWv0QLIahgXirAc+hPXQHcx0TM3LLkTulaaIhA03o7een3QXe
+l+jzB2zgVaPQD0U+svGztaeKnh55zaCVqVqfgG/TncYmt2HtxgaKmLiGlGMSLig
SUkech+8b52aKCgK+lxgcPcJJ6JMpMSrOaCuI8c5UUrhuAPTqTG5Vqj1JaxRrxMF
W08Xz/KTaWFYxlbPnXNZVEOszXUtH3KHzXmIk/TKptY34Y88RvMAlpjCI9/kHW+w
D4DoX9CPE4ZgT1PLjLYYDP9WlNMfCOEPoZpu5xLEgXxQ0a598INc6E/J/P/JuYM1
AwnSEsf8pgzwQDxYHRTZXyAxxdA6s1WwxGyH3q3in0RJqtQQeoEUMM8exP94FcoF
JQWY//A3DYpdoS05/tjiesAjdjr4eN1ycKHvjJkc7BUrQdCcLuS4U1HS8tA6DuJt
9HppB2XTWQKyXdoQocS8bPOFcpI8oRY4zYD5BuRqJDH+9WYegcLyIEa2noZyPnI2
4JaSOeOWywpudfs83UIpnrFSv34H2DXVtG12SNu1rfOzMIT19dg3HTPWPmIZg7Ny
IZhkvew/lRcFMI5gkflZtDlTfaGYDIXFyTWu8H7ycLauYrWvnimgMhc4Z1CtK27A
DsyYfF9X8skWPFFWjW+JqvmSYb+qdePL59iFp/cSXqxtOwWnVdzD5TL3gfQIOG1f
y2x3lW7zpG2CoDjaxuBtojqf7LKWRTKFM0xv2p9xSUikrkFAUlPsQDVeDx8bPGUv
f9frMhs4XYOiB37QyJH7bbBaDFPZ1z1uY6QTEV9JcVBwobWF4Fh1517WWv13xH9v
9H/KMKQE6IC19Pjvlz3VrKkkGHFUw8m2tcvLcdUePoNXtODiK/AEGhZQiAnY677h
IFRnNFiWKHu4u0QZRk/G5tnWXn85/nfycBwrXQgmby6PH0Dj7OjkJjoVJ5iBM5IP
6YAqBpVzaJ7B9uKHockQf/XySSek4EP8tay3MLHMzH2Rl2tS8nlrv2lOnpfomGeX
nMz8oGPYHd9U5s+oy6jZ2qx8tvcsRxL4cCDsM4bkHWf6TjpsgM4OTq6DvE+rtXcj
j6Ssn8bJzMAqDizgc0QyKSI5UGHpYH4H8x8hkbh3rS94UzQaGe/U6eyPT3IYzPhF
VDtDHP7oegLtAc/OmFAf5F13M8cXLCoLpDbnTAUlzxCbySqcVfJnS/yQbCbVLv9x
GPRLc8xl+1QJT5rGhmkfAOzGm4iYhx7wq8ug8qHjzrnSocJzT1tdC2Fq7FiBAlQg
fEbrjIfdUSegvW05PaVmq/nRiizwKJfYdJBsISDsL9hIjk5JR43ggnYpzu6LVBPc
O0xu35sOKXGfxqUw48NE2LuofkRnVDrHQJWLKMqlHUN0LG0Hoq90JAr6sLPyX8Mg
iazak1bP7Tg3CtW/7Qppjij8aP8zU0yA4KII/YSbb3GFGTX9nBjMn4oCYiBQQmqY
OW+z+FgOBpxaymg8dB4xOvD/cDRWREatIFfYckNlQwpYeKFNaK/cnNpquW5EENTY
EiwATQcaT/Wm8ZmjdtnEjlrSQ8LCWHW6GSKwMApsZnILDZ0knnTOVRvFPzEMjcmF
3mDbRGI7pwz2zY8xVI4V30uQFjd2rbEQP7ysHCXMREvVHv2KtfgCQ2j+cDge3nZl
DWabmycyG4MMASramndWk+FgLDZjH4hciaTute5gRyyE3QcQo6n/Tf1LyawKOMQb
Sa2vW3d//rGeedS3Ba2mwIpbhUgRtY6mkcuS+h7jemf9WUbta0BB4uNXe3E5dcP1
JmeF548gZvPHLYqIDka82Z2BsDnz5JItn16T/dnmV3HM97zs/pJhhQaPGE+IVJU9
nUkU5QqUnVfXNuLEXnS1V+OvMyKqM2qD9AixLalibGrEZ71Wrs11xlEP1YRhLWHW
VeWUh/37MBxwAORv90OLKjc4Qp8SwQBzU+kok0Av9rFjZTUxCrDQsLBAYJ9BM0On
YIQsGdlDNImrW/1nlV4uQc72ms9Zm7frOLLvJpE2BQAlhdI/c+fWP54j76LvL0/v
xR+iQ03pIHvO2tj/EzjBoW6ARr9n2Vncr2N87ZFlLQRiZ3+j81rdmV5qqUBjhIAM
CoLdIoxywSzoHY/Znvw0OguYMnq4LqTwjtue94asKZEDFvcmnoClCUPi6twASCe8
nV5/mJt85V/SjedbR4QVtr+SIg91T7L6xbltIJWMZJWUXz+pQKADckjDY3VQGeuM
hWt7v53Fvfi49OSTZ3+8MXFiRdBNiRqObRqVbkW63SSqSb+UeziZimJwhzRDFZtd
AbkLyr7RXLRvvdPVe1zh91rUQXjV7FTUstDzX67ypTHoSqKY9mwz9zhlp1qg4+Hc
LHgUzItdnbTAiQsODCWVrXjvA+GHyWGZFIeymHQbzWGfWHuygSpdHjtEfpAz1wsq
ZkCfVbEYXFACQe+BnRQpju73nKTyKcqtsZKeeT/Uh3ih2Cs5sGiPEEuu8iqNyicP
HHm1k8q33AroqjPzfKhHqwJWAGRCK7PNLl1BGvS+CO0zAOD7ulZ3CxfRxx4oP/8L
wjq0MLhji5J3kgH9xFD4tywgPxWw7WhbTjjP5nW5Oi8HvYojZYuG5ccRg2AqO9/L
6Sa9WNBkuA11loMeVye+DLIJVCcndW2dfGWYqileljdQBtJzcCT6rwgtTeucFtnl
4+cRFCt6gHmwLiv+J9OgxKMj647Dz+OXJJ3+fn6VgPq/vGiHsasEO+qAyuoc3BrR
u9yj9TyOvpV5zl1wnPjq9ZOziByHU9dS+j6v8aWwQHkL2SIM13AQev5Klku9wHlW
eAuArzsyMsTWn1Zj34eIoibBRuqDJ3lIuoy+qyqRURTA/FQNVnWEVJGxmmHNnmNp
BmlbPPamtai/1FHnl7PAagfFsU9ERJ4XRuP7+KmoKu+aYenr2hz1AEF0yptTqBHO
0SpsL7BM3m2FunlMwqVkn1FvMhipnGkegKzXdTe1EFNVRebL2s1dEudYNAtwXQbC
gK94tNgmsdO1reVYcrhX+rjg8hOMIkkMYbhd3AJpSB+44N5Klhr4TBHKts7b5kgy
YImxb6E6udP57cC3j05aPZVtweUGhO4rnaabnuEq05Pd/4GOOCAJn+dKKWAoApaW
YpgPUGDbZxEjssN6iJ5km4YtmuceHxTr1wf+HQHulOBN62z4Uxi5/djIm2M8IUnR
fpezdQnU7ju2PYbWzr80nW9Zm+ToDwB9UrJ7NH7HLocZgK2n7VXgpBfSVx4cafnr
pOaa/cShZ05xCyTN+H3X4UwcDTjHnqipqp8e2Yew3p1+pP0Y7JoREoM+xsNcGEIq
AfbUCmATvhM1pi+FPXdZ20QtMGsDeBBm+NxN8X58me9mVzWAYXl10h+gadNp2oqM
P1H9RPfQQ7nU9jDtK0EvHgb8o8WhTQhM+Vrwe2JrdLx/t0j1Ds7HImjxHvW0Rdb2
1zgYA+WB/gM8vuTIYyKaRtpsn1zbxgrSw6thfL4IFlNrz6MqfyvyCj7fYk1OLbU/
7sA/n9MEt7x/zrYrWAT4XUjwMfiL1vD6LFka/Py2ZmFqvlWtr4uTBQHuhhxzBSEl
Ph9fB82oDJjm5URgDxgJVBBfao2VD5pnRtPIIdroDi+ecHy75LytSLQk1HyMOqe3
VYeXOE7tHsTVxkMueeSP87EXbpQYb68TeP01Tvs76rb9YvyHMeAnsS+GR6wDxyTU
ZGIjujXlc+jhb85sv8jOLgqK311WUYoF95fWxX7eQ19K57cEjetUcSvxb3dkD5Ok
sRaP/Ej0BLjJaosCvXWOHA==
`protect end_protected