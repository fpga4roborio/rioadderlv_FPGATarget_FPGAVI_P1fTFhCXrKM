`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
ddtXksX2+yylW5zu6QL2Lhnb2d1sD00763mmSITNX595NcHTEkwn0zB1Dry37fOW
FufOhVzEJp80NC5qZ/+F0Vk7Ik02dIR0elf3clrjeJRK85K4e3Hoo4xn7YbFUIms
l/8VZSb14+JVGURjfswrIyCUotIzlzVYZ6gzoZwDXIi5gQIBf/gI+KxNXPaKV+PQ
Ufys/12rjO6aI/pPlqSm0hCvftmBcnezN2hk1UeXgOIuKZnogjOsf0iJVX2aOOWE
6pD/psybjbnsNB6kH5uFTA5frkzIzkzl5d9+YDm9OyC+k84E83I/7/j+rk4L2dah
QJOvksSIzN867/4Qt8qYTQ==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="MvBXkzurAa5VTw+1JJ70nePUfoQXBvZOku/SMmg4TwQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
oRtzZL4VJ4iwysPsC8SXYCzXS8Fw2gtZTOskLcDV+1B9Nzn1zTyNtlo6lNICRmmK
ZRVu2BmCc2G+fmzynYlNTnSa7C0Cuel6FYpxCBlOuk3OF2tzAmLAuDyOH3Z1Yjzk
a0aHuoCdIRKv7BrZCdALt03JeUmXKPdOmIlkVGFl8yw=
`protect rights_digest_method = "sha256"
`protect end_toolblock="Jn9CQpRhJt4rnzZPRk+dOpzAubz7omckX1MrFd4p81o="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 28192 )
`protect data_block
gD6l00tciPUa6pDNTk/+t0OO0nC/UTtBwLB41d4inuAUA3i/ALrNyoJVcBnAmEQW
ptbcNp5fxEUJjnOxnedyZEuEBxWRieZFQnkRdF269oOgd6KaoikeSr/8sD01eXAy
Qh4F+KzlhqBTBcPH5AyfEcKJY4UW3YB0haagQ/WCv4wSSADw14nFxKu3DLezUurb
WogzjBdd/0QfBs9Z6C6aJ1TUJeup74hCCsvdTxem7+UqEWMKT4v2MPTDvkThyyYP
RKEL57uH9Y8Xy9dDtil5jlAUoLyZbjlaN+s/mVguhw67t9vMDGdmzARy1pDX3Z0K
w8EL9qwNYP0NWWC/Tbb9f5mQEtSV2jVVn/ewoyusHQzWgl5QHgpo1J21ILdywKc+
+hmW3lCJvgga1ZIM7tSSdxzh1U64ka7Cm7D//TO5SOkwY6uYVTUwVsHGhsTOsMUt
S8OKeh0699ClLDL3JRYu0DxulphIs4K3WS6sGJ6ZisXu52viP4wccJ5gJWebeUo6
Zrh3M0LaagcL2u723GhCnobwbHM3h/9cFaZrGg0WZCPv5+KZFxPPDkSA/Bmq8YCj
pEe+VFN5kF9eF4khEyusdUf8kq8+lYklV5WS+y/vECbpPohHpcUjl/nJMZA7WegY
hEX1wxOZ8LVu/y5XNA/QgiMkDPXM01K/OC4Srp0U/ynwtOFBhBrKlrf5KRHZi9UI
HV29LwbE0TgfVOrhMxOR86Vf0BJj5ZASUVRtsDGgAGnuUcvnCpJtG1pHW4535r2K
TfvXM6zX1awz85lFH1ve+BgI0klMdw2W/+s5yoS139XHadwmEDcYxA50q+0DrA/M
eEbJo/s6Feh50KLcKWzkPbJu/l4xK+GGQ4B6EbIHbCE0l6g9k1S/iGSPfary1+//
GMN83OONTcjP8p4vlEHlThf+h3dmNUeFvUvmhiepKMlRmPabbEp0sOgHuMQXqlgV
VieAklys50VIzhXndYUJDq6JPqyl80RG2VFBwvMQ/uIHpLk41wCBNAiSOYx0qLti
4iEkemrim6S3RytqGti6apYmgdUTxVaGla9PgbMU3aDlGuq1o3YPwb64zRDQ38VL
I3c1+dG+cefALXKyNYk4mPAuy1D8tSH78BQ0X9Th13Bv0UY92DapR0P181Zck83o
CGFcsz1orVmbf3RBB7USnzRJZURm4IaLJwuFHEw7ImWP3XdPBVrf7hSkvENgCnkI
HsgKaztQiZjWUfUVxdOIAjV8ba61qXluXAUZkdZPVOCLdPCaMhcc3RG5TfL1J8tp
DvJB/J1IpkhvVoqAFJsUfcpsYwxRIsNRKgUQSyZdIE6q0mOJLQOqXAHkp/yqjXb0
e42EPPxOJdgfdmx6jzLT+ziEF+spp7tYmdPDQ0HAhv4PTn9qXfO/yxGTh3x9sZ/F
A8hg5CyO84CoWWriekRD3COlmvWTwXKTIxp+PHSUJXyDvHuJauZkduWHDrXH6X2U
b6b9Kd4fecqzrPaUdy40hI8WWFk+Pm5VIvE0F0n6kHW96TMLxa4LG8bg5ZaIgzij
DFxhHqtMB1bqCBTMc++n+lHK8I3847aMGh6oFsO4v1zFYdf+d71cR/GMF5hu0dLu
yb+a7/BPT0YNadZPL6PF0etgxLR8N/AH4e6+YO8BPBYE2yy+uipYlJZ2EYkH/KxX
0c4e+4aYIfUq2LUwQRTOuohYAuorZ/PF1XjrYc6oD4lEu7Lfvf7AKLnCvboPdkGA
3jdgYpmypkB+lrVtqRyvhwOPhaPlzuFkPZPkoZazWUSHiEmN2VzUZnBfjuggv5lD
XUHHVLql3ezGNZIXUG3+oteHDSvsHYzCGOVgl2tnkUEcXNHNen9Wp3lEJU1Rlc46
cm58xwYIeDUjX0k5yoyb1W62nQ+PDTIfRblNIss+aLZPewvUaWZApKR4oSgbaDfq
0jt2EUiStpvGCU9VjkNDruhp7xVFTkyaGyYlEiepjk+wcY23/GrVgsTbN12Z73Yf
YZ7jkEDmEXeNIDn8Z9bXntEmTG6vCG82ZM4Rs7CjaokJBm2NLJtDptHNId57QnJv
vbiysCx/9se9Wn5sNkvWOhfp951HK8TCwApNbzlDTCtDgY13uoeGOmqDSYdhdrPX
440sWJj30Bq1+Xl8PefJ/xfFLz5rT9ie8t6U0i6vK9tVPVPNnFyhCHZVko5nuS4e
ayjrCcRRhSFziKZsMZltJmkqGs6/KTmzjPLVvhrKL+piswUaqbKL+JSokPtNp59m
LawFm3XCVjNrBHnBqPWtdDkkHDSEzaKvyIOJWQOB2mYT1aOqUfZ2PkdhiqGPoDGc
T48J280i3vTsVx+EvII9Upqq1sLbStrzd0uShpJ2Cp+zHEIEubCji8t40ZcC1Grf
JOShM8zksMWeHJjDBiOMpAhhrRwdn2xBEXYWPst2FoioQ+O9CtNiKAGki6oQd9Nm
hkB5K01ibf29M9+4Y26yZ0HvjBKW/Hrme4smbre6UGCzADKTSJpmplkmR1LrirZB
AO60wP6TRJlH4P79MS/GMzc98ot/2hruN0Oa1TST0aQMRrNJ83Zdc1z6tcTmmws7
c57WQ03ytvo/NkRRsvcqRZM8DcwyIJpurBWyFVLX3ffO2az9MCMV0Uc2Cm4sbc6s
Eu4HOPfKcLUrvSCJS91goYw5C4QALK990VlV5eOkSog38iFEwoLIjXz7EziaDEhT
g9niklPbA7B+evgsLXAyGQsRIoP2wY73GygLohW8lnIS+iA2HBoi8A7Uf90irqzq
7azih11xhtw1bcaB5c3slu0uN8OAiXYRsXFk2rWaFxheQ/ue4zaMPAm3Y8vwg2/4
1HfRzNMwj2AAKXgYAt4NKN0F1qPsGfaQpP92g50imBkuRApHCnewDPiqkF5kzMwp
BfX5GyLs37lMpp265Nl5qJY5QIFgWsKoQdXRIf/LDao46oqocc8SJpTotaayNKMW
ShU+bFRdGbL6OUb5nYmTmRkp7AEwo2H91EBQonV4U4+qU+XQQtUTDnc99W38EZuk
C7td3xqmZzzJUpymX6TTB2JrJFM1OGlN5aL2/ApwxbHZx03C1UYaggAvJWhXUJmZ
9AE8sXNM1yKDfcwsCMj6ixu1w41yE9S3Ft/cmnDmwvxlLcIQfv+5drKJ1QUf2kDN
AvciXkIL8NKeCpT5PaC9bXt/WR2W4uZvYv9/8gnKOJAkg9KlbirgQ9mPCSCCg2K1
isJgG2RDW6RYqjDCWN0XwkwWH6x8mScDONcrjkCFVJrZvYX4Ymnak6h488Vwm7gn
GzqkWRr0aH4Gc8wzVeNem3kCbSgCULmjNSqg6VLqGKEUrJwjqbubPE3qVOhe+tiZ
UjJRBT6N7ddw9aLMaddwzKq4btzb88zSgOxB3H1467TGTGQnZYam6Goayil4LLSs
EfnlePuFESv0vRcBtMotoI5BrTtw3ybDx7bbbqxVuHIX0nt251koqzPvlQu/NPGQ
RFsFCJcKChJcqcbvEe/Y0qoXPBeFHXC/Pk2wCvukL9AOoKAny4BV070SD/Ky/a5G
3Yl/qlvlQ6bOyIc9TG5BWZ2iYUM91J9m5CH66JGKxC1s58qGLLPuNdvnv63nb7BU
/tpB0eIaQMEzurI1YwfrU+9vqlpG+kl22nTFxYGJYPPg7K5XrchbzWhwOPEpiHHK
BSj/AngAzthoZiMye7kSjmHU8B7zLvldJxcZR2VYFB72Y2dWP6HV5yL2IyauiXfz
ZbOp/gJn1vTCIuqeX8gzvmQ0OFpP/lrj+kwwOQ+693va1+8RLZsYNWRdH6BWR4XM
yNuDSr4oUNqXw1h/oR4sudcMeIZc+YtfYYgsuCED7QjB0r/CCY2LoZ3oiXnTJZGC
CZ+eO0tHHHoybIgsR3OI6v4v+uhz4gYFFAgvU1hJfhvctf3cIzVbVPCf8q0MLhwV
VvnpEN7rjzpHJ5uObMWDv1Ga1crw0qlFHmPZTyc1ZNf1G1PH/1vw7rjYoIx3X8Z0
AKxpOb8rOwIs+mMuVkGQtfJzFKCwNnZhKmfHLLm8VTKEBkIqm/ZUzhDIW010l+vW
okxYIkbHyNVT7q3T+jUbu3bZjhJhxfrFhhtLEHuLBwfvInkdqrTR/s9n4nMmqUgm
lr77ztSd21frdXZRm+iazNb/QYAdHmFCgXzEHbR2SFrU7nQ/UqYb5LysD93KySAy
9pyq/FymiD2kPphABEaumURWpwmZPqbBlZf7pRfPIaT/sszGR9l5U96LmzqdBa1n
Ax2WxtfnSjo8mNRjx49DtHwWzeR2J9e9Y+FBhTvcucqCf/uwTUG5YuWhhNw+L6cn
J/IQuQ1fRLWVtqTrznTiXjYRdo0vrmxDCKw5pxlP8QhNlJENW7/jrWgSxIc2HyuP
j5TX8r6jvtaAHCpiHpjBrzEv2+oF7J1hLZq7h+3RJWMiHvkt1oXVR/6J57Uc3dP6
CF1Iye1Z3ahfgcV46VY7PUCvOhVWUbdGdmW7ct2X0MBPT1y+Mpj8NWSOh8oYS5rm
P0zhpcmI/AuA8IF1k24VH2SjWXAS1ceIuy3gmF0o5T65yKjcP4OrGFRpm9EqHNFS
amjPlImshQQNAiaIliclFUyROZSoGfgpfMgmTjn7fwS7o5dPYXWKOXy+2HCsYses
xRbheq7rdJVPAL+U5Ykm9sTF5X3SFmDFqPbaeKLlPCljsNJAffU69kClD6sdexUf
nFpremFiA7YsOEOPYvFrNg9GqdxhkRVCfdEZsb4uR0dB/jmSB5UTsdZ3db9rCJoy
rIIwm8uUAlF9z9ZFCMpft6MM4+KH6xKEBr2ubuZ+QD1rJL/A3cK+aR031V/XoyKI
4GBRK2o0vfwZGU6L/8T4pedkpinpQaocTvmUjsSFoXKlbk+/X5utpvzYjBAR6R/v
JHQpWHs+IqBBrU6qe+t4JidPvQ1BoCpqQEDsCElPeAF1tyTZ97MUO4pL13/g8O6X
lF59sH3rAVQWAfKiNflPnBhkHJeDDcilsaaWTL7DLEzsArsO+PyJ8/3XvF4khZ8e
9Dukqm58OIKfutohd9VK4UcmP2xyD5VD9/Asj4DPnEG2kht3CI7T70niQySrRcAO
GiBc/w/RwjQN1zmqZsa6h9x8tdGbdFe1w1PwFepSmTE+IUfaavS+fTEX2X6XnKnB
Ov0wuazqdons9rId5k/ktDtLhQTHBiZaMIA7MDZBkaTfeeahGQHAlFn7SCaYJWSB
J7EmHlwinxiJllEP8LK/pi1INrgnRpdDhEJR/zjyqiJ+mqBUN/OA8WmigEM8ZS8Q
zGC9P7fxB6QECyftnBrGh5oZXvEf+ONy/lmW79OvXSitP9lVQwlZxUW8PR3MJSZ7
L/Tb7FeiJ78ybXP7EaX8Oi3/zSnZNjQOyA/kPNDL/3sI06KAlxN2NDTnNI8L5y7w
q+3VhFBKokFAa6KFJ4d43z57g48gpUMP68DV8t+JLDc/GruOTXO8T6zgr8kkVNn2
/L7Bo/7Uwti49bJjUzVpTYjTx8KcONAbw8wESoYKK5p51pXUzDwMdOznOLWtxsna
dUbKPX0124wY3DydJGsAkdwnXEusOdkWcdkntWuMNvFcaRQHeViu7mMOAZI9HwnU
N42Txtfb8U8567gRvhQvOg6gVkz7SWjcjvM+JjgaOXL2IvfALU6+74LY3Xpw/leg
IIldKUTg0WBeMShspillWMmmIe5LYZ7uGhD88vmcigGOIenM4PwJtm16zQVQd5mY
3vs/2Qp2RIZD8jFbpAcetbdvQCKY+uLzublaeZ8HRD/oqC8U1RN0HG/JCTUPYVsU
bsB3GGH0H7POcjPsMm/+EkyijvP9NO7iBZQAtzIVC/sPtelyBGSaKNjqnnjc96+5
xT71nwOz2g6r1VVzEzR7LwLQHlgp5ASNfq1LAyZ2cXwWMpRsscrhRt3NXyCB/I1V
23l6cnJDFRZGTINqfj4gbzPnRhqZMf3LPHvaIZkuUc6eQbIz800duhmooyP0PCt/
GKL/5LZVTusJ8QXf78z2qLE0KYlmYnxMK4tqi3qm/MokEJ7YEyOqkIUhFvaoun8R
6qyXzvIjb3rjh5KsqjdZb0b7nRa4ECUXFVIAl971fojz6y9VrEfUsnF7I6VU4lzP
E5cCUQ4RsnCvZ5I5sPbZfcDwCWb4kSaLFde07Z7viH/Ta1jjDI6drFdXsOxPRZH5
vjEQz8HiSHIFdlwA5gIXj1Q37doOWLn4x20syXHVSeJS/ViLs09Pmzzql5IHTkCQ
tn6czf7G9XwKj/fBtAsasfFIQPcV2JaEcEyGLCg9Kt+xrQs7/AlZTWZj1Z5f6AVD
6ZviqZv5XEPoBdROe8zK+bnnwSN3mmxSX3n+HymDQ2jGJAiHjJNbQKG+8E1A7MqI
rGCh5KJzmNdrEZzAKppr8OWHbIVcaiIeDW8XqKinVDBANvmqGtwPXtzm4tTNQSJS
i6BYZV8PJTv5QAvgbG52n4MIoQMax8ZG/wSLZjBYMa4+7S2BHI7vUru+azI6E07F
HQ/qTzwN/fy+onFGMkKtS0JQhlRs2/bM00Tn2Le2+50yBpe4MlqZnyEECtmUOYaz
lMZxuL3CLTEHNtzTIgFmGaw45OcZddgDJKT2a/j0NKW6jzrtTVuSC82Zyn8mKcO2
RjjfEKV92EGVCpylNoMH388B3T7P9rZI0hOqGtGjMVdkfUNnMOohnIyS/tUgT7He
DQDAlJo301RPR3AGS/zs38LYc4u6U4Wzn10pyxSd9O+naiPTQnO5o2Aoef3Hew0L
t3YSj5HDz+ol7cQ9kdGVER1qvAVSShVMtKBcrDetDHiUn4CzJmAzWFHDUoQty2pb
eiBxDhoOpIk8zZ9sWm8HEIWFE5Y1xLvGEuZSp2cxgzu+hKRzjgQbjve3Ho4xZyMZ
Ps2yAeaNsdsd5PiiXHZAZzzBWp9zo59GX/rb/WjAhn2tomkPw2oFIsHTRVcmmnIr
xW4PPuf8e0oe/1aWKGlvm7y6wm5Mc29WqiFz6nWQ5gbCm5Fs3JBkR6zq2T3p49Rq
yOTm5JWBt/k9ofMYzXqXN+nu7UxlE3VQ5gQ0eMiDc+rl9Rp/ILHDVJcqEUnzZ1Gx
lJQLwae1E78e5VP1UgGQ3PhKUO9shLE9D4qWRwYf6Gc+zGh/piK/becCN+U4Ix3g
REo6xFroVKEevUFWnQLYUCJ9gAs3/xgu/rUzPuUW38DZNMZHqTqoEvgdeuPSxWyZ
9a5HNRRH+JA9CwXEV7NaOGruQsch8XCptMq6dwmARrukb1AEekOthOHpEl2fdibG
3aXgDoejKxm+p87wNU5OHQ7Q2QipdjJeQgyWYaeaTczflmuQThuQ8e8LYtCtwxmO
01Gm2ASCvDChiPtxRf3e9wqjLJcJL7PtuZkOKXKXo15P1fDqbrni/Xf6CzdixBOD
RoQJ60tROxRNTUT5Hkil2WUyIEBB3e0K867pRS+VcahqBoD9g0QPNhToJGE0lY+n
l5d/mUEZ99tDOnCHEuDziGk/0vpkWIIsI1W0VX6X58yxRQ44wfcBEipjozicVXhT
qLdEe0isGsVxW3bRy3BYUl9jMpKgJxnvevw2UkQemThHb/yMWSG+wSmZhfzi9De/
cwQfyHVcGrVWhLocii9GVRCuEastWTsugmQYjqNYI/ITjCQTDw8Uk7x2qG5oIyXF
oqrQs/MRafJrgYIcrmqnzwcwyZ+9visL1tTwtF7CZML95DawurCL6RIeyymth5U5
CZpL4WQ5o1NnttdQm61sZgpc0E9e0Lb8hg66uY7ZxnxTvu+Dlljq3tKN5Y23eyMj
HwO1AEAwL8OJ47ymQyTZ5zfCtdTgSHA1xLnCyfr+VJWQ4QIepztJj9N6MvzGMWYU
qFlfvhwxSTz5/NUN6x3wmMpwYsz68Y7HBBhzt1ASC0LzUm/tyfw2zADJHVHClfcj
sAQua/9liLWQtJFXORkNi6cP7hSvQ5lAoTEkxgufr7dDmON+prdsDjYwoJaD/EOu
yT4I45t/5zHZ5ws52UnyBqecx7LuplDWP8DYep9vrmrPAG+O8RmAaDFr9VFR656M
QTMj5VUI6pqrHVumNFQZqVlEn9ptSp0CCBah/jIbypYllmXPcewfKADKKE80bg0j
dWiPIL4CrtrvC9lehHGdjE08/O9lIwMic2bR/rq0X9a9CZuhbMyjayIBQfWICS5P
tzSxwgcr6F6DRmwdyRYgNbraH0618GqQcXbj+0eUrBlKq0A9ZmBRD8hbtwaBI5KA
lXHcwCWT0urfjZP1dmWiZbh5oaqHIpcZXSp/Ua9TiH10OO6DuT9cjKjZMt58duKw
brOHVihxKeX6prCgW/aZRFtAicnqKFtQh0m17dWQRkXuuRaZgCnXbuZa5uGquIe6
sg2GNW5qFJdzzZ+GW0g/MzuY+yc3UlbVRCZZ/ncZokElnyjhSdJZT7auyYZg5B3o
oGshGI196s3zcyatV1NYgVZP1SXOemPyw+J12xvoXqmCRLvpCXptJuydwSrDT6qN
qrCSIOajlIzAJnMo7DCKIslwN2hAGXf8OGGGgPQBpqF3JtepoJEVQmNZxrJpG6OU
j+TjCTZOS6tJXRG4oBF3VE7m3kJ4kKxJaq2z0MkU/Y2mnoY9XTM6KiF6J/AOs4qn
H49Mdtd/b5IoeF+uMtbsXHxnDGxn0EIHUxmD8ttMZhMte7VMTKkPOfUh46SY5LCX
f03sOnS6f9mpTsmmneKU5y1EWrPGGKuWxNv/CjMUBATty8jYlEOP6pfkPoOAm11Z
TSHV/W1FGmcDiwunDOQk/6lMITzvb+1IMogQFZ6y4t9FAfC+OH5f2Bj64QBMJL9c
iKKf2regc+FWqA01Tvu78HKsCl0Omd3Ah7E3yAargj75Vs0qAC2UfyufISkR6w2/
35hRpyzlmKrnHy0eRr6c6VlpEi2rR0BmqMsdmQdnSTDxu1ObXiie4mh/rfRppaIe
2ZOcEFR1yF0lEykKDda4b/ZBc3uoHdWozVN2QY8+h8+RLvkxGEeHbz+z9LkjlD/6
E6C9r5jEss6LuwFFTA2AfFiaexYS9Dnb43Uv2rwrK8e5Vwd/Kr+/BAa+X68hvI3F
WZUWQPdHIorAw09ASRdRaaERiSXYfbq/cOkYby43IYHvHbOMtuJGAjbSrwoiRpXh
FWfT8dnAJlzqFW4wbWuG2zw5E9S2OE1TKzwOP+89dVFvxWOafnHFk/RC3l6PErdc
aLH4AoTysaFNcyc26hGFRzDVA6vgrZb4JRas0NuGYylULtSjB6bYa5ONCIiNVzdu
sipx6tvMw5FGddg86bCZK9vdYeGkQ+v4QXoUphgIraFSMhsE+IKBpchLj/CaPU2X
6dH6hdNtl1vuRPJZlCM5/Zyi9KhYdwi4UyEYYEYMLbBAkoS1bYU+KFSMxftlNW7j
9qgqwrxK7Y088RUKrVt2hsM2WYSNCW9ahIIysnRpsCTKMDgHQ+h2wmHphYCkWx72
ER6rtjJXITdTSYQoFL480VG6AXErh+L9LtAhOLsjghGA1QzXjv0gcwiBBBYICthf
M7nJJXaKSJQgPZhJWMzbtqdmGG1bczkBzrpwJDmGE++9jBA6fszwAF+qUxprpGVt
p3mYNyHu+yjRIug3UbOaNkr0MNOQZDScIauEBhZ1faTk9rNTdmHvCt5Mtg4p50Ba
KfUFvbh5o4aOroW01QPG5ASQKf6Y7FdLiQgTkQmfrfArTdmhMetJw6rtyA60Ftsc
O/VjwXjRLRatSnrAi9Tx0SwFUimD5/TC+BKeg1yXta7PcWOnEYHrozKU3Y471uw6
Pt7q3+eOfMO05I+tX6P/aXW9ou8esUOhPs5T8elyXFf+pSQv4AYECwY72qB9pCvY
nfFfHjLlys33hewEZ3KnbNJIBhsc36ElF/tZdlXLmmSI2ZQEwXDP8g/M7RtTj00B
ZvaGZCtR2C5/rannZVuNCnFcyQ42YaLvhgNdPBc7Ym9oSl+9CPwzcTdWeI7dmukA
wag+V5UGIQHbRrZCQzKj38FHZ1hcsKso0NmMvVi6IXLi+WT8ckKU4J2Le0Ky2Gvx
zitwco7WQx4MYBDWgWNURUYLphE2Ieo5LO0FclUtKKh6aVLadZN3FTaBTkZ23JZp
6FA9qFC3fxGPvE0wUv4PbKyovnPAHItoL5hGhoUalXIOQ/mJQ+cuMnYfUDhDTTXZ
jgQyCdVieiynwyPWcdZrPYvEu+YqFstg8h6WcB2cpRMgbdROUlzMTnQ9He1fVAGx
RqkD1HezpQmUXUbyeUqulC9W2ZjCPEQ2d0c0Wb+b7cQo7Xwkf/jjtnvVbSQDXfBm
pSU2WNLI55+KczR3GdTCJyn0Resjx9oK9eSPdfa5M6YMdF/i06FeIT7NMJx+GJRK
VssmvagmfTMj3XSETNrPF6EEPqT/wrS5A3Cmwt8O+cQNpUYuVceLdWAbFtLjPQav
5HAlCWbxvpDdFOZq4dp/P9Xdhf1cI890qqO90rjH8ri+LqCOwgHQGzLHoRRtmr3F
qSuaKNPXVKd/ab/l9/h/bgj2CN4Sdy1XImyk75KDqw7csyJEHk9q4xYiQGnOCQ3b
8wIOEUiUYpB4kKwJrja9dnguHKAnMoo6DwWIVjfRwkgg2iqnpdaCOwh/IuBm5iQm
ybclmCWxqQrl32e3rwGo5bTMeDfXW0CHmMBReXRLk81/MW7KAjQu9qWmhihGyYuM
B3UryZ48xvKmb/gxWasepLYHAObADD0VMS3kMVh1pfJNIdQ+MaK/zwRNjUA/L50w
g2caP8hI7D+RvvYcOE0Z4MWtFURzWcXMdw8Q/OoNNlQQUtl4aikhLlw+TLlydK68
ZtDsU7iB0cQ5yZFPDG5lgCOtSrW663JzBAXkzxgtXbiwTzlff61UE+CjOo07rBh9
oPUO3m0Fm3Rwf0SgAe2DkuNbJQYkw91eMv0ggz2Zv0byjTZrR2/5eY5Rob+q2qnY
c8TFd4Bbt1CcP7nGbcTYj7+D0ABkk9nbhvQU+lTaCjirVLUHE2c0wW41s/49Smak
3XW8jHyrph+8F1oFqzlQIB/apPOHvbWvlJzd/w6yg+6Tf1Zvhd1k3GC9oXJmibay
SycPb8610w7VW82iAJ9fEK5o88vzJfkES0lbjfGLwokP0x4695m1KRaiYM0X24oW
Y1TPJESrNofpIlxii5SdOpGSQ9R2IlMHaq3J6NO3Rboyvk+KiyvND0KtHDOHrnEY
jx3PL8eUH1VotviZz1+H3+cmgKq0ewFqYjW3+lSOKYcBMA5sz7iJ4tb1chdSMSyr
shqo5W6LG8XjleqL5NYQWBe0uxLUZ4voi3XNkQHGy79Ot2xCen7zLg3HPSlZJyoU
AOcfgCkq1H772Sqty/+J7F5V1GxRFkdsvc6BMVnFpfyw/Vb70cDZ9wXNC3f64RHY
RDYy4vvMmfn1gPbPF9H0ZT2a6S4pAXM+G6jyL6zaYbTfxy2L1IZhOweGXOUEw7aa
yfncq9/eYhU4PshUpP4Z6kC1Ni965TWKkSAs7hzFjTsUASH8e53jp8GnmyVAXbPs
RWT+zahh4RVS93RxvWhFec4RfaP5D17BnhwxwNq1dRPPqNMKffs4FNDsh2+A2eUE
Uv2xE2Uro58SoZeKx5l4hQ6lHD5LcOAQvQt+4eyrW8Npiq+OidbXH5/4KalUIYja
t1TVGfRSgnsd2SNLgQVaob/HWEpcVYrI2AcyDCoK9p1yExw5igi8ak9kigrrrDaQ
xTGi9jshn1sPQHo5XRZnHNGhebTQ8qtagqoz6g3qxp/GAClvprpcRM7st9BdqFCy
5U0hSVbDtLXLbEoFEQ5HJv3M8AItKLLKBCaz3KnCr1vcvBGWMrR8mdogMC9IcfIG
Fx6JJFPFgeR3vPOjHGFiI4TvbbfO3C7BvEGUQK4cRivSgfAJ8dBB4t1m2ZTHIn3f
eFWud4IldZ+1f9oe9hsZ2r/lXjJrLSNC/Nk+IXVjcj9+olW1vMVsbXKWhz04R+6z
FLkeyIpXSCc2Wt4xMaCCvH+L+8G8WdGJoUHt/JreVGyRSrmmX5C/DIXQ9vGqP8z5
upw0+NXP8VGUYbmd6pV+3VDMoCQ9ktQNQpZrB2KttNsVsfNFCiO72etpTbIdnFrz
nNhxYigl1512l5aN4ZLOvkIO9SPk1C3VPrFz2QNq0JYewQtyYA4/5mDdiJxiHbTM
mme3Aw0ZVjBjXZoMf+1YJLepOUL5HmvBwtZ62wmXR1g5QyU7/ja1yr83eTP137wq
KrF6pI1Pv02qpG+7LIKyYMww/lm+Vendb8j/wx5JCiTQnb1l0PBkDHmPGMz5M3yT
nI96gmNxVmZju5ZpDjmWqIFVcBuwugDsYOkTHqFM9wDmBigXXiPrTmXWPkK3LsiD
MjfCpCABNY2nNj/eWZPAjKzg55keQw6A9/xWEMxVq74kOSRYNjcdAmMFpDDkYjri
knFfkLpXNIxM+Mue8Hb2ITMH5jsF360/PX/sTOyPLbK7hVFr93h2n3Q949J2SeGM
OuasYzMOAIDmm6+C5Ov/oBlZNkhspZq2jJreceOLQrhAr/mk2E6ZjxUKEY3wgh23
fW35RPKEFL/+Ft29x70oLjfCJMJEgvTNXLn7OR1rxmbafRU2NOm+swZHoQaHJCyr
pmBTK0egV4ftop4eAXs8Pe/J6nDkneDWwc12WnzUpDD60nxshaHLUgDMHtNbKz/4
oM3mDnmSelpbRaiUclhLRTm78JMd1feK1FBBiqsT2RkdjfMGB94qUPwxPGEbWLyR
/HtUrpaYAWQVsVVvet+g0/XMW4f6zJSjhx0Re//nGuOe7X7TfkvcBvFLb4nqcXNZ
C2YFfb9aPRbaBNtmnkCO8gT9Kr0k+67XytzAc2mU993OMaJ2NMpenmaUpuxJ3K0X
A9lnNep4N7GY00ANs7Ts6jQpcVbsm3DtHw7n/MJKXIjaLx+B2Ecf0MwPi8ioexcw
Y9Z9IiCGi7Yq6pYUYBbKCnZyKoOflHKEXv30NseAUFEr1WF1t4Il2kfezA1/7jN0
dLMA53w46RigR85TjHJiCpWZ2i2BBFnYV7MAS41LVL5iH/umxY+/qQBwfN0Ep0s+
XtHUng9cv5Yq1qToEqfPfuKo68ZcfcpRY4IW40dnFcTkuzPo4Ugs6STGoKWkEtNJ
IwZC8Qckpq27PGyrhY9hj6tEWN1fxSU8AZWOxXbKxjRT4h0uPnxIfwMBmlID97jU
bMhFoSwgooDYU+yZqdKQ8PtqiKthYtiS/woGUwaod2ioSTEE+gHecGSf5uD4HG7A
jFAMngjrjvd7NHQL3zy24tyBMhYKBZKkIWvoBVL57JG7/gOjYfHsuT9aoYm6hqh9
7h1Ka4YXnszmzmFF7894KmA3Nb65kESe6RsZzAoE8SSAU96fPc8uJyMh44TREFkh
UZFKfA8SXt3FCDfIB0ESRlP9h9C0X+EA4A2SxAEXOQYEuA83WJhaGOHNNolH7qxL
waxx1U085KPl8EDQLVvbv2FvvgyDwrQsBXlnB1l14QcA52KZEAasJekF4sIwIGKi
xXFLydbBlUx0p0MZyrsSibKf223EUYArvGTnDFc8BqtTfyK2SlYYVu62vBpD/5vx
g/PHwm1SB/AEul1wzive7zObAasnfWCNZNyDQJ5hp+Ud+2yeNfcLYh8B2u1nnncv
c1zJ1y6s2vwrWHEBLvp1x/NliVmiqxoaQshCJWdik7OCf6ZVPS8L8rImF21e3RUL
t+PUe86OReetzspO7UTHqIBVDpwT5VmMq1KPEJXI8ZfAIHvQZJDQSrgBvRN/x8Pn
yhE3wsGKG6t2sxJiMI11fNJMvvTJfeeOA8NoXSggj2IOMK1FZ3jMKUjIlRLKFVJe
/Lo5RMf47isRO7c1pwDcW9paoxzAprhHPNsXtYXrgYKuVTLZOg11B/e/1UScWgtp
0oVjSJIz9k/n6iRNjUxiNyNtWhPldlk3TTe9kU7wY62vmUJW20/eEbmhLbsQ45sj
qOnBUB4Xpcqqhgc0DzBW0W3eTGJ13TtnnTo5Tif7Nm95GE9eUVSZUnsQt+SzDBNM
kkXZ/Hc4FUwSw4N7U8Axx29CZ8tx0VowaUl62PS0WCtSiaLC/DY5laFZ8eQGGBFD
nCE/PQaD2OXtlOmrkREk40tU+P2CTQIdQwTakhvEOqua958bXJ1z/SRjb3lp8rlB
QVs1HtPpQTMdTyCsh1FSGVZAjqoguRzFkeaAudAm6stTNVKxcPTkoGogLlGp53pk
+Qrx343JJP/Bev61wF/reNOkl1jNQCn93d3oRP+uQHXIBGsVlkMovgpQG82XqWt3
vpoekUsGRbKz/y3JF/jL7flfZiPIwjSNNMxa1K/EB+EGnc1MB7JPiDdVAtP6WpcS
SmbdYcwABFEsAh1/alG9m1BeCbyLZNKuVXOtcHpzdO94WoFo3C2tExoqxjpkgdJs
YYcl7IpbzWB7hio0qAh+gZNr30JtpxnNzv9+clFj84K+B0sO3no7AxW4OyCRvN8C
rY5MVKFBgpO9AINYbzF7tOB9faMS+kmB/UQl7G+37/Xy/K4p4sxsSth3MZWUGxsR
tbg1Hp1SbXuPDANd075ZyAmh7RHmBPW/OfpUODON1OASYosjHtFim5k14EmE8OGI
JXhx8259HKwsY2JVn61VX0TTYD7qHgcg1VfbIUy8/j1hEQ/gHlolk1HmL1L7yEku
8TbsQLaVG32V4po2QRloFNLFQ0G20L31BHatCkGX3mfvpAUpSodM4CpeSR5Q9bvG
ut/5kIsmmnQzEMFLOK7yIhdKVKeIdvRxz41vkgF63J2NSIaTtUtm+neIU5rYPZtZ
TDLv+OYaDX48sfSm5YpnHlbL1GzM9170nHF3OZ/UyzjKAtxvfH1HzJkNqE+NKbca
K0Js6brN68Ca3DIxFhCAdL/RBtpH753d6Q3M7KYetIEBlsqq2FiamX2oY7DB2Q3q
OG2gt56ol1bAkz7jXyTtlYhMs0nWqL/5/fHfAHp/vG3tssS2vf+YHNoscO2fjDoQ
qd+ca51TQxQsg6K3h4YgM4poV8FBf2wExeLq8I9OB6nMzJ2SfGBaDtG9Yo9caxK7
dl4fdUGmpwIiK6JlgJcuDSD7N/oOuOqQ3FmyJKlaA/s0dbiiLRaYMFktotRQENao
hxBLiVq/+jcw4tkj4NhFYvHqFOairr9FnZRRiB26wSxhlLdprNRMLEP/ls8Pj0wk
Gx6/bTEAwFn0Uis64xkhwMenYXlYWswOF78zvdG14c3CjcX7a1AkmGfMc9Y3oyZZ
DmAIMedcbfnAM6VLH3DUOgHVImZsbLKc68bbOL7tiVIw7ASYmTJFnGdwpkYGuGSH
FCZ6ciw3of8nvh7kKqk15oqmSITumkt4DAeVGMrQ/aF0rj6Q7DEnfGE/cf91T75w
cV/YUzLA1vhbWAHfwc9XPN8nTtk++fe+MwPcwDrTH+Hajo4BgbC0UsZZW7on4hKs
QhFrXDd+NCOZpPwhw6BVc0p6UkrF8EKLf+26SHZxZdG0/Gtkbirrk/kbPstCrS8u
mBqNSvhXJeOyH9GpX3PkQ1CffT37aCzKeAyTO1n8RBbtTeR9XvDzQ+phaMGPBhR8
1anirm9iXg3gLH1wkfAXbw+uYUBru4yA3DQop09SvLFn7J6OvwGW//52yoW+g4XR
yGShEA7p37Re9Gfah5iKdzfmP7RLmA3UktrXfnQUUpP53w/6atmNRDNGU1kbr5a1
LLrXR+z+LmfVyFoKiMtW08k0MWyMeUUCAkblLFm/6Q+3lNQ+OgwtalL0JCwIuZXl
HMrKSCu4kxOnqya3Nsu8RB6pbEkvt9GMqoLFucrHNKTUuZl596TiLPtJDOzraCam
SW33xu6FdCoFK4AvfzqEH+AqGhPvBY16gKNEzs/dU9okHryjDbhqK9B9Ct8IE8vL
Vk6DkcTIBnSrdRXCmYrUyGpVnSYcxh4lSnWX1+XzJ7Y9HG5tfjTwxdSDv8B131KB
woRxFQ6Iq6KYCzoJgsFshDtdE9kKeHmZTlB3BIDza/7aV92q/h7JZsov0Fh/nL/D
MqTq3sHWZytQq3mqzx3RurphNDrPFtysnctqy9ZaPG4SVqxOOX4d0Dpzmm6DUO8L
UZXaQ6mVH3F2T6PQEI+1Deg1T/tnhihWLyeyBtrk3zsrOtJZC2Hyk3xOc0VZeKNw
g/W5eT1D90hMU4CsBwkKPofBmAK0fRH7XWuIawvSQfSc4P3O8Hr+YXWnX+73QnEC
cORJtXdDmlJWE123lG+3eQk/B2bV1Fp5T4PzJ0hIcNqOMnfoems8RJcde+2PbrI6
KgpXtmYccS/3nmMHxUkMzmzV29KZXUL5FhwVqDYJD+HDNaIXqE4NdLnriTvdkFnc
SyFbI+cojlPxhy/E+2r48fhzQHXC7wD94ZCr0QKaQRhORWvUgix+uKzaS/86/g3g
+CHZCTN9ZZyQ73A/GlrIlJlzwfoeo9U7Q1efCIjPLjt85Fkc5z4Zh0V5h5C9b7Vf
aNGEvARLCv+a4v19YfagbQ8NSzDNbrsEwTrJ755wvB36z8dx4cgdvl1f2v9iECpQ
gklwwRQkSeFIZrehPqL78hb5TeGhPWwHRA/SuZJ7/SJiI3xmor80ckenbXa7ueHu
c07IF+RyTgQeI8+Ha19fZ4ygHkbkZQzyqUzDI4Ke+pnhsyaiIwWHR5aI2u9gg2wY
icZCnLAp5tHdMy2I+r8c3/e/rPG8M1v88gNPjadeC/Qz9vsy9aS7WBQr7x7CUjnq
pVB9g4mdRsY+z3qjOs7/CiUOPRz76jBjoUHbyK/wDf39OHdtXsOG6xbdXM1IcwHb
bJ6mMym4Fe435/80qE2t/uw/0yPhvNUpVE6o/1sG/jdYQvuvmaybHus+8X8KtByB
/CPbYwRddYL5jx6Unqf4EZjOcC2ISnT0WAFVV/eAsZlwDTscxHiiEK9iC5hXqrns
IP2j1X9o305JC81eeWqn4JMdc2RBkfRdppeG4t7wFloYYF+ZcgFhAvUDhptiXuoK
CrlVH60L5iSzkE2J3VYjPZ+sWRlOJZuvGANDQzRkcCDLXCJi6ZZxT2bZlm954+aK
yVyofbB2+jCUxOplhvaimdtGwTHvhpwxL31vM4tw9hrBHEDiH76bDdLgXtBGiByq
w7l72WNeCz5lWpkjV0NhFWeTPWjuyfVlJv3YRdK5TD8qo8cg2V2y9bUOPERfmpMh
HuaNr4mJvFYb+2s0Bivn/gA/RwpT2GKwAJnqJZ+XDXQ10l1sy33UMrpOIC+FKMLv
5qOWHpYLnLNDWuW1ZeFPxXCDKYpQxTVbm+M7LtIa17T4xhxqhiEOIHG8/PFHFoil
/la/L8EY+OgG2FTC2DqOO9sNPhLZnaNURfiUrAmEu0j+ZQJRqXRNh3tY+qpBNbzx
c4M0Ubad/GuTTyYL5g2nJI/pwLrppjYEfUHqdvuXf+KgfsFcrrwikcoA4YAYjZ8V
/R1gF1mZvoK9TVi1DQT8nA9wpdh9YEewnJCIAekRUv46H+IjWixwYQAvmMxoK0DF
dfrzGXelSGMmmRDLNX6Zi6Z6L++oyAbMSX/WZQZ2qcF6HgqXcGwfbQC74z9LVnET
4Dyz1Lfou+YkOI8CQT/yrXdMNqM5eGUacsNMUhjLe9BF6rqaZe5pKtari8EVMND1
q+mvM70QCUIpMaqGrTN8xMNMkT9CGMqDnXd3JbJjCunXtWooUN1sV+gfIERDmpAU
bRfmkBUA0cs2CC9eKRVMAkh2OUH/S7x7xHJyyRCjR4O92adrVT3DY5aYO0FeYTnd
s+0JXEeTXZnIrCJn+kYEznZVc6OE5RJxWtr7jQ2CfF54cbEF63HLvEtVV00hb8Ew
J9f2bS8tRwOAkaaQXBXqct/rHYVkTTIyCi/P9402EADHIj1fY4jvxj5ToRhmgE05
sdRKDujHYYM1Ipmq/vHEA3FBA+uMDBDwpn8F/Ry/PveYUvSY7u55Xy8vUmmrjG33
dhFPlwl1YmFWCINcdhQTJ1V7jS1kVDIWIVhGMian+4iCX+2nBgmD0fVOOLTgYXOy
zdHDb0o9SvGKx2VQ68PFQbAaDPQ1pgNDLGFK5rYaP4xNEMLWhTHNv0sxs/jpz1Ms
O37rkIcd05Am6lgN80qomrsYQVHoPSof/d4loV1ZOreQoFg/V02OBzfi2LDo6cua
nqcWSMBnsTO5ZTepiC3e5FJKCe9V4cewuHBigY1w6j5VO4lDXKGiODCWmSj0mcOq
ZweYsUEHKAN+tWkCVoxBdAKgi/CxDbDSNL0x76B2397NpgGkK2FIyVVrh+omQfI8
7bngTxORQDb+Jb/WRmJZ4VVKfrEsuSzrt5uPkkvfOFRzuzgupf890UC8T+JPyIk5
pS/nasbK6deM+omnZJpfPWH/dsv3XwTGLDb6VQzbJbsowe8KiMxGy673hmpTj6Zy
bv0En7r4AG1dyBP8TbKL+4fXl/Pt/OhKqlayhRetAWZngdDmQ64TWfnDeo9rjLNG
TMB7ilgVZXrTlfm6in8EskFdG6r+NolYX8nE/L5IGjWpenUBoAdfcMjAuiZKVjx/
1bTKL7V75S/r+W9taXr9m9AHb8dl9drT6ONKQ6y03C9sDXHqmCax5ONvHfoYWhPB
TVs6/t7uXawGqjiQOVi0kHHPlxzyJ2z8oEzI9doC6XHlLWGMJSHp/hO0HSReY7G8
fmirpPiRNknqYCSu3QvIZlODKGlfwWpR0GTsPJURQCkWLU6vWPsAPJXvTNlF3eIT
fChN2TaUDNmKfCQPwz8q6DX77j/mj8jZTEab64OXkvQ/7ndUhdutyjC6ezmSTEdd
CNEzlKBO+WseXYwCBeiS78TLrfF1eYB0NtgktCvsAl99jEGTV7MyGLPo8C+vAjyy
DiObjkfXFcSdnbUIVRS9oVJSTqaEA4OTjtBP8imgw8xOoq+v0yq46lT68Gh5XuUl
EU5XLnghCwadMdPgRKePCJrrLzf6gjr55C3L9Kc3oetU9D+lnFfM1Clf+r1D2Snq
Ogtn/2YkHdZcyTWTxmeSuilb+ysyH6TfBupubo/wjwN8MSoUbJi+okQN1rVbUfla
NYXYYPOsi8uv/9Ob/SsOrTQ5TvLQYopC0hrddBTGLdpew+quKcEiD0OTWqGKugPj
/SLdTM5ZbQaCBN8yVP0YHMziG0R96D5SsOn57R0tLyCkNUzlaFy+kg1P+2m5owQH
YUt58jvMLv9VATsSfteX9nn55UYDBmUTB4NzNLpakea0wtXwf46gIVqkD6VgrEnd
eMrUr3W/Bz+bJb51f6VeEdYs8OMyvi0hA+rfeAXvoBxIYptdTb89Liyn9g4wmmRw
kpzfNR6Ij5bIZd8xOYjI5PB9zND6LuoQqDS2dJedVx/yNoyGPf+70khu0pJ95RWy
F5Wc6lHBpDZTWwo4UhVefw2GnL+HNKkLBTMZIvDRN5y4gapOyKsWMKD1FZTLQmGB
bZmOPMF/H6IP+YbShMmSKQEoRunty09nAuZwpvs+To4i8So6XVAS59lDjCW5ejtq
ZmNv0j1G2yBh5nmc4vkSZA0hvzw4ENorJM8wSTz+l6sYiLtMvaAFpvi299nm7Eew
cIEgVpc9tPyvvGSmQHsw71KpHdxLG3jdaENB8P+qCNcThY1vPrW0OtmNdZ7fXRWT
JZ6yUKwFQ998ZlhdC8+dwv+LqDaBi3vnj1WiAKX0H9QTUPQJDXuITU2m+hZ8Q3Q9
LG+XzjW5zsM7CVlMUuWwBA1/2dQSgF+ibAcbij1Gf3HbsQA/faqpk7dxk1vPSHoD
xh33DWvVWQiE0lT5fJljnkoxJ8R14mLM+q4EAB9H+Fdsg7UMa3/92ESAoLj4hhuA
EgoLLHjYUQMSpQelWNoeQUAnw30aL2bDwZcvMumVIyait6VVrqfWj+NJUT/whOEI
YLq7li6yormjLW0zyrtyIqrCDQ63B6jZdcVco3SY5Nn3LH/LYq+LUceXWiN0qPto
gzGWHCzPdOtz8bRTz6tsEx/O1/AyYGpxtssQnxn6MlDSfM5hE6d+i5uOzughIVjW
ZROT1oiNZ5BsSQL4/Txj3AUmbBGMSvvECCztz5TRhEt4dKfVoCj6E3c6YuKJBN1V
B7dWbp6h0hty5AW5Vj3dd5I89EkDc0D0xPPXePuSATyWd+WV6SKjE8ageMDJiHkP
aUUb3zh5nntpNu0X7/8V4oOhjj3RNpvboBap7uh6SddmNaxCUrJV5Ru6//IwYlXI
PrpLBEV2vWSYp7P5LX4fHQo8ndmMMEohn42UEDMceseWhpJYFx4Ung43yeAJ6YxB
0oWyqWjpB6wI/6VMdvbOVLb8Y0Wx/ghUjILoZtZ8gcrKRoe0KyQ/LDh1wk6MpbE/
SHREsBNtfjkYO/0Gs097j4bCNxReuqLjWJQ9OuootA0Pplp3ceYoCg8x2kBxN1Vb
8feF0GNNFzHwWeWk+eXBZSQUw5FDUnfiXYLgvZX0El1XnRGaYT9S9E3uNb7L6XTJ
VAFOhy59PP5w2qiHhhdUp+enaOYAkzvtWmenQvCO3IMHGas+SJ3WVF/zs2Q7X/2h
c+YL5CEQBToDzLSeDdeU+T/LkyUgEGRNmp7vQK3xLX6GVPYKQ7/c1557dvqaWzqh
4wHxVovB0COiQp4EN2gFCWDfsEUCS3AaOnZ24veCHzQtFFNw/p0xgaH/5bZp/AnI
TRz3GsYQAClm2nunUORD7sVbyRx748cRhZUuL07zSvbrSnTugTrTI/p6Sq6gKWPc
GXFDFNixqwcCnjGz8z4fpDBzfq8fkmpqYTvKXyanRufjTntzuoWqd8moe6khTBdi
2sWuvh3suTUZ0Q/Kizk+zzKO5a9VVhFMqWMug1xah7r8iQw7dh2hwbNGSKR/GFxe
PA7ZyqIDdz/wGuUoTabvFgkaSHWVDcp6Ax/+Qs/WDeOPki9tyyK04yPg3XE15Is6
Ibn+4ahis6gWE1A9Ywj8IiEGCVbcQOUJkIhvOsnS1JN7SKI+mtTiV2OlgOXP8HGs
fZRUv4q7F/sP8+Dn8HEKNF2uGxSZ3xlOoylxM9wrTHg/eu2fiNdcMsL0qgoYqieU
4ybelWAxGJUEvWotj0J1/6TQNUtt3Mz9oZuNq9+HD6id4Muf6Xx2VAp/Ah2ofG6E
rYk9NyIwE0qsGKWlOKQ1FkXLNH42HFdAEcNY4PUIS3dTSd2A4OJPMZizp4xokedx
10409KfJdPwepUY70xTBRe6y6uUIfKCojOdFZHwymKHCrDEsTrsY6DhslXk0z0wG
fxcPdsA0ESBd5thpiXEz8i6pfz+d5opX8PNJVRK7LWJiqwbbcqlZAS9cSKZNCNWC
9SKjEMyHEfaJwJF3MAmIvjH+dr5SD8aOGuPip4gpVkwSBjtzvaMqoge8xhoRE1qX
oKNkzxwo47rEl+j+ZDGjK2lMJGO0FHMQkZyB02q4N4gOyKcm3/fyIYY5JEEM2ds2
/APJvf6xcAemqxOkQ9zGTwn7tjBmM2gV969qiTHZziorF3I3cuoQqiUaOOGiI+yj
luy6qbSDJ/5oWaK5m48ydzCwr5vK3d/1aHPcptMXU60Swx+uB5MVpqxsaJ5mcyWl
/5qhoSbTX/Lh/Ods5TTmSjw7HAV1DXoGGzUR70bE+DGUmm6lFkr5+j5k3vQndfN9
zfDpUgS1jYAcOqQXhbdU8Gk+vd1XE39F31R7O14/Mv4kfRl7HQEzLJhbMbeAc5Aw
3QuGaYVXbJDZK/ol6zusY4/w59eAEEdeQQdQ1mxo9VVImbN7aeHo3BymfsPX9oUN
fgV/ss4GlpyKmjQ/t6FDgRV6rHCRbDWOwbUe60bRAfz1afHMYOopLC4ioANkf6/d
y0YQalWY+NODPtnwr8JYsyi8GqdfdhXSvA3tWHz/0vEKpm0D8qz2f5NDiWg0rcL6
UtR3hvj00iAL8zqVj5yQ09nMoRwTeoD7m1YbnbhpjRYh+MogmzgVL+l8QaDOuqRx
MmtiDKaxuBIjJqBmPU2Y8Ic/dj/J5GhvL0bu9NFR2ohO/ev62O74bfZILMj2RcU+
Uj5bD1lFvhEFIVvXB9Xa5pA3e+p/4xtsLQdT/aBVJfUiytih8hp7BZInS+TmNdo7
DkJ+R1NxIdNHuXa/c+3ddxkuA2R9trcJyYG5HqzmR1kHFQGNehxedSfpQJ0Y5tdh
DVOjDF0Q38eC+fMBwHtGSoaKI0p+jvsD32gsiiMaWIBxmw0tN4Lw4DC+B/1EI/WS
sS1lkis82I6p0DV/YXqCmNRa+gli3ciKperte3a8fbme/Dk5q3TOK0dVzq1VTI6t
LtvZdVD3c8LlgQr9sF+lI6IFZZnpMFXpJTrHqhlIgaNj7lrIR1leJio41H15OOw5
NukI9b1/IpDyI91EBN5vpF5Iu3zpB63vBmiXRErFvQPVmbDMAuq0FFg6oCv99EYt
VnzlyyVboMooI4Cg0ZKNtcJsRLjZXvAMp9w+SvVxnAckGtjlUODUhhauL2nxO0CO
pi9AVX98FmEuqC+Tq673dZmIKM1rVgecTS7OrNJC9hAmIoWWBMw0GJrvRc+Gwamw
r/iEXzOkxgJHfP51RCDDOKdFJTD7+SHS2WteuWecq/m2d6lmloxK6kZ7ouNoiSHe
j/NnxeIl1vSH89OxMAGdFfNPN+SBMKEhkMVOhAuUVruZKo8zWG4fj0g8hRt87Pmy
52KEgfKbmfUshXZtyjoVWkt1u7nVd6T21MdWLwZaopLXMPUJuUK76RMM+rArzB5k
YAE5f6bb3/akizrwxOtfXAuxbygJo5QgJOsefaHmgiS4LyWsfoj4kM+VfzUo3NlP
LpzvJEmD1Ry7qQGzeBBnG6t3utxyJIExhliXn2cstimEBiVc8nl4dX9xOdmOFSJU
9UTuPUV//R9egPVGQwpMJmb009tYX3bWIHL8O/IShRb11SeqUpXr8jBC2FjeFQvL
DFTK39waUIQIyFjHioDPMbgZqw9aBAf3slcTvdXvzB9kB0R/szN29Z8Xlh7Q8qF9
KIuVvELhXBvH7Jtrwzli6DIlEz9m0mHKmkXAIaasItnl+ivsWR12zjBlLec8urbC
nT0Jio2yv1cJUKBdLATFWD4kVbFPZ/AowTZkPt3VxksouANlouSWejlUVwneFspj
/fAZ7wCsEx/9TGLnFIGolO7sKpaMrqCswTuZWLGo7It3K+FohRMNSu6jytNO17o7
nowaAlRt/kMzru/Iqh5T9ORJn73BzN6oatgaifC/bXNE8oHTHq+lqXgoGoHOauN1
vYfRANTzn3BOtqSmyPsLlJRwyndoc2Dq3HpLEG868rInSPDXerF4W62tg760CD5A
Wl0DHzsz+qnyJVvB5yWulUyOE4T13oLuhydCpG2ygQ56Nd/rhODcG1WhKk5wdU+0
GvW89/rZjYc0rgsGGSEuq9Bf5cOlef8Qwuo9roeEtpLchej2tC0KfX+jpfS9eg8i
MVnaV004zLKiU9zGQjkMbZbM5c5Q2+5WVX5YSWNj9a3vJI8IijJIK8obe6T+/gg7
weoD+gDOJFhjSObMxjIu7N7KgvdcHKgUi2JXgFubeD7oU8D6xe/YgIa/bi1hzOtX
mawSaDxA/7JxVrc/TVCCPk4ub08iHYZ6fbjqUO6QIg2tghhmkqa/C4s1lDNwJ4j/
oCRWHZNwRrfR8jVIwNZDo+fVEIS35vm5WWeF8L6GW+PoKd8REJ48Qvjt0ovZtVtJ
2pChd04MxnGhv53ZQhDAlPJtwEiGlhrGbmU/41lXBLsSOdprlT9ZyA9UYON3rPtA
yaFj10xnqRyWkPYnIYLOnhUU6HyS2kV505njENyueysKd3DRQiVB1uxElhqa2l9/
zR12NV8KhVjem9yEywekDgACJ2/djCcxvFtko82Uz52BsBFb5j+AjrVMH7KGLfEK
JhsyD2PhvK0dzLkhBfeYOeNls2moVT9TSNrJRgt8Hyr6ymoB47LurfHTPyWM9eRi
6sT9EjUlZlGdEaq0StpI79ieU7TS4tzwFHKgE5XS9w0vftQK5lTM28J21cTtswqt
rYKD2N4BvHCirQECKtlgESkItpM79OAFN7JVe1JPO4coTLm/jk7bEePM1IMKr91j
qWjEmChDMaS/rYC0RkFxAmq8V4CbINDvy9LyB0mogtk/vBHuJAWUf1r5/I0xJg4g
p0RQdpgmlVC8A8QIDB3OFVpoR3LeGwbsHsawOwft8gByJBN6ZB149T6YNxUmJLzx
o0r1Gggyq2PwXwOBELfupiHSbzz0gUeiiUURPH+aSDAcHbXPDubxWmEIDahbqdXg
e+9qREugp4EFheVP4XexqZmO4KLuZ+hw/zGIfu6kgwJd/Mdyi+6HSc3K3sZcKcEg
FBRqgT09Dsu2QTLPIPT0zWwmUlFROANsUsFM6mrLhkMa5PcW3KsC2fq+tSXSgVg2
iWh8duKx95sp9r5nus2LiM6QTpydSEaXnvSQan0edi3uRUU86CDF85t8gbhyloAZ
LC0tZDFEPu9ULZuf+ZSFbKHn1Vb5cQD/rl5smQdggtN3vzInaUSO5Gxtl1+CwCZB
eXK1y6WmT8zTRWKNv4haxoAnvzjrIu+LNilviVRd4bBtGelzCyNZrUss/jGXccOn
giHWi15HosU49n0EPUIiTP9VzPaaj6gm8KvDoLM01yuCdbqR2HOuhyl8OV5uPLIE
J9PX4ypNCNQvjZrAHoh2C51goCFSGu54RixIKXPL18uDpHLYuvTp9hkVuc88b32B
o0OtLGzCNUnwsk2kILBcZlA1dCllKiWzK/J/bZAvhhPRxfFcH/Bto7XJ6GTV0vI9
0YJc7WlPqERPMmNYiRZo5R84xvMhp+mohOJ6BDnsHToqEe7G0IxBAx8ksnZMiDvR
nLp7oixVaxO6O/w+DUv4lwwnX+b7b4wwmfGxJNW6qoc9RgnXy7XIAX49dgUYVm2k
O5KPzwk+4DPH7tIkeaWR8WpF90zt3aIbATaqCEDOiYuaIHKH0LMK11UTrQSsHJvV
u1JxN318dr2IUAXyKbLEsjSMjYkBpnMA/1Y3j59PPgZ/C/oVdxHPK72IDdadoiQF
VDL4/t9w9dK4//dXhS87mzOPOv3U0mECLi/h3FnKwKiqqQKsbHlK6a0e/kzb7wQT
LcXRlEp8wafSGWCrzdUPg9h2lfwtib89M8WOa0q5vWcOUL9vddpOUKI0ulUFwTO+
SBBZESmSqOKiDnRj/bS2PvOn4I02FW3oUZOwI/OqWKrGz0ZUKRpTVDH7L/gxC2T5
nI7vRPjTi84NSD29ec+4i57UXePy4bzUmwgox6ZEBrRA+3kC5DZ41AaciFe5qNox
bNQSqg3PnhRxJmu8mf4e2P+SOkz/Kc1FehskKN1XhlMQYtQxBLty1yxWldH7w/R0
ADfuhFvHeAnmsCQVPNr5FIqDC7mVobxF2Gq7gxMENmuGKXS3gXTCttJYkJ4Hb3tw
aHWFl0K2jpubqudYnU+0s66vE3/5vSY665wx9YcbTResfbGD85GWE+C4WQNtH/XI
aoERuTWkcUz2CMs+w827Py6vWQ+xk8lCDLMzqXqQWNKRO6VE+5C/zmgNe+nkqvUC
281n2FqmB5wYE9fPN/VhXxXZhSWXPDFZIrLCEjsw/307vXeW7VNUp890FdtA9WBD
XrgV+Cg6uQXTa+RoV8yWzrKNPSOA/bznPCiaL5cvuiGKdBDejhR3NM+DxdEj7SqW
USvr5EtoH5Vml3FbFHQs4eZuUbz2USxDhxceGrOfvVjkTUfD7BZnkf+fLe3C3LkY
MI6eHl5y06QoZFAbCRcyBKJYDXFfPBG5wmjyBWocfrIabWSbNPuWehUasMC9umKJ
E51BqY2O5Af9WUP7s0PfzEBy4rlWxeXtxvyCostBBbn2bXLhdKBK/GONVWdJfbm0
wfy1RmITjCOfTnefrCtm2abXs8hOETZsJbiVVreplK1eXn1UYN1eByBcK+xnFWK3
oxmO6S4xI+24PQ7WtERzBWMOVaDFSKaETgPxk3lSlLG1oqfZXRgIeA0KQ4ZokDVi
+FfEgx5n0OU8j88/u7PIfXdZeaJ1D/Tml2Rd16nBu5jEpqDSBIoSX9EhdRTticpc
/hc8VNJfcI65k7ouAwKLf1EQbpeFWPFwio6iGgorEwiO6h4juNoQbTN/uk1zVk3d
sSJgkHaLdmzsWtDT3nOSvS/ZyL/ZQ+FInHhg6+Q9XhdvQnixHeN+RlZeHOOERwrv
PZGRZ7bYEFs1Fx/NAcDksi0O8PsCycZZOIYZ2XXb9pBwhKWQsKHrafZsVv2hQpNA
I42ub+rfJAM0fk66Gy+bDfHCv6OGpJCDKzcZJhKX3tClPeSSQOeuvREyBnEg892E
2ZvawVdTLlJy7RmjZomVlzIWwcBccWMLPbC9Cdr/CKELB/HNILhVx6ZyOEKyT2nd
bED5YPToRPPYAoKJWL3YTCWtPCjHJg4UYzzlYjRujW+a6BYQtcrwXq/cBlfBCejg
cZ3pXC6R3IMEIR27xvbmpAoXdjdpkW4SkNtNOtlwTo/cHOSfyZpF7uzICb5bXPNk
VQ0xC0NMy3apmGNuwITWAuiVvWQIaDvci4uOGuLIQ5N2S8uXaNRE/6p3ysIoArKC
+9f7TWGwEWWc3y+fi+B9OfhZ3aj6OvL/ThKh15IlnwpuUYKDmj1ng1SzWFwDgRw/
qfbkAUN0x3zBhh2Epz9ajnhxEkJQsxK9k72kZV0dRZV1+CZBwc7z4GJaN9dSsw13
hbGZXvXMc4jGU/YGZxNtBx6UPpnc978YtLsBTlhxAfo2X4e5k6jCK2t94IxaktsZ
jSjYslyjlCVNdVXDHDrzhKDDYQBfVQk3xhPyBrWOMhm/yplk4XYAvUym2jOuA2wz
uhk8zbERJa8ARAQ+V2b7zoEvcz96PubVzWVubDWxOf7T/YyIF0A9LIRgffg5HEOa
N4DyrybsPeHmxE3TmhAmq+lbnhLLnTxuhy1XksS6XM0G61hHaMBO5AuMdHO3O4NG
jCElJK+yO/WPeIYGunDC9HR+YQ405Cp7SUknKB0OXUV2Cqrfp5pPDBy6ZAJI9Rga
2UXDw+J3a7t/zkQZ52qQ8bQjGn3IcZWoxogNaNFRYUN60x08L0RNt9hQqREYrXoy
ouv2NluWRa7esHp0HQ0lu1shNbng+nc5hnzc9Rl2msToVllnwPSlGiMGMeDhXpkS
hKRks0ZtsVKCl/QB0eX+FMBFCvOwGIShipsHk1ebvTnmaVM4pRLZ1S89sDVqHD00
XjpStXaxLrrXXiYJb2ZwqQzmkpK0f2m0fv0lXvLQpzZH3RGFt9EYGt/b0jhsbQwm
zKt5uoO+3KrROgl/sHp8mGVvM8oI2imLXTEH5ONNHkPrMAFGEDSb4SmL4ItxK1dk
+9rSZ/L8hPFQaRY4//MQgWWyd6OJuxWg2Ol7C1an0aR3WFJwZdYqyK5mQhrWhOtV
UbKN+Bx1ypKV45y/M4I4hy2cNNCja4C+h5gZtZc9rOfYmHDMCw1HC3ZAvz0Ckyme
EgdRvYskq1Ef1uDXE90Dt3Fy9gQkeyUOyB3dSD4uJoULbtxcktml3EDfBe33Bv9X
k8pSA8uVSnFAhDqApM4tOnhvp8+cXbUvSTXynlNBNcIHO/ckwDalAIU6s/XCi09q
AnWudQUplKMRWy0tCY6Q/3t458Ly72OyHeIkfgGOW1IE+CauAf5TulwOoErSlfR8
F/vmny5Q6QBg1dtUTqWE5BOhzC/Vx9WCY/tx21bbYkFZPcniiAP9Ik/Twt59KGBo
cEpS0ehzZSJ2o4Kd5LREJBLcaEq/W22V4I+93eARzziH8KBskA3+x/wjYUhuKHb1
qL8oLZVHnGztySB0HNkmOoiZpk+tgvlb3m352KuRBNxlTnCo16BOcWf9PBT+351p
Jrd2ROtsw3ooa+E9SfV6LoJJjjbAC3c9TCr0DMT3gbT8+hzUM//OYS5IUhdJXq1j
zM8d1HJcaYzYPzlpKr/+BhchqfiQAM8O+9V1/k3vJEAalGtvH8KW0u00cC3nOgRB
bbUnSNk+IzfjwRDpUzjIavJWqHTcfVrhZQrp/XhUS0I5f8xAVK1zUJXMoAx9Vob8
BtO5s6QEaxMJ211L99w19HBkcYWlmgzUCWcXf0WqSQcKuphjBnfWQLCHKhvcwrLu
BfXYQj3vCeZ7SgFs9++OUFhCFnSiSqR8Sxsx0ww0f+wnPCIrPfZPW9ac9pZn9rDH
M5U6Ra4F95TFkZm1QXr7EW5h4P1hSSRiu/zEhGSAFji3M7x+ANsbRebRUWh1NatN
+iMgI8SeHvJbFebTj1+AyvaWBT4YHh5/E8PWUjWugr1M3sNUxZKA+5d/kOch5j0w
ghiGI6aNYm1Fny3phFEzWVtobx4MMhzJD/p9TG7s0iVO2nNiO/BnolI8sbQi5BZc
KHZJnA4Wk6qwi5OeWqqYtwtdmCRUqsHzYTr4/MXapgbsTPo/7eJrY/fIx6vXNbb2
9ryrWNi5YqEM9OCpeBUCEwfYsGdAiycnV9L0YxBhZnsC1+ogymxcBVBKdgwWbBVM
T3uqngPcwKdLV8JjORUdCynNEd4tv7tKN5uyXkeb1ZQliQOtECZLK3DDPpoHT0wX
Up20Yl4STu65nnDd2+JFiuyiHoJyGG5EZwORMKWCXTizuTDwZIpr5OptwxFkHpFZ
HPpOs1g2/DVdfiK1PbXUH+ph9s1BPiXg7rEHJS/Qq0kiqb/r1Wu/J7cwjaQ2zyKZ
6CN17t0QwqGWGilNsuZox3K9YD89C+zwc8TEoFOC0SHobAmymhWNmeSv4dbf01JK
ZgljzmoIXsntnYsTdM2lNLMmh72eXD0NVxhn1KEyjdBL0YsdOQMJ/zPrOvadn+ql
UF/liUySPiiqbDUbfjy2FcazvAUqzzk42VJSO4x5FulDIfUba3bEUiAjfm/ktAfB
IaATeH11OKepLjZGC2P1AdA8k1alzyuOs/IGbLZI+E8qDuVHw2Rxq8Gz7ZwZni6c
JYK2OoiSi/kWGiEHEvREpdUkwiXtYczowLZf4tAOwbZesC1EGQB+8nFp5pTAXzdV
cjhCh2dGeZ4Eg03pf2MVbshZWfk0e6CFEV/w9KxOlfCyYQ4xMtbSPnM7200ahWeA
S+fJvCdu1+0L2/KwQdhbJdQUm95EwWmudFOLiwDeVgbeEKZ2cUwwZw4w+Qn6TUoZ
aoFFsFKJ/5vbAO62imW6jvR7AZYuvrhhXdqp9HkOVkhaI9VMS9Gf6LfQ5N50CD96
0puPdHlzmxGFB0M6cubOpbM/7xnV5aI1bACIRssDLo+0mQEg/Ro2SmWLRUlwSdBc
n1gOVK5I+NcPWJ0t28BFDhE17lf7mSo0tgHYeww87QSLIHfnL4gBV/Lb2Qwt/Cok
m3Ah//SjVxm3cFQd4vB516OBHzKeAvgZN6DMOSQBgJXwg/vbRQh/LHu7Ec1XBHQB
mAlsEhPWjpBU6W3vXFSG+7nXMCrcd4NWs6Y082PVdThJzkuUUWbNePEKBckoV+CU
r6kwZRdKds8w8PNIctSZz3n6RkOz2edtxcWvTJTGrlUORp28o4V2htiW/oyNj1y9
AN4N8wYRzSgcF9DfByzbCLB1ej4TwhHjkTzXLg3pgluXDUtcxu93Ni2iCYBW1tvs
QYtKXgNFSa7McUfR0oxgloy0Fj/2YCt+hajpNcQQhUIQDq8Uon6HPim7ZxY8dBzm
U/cSkX6ZPuWvTaQHO2W3xlPbtHFYQZvDu/ZDxWBcx/mPOVf68UVcIkaGfV4DlWNC
QiZOmzwm6ehFOofXCQKf6l0/4XSrsjgwPlff8WPdXaA7ZUF+ixv96MZ+6K+wO7st
Om8/y18liTX6ElsPFAtE2VBrsZ6Vs/aVYJ9GtgNSZ6Bi2jKruK7CqS3s8To553nD
wRky/xft2TG1ykG/ny1ZaYi09xinbRukMWGD8xPD4qIfFVnwTmYti93Ll2wFA+Oy
aOdkN6G5obWRo6ElHfxxFq/yUC6CO0g2xzJAQbvT2OzBxjj18AVXswmwNV4ABXF5
DdAEZplN13WlVgjQGSCTIzZYWqKpjln7ICvfO8whJbxvZlZ5Ce1En/al8gt/8Q0g
d+zbm4tEB67TzMtnKEHOLc6PSHsxM99tSIaJ8rZRD6hCdoFW21e0uzigvi63h4Uj
e2H2zJBwfHO/g/ezM0RefTTUAgeTVTTBSC6nA53wkLGAZO7ZhfVOBwBWiFpSNU/9
WpfefPadd6EA+IQMU3PKJg4HOgw0F8Al5z+ndAwEudsCzyjLra8VaWr5QMRpA30A
I/+s02RgmlJQLu3vi8XEAAcfUVZuQgnbRsMlV3lwUSlV4StuaV/G7KFSQRnz0XVV
TT633iM7fmI+ZbwB9s/CYq2ZLYfslsUss/1QHNdDUTSGQiye5tLRj+JRZJK3Vf0F
MgJmouAC4MwudjUpf3xCi20s2BtJcLIQXs7KtqcuEcNYvjNliMHmsbF6/MAtaLzC
3UURog8XLVLOrzwjzMrRBiHj2xutV1JxomeLfBzhY8ySoS2rRLnxUPDw4OvqDFCa
EtNASUYTru6bsBP/OLPwgDREeCxnHlnQtJVwTjCvyuHlQe7gxrxbZncERsI7+G4g
q/gKHOC9teJfUVxzUjIu0YodHfzqKdlLFD4wvK1FmW+oyz4iFTjHyntJoTZ+dT8t
wELxyds3nJHYswgBlmTcU+mjKtoBpkX+8THkSGfFro7vmzyIaFU5FlXtREQxcnNd
du7qR1NoahZ9FaBRA1EMTB/UAg6wILC8kNGus0TO4q5Y0ecWYSS1iLV+1c6hyH0D
CQGLIz4UM7Ci/9cme2Yd4hHQCnlBwYjBB7lv/uwgneDeJYIwKNvKGhfIBrUjvnRq
5H6/O1q3Elw/63oaIfwj99kprFMvlTQumnJBbdYDEjFtR8l3Wtr54wUATWzuiCdl
YFmjMQWPEFpXARvQ2aiak61SlUaQNof9Hk3R7ec+Oylpd9kkMGw/WocTVegAlJdc
jVNyeoCgrjiU+s3Ay03986RiBwOH+myXR9yBR5E318TBka0dBGHR2zopIMkr28OA
gxOAs01lWyyhxJKLduojXwi4cJoEI3T1eum10bW/xeW2lWWry8jVf6PSj2dDkasN
vZz8SWNfZj1gx6Q26zlce8Hp8gGLPnAI7KtvRBx/3TDnEsXGh0GAY4oBfBRnmTIj
qMBydPPb7A7f7hrOpT9nR4O22rBQ3RE4xy9+oBfK5RSXPwOc4hsZ74DBGAdL5sKU
4HxjKDXUoaMFWpL5hHsvtj5b/FXVsgvU/ykGtYrFgAX3wRskF1WbLwjiR7/tFkxZ
c8F+tqc70sVDiNrDcDQ0SMjCa0Wy9oLLUfLQlBlX+BokGsx3/rpcf165INePW4ti
ZEg3gD/cjcDzMeUcBPXpoz0b3INpRO3v9i5IXEodwdTNQMnigofY1csSlKJBm7V6
SX2CuRef/pclIBa6wUN8JpXeO/4ZWUSqLGxsvCpHuezHNwQB2dOpD5Ycl8nsoFxD
zxuP1sQErXH9AlDDgiu13N+dAt97sFMUTDiOE8OJxvDFhPg8BiRlxh0y2PfgXzLH
CXeGXnhBVv3jis2N332FPoLF9w4nD5AlGQULut2Y8l4HP3uItJI+/7eDXet0sy10
mvUhrvgQre/3YJHds7zMp+/2Mp5Rg9IcE/Nuhbx/n1dYBK35nbMcazIvqfA3ck7o
AS1BI+Bt6ApRzM5kvlEe6aCNWQur4d9wmJcpYWPZRnCY+jLsDnSMq4ibYfs4Yymj
Psymwz4Db8KqPi0illr1xCUumnq4nsron2O4L3ByJtw9s+vrz+QJCCWjH745EVaL
YGw0n2nEGBDuIUDKsVmcQelzDJTLDTt0916N6/wqiSYvKkrdQ8jervq7kVtwhhec
zsxMW9nDhA7lpWbg0Jnm6ksIx8Ox2yFNJT8GRcrsXy+Vh+p2UNQnjhUvN2DLsurp
6QWAnTlJpxohlYc6i4wVnMWh+hmnofz/mRDcDB22/noRs9s/dUUpW4Juk7mRapIs
sLvV7d9Quw3Xd+WE48+YEgPxbK2friiPMSFlbajU3wqw6ngtBUO+4cSAPt8Cu2SG
oX0NBst3yOudCXHlvKTXyZG7ZbJ+c2wUVNSwEGk1qO4uWwDwF69bPpVaw3ds8Mn5
YadaleWr85HsQaJyt/PD6d08mdXWwPCi86qynds4I7nvezntWWosh0amnmFQobao
PUZjb+foykfPJ+ABQJLTYB08ba1zeRLHPWp035fJhd7ol/ulpAZfJK5gHZxZAeo2
57IOGaA+nbZhzAjLZZ7NqTYVuf9uFfae02GX9vXzGbda/xTnp31qkHShs8T+WWXx
k6jLf5Nu9mPiVkm2OHbi6pskvWroXJ2PVLYZn69Fq6vUko9JTzH5ZUiHZaw2LH2E
pf8wxTL8y3ishssJUCGQj5CNcu0HNcPABjY0DduIcW3202maE1sQRBftzX6slo1I
T5ToIPhqca4az1mqQl3yyzfJq1tEoKo3qpXrEQ/Nt0kNAAFZEnfiD2TgaPwsIwzD
0GPqvRoccv5rkoJwC7dOR9g7OPs9X6U6zs3NKURgamodX9p3BHslSIV5iqls56cD
1MrhlKi+hqbEhLLc2InAVUvuxyLsvotn23yQH5UPMh/bJeUJ1MDKkCp3Az1g1TkB
Xx3IjeW5viUaURwwGVhoVUAEuHn/WSFcajwX2mi5c7sxa7AQoXeDfjHp2m4WLdh1
uY+VmJfU8a40hQineICNSQsZPoXsObDCoBRruQZPcSypBQv0Js6heQz3/wdZpPHR
eav89Qk3MhD8V0AAhw7YMeep+IIBmtuE1qrin4pbfJ0RvC8fID6NVm/vVrDd/1Pi
NqvLMHhhscqcpNVOopFc2qQqCs3y0ymM57pmyWd40MsOjHUnQBn4WZbvL60SlL9V
o3Z8ZtpURhY93JPc6/T06j9Q7BlIRyzkKY3FvHhBwn8HPs4Dv0oyUmxzezhg2UVJ
NqSa3Pd+mhU+aGDGwxoziFavpyC3YY3q6SaQk6vYnSlhGrdeAq0xjRkRHiwd1ldP
0T8fuZwb04NT2D34NjfyN+FUDc32sSfy8283VXVGCSCdHY522cl+7nC07u/qJrn9
6qHOjsyaQCBa3/9IYCeM/7Vwbs+GdH6UHJH2Y5LtXOOh/+JQS5NMN6v83f7Afq+J
47RjVTe+ThXEqIY5D0jtTBiCcT0Jeirt2+goVUXU7SGLlxQjq9o5XnOMt0g+HzgK
5BJrmKUOSIsSigBblY4PFMHSU2WsgET0VE548XZ96UHfFsFoVyhVj2h8Is2a82eC
VS22X42HFlP7avvlyRAlEOCC7Q8Nz0Fxgr152L/2Va46to6tc3I01nDrHaTCZKH9
DkMLZxx2tNDMSiERgaHaV+Oix4IXyQrYYMZAYnOA4uETS33kNnGBQGAX9AjFNO8X
7WpnONJL5LWCDLq84GZChxZ3vDrQTnafkA8hBs+4AvzQjmU8JnjX7pkeBcomi18f
RtrbWjjl3uQgHkkojR6gFVeqQrIx2hbhdI5DbiHbacq2aOQ5+M1VmxIIYTe2oZYB
sMbsdwuj2/P4OsrHznGNoG94WsBVYdbOLOBg9RJFtNjzsyKA20R/Hx3GJPWiv8+R
aDfKKQrJsSDwDH9HYB2kcqmFxDX5/zsVqnz9cSF+sXmCqCBhyMF3xDQgSOgV84Xx
YDI9NNooNI/2PYkcCnYQrUPxICty1nrF4bQalObeKcisEEtGMYlcp7a2T5ARcVqu
7UEUNXPj4sHTOt0O9CNCxgIPuco2D2geSe20gg4emxDfAv75z70Rksx6aE+3uzLs
IriWyqYsO5sfqRlA8pxBbk5Ye0eG45+0xQlTdlhH3HskHzw8khbAQcg6nMsgitd1
K6zm5XITM+7HiR9s6FpUosXQVcnWnc8KNVGITgSN77j2vx0WEtkOIF6NovcPKn0s
nW5nuRRLB4RsGnCbE19CEx4Tfzp3Dp0Orlx2uVQsTCU6ByoGALZAF4nAUP4/zZaC
mNWmbs+OerWb91TSSxyGUDvS7NF0ywNznn+36pw0L1d6zs8S312dDbFrx8Qrmxq+
vND8QjiEgx2hNEwwZ4tBBodmrWW0HyXw85ja0IcqE06gvl36/xmaa+nyIChvMNQt
Yz/xJJUchlGP+Cw8MUi/GBZhb3a5zZSMeQcfJQCZsEnM7b9LpukJkd9pLQGiX0HV
LaqMgmra5dyvXZqMlIQLX97r6+Dg/+72GrimBirp5aQiqCmUUvm9Jj54YblOtA7q
iNk1LAXD1XVA1Ud6kijTjR+bkyPe35CIKayEU0iozIQNThecDRSPeDjmDIDIsQPU
oVrIluXbDQHW3PO6pH2sDQUcAMfgTrmoxbT96npvXL83S46DYnQy4Cl5ep8a3CYL
1cufEoaB/YkEiuZrxWiRsmboqqLIHHlZ71Elee3t8/xjvGcfxTRW8yMCcSlEbRwV
TV3Q/YazCg/eSFbN0bHx+XgNnT3CJokcy6d9+1d6j2DKC+mQ/P+8w1rqHI5WKyBW
P2CCMUvo/6ck+GxU9Rt8zGQ50pagg7Xkl5q8olGdmCDo4LjyIfFKbQ8QBiUOFpli
eo/ZJrAgMl12LuiqH4y7Yu3TzX+88OtItTF9Nmkf/VHK0yJaB78XxPRUFvo2VfQV
3dUgz+/hoNtEOq6jnNvk/3O+xIM+csvs3CvTZQf+lwKS984xsYe8EdyOoyYkfnz5
TjfKneeOAdq0jPzSw+1ikyQGz+TVacUTYjcDZd40YleDypc0QJqS8oygFDHMmU95
uHtYikxtAf2qu1rgXmC9u0V/vM6uGbSx/a+G8Mub/nLq0T99DGDkTBpOy+BXv3QJ
WQQwjuds6H/Y2so8CiriE2PVhJS8LOTdtzwuD5gHYM65al+SKzq9/RhvQFreM1Ja
R14LdCHNSrWUqbpl2HsPond7m2DTF33pZhQaslYKbX0oJ6id8KwLnFfJUM1ap8Ce
svBp2ft6FfjZOYE0A40IH8HYDTE5fIkTtJCcjB7hkPrNMMPrB94eOvsaMIB7cTEe
KdsMUPdGxzOenVK2CAp61+MAy15kdMa/LwIcedBHViSIam6JZcp2fgtbp4XOcDyX
J5rr2mdzzEs7M/DuHLAklaCpcwv6ABZTe75MIyp7F/Tk23ucZp5GBoa6cN+TV956
SF9ywmUSpnDlIy1xaNj4cByP3xDlVSVL5wukXItFAWR0chEm3AHKGsuvNsBzbm/C
D0M/cgZcgZ2ECYK6T23IebjH+qQqB/8bOtqfh+zmKohP4OQP54x1iDJUiPO9a1OK
sXynbksaVMup26qsziycf8RSjyEYtrHazIPnJ+YDH0SdU671wNvBmuU8JS0VUkgs
pUFdm4aeM9NAPVjkxcnmZxbbUFRFPY76SNZcSsgwAtvQhHBq1CCFmYafsaVHTllw
nem4jptkfGtSZjjM/u06HZoiBE4H2kHYwvnHfj+Q+YrkuNkqUIFaTWdWFjkG/Iui
fjIKbZV7bktO/95w6Y6RFcAOHQz2beL0vBvOSD69PS+9MhhbEPTVFgWGkqSMkUzH
1sj2ppUHZtvMk1UnP7zYNSLAHrvh6aBwSBQgi/Shqm143oHXMPFbemfBjxOtIUDo
LIkGE8vJd5xSxG3mQgtH7RbpOEibAEU/XmynnXO0KvkVpBmxX4CTDAQZYuZyawEH
AZKQNIxTOau7vzLXgKyOX/aB03MIsO3R9bzshikgyvWglXSmvqLpI4XcIi7IilkF
Ml7Ax5XZ5XWx8fGH9djC025f8nBxh51cLCCHGM8pGOOb1oCqL0xmhxVxinA/PPk2
1w8oweaYsm38HCfCljn9bOn16shiLxdI6/Jfx7JHRAwhv6LQBSOAIGuFQIbztawS
uIbi7aD6Sw6Ws9SkZps6mP7aXiFBpsORe8WrGo5tv6BhedGU00T8txHCjrLCeK8r
sgtEs5/eKweLMCZqA7KI5pSNjhHhY0EM2gdJuiaq2htOBeUeX9ZJW2Q/+/MYkMvG
e+DDKydZbCDIgy8gsb1q+TmsntEbCpmwDZPj5a/gXUdL4QW+kN8o2+ae8u7qZ6jc
mEm5I6R94yFnCEJq9xD0GYTyFgFgz3ZIcBhNVzcDbrm3e7lezQQZJ5JPftfVIOik
UP578+pDanbFW26ksBREX2lHxFUxSnbnEtGAANlcJITUiLIM2GKxCNdpxB2jbQ5P
M8JtT7y3HWHY5i2+/eFIyBu4OWn/wkPOWoPuUjORW1Xdi3iB40j2fD/W+TXR3P41
wKWDilPuBIYBPTPP4lN9G7G8U5V5DGUYSf0hfS1OfKtZLahvGYNYDzVZBTKUpTJl
Uz5sr0Pa6OkDY9mf6z72ztR7x9zYh5z8q5UOa5GUgfxdSGZxouoT5nXgh3uBLVNb
4+e27+/9SlKk/id+byxyxCTOAVXWqTU2e6CqEThZV5DLtbbRPEGWIwppoEkA2fjm
63f5WbC2U4xxDE7VySIDgIH/bx7fE5TN4Fp3amAUFOh4v+hUjeIpjpvAmm+ll96B
Lppz/1kDHBXZosUQb1dmGSt1pl5lNk90+DL3e5aMTyr9piruyKwb79h5KnSfFXEr
9/FzkWTSIHlli9PfROFa7Y7YqVUPBD7wOGuZ5XTTKOLX/x3bpdtrqne6iQfIp8KT
IubziFBsTcUnyr8FMU11mGtlhQ2EgD/dUOJJpCfFEZc91Gn564opj4xQaXgvtotY
dnDgVh9kimYA9ZUWEgwgN8mXdR+SjaDrGQyGvbXld36bqVHi/mLMvOsh7/Fz88mU
X28IoqsCIypA4QKDpT2PYUL5Wvg/BWTs64JT3l0E4M2ZXwqVWAgWpGCcCJtTAYB6
BCKsuelVzw1oQhatIVsUZJphcrNr0s9EwtBBM6EDpoxt2DkuxDLxYtYIUfL7STdq
b0rAF6vYIqncmweVPvlpEQQ6bGssilcj93Ed76gEC7+7Cy07b8P2znWUEEEOsch9
lbX/UbKnnQNf65ggXN9frEzd96DzQ+XQ7mlLSBOKZKERShobCPdskRjQO9PbAQno
XQ8N4tGSb8r73JjBk35NRV5gIWj6VqQ9DJXEqxEY918i48f7OOgTYvZsw3i8iZPE
P3iee9KH2rU7v8Mj6SKO/K/miuN1TC/LFz8GcOzobtRqemI98g1Anxwj36L65sCa
ADeRvjkmKzgI76EMLYyJwf11dzA0xLujBqa6rbbWyMXf7w9vECuHQCbY43S4Hkud
+vMdbaudVdAZoLYJS0qS848JMUVYQLnjTvdqoph1yFnlcFTsYN2o3HoKywszkJqY
600MqH3YusjiQYIV3Ze+QbNyR6esQUm4u8QRC2+BU1fE+JEJWMrfXb0UQTab1CCk
lC/pFzaa0qjz0uO/rGZJAqhvVtd1WK8l466cGnOU/aM0f8F7Cuw+uB/doBY+X9pp
4jMIVcHymho+zrDYMhBFtN1L0IZEs5eTp3kIs5Bi3Ktg9nv1oU6eMykKRKxYNbdN
TJrwxc3JdXBj2WYqVC+m1TDXQvpO/4RROs6orvZ8jtWL4+M+pdnuAr5SjMUkesEs
1jTSW3fSIGBSGhA16o/TcDg1KUaz3AeIlFdA0Am+kgv6t4s7tIi6G9iArDJfP6bI
a7N7iKhsMaUXq3dB7LjMi9BSAcKjzW6hEJXvSJ+HLKYVV9RQszpIjnzVOKzqSvl2
EOndJiqMQ7GRGgoNdkOYyIDUKvi2h0dqOkOnBl3mFn4FetxFqymto+z539v6//4n
iCtfMSI7jiTGTD0o5bGtb64kQPDO5GNcCnmTia8CyqP1RbLud8CnLz/kTLWEwFam
Wp6v0reM9Lk5Rb4D1EMORg==
`protect end_protected