`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
ddtXksX2+yylW5zu6QL2Lhnb2d1sD00763mmSITNX595NcHTEkwn0zB1Dry37fOW
FufOhVzEJp80NC5qZ/+F0Vk7Ik02dIR0elf3clrjeJRK85K4e3Hoo4xn7YbFUIms
l/8VZSb14+JVGURjfswrIyCUotIzlzVYZ6gzoZwDXIi5gQIBf/gI+KxNXPaKV+PQ
Ufys/12rjO6aI/pPlqSm0hCvftmBcnezN2hk1UeXgOIuKZnogjOsf0iJVX2aOOWE
6pD/psybjbnsNB6kH5uFTA5frkzIzkzl5d9+YDm9OyC+k84E83I/7/j+rk4L2dah
QJOvksSIzN867/4Qt8qYTQ==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="MvBXkzurAa5VTw+1JJ70nePUfoQXBvZOku/SMmg4TwQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
oRtzZL4VJ4iwysPsC8SXYCzXS8Fw2gtZTOskLcDV+1B9Nzn1zTyNtlo6lNICRmmK
ZRVu2BmCc2G+fmzynYlNTnSa7C0Cuel6FYpxCBlOuk3OF2tzAmLAuDyOH3Z1Yjzk
a0aHuoCdIRKv7BrZCdALt03JeUmXKPdOmIlkVGFl8yw=
`protect rights_digest_method = "sha256"
`protect end_toolblock="Jn9CQpRhJt4rnzZPRk+dOpzAubz7omckX1MrFd4p81o="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 44576 )
`protect data_block
gD6l00tciPUa6pDNTk/+tzLxvdHE2s3DQL3/JqqujQBC/Ei+vcAB8wM3doqg5vTg
mdfn9XB1bLOis2CVSfu295W2DNwHfMSTc/8BhCDRnTlLIX0UCJs9Za0+LoM0rMrV
T7EjVWppbP+Em6PkVKCwlmIQ7JKaifJ+Y+kjw9HCGboYo5074hY+K/CBbfsBQY86
DFekqOo2vgag6ud273wY6zuCqJxhIjW3yna/C/bfxdMe7u2fPOuJJsGX2edP+NnI
28pnXjfdSdy5Qu5vQ2kUAB/yuIuy8Wtp3rRVGrGRIY70F1JSxiy241uzWgEPLbQF
X5Umt5G1/dcGMppi8fXFR+croVFHLyC2xwH2F+EiIKg3bVCzTs8LpXNRgU9Q+9R4
4TpkMSg4bNgfUt+ALEqaUiS+z9mSDRKk6nAPblJE6rWBs063Wa+c8EB3vPk7cyv5
j3TozAjjpm1cbt47Sfi9lxlG/uOxLP11Go9sUdkZN0nBRDrCxQ/dplueG6jiIsGv
kq0wqZic52qdxNkPX8Qh9g7FToRvzPWInKb7Mk4n+SVrcMHmaUOiOj1lY0GSy7ib
hbihjE+9xvEFTKAMJb9noIrvTgzA6+CibDgvGv6cqGvuHVQ6AgB1OdgeFG2NMeBM
qW1omIMHVxk3fOAsx7274Q6tKAZp/6Sds46eC1H04vFBPSNjhv50iIR7mE3uVLRg
1Zl5iTU3BIgPa9BQfHX3IDpvHejcO5Fyc1zsTn702VAezKLq+k6bWDkGh/6cpeE4
Xky8Mt+Cj/Uack3XZSA8FmfHSBgpP4AoQwvP+ew0h87criD60rZU3VnTw77znFOY
RYp5SJC81W1aGvhUYxSIcyAHUB2uO7rpptch0BKL1zU+SOviPaT27HOblASCR4Jp
nNB5IlGqW1hZtN0u6eOvIM+KQgSRDUF4XMST2Dn1OxNrLPuC4jYJ1MgQ4KrDAMUm
oJMgoAnyOQfW+TBqcOEsjm8oWXkoBS36Xap2h952BZaNbCmsjQVF80ZnGx2v3kXk
aHCHhYmrA2U7fDCcFMMxIKPSRAb27YraOIWpV18XvICfpKK48YYcaXo7travG8zn
TQij+Zid2GL0D1akPaac0mZUtUgjoLz+jnPDb3kb42vYU8y9rPlEtw7fSp6gZHE3
nx9WEP8VO/utjvqy8OppV+xzTLS8M494BCBWreBAWz943HumBO+79djo69zyCGt1
ptxLq1yvDarBXCIbL/EXbpZvQxZ3fo2vnvkzNAHXZnpxHsJUYrYS/ge9f8LE00y2
50FSjOha4kI1T4p7z3xIjkWhm6reE1tH13mjN+HTLM7Y2Nwur35B0BbqGOdwcPdU
FDF0uWvV+KjY2oPVmzMYYYwipPFKXh2RxY47wOtPjIgBjMVnGiCCMJwNEH44d9WM
ld85fg+RvwrVeAoCO9tQIRsM/U5P6SxVgd3dKaVbdYhJr1ivcGAAoG45b7/JDLI4
gQwEzQd0c2vbMFAmKacYjKs/J73T+NcKBaZ2LQCb+rUrqf25zDWwGQOQJ6hxB8sZ
BIWyd22Vitpl7dkIO9jEJ6BD/pUzg3v1lPSLQeEITr1tiF71AUEeNYCAWiDN+PCa
/Zowb44v+ts/+z5qcNevzpypiwq/6aUlBKJRn3lK6eX3xqQyQSvM/s3ndoLHE5k5
VYxtNUiI/5mFzRa5+irYv7lDfZciWuVld4/RMp9FkGB3WSZe7Do1JOF7tc1D2C+j
NSgvrdsF+8k5hmdav9dDOYqBQ4mUuCKqRl5z9C7Uo0fKsrzmqHo7gXjRMMMIvmUJ
zm65lxUJczDKNm/ogw4jd7MtM0nK3tlcCQZrvIY7tZFXWOmwWOv4ka0zW+SKYotY
QiodI1PX+9d3KTHSGHg9UPavOrzpCD2M1h2vkqxRSc/7Y02+plsuX1I7QOOnmie+
NOSe75cRQbSmk1FTijQRdjlSZDEnOd9fVmALfH+6riEjJ4Xw01KEpqdPaHAG5DT8
N+kD6he+eOHnAfCCPplRl9zC0X3NJehZmfBEUZY0prKncEK3UZ4L4z56kWyhmcwc
7aojcF7wDPpWb9OAFc19whfh3XosyZcjln8Wb0kLJot9EmGzsAhVEN/XGUI5sRxA
1/jTqgn38AoPEsW6eHvQggpCRQPEch6Kr1yd84ZqR18sEAfY6PT59oGQuesNFq5q
ZxmCj0OYdJlagPo3u12gACejIJddP8j4INsjDK3f47kRITJFIOm8BRpT9NqQpBmI
9oz2vEXb3RmHcM7KegCbkHXYXyzeQ31hb0mlutVo/u62S5orsjJRPNlHdocfBfEu
FAxj93tcVsuaIq2DRroyY+sBnUFOt3Bq6B6J6nWb+/2USZjMQXaHgfVlQj24JU0j
C5rlML+B0InnDtNsEl/RZR5pYhz1J7RC+dyZ7Pb90f+IdYmt8nzv/hQhpF+QpvQz
JyZsrcaZ+R4SDCkVPy5KC+ms7VF8LKx4VT4f3ozB7EDUA9y2OntJkKax9ZUTrFxp
hgPScOYwt55SQCYClPWHdnxQ2WV+3sY3sCTnvc/Y18glVn1STBck/4fl6jKIz7hL
YQ6Pkfzpu7moWRAgyjxRnwGAHKbLtqwwoauen3gbWAZF8QjC7dwDboj8XA0oIj25
+kvTf3Q9e3jRQ1T8QVIWV0NPsHbEQ6eQwLjRyKpcnsfbDPHtACbVTYARKATIr4W+
zuN963xFMyi3jT2eT8isAmGKLzwzNR4lJQuZ8/rcZd5UcOfoICsyIaXg3+jVlOGz
rVKnXKRW4UOcgnDAuyojYWAbnBBy7YbTdO83C6m3OSI4zo9tplj6zx+V6Wau3b+h
5d3VMFH9h+h/vK31NJ+49lwUzscU1a1+ezqMFHf0DHV01fVQ2CbrA0up60UDMDI1
2gg0xaVrapjvQ/3x/SdOcXcqpxnzIDS2UrquZ9VRY/SXe9LCDimsIh723jlBd3ud
H6kRGK0nvUrNFmFzctUwlxwyWARaqzyK48z4OQ0mQaglhyUdxEmH3AAffGr4I3yn
s2uUmDpAeX6efmAWQhbeKHif4+mfoTY9V4gAl3x8PV40A7Tx0fpPAooY6Ec1FY/E
ed7RF6S0lRYYuoMsLH5Bfep5oFGi5svxivxljU/B16AIau6+XAfzPagOHr+CrKV0
UsxjIgVW7vZVMcah1t3sIf1OB1XWMxIrbq7pVJ7YEJrZjgM/2uNLzPOdst6UaWZN
3HLbfId4FechGgGMgOYTvn3dchls9eOQEP6U9pdPqfbBcFonuanFJEKHkZyNx0vR
BMwV9O4Cl6oiK1t96XqmrK4Tqd8/KR83WqiGP6apmEm7sdCSxrZnUGmtB7FMDlmk
xOc5bYyiaqpLi58E8RVNA82kd/QMAXdoR3meS4E7V9p9nM34y2H/xM23vx0l5c4j
Q1GDbtoBmdTQDEHO4iw+UlKVK/Urdx54AW4xZyagtIsbWTDPCM/glxacRYXNVEVq
+gT98XLv8PNK49bI4+JCoZBl0ev1p4uqgrDf0vo7jfkhIgwz1yfZ9cL+8XaGekU0
PrGkGnNOovTyj0ThUeXzosNpFfvkHG7TdGXEW4rPV5rDAeS3DqTLxgXy8/mHGVFI
jhYZQP8+XCkxGXedQmzfAsLFzVX+InI91frJMgNWRSI9at9tQOZ7VYcIvvAePr7x
/+uDd7Ty23Ks5b6oG6W4nTKFL+u4qKBQiXkI86iSdEOS2MfgrbG8C/6fgp+6JOe5
4ns09NdZR3tMJT/DJX+YnIzLigA8C/kaq3ogSXDrenCjJWlpBPl3b8zzGSTx+wog
+fIJLgby0DOth/RhfIoHwfNWNWpnerKHJi1HuuOiwFsZ4atDcOCuFSer+8uuGLSH
BIhh4zcbOarZ2WglHhEh8Ebnr+KjahKdSx3t22e6Gt5MIs2D3PIhrQr9YiSopRUk
mhPElEgvwPGd6nCcfmlhn9QgsvxotZtAvkD1+BqtyW5nkfoLH0X2LLVtVuC424BP
zlvfJWXvDf0/LTsRveHLIq8RxHwgj9IKK8NMI2SpDuGiGy0dVcFhtbSMg1oBgYpw
hIQCq7LtqUtcy/wOCjroPM1PAORcrnSSE7pcBqAPfjYcW7jYBwFiFx7PUYVLlLoo
LnDy87Ub7YYJXH0Q4sDq5yIaGhKJ9QMKyvzVnuHNtobohiuUcnyCCdr+XlEUyo0Y
QSR6XVzGxWD6h35GDG/aRJJd0EmtDX/Bt8Xa68Hqh8/mXMheGqgmDJgP+wVM6IDj
jm6qXMv4CWDOZ1FdTRz0AOsEBTI5Sh0vGAkp2y7p7jN8OJx7CYVqZ9M+PDHE7GG3
h8M79+lkl/qljNho0Mk6BFaV8PPE77MbmBsOfp0zCEW/8ULW2EYQjoEtJgk871wS
0q/3my5UJLepuCRiszo/+JTANohBvOnjYprmurDGgsCKnSh9XTW1tO+++EzfQRH7
QIpEVy70XrjeKjCCYUJntTSnuXf2Qf5q7j87enUQLRHQZxdV0hSdjXqrIWspxea4
McBKCH3OUAzcz0kW5TiBy51yshaAqDAYBHey53DB8wo4uDxo40XQK/NbslUzdEsO
tBPIdFhwqK2Mazz88XJ4/KHiyA8ESvJAyxvjfI1wsn+0JJY/hKbyzXmDCRmwDuWm
tSyg3z+EnoLbo/TZY3prwuuF5lysaYjQX82dOoPy5m7B2DhdJ9/kpSK7Chnsa6Go
VttW2hGlwBsV/HiELVUbW5qwmxkOHzcBpZGg2krL1bRhwqGQ1tSEw4LrUkspk9Wm
yVGTUcby+fedPs2fPXW0qxPGHgXwBLH972mBcZZIT8O17QHLrixkTujKRNVpKsc7
JddDbbGnr+hhN7QRuUzs41yBDNjO1DDaffEA/lzMmuLEbj7zc/ILGxFHzCq7g1dV
LgUKodK29JUI5SqnSSB/wN8v+QPe8eGuqny1SzFDttwT5Z4SfbTJ0pyGLazRHl9f
TB3W4NIWqSeILrYKwS0dTU97peqYqINyz7DJVS5UhVxPG8sffXiL0CY6sRX++mD9
okrKDfyb14cEAQzHvDs96L0Bh5nI9FXG0uz0Cqo9Qv9rOejBW0n2bYHTrQkt7M0C
4si8979W1TF1alAJj4uas9MJttrYIhpMQIFhnf2/NF+tesYgKx2evhNLG/pUypE3
MgPjV7ne9H0I8SoC+J37ZSEGa0af+E6QuxNyX53r1oo9tbjW4dD+j95GoUd1fO1n
wxhtfvQMMv1tKmQi1SFFlfZcpdVEvEezXkRgrioAvAEhKVjlIFB5S+ZFrxYFpNJv
/RXsmX5vSfAF3SJqNgThYf2zazbAKQiZJie62l70/PoNk0JuU9w/G9GqUkbmtr9q
Sgp/xkQ4qsMWqpaunipbir065V7GIelpbA58HZazZGA4JP+jMD7G+shjmGTZ7Yx+
K5Jhav+mwzsjgKAMrvij2BtM8iWLpzFAV8tD4mo6HD0Q6YNfJswMY+5zm0vP2Dhd
k571JZ06vXc8VOLzUV9Ass1hEVswjGaZIpYoW+9CBttqb6fE65YM714Hr3vBnZN+
TKPBzDnUPoDfaV8guNhXsh/+Z7M1m1YcXZegzZkomvWAZ1pef+yMBaqcVvmmv6b/
Rd0FqdJBknPxoGuRZ5e4ZMrlH9HThgOcwdYpYcVGSrLfl0vCeID3fWAxJn+d54mI
YAWJ9arFzgdLoZcuJXiTVfqttQXVMaZ23sGebah/U/MQkt18x6GoGfM5WtqCyEjD
vZV6DS2HcLFPgM6siXQMyAs1lrIOgagTjVDegdrxQVdqYw/0XCpyn8rjxBkYR4ZY
A0EshIQgFidDU+CBaCSGsadjuFN0R+wQDpI2/87VxmWUOX9cKDpmj51j8DhoGpB5
v6ugUGVVA63FRWcHchO5avi0icPJrl0AMCYlklpcIMpBQX51Q9f1vWdKs+0twYRs
DWk95hZbuvGGh2oNJOlF3IHFKqQEZgyrv91PJsmyEvgVw+f34UmeAvptEOSpkpq4
xlYwwnEmxkBhvpgVFk+sNoelGE5GenU2H1Vn/P2eH+gQ1wfRvo0fpu1QHJn7ot5I
ZQPGj0na8xxENQBQlQzXjNHAhHd7YXSUe7ZlYOwkzml70yc9H4W0HtmAzjlrmsLm
PhMq7uuT41ThSB3zUBIYYT9eJ9pJaOweOFRArlCJh0cASGK+JaNkhlrGGDOTfmy8
uYSVI+8ipiQSr8T19GYDzbCkwlUU4fVXctefq9Dlz7pEWpuGNtK8qMkx9Vxs16Ts
BCETHDJMvhEM1pmN6u65cI0YxdQhMvkFJsUoeKn9bgepobQN1ro6xlsJy50YBIhF
aPS4vJlMZLJgXf3+SjQvrzaxd1WtiOamRwzLIrI/ZX31QiO2drN0CQSv7uqUEC9V
pQY8a4+OOB3JnFoyhKLSPgtOcRiH77/939k20sr4YCz2pDirUtDH6Jg78/B5OqxG
k2cJ9eZ8J3RKAsmU9dk5TRarK6wJ8tV6xzLQ2iFHTmWWTrk8w1VXW1GYUIgeEBt5
c6WScG4c6SRMOLQreMMF/KhBInvvfXJIjbgiOr7X3q+e3v+jDqpWwKPdRQLTZ9dw
cget2NbEEA6YM+bFUreukZN+2Ua/Q9BNleKR7CiuakpNa/JZUjfU20ALYEG9vOle
RV1sQ81l3IZ8RczwBa/6MEKOoUeL+2az1xv5xM5oSdgSyIH+ukPbMAg9HbhRYp8S
jtw5kIx1tFNUHWPZQxtrLNx1ijMyGSFWgM1PQ28BVHmGe0YamdRZzuKx5ihBzjB3
MbZ+/aG83VYVl+muSarES+43q6ccWqpVuQdw98lBC9/jScTESg5QjFJSRVG2nSv3
eomCmEkqSXjmTNCAKpDCYsCLbGK39F2jFeUQROh7TmHfM4fRkSM9KqtUYIu1+K0W
B9FQwIRoAbWGjx8Bxd4xEozYHSAufwEEEV4K6zmaCb1H60ekqEy7WyZWyaPbp8mX
QNzYxkm6lHrs1ATeqvFa97ewjTMgbydvkNuoP+NUAJVm4Fv9OKnbgqS84a4kuabZ
wEIJQ8PeVKR26pPsPdTBLEIT3Ask7i6aW0Yjw8tcyPgZp32ht6/xl9nGfKD0H3ol
rDGNb6Gxy0Nusp2gYaGCnxkhaCeOpVj20UTUBYetv0rQdbzQFm2psgLZ5CETMYOV
Ckf/CcGKqoUYgY0yn0lamK/ZdWtd3IOwtksydpvfYuUgHkQuPz9rBOoYCH6m1BXl
kfFBXItuw55dY67xt/XHSIfslJDw8uMsnnE8GNgbd982O+Jz7LE/r/LmiZS7LQ5E
5kXSa53yR1Q2VnVz1ePKZvTLAwWSCTRUOCzQuysjKT8AcUX3PUBGFLnlk9Quf1AH
3yxxb5v516mEaLOR7G6E55Src2BK5aAvRCtpJBGzXfpZnofArrvuer88RslbajZK
tr2OgX2EWza8ZlUPdM3h4VKvJJVhlj+L4a2lLkz6rs2cyYETTt8lTvtrMfTo7FTj
tkMrnxO4fi6Re6BPD0J+b6tu9Yk8duvQYrj5b+RtS3vcGDVADeq5Xw+cdNfdCUjs
y9896Dn2OIiPsnpGWmqhoxZpQXo8xP+GD/gfXEOgAoDCPjgEYRAa08lSwLt7LLtl
jfnn1mvLWT77Jp4y4ySHoOPLjcu418QkLCDQsEu/xh2rFj+E/5pH8FRm8J9VT7nj
ZRSOn9+G5RmaH581BqkRfTGViWuVrrwTlG1nPu1GfHT4PD5m0yX0IrE7yxkC9NBa
xc4RaCOjuXLoJvGsg70gcoAfOy2Ohim3Mf5Y06KwGRiN6l66wwrCEsjylnEiUcw4
IMzEGSJM0KuRokCTBHQDBGYmjVItQRCT1UcammEMFgZc/gYUD1Z7hIOrkVhxk/Sj
oxteEs+WxFbjsH6LEgq2nqJ0+1+zVe+edelZsLqPLcVeOJe28hzOq/yPm1qMfvzj
ugCxEGqYx/CDvpAZhRf+rb7PAMmiwVeYMyGHuV5UbvR4QNX+l6xA7R8E5Hkq/fH1
NTly6iDUEkkAvcxmwPD8Z+IhiJdw7LMCPzy5JzJE6MPO6cSNiYFfanPb8CnuKhxg
FgGIb2zfvwO8Vok0gvKyKSxgWWB9wxA05tQpIMO8hjLVgzha67+5TUJv40kdzYT5
fVr5moqEdlXPK/J0Qc24W2S402ziJ6MFhVkn1ZvJAncgtjHPvko+kdysKz6CbtG2
20Iu7iEiwS7G88R/uAYONlh0Q1ZDt1EigC1UD5jDhJ2tNR6M/y3bZb/T4bSeQa7X
bCjKYZm7PnoCsCMeSl928P7O+THC1zrdQmYhelnhBr1wuqAXwpC0/q9Lh+zxZbj3
ITf+J2DxU7Gw1XpQFuffUMnTbrhsAkXd97FicRfwtTCsqAMBOe/ZVfbX1nsk0zoH
9XsWD0dSHX3Kwb0EmMd6z+XNdTN7n7j2w2RpY4b1I6PaBFtcYAPk0O3OMJgkRj7Y
AW7w/ZHoYGw1PKS8ixEOW5s6b+RgPkhHoyCWYEzW8Cu0daL3FnZnfI9GsaOwHgJa
eQl7bDTHEZ1fbzTwpk26lm23dhyXUtyJVlHgCXUj8rIMNN6GBL3zSdBq+xkBZfmR
WQxWCoHaGwx4LlX4IXu6YcBRzSwK/edL/MCzHo4UIW/pbPvYIBkeWc7ZiVCu8W/A
fncdnnPexHQgDNseq5xcc0eXPRn+D+5EQYHMSh8hy+oVSlFtAGHqvQ/R/CoTPy7B
gNMUN2wNBjK4uOYDkRgNduZDYvFtxmb/mMjE+bLamDJ1uYbZjtA7VIZ0CfwvTJSR
AgFw1qoRPvyShHTS2QsMyNbEDIY8lFLfc313F/4LvDJs1Oh9G2FOLmcwKvtHMHNO
Z9+fuUnYASC82WIzWi0xOSHSlpa5l9AEKFgI6KHx6JJITxk3gDquokSMt9h+mxnd
PkFqrehezs8HwDiyLd7dgdV4QGpSXqIXjAmQZsiP2vtIokHCgi2nqb8TVdS0Za/G
Vg8nTk0LsrJFXFqx1QN4hbwN0Wj2aq9tWLQ1iypFVHf4T05XGU8ch5QMuoy07NC2
3eK00PAD30Pd2qcmuyC1MVX6LApR5FBOZa7Sibn0o3EOTug7/UY2a+IKyK2iwa5p
fj5lfHZxLMqDWK1xNWp2NkIiZ85R5s2d77YlDGwqU87zvadWLBynyAh7eUSKRCCz
K36YGUnrC8lv85PXR/aUn5/q9SimNUCFWF5Bcy85EBvF8S/FtghN0lreczYXGjeY
YbfHJ6UDTgHBRLXu/oLwekrjr3ZS1Jp5TeSV88rVgbkgMr/uR6k7wargASVBO/Ua
ZipH9CpZmO6mUFM7NJhIG6eZdW2VVUxF4iVfTbYkllra+G3R6q3vBewodm0Hy2Cf
ThlAL5gm8nX9HIILwc9ZEtsaEx/9zkLE5d/FBuVPDYNG9QShyPp6HZfmpSsvCK5h
7Jxi/ly+Ie3FT6r64inM5KncPMwV+QBePbKqFqZcR+eup6c2RwRNUcGa+y+QUJ88
nlApc5lWV60WlymSKWOT71Rd9sUGinoNRlwHDhR6/v0OM889aasH8KCHiA91AVLG
aPKImdVhp/eDUK7EBUA+kq8QhLrErXQ9KFJsW1hAmGtg6bI1UhCDcRws/61zSzML
lmCCKHJ08fZqy6SVtxswViAM5tNFruRnCHVM44Dzr3PEocDbLX04mbFVQomMIUY5
QbFFznlaEAFI7CUT6MxmDx6X61JuPj/xu50WKMlYnTy9jVrFXiHj6ep3VVVUVdjh
kV1M6zZS5A/awVU5csh2vmgHORACs2IysDkP574Zb1ogzyz+LY2KRY2/PMydSxHI
iEqETmdOKWa0JIbHCdr8/1ZG37vXR62F2wk1yM+QmRVuT7+Uh4XykgndteBTDKcS
6nddFD5jBQfDI0/GakHw18KxLJ7ZMeFaVwojNTTK1Nny2mMgIw29KoIc4+PjxBxp
m40XwPIZdtKIunG7s111UFk4LtCD6YzwvypzVS8jm7A4GFd0oGlFzcUUueHlninW
uksu84I88zyNcKHp4Kh1+x7OKzwGd1zqXdCtqKTbPU7h2sW43uVIHwm0c+w8YVys
e2eXLllFbwqCnjkn0fCJ7JZZnTlzHereSqDqlc9/uvuyx9Ji1J3bFovLvDcmEDOu
TCSON2ZauxPH0GNbVVqo+4PHjpi0iR0te1Ypq19z38VBpxCEmGEpc3NHr1jbKZy+
d4/UJHLpbi/2GPS4LhkawOKVSMReWL5h8QeqIoyl5HqDv0T6HDnJCqxVK0NhBOCn
pg7qIkqyHX6J1cpXR3llUkexSMnCAD0p0nkDJSf46WZop5IYqmFqw5f8HQAhprlm
hTXzIqyXcuOqvX5QI2+zC2GncQa0VEVjg25WJr0aqxdn7OSPfffbjEqurmbeHfTO
l46+e1Zvt90ER5+MPHyVNhihBi7HDEqQfmTh1sGl/T1NWx05VzmXOMs5YoJfb4Fi
TDntMzxmEAPNBE+FbckDgs8o5YIF7IJpBW4h9Gj9qt0hsNtYK5zWVpmWYhT3DuEp
1MGJ51Jzdi3DGigsCfE7Qo8HUdroEwFUjQ4xdC1Itq17yeJj99VOj4Ni0PZ2eRuf
bUxFdI9uUZZN8dMItO/znLp+B/6Fc5SS1fnMUZFeImE5ndEO46SoJReIRmXNLO1t
wWRTfp8keZUslRnrEV+WSwdb3Q7DQk2x3rNFdAfMLsD0m0AFkcyIZSPvvKlgKEx/
6dobl1eBK/KvQepU4SEUpYPzaoMzhnKRDAZALteVLux8oHQZ6v0yMDOogtZgWwoG
TT4QV6TilCbzGuTfz3EONpMrnzs7wIqcR1YghO6n4g2uuGacBFgDUS+asZfvY/oM
UREnMKjqAmYyxTT7mNrJ8Qil//PviJoD70snnkPoV/bM+Wt02bdnViIEem7Jmwsf
80hDQlDgYhlx4tYJp2DpQeZ6nsGfXQFKLkMSoGV1DvaIJtZRM4d7Vq4SG/kOmWQW
Z36qjGb4VoGBmKjRI7kiIdKBEbIAyeMUS5HNX4JEcIwQ6mXaoNIMseyfW6azNuZZ
XHmIdjNXwon2JUftX+CqBTyWdQk0H8ctzfRnZcoygo48Pln6oFGiIja3ER5vA4Ou
CgmcbqmHET83GlC8NVllaZ6TQO2Qecmkn2NTA8r9WgwNZBFOADjhs9ng8/0Kpnjt
gotEyS3G8kgWa9MFOWZZxNJD03tIbrjyrmH+bKuTWFTd3M8tnBdq5Q5fWjiPeseJ
BQyscMtbhgEzZn1Xa/3DuE463Bw5RRZ5/b4srAFUAk0ISGFHgFCK0xAFqBXHmDVK
Vnc8pjBfycUR3F05Z3/68BDOL5/ySPMIBjxVEeI7HFfUgydMFdSofWctDeG2nWqa
4MB2hZ8UjTADLYtleHhoQizpjeZS4vLNq5NhllqSgRsuc3Lv36qlrKH5ZOTHFi+W
mpWDuiHtMsgWM6q9m5VnRwe1jEnmXc51st0YCO78pPR8Ga/IStAcUaB2dZqBbjCR
jgGDYpXHqEgfwEq5pDEV/YmBnVKtTLTrchkjqgdQ4n6HlY/3PlaHDp+xWdaR0Ls0
DztKTJUYWogXYkYhEE3lZMzQsedUSoU6WG5hqKjDEJeHWMKjR824yKanf3Z6S57q
aZIFvNtiron7WWFwFMljdqGZFeUEfKS68aybysnUnyFV6DjNMQbol7j4KEVFwPox
IdbHCuUiPFIH+YJfxdnI2uxwdTyu293JMSZDW/37ZyuBMAUmzINg3N5eZRTrpLYc
UavKteS7Q146NSk+LNXlAm6G/e5ZZcQB+8v8PCp8zn+3jBPB6JD9ludNx/NSj6zI
1v3pxsqZTMho77K9NiOQsjbjHd0YglNYF9O3HfjKh64+S8Uf3Le77HjZs4s/X/8w
lGBKF2OlbAYIEj8PaFYvGVgQLOh7CUyzwELOtdi47Pzryqw/y80XqZJ4OPWpFiWa
vnT7DO/DUNBkLqeHVThJK3kHIwrLvZdwWwtj9/4aq3TVINXZq0Jg4xfRp92uhqnY
qvBdtRki3cciHOo1YgXchptuFq8pMQJBOvdu8g4+J0lZpdc3OvMjZQoMzarezIop
bPl68f3qnCeUKr7Sy08cBiYL4OoYRxH/S4FzuHaacr8b3KGGakTt/x4EeHPqzpN+
AU1b6gvZrRnHbvGTD1YbzK7NhMW0HpI8lxZQzE+UVqZbW+0y3hqYKws1rFnFya8I
9k0S/6OU4iZ9EhPLui5PpP7ydrJjgksT3PR9bXltbJ7uEzhqZxa2utsengLXM4id
ZnFHIxWrTRHK6mp+c5ShTTp8+R8CsQ0q71A0P1y+jwmCrLtfZ+CMD3vv0bi3BeEj
q8/lyBlzpEMbCOGHO2cIBzG0YMJFwS9XDs0D829Dd8+QUbdR2sbWtFWeDjB9y7+3
eSt1+IthS8Ogga2EVrNYj7LY5zCxbhcyfGyTK99e9LZECjRrNgY/O4I4dpQq0CTp
+psFl3cdwfzormfs8vCBTVY1SE0v431TkHWNvDjAXqG23lPNewzHy12yg0ECh6yp
EVmQHHhM7Jr7h9YI2iHYxelvabN3wpVZGjfC0q1LuYjUk6XDtNHPceL0B8cKZli6
FuZdSKfG7qXauYsDrJla+KRvA5sSztwZ1juWflzy4n+PCPHNQU2DKD0jdxurD3BV
S+UyciQYEmNc+t8pw3LylfioE+ehHzTo81LyCWnq4JMVRLlDKazeh0kypXHcmhwx
k1xUquMYtTugGQQ1kn6RAEG9KFIpYltBE2FASnGVT981qqKa+JHLDxrm1DOuMr28
TaHHQZtfAMgdBEQAjfAtY5hfEoGK5KYDWjDlf09KrSX2y5BkhRftMPoUdVgFcgMH
ikghdTgwLY4ttCyFUelfW+7M0u0Nb5TIoBi/i8Pe28w4VewjMYzJqtl2owiHPzwJ
VN5TdMb1xhZVpk5595k/UPOGU99Gt4MwpxXpfWnbhsy5BEC26P0pKX7F7mkjJEH3
dM0brItqA767uZGa+JZ4eQUwWGF6E7QvowyGRw+Cll8rXkXa3k8XQ0tXVZb/gZRv
zEaXr5CHhehd0irsTlLvers4pINUr0OVuMUmmtQpwRDThf0m2rwSI27sVTjiw7Ok
AtncxOnelUW+Pil+MI2VUSwLKPcz2E2xpBP87orRUnn1pEsQ0eTWOPQRNC9QneBd
bY7SPZU6ZZwuohZl2b1m9x/Yu7dzGr6UGVqKKb5iAhmOX8uWqjUJ2Yf/xhMKEJfY
i7yqFPizguZy2SK4YLfFCBiqlLiETUNzyauUNDuAqvDYOl1m/ncJp1H6fxAVD95X
5UjHDJyM6B/mEIZd7hYUxOwxhgxl+t+gRXDKl1h+G+QgnhBibvx89hr51bg5SAJ2
wFS7uTPvUPSX/pNh60ve6X5Ed3RCplxcBXJJZh9Gg9+aKsGLt3YIANrrtyYWZRpp
G10X6dHdgSywvlYJH4IPe0PRfYY3HNXCd8iDLrIgCbbUl887QT1AR/OwZ6AYcrLn
PMD3fJ/oJNt7LM/BDooLvK5gENDGw9oQeMwHVrJzejiGidj/3TXOhY1l2HVXYjZi
QJ1vOnVsN2P/gezyBPSIo5/e4LcjzmqIvC9gWmiVOI/0k2+QVjl/LUCyqM+FZV6i
ZSTef+dgZxc9D6p/y/gb1sW1gBjZJ0RFoSPnR4WF2eraWTaQ2o8uCI1ECrmnN0uD
ssxGRqusBupoqKEhrqJjxOiTm5LKuI4e47Rr07LTvHSSdbcRravaSvT4hogDbzNx
NZhToHwYhvv1A6coRh+xozG3viWqn26X3xBPReZYrnfQRF4lHdaZTyumgolDbCKd
lSbXzzeJXvjwCEzMzlXMjwEKEc0PAhpOlcrHiVTUiCvQeECzXJeyGy0btjhsbi9W
MAxuNWRWAavWMxRjQvWTrc/yYgj7fmrYKmHs/nXo1wTRDBrXOwwQn3jtsykz68Lx
PWJwO0wUW6r5F9LEe4zlv1LAoQYFkoEhmQ/hWzdWhuxonij8jI1uAFRsAmUr7/g/
If+CQTP/sfo6A1F1n/6X6j5SiAYqXwbyaempclbKL155uqtEip2lcIYSYCY/+huK
tvL8U63QxOsITMq1KQ79pJC2fPk2IxN43z/WJZ4OhsNGKCSKU5meNU9pcY5eK81n
dZXaO3FeHC5kk90mLo1eblAQr89mj1AZa5S2I0e1gkvMH3M7uSZZQEsd9TVSnTXb
LMvMAk/G9/wcPLlPH9IZqtN9/JvW4AEf8PB86copLFX9Lr3AePprguQ4+Ao+iDAF
+xku0j4FOuZQ30NZF5PuA9tuYdbIsL+iK72Pjvi41sfTipVzU7mm3tmGdH4VuRlF
ZJ2ixZWc7R1bFdp5hlGhXQrpLTdr+QnVMlj8ooDija4O72O+xTLaOoJwffSQ6JAm
FIy3MFZHRD4zbcISQUxHyqqqhqcl7hLHdEfFuJqJyu4jY5vveW5e0a3uL9XMKPkR
mSr3KpMxivn6tg4ibWkNI1m9vJYnCK7XyDyy9hyl23paIFf6C5ByPtA+mex1ap5m
CsApy0XZcKP/izDSYbOLxIgMd3fdPonIz9I53uC/n78P58aOEo07bf59EnBr64sK
CHF3l49ccU2qstXoFrZVEGrnj9J0b0fqLhfc8veKommuIlS37lPhErNYCHG6iPIX
HamRwKPul7tVVZ+GUGwmscrZ+r4Zs/izM29ANigepkeUbbPj37OevqYDWkyWnoGT
CTKhxNURCPemSPBn7SicvzNCabTNZC9RfAE/DzShAP3zqFvOO5500nryyUBfswcl
VR++c4U+LRX+N3IiuoZXBCwdzRvVxvEn5ptdDfvhcOyM9nu9ih688LlERCm5ajzB
GnV7gGSbfl/MmRYWkd3A+sic2ZeTd7y523E8J6mueBCfu25i8jJwthrEaI2h43rP
XSVkonIHpFhG6INrr4uXF0s2cwMdzUW6fcXdFN9vE75HJL8AqB7MfBix6iAyorCj
qg2IYwTni0Ro/5JDEV5iwmmm8t8NxncYtluYIACqM5A6qYqGa6BhhSwwroVNmY5v
4SHNUPr6hkPSl2QlV6qyxKRNYadF6B7D7bcnbhEhrsZIsMkJfPAYHIE71S73dMmf
P3FyDalW8xEUGLqpTR4p26jG3TMwzLHZCxIp9Gv2vqxgxiitvrtR7ZWYtyGPjAaT
b8I08SOAwcfgMr1dhA/6tzRit1XtgW+sd1OH9m7KdqD8ThbHKX6GS2sxueAAsCv9
hRwaKPcUmQvn/O7z0UoBVZIf6nnfvyOwm9Wh4hzWmmXufQnkPpQCRX5nkOg7rJZz
QbfnCL8gRR+n1A16iAC3MII+e9QaxMVZxi41bV1o4/Sqih3If2Bp7mPtezJbMtr6
+orUWKFE3mOmJDhfzPe+mXQD09Pgam+6tKi2Xw7LgfcDoI8m+2x/RftM2Oa6flj4
aT3+iyD+WMstJV+8+H5j0sXEAXGX2dUU6vRABUYEuccuTjI9EYm/SdtE0ORsYR/Y
nRmh7GvR6dz/l3OeE0AuiDs54Q5vQxGvwQHjOXK+yYEyj6HqWhsEuBthtryqHCll
5/9yU2etym/6ALPP67qOZ+aKaS5fmv9+66tFyD2tuQqweVYqAuBrT/OSglAMW4J+
xvxByZ5pWqIWpZ7I6DmjlllRL/5tVfmJ3bIIXDv+u49JTkKP2Ms3bow8Ca6jVJ3+
kpU938LaL2L+A5AERSYrMa0P1De0uD6RpAmoB1TjCL5TTVg6e/9IY3WtbOvj1vj9
BKCOFHcC6lKS+yA1TAEh4BOwwfUHBrspKZIB9xgHSjE0BBlCJtIsuY9S0rqHnAnM
ShLNFu+0CBLnIZ6K8hXykSCwEkQUH5GF/CTHuMSigIM7gZi8IBAcIZbMjfh/1wsA
bohnVGjwigkmYqFhc8ioqmC7qiOlVDa4RoAudsijBtWOYYg+Y4qT2EltqSdHINta
Co3nVaWWxQrxnFVEZ5oMkBZG4EN0oF0dX2p0cmXJFUkIRiAZYEnc35GGqE01XswY
PP5l/sLfpxqC6wQvGYB5OF/mY5Ujb2lylgEQEXnhTQctgOGBi2GQyzmhPV4NBwbM
qJ2jQojFfEK1Uj1hS57vJy7b1eCCp+Laszc2j0U4eKGBeXVS3PeynTAVTbKtkvxv
YsvY8apeoI4/TtQ8BYwkE+gwa+fMWL6vkLx6uvBLlDs4wjr6QmIZqLLH5Ik+iVhT
acjzr1BU0rv/N9VQItWpHEzZkTtks9KYX7KLu/7D8bgFVD+YfO5+a+E5mYP3TD5I
Kl4+B7WnJpaTXb9hgJ9Y7qHAkhD3agP4oipjzBbE7oich2epLDLxRUwYGzUe4XN0
N92Fv8XuN4celwt425SZkWnmo9vbAF+yIL5dnKD8B6BMYsbawUSS0mH+XxhAhk/s
YZQYNJqEWDJvfJaMswhLLxcknunWtWCFW8z/ZD775ClqBrYHM2DzGCoVTk9/ijqC
LJWCrAkh07Ma1iVd8LxSJe+cY40L9LOT4ouwGRrmF6CGAicijrNfPCNhReqq6289
WUDHjKlWnGasQXweSsxyZ+ARFsnA20ct0TjdmM8lHJnVlp/CGCA7vL9ZfgmY2/0Z
s0HwaHlNdukM7cUck2tGCNPcIPgwrpciossFxhO63kr2tiR9khcMwHb7q5RQjDD/
aZ1M6gj3SemNwKUPGT5xF09zqSELwdKOj6FKf0qTxKPJdVh1dtKrzRCyO3YPBOKF
GQ6WZdXlzFQGAZFTN9TvxeD26R7YX2GwPkt6KER3SGTbK7SpipSeHO5uoCGu5zrb
aymDfyJWT9oQ9+dJRsl2gWVi5S57hSwDkMcS+8TJ75BIxS5Fkv0pO+ePK3mExYpo
KSsfiWnduHq8do5U53dXF5ushL/5Nxswt0KrlDKqK/IDCoDM+ZZX7n6s7LE+bVik
V2tXE+phxcVOlhl+iiD9FdhDbVe/uEPwOEO7+jH0b4EW3r8AKNbPTejwdMaUqvET
/WLnmnzmqf2uFqUwaaP15CzO7KxKXFEVla0V0z8eW6p8Zqcu2Efoy45958NLjtzu
hFa9or9SuDe1an/6uTYQYTeCDenn/D8AOJ54pxExXQoc2cYAMkLkXBrtmKX24lr8
BUJUV8a+iQULkGcoTIgvLjGjXBS1kd2Gejp91FQ21EHp58j++TxUbGMy67upf6LY
MUhHZ4GiJNCrlV1AKOGyE9dUyN/S1r7t3H3CrJZiPuMI/06vp+2tkdMZ0KotfB4N
UEXRbGTmxp/HV5UXXgerdH5JX5zjrLk+ZrRkYC/iA+MMEdwYpq6jte/19vkJ7Wc8
7anTmux/PaX6uUL7K+DJwSgNyPS1oUEJklkjOGxljFkBTPoShQFpyocRR92SVBYO
xYO405hxLl/Q0kUGG+WNdl/JU91ZHabV9nUhZnAidR80kpyzUQK2BOpOinYBbQDL
KlAS9F3n+n5Gtes8QjgZv4mu27wDm+TveQX1iQY54zAi6NcIkor31ITlgrR0c9rq
z4OjdsjMQRRVG9w8gCQRWv3LXQAiy/6PVMgWjjkJ6edHTKJUspuFI8swyqnb1uP1
Cae2SkTpC9CGE9H014h8JZ2vfoQvZ4/aTA2uQeIzQ0CQU/xZxWMVtbZJdBR4Frx7
jMOUxxCOrQ1FDm2yx8cmN1GmdCvDtwNpcTO4omeRQuZ6OAK3p0z22geborf0vOML
inz9YXlLhtZlDyRktla+oCuO0I+036ZVasTf1JfaUN106ZeD3eUcnNClMHdQSpsB
3kIbQj29YOwiRaGXpkjBqYGwce9oNNCWr5wo+fMhND1hLtawsMQWbxtsJo0C7Fbf
ntO0PriSfCsqW3/jVRiXnYlyJ+nOpI0yAPQn52lVHm3Wr7HhWg7Cx2l0g8lHneXx
jNHEOaWgpa9KnxzUHAICY1asOerlqjGeyd6jD+cxnqOOneAQALxxulnEsxpUuZM8
C0TCJRMMHmDMgR8GngAmKPhLOEJnlz8L4AvylTLlRJVVAQlF6JNosax4M/YiQKXC
+OiW+3xgivXlJ1fLozyncDM5kwcFxGnEh6tLo7qt+I8T+bgXWv9+l+TSGb5UmUm6
XeP4fV6OLacSNCq1xGDyzMlIwDNm8mH9la9weBGBUlViAJz07kVh999WEe0HBlXl
Hqepw5Q0GugFfNb3CuYLaqun4rrSWAP5IT7YsyX7gr2JUASD3wsFnrAXYdMCmqw+
OsKp+sr5RqlCogUerTE1kl3s43VuZVQuFI9r0FDbGm2Ru55XizouKW628N1A7nHD
Jdk+HULhi1P+DTZ8vozt0hWOVTqc5mnCBqtV1Q6V9ydNtkWehv1KVyZHgG5HDwxR
ulQja5kjsz6SUPe+p1tTvpCSyeDenccyODIk3GrVVsNXn8LYMRwkAgLYoFOjLw35
/O7Wc+s4LbXcs5Pi8lVqdYAWP/aQu6YvWlyUWM/dxawG/hZsDpyLy3penm7Fi5F1
NZ01yppqCabAfFXAbbqqPnnRBtzZbp/aF0MDxVM+qC6mlpY6rNan0jxCIQHOV2cp
JZdzVH5VaivVOcFFA/vKypFyKRyXjCt4jidazo0cXWZAM/RCqu4UQ85p+Jq7EKEZ
lX97wvZK79DuDUvsjwufgyLvWU168JpmQP5zH4Q/qsynVG+zuNMRtMJLFVyIDRyD
ub5ABHk5X1ZBUGGuLwDOsyxulqkFyiajG2YF5MK42JUv2+gFi5VUdVTOW6ytkFQX
PvqDF81kw5kchLw8xT0MtVt5qDhW9jKBgxtkX+6nG5RX3/kHc3WTNZ3i+bPLzx/n
KeHZQCW8t4EuomN4GbQEMvS/3WyytbQyRnbeZyDsFvA/a2aYsNkM4NvO07g08E7p
/pBqOp1pg+x03tDg07mtEhzVxwoYDzuDTJ4YgSmBK8YEn8+P/K2i5Pm6GsLj2NAo
nPqVqcoKqNTJdFLifAIftIn6Xo7yPBBPYJhQwku7zhWPAGqW+QQtZK9AIVkJKFoW
nqBUbZlLwgsYs6BToICbudJE/iApe4pSscNUTuDviFBs3NIJp1Jjpzmp/rdh35x1
DtvIGiIkTr0rgCeonRAkmbolGxRi55dk/OkAHiPLCO+sE5gwarVTuIujajt4zr0f
shZTwRQ2ep3b2HxA8ojmtkVhqa6KdUWCJxOHUmNT1DCzWYx1SAJnyZXUmaUkdut3
yC47i5Nk4ycemLysRSYkYykqMvevGzzfV0yhdI++Q9+qUunyU40IjssGgcXfxy0H
xN/ctvsz5AkJBEfOJWkUhpaM+ZEoQb30ZUp6kSCo42PArjx2rMMNy2XTT1HrmIhZ
az283DgcBfSoRAQraQbFZLHehEv97vPRUv3Iu5lEAx4K+2+dkeXaxG0U/MBI5ihI
CZZhA/8/YQYMAqFcdsBfC4dV/bVwAfOFdr32aTN5jHQ9SqYENmije4ratXIRqujs
OMbnIF6vRebsgip1ZoSrh6okSfKGeDTtZ3C3XuYROH6dhpFvo+LeYQyp3uvWFdFT
R0vB/nL3cOxlHA2bShNASUQFkYx5ubDWi/mCPU9cFz9ggZka+hiqDTsIG/JNqD6o
BU1jLBhtof/yRXMJEf9LTVkmRkUyceo+8cYx2/X0mnGJy8KzJJB+LzTbGFtgeoxN
/kiI4hYTxXTXEukYGMHgZD8dsr5+0Z0UyXDCZWWtBvCbL2KSiw6tiLUqLSXqps4p
15PLSbIeifRn8+quqeXqInl3rs7BGmmjWCqNRAQ0FQp0aN3mxErNJcNmkxa/Or61
FfHbN3zt/X0DdhJ9vTuPGb5LVMtjDNoKn/+IuP6VZoyE8YY42HmRoEUxIFg4Psog
RaUZ3RMZpsxLNqMY1Y0N8Mx3KTzI2c485Kqh4e3gDPtI4BkfzXcgulWIA5LLjWnG
PPq1NITxDP22r4frgCEquCI5I/SboOAf9bpyXvz0vxtIrU+tLqq907kW3JZ3ECc0
shE07miGReh4rXRtbTEcvbGZHjl0yskbdGt2GCQLHPzlx2AMtOJba42GQT3XQkOq
SMfI74Se8q7mkq49mHfFRSHrPOEkbfpOBcpo3UefosKs0GO2nVkdlaKw1ZHwRTXf
4/YTXxuCpTKoERDEZKKVqHBEOFN4Be0ghxO3vFDz0ZrYzPLJE7AIpbtZg+CHtWAf
O0Z08ASW+kkKAtTxz1oioZIHDy7QQN+oPV3O0YdDMIMRPA7QLMfI8/Tef7rtbM+s
lbooOUqm2bv+F9GDPlor3xjhwiUMfyYIZNbKgthIhUS/bbRP2HBfHb3hTqanxXNi
/PrWsuIJN4Jyqn5Vm+7DU+XzYI8cfKTuRp3e29dB6Af+mqjbn45wfsn4eyb/0NL4
k7CtcwOE2WXikPfoFmkC8ETvEUaCtenrXe5h6Pd5+hh/j6LCA44THqTmo0iLuEZX
JUQp6ZIlmO5m39OdCqU2VcRFU3axOw0P8zP5poAIx0VBK4A7Df9vD8O/IS+d5Re4
HcVmwyPZ6ruXwMFDpxo1d7nPWwg+61b4FVFOLQiW6ma1ZgEeXhE3AejQ2+udNRzW
0QusyDauGK8UiJL8oxUfxl2bOQxlxWWgb6wwfVH+zx5WiXCfyR++tXIpYjOTaSqh
n2LJ7zK+ATA7ZR2hB89YpqESXTUViyKRvGtP/VU2/mTdbtxxEGTbkeW+DKepYoo4
rkL+u2l/6nA3XgItHuzPL24aM42RgndweSYCKIlvS8krX0P7EMfW0JtZlSqBmj0I
C0y6GPsLUVN9o+hiNlDT/dxwIrGswPvmi+uk1W1XK+iKq7Io/RjMDph0mQ+OLw/7
i7p6G9ayDqXoLW12x03/PbuNZDpBZzUd0lO0oFYwtpPPYXdiXEplMY8uHj553WOF
bvgJc7ci30LrCQ1OyPncgp5DN11cbbqDJ92C1mQ7Te+gV3sVo14G2WrJPznAFTLb
w/bbRLmC80/I3zuSWL06Nc/2w/Rue/abllpBP0ZtfzsvuW8f6qcWmWcNDQ+csuw9
uAdHJCsy61uo55DRjgBszrF/F7cVR5M5ak7E4W3LIwONuTByVPo/g3PBUFJfr/5c
Ia53/zcgZyYBVtGzND/n3j5NX9Ep3XgkCh28c3ys6iCcagMQU0SjI3wL3zvd/Trq
6n9Y22wiDh9NZWyoqtoFImwEbnR9GkvKgRHBRSUS1gOIjfoi/J6b6wRdiEJHLHeJ
zXot9Pw8VPlu3PS1x/N/w7BLs0WOfB6hIn2itmMYXcbdQ/p+WRyh9z09x9Jcy7Vz
9n1EbBOU1iqqczq7NfEns3yKDo+gyldbRHwPj42ISeDAgGwVKrBsIZEdVD9SNNkB
I0Knwdv569MomD1rXgI0ffdnFJAEDwNW+ozVO9qOqjb1rrI+jd1czn9+abCkSSzQ
R/YRQg91xvS9U0NjNkx5UAyrYXgi/rIcAsgObF1GBS81eYrXySQ55E6GspTW1doQ
X5pWpp6W2R/SkhIXUVOFJaAtcSRLP86Ju83qKnLlqaTJJR+Nk8pLPbYD8rJAg7io
opdpNPAhuz//G8y2+0mFMHrYuopagY9UpPjmBSwg/qmmHMRaUjYwPsJwaLdGAk++
4m//QLh+sjxAF+iWzUzdI2erlIebKgl+JwrLXZhZHX7rNy1Ns628bFoYCDisL7DF
TmEz++KYnv+3MhYSqVLiQJwV/y6ba221UmKVh9k/0/oZcBZFUjUofeEJQG8BoCb3
kNJLuQn+TzNCPwJ2m0Lc/CIJIRJlUd4o/fBIm/0MnnlkAWQTZivHazRSeveP/Wze
cFTbGwp7Tp1IaHJS018XzWchAn13aVikzYZibvuzS+O6qDjsj3/aoi1Wdd9g8Mv8
7x4aP9XwQ02FsUmdqmSXJNZPUpmq6fbKzTDNnhxtRO0OemYCbasfjZFGHFIIjHOx
AcUbUB/WkZi34Cpuh4+iNz0LOH3+tlpww+SBkLLicsKYXVDAWfyA8r7uihmilJVD
LeSJ/Iz7xIS+j/eJS6HUUc6Rbsja0xPggDTTKnpd1ERRSYtwBBqdp0H+4wshEAHI
3Sh0vr/aSAgMPpIoNMc77QALfus4NVzfYc5RPxe8LvnvZeQJssbDpGk/OxyqmtZB
DiIOBbQGy5aBB4VLrV9PhG2cqHNp7SZv6egV2tfol2rvQ8CJPDCw7Gq1rHGgPLg+
Eh/l6WFcUDqOlgkVDPxlUtgHRudAbMJFzvxyXKAWU0Ge4V7KfZ1qcO68yIQYwJGD
r4Sbh3FqX2XSzAqvq8Gfijx9hD3MQiHFjhEkVJwkeFcetlYi/WpsgZ/bH9ZV4RR3
8JkK61K8+TGRdbpcMs2XqMJS+Bg34q3nu8AtxJHSKyXfzUcE3NyPdWJCBE6PWMIy
9tDyigbjvpYfTy1T+ImI08Mi/Xi4k1/Sa5Mcfxgz4DB1FrVjFpACXsaNu/a7jpuF
ID2CIiov/Iq3wv+G2Iqnkioe8NQbQFaYN0HlYCKPGQuTQHffcYauh9iTMGuK2Xx5
LR1gTuH2TZxv5t+SvpF+l/HrP8NLNo5ql3HYyuq56SZi7Y0orHOHuRnmxAuQnHdG
jf9/kEh/arpv7DsvOWvMe53sjwRK6Fhg+03vdQVBlRwgnG/P+RVg5WojY39U30IF
tjoH9EMb/y2WxvQXKXtgN7e0OWqssp4eWeAPB5D4nFOG1AADUSf1VIK9/dyUxZwE
1w7FpHkvTvX3mdyu7A2ASBoLTKUNFqA0JfEATAY4xijYwHEXh4ys9Fu6yj+bp/8d
bWFTdBvYTL5IjBpboVlJP3LjLssekZ2apZ4GC/p0SLzjkNJIUmSZPFBCWGS192Hv
VmuihXHp8TdPqY9+FLVYKehPMztnhDW3qy/mMw0+IgnPkSkW2qOwHcSjDYmLwdcF
ez2wtVn6S8YkWNn8Ju3G+e74qSLPKhRbwDrpQ+H5uMLMcBrcxbq/7Mp3nw7WgdST
zH08xtyWP0logolqQekDYMBayDH3/jfnvN5OCMtXd70KlkFu5Zcda0ubq1sndzqQ
+Nanudk6pm20N0GnlGCoU5Yv7Jlzg0xao4RmhbFWVrcU168SGv0+aBe9RTS8T0Yb
4GuqTxDFa/ohA5ziqrxOWQtclX/WtqTcDjsLwAJafNp3RijXANfmJCDrd9uaTphQ
3psDoyIOrjRCGsW2m6hRAy4EsuWMAUcqp1xHK7Jh3ER9d85VNvK+t92LwM09rG1U
zQ/XDTcoHzD/EvX6HSqAuhLZR1DLE+NsK6FqU6nFf34aHbGJX7oyskaiRGFCoWfL
V5zWRbyOnYXXb509MqkkcGGUxBqD+H7PvV9CwLgngjAsrGC7oAY4y4ZBP1VTh461
/bJVal4HCepLCT8pM1hqGc2ZnQTZUyAo0sMSgz8D1DviQm2yBafpNX68jilFM7f2
5wgXLOz2P0n3ZPkEKaKo4ttVHXtD57x7nc9Q3xdNgMUVTr+JHPWsiA++bQJ91U8a
hXJ99jcWiS6jNqAYrEHH/pbFg9OUzTsZBALBuI6HjuWEjHD4dAWhvJRv+sO5mVvh
/VrRVugm7UC/C//CPHvxy4p1x/OustU77OMnvicAeDgrPbUJQVzfkhCZumA1LiJX
UB+H570ELT3kRS2nATJ8zfMAkLtdOrUYJNlceJYZapkAEDepX1OIfl7QPEUlgcWe
LNSs9cfrDTHQTsXCWIFOMogqyKlQj8g9Am9ougWNq8b9A06+w424xkQ/QZGd2XVu
ddbgN4+K7dEM2bM1h5R7SFIM5p7y+Wg1RdaYyNMtc2hgsMeDVSmIbkfxY+P41nEZ
pmNu+wVI3Emf1qzUL9R+Ju/w3g21WS0uOpN+vk64wtJUOsESSkzm5+jJFUu0EyeO
s+shtuIAQ1YqSMuy4nO/ASIO/J5+veFTlGDS9zsemKTJrZuo2UAuGCm1qKY1wUal
WZSOe/wPNzXbhwIQjub+m9KUf5QKqBiXCQ8EJ/xGfBG0KTsaEleGMVsHMfKZdtYq
rh/sd9mI3mFYXY/AiE4wlY2U6jmhAUYYh73wgso8SFSRkNBBlrlv9TrQMYEi3zup
3ducGK2gjKZ6WvGanT79bKRUoiwlU3L11BiMCaFUNIR4Zn8JhhKv7+e8w+ZRzqY+
QYgCqCr+/l0Xkxhbwfr0TkOSBljizxdB6y71qdy7UQwhd0qO91lKWqnG4gwMQ8/E
sN42hq5qoK5GKZmw8itniWG1SIndlqAYYYzSgOmX3abgCp++fyzCVXfB9Lrh6IUd
DTEdp6jIHkQltaJVeSfcTkDN3AUjpoDVCOn2377rBD47QOyAZw84pLTExjy7Ld/O
ldwa/wNuwyTf3pN1fT3AEnpuA2jJ8s1nx5hnyQEKz8gUcxJit1kkIae9c8mzJxIV
nLEHCgcpd/4gHmP6KnzJs3POYB9ZqFvmp5qJSVuM7Ky4zzlv181Fq+8Q6jcICpOp
fvp7HUTuUPR+VDKmBglJiqeFHfUsYcdXtPa5UehxghTZOCZTj0LhRFoTcSH4gxqW
vXCGMRPH8XPmOvQz6tdg398H24xk/sK5bbGRw7pJcKlxD2rvv/UIUPYmmqsIfh47
9sMc4iafoBi8CY6uJP/2ZuAGKh2rqbOaJ+ON2UgTQVQGz7NS2Bwajl0O/cjAcVUr
vCY0cjrICNMc2a80U9CPn5EhVIfjUlm20023xObT7ursFf5nYivalE99cIgogF+g
/pMvr+b98MzB0DGtjdh87Wf3cJivVaf3nPoBoSAKV94iz4T7K55FE+IWgBsnWFvU
hWV8V0kgRdULs87GvP4oXh4dj3y+bCkN/lpywvnaVAQkJp1u+wBbEh/j0aoDvHZ4
dkjszmdDmDs2t3RZZKuwWseHMQ8rzsuEz9R9bovN1di81Np/kWfx0vcr9RK99QPv
rUielco8FkOov/hLvJIooLmw5IrsmS2ubSYUEucNn+K3CYSrHw5cq6YcxOZbiVp+
i9mb6BozlFVGcr9spCUFKH4VhEij1KAwFCKkPKNSGO1Y6Vn84ZdBojzJEldBJ2yU
JdATawUXXc/ihkLDZ61UmmrPNKHdyXXRgYEE5qhtC/TUtX+uWYDKw0xNq/wb3tel
PItPuvkCVJHnD2b41EkMOZQo4T+8pastnbUO/o6L/bOuXYGN9ZpPPCrjQGKwJJZx
OsjFe2a9DYmFzswt5/ZG2Lip97S7xO8HE7Q+szjRPKbENVc2tHlLVHLH0/o19ONg
iVSdR8bKRDdVdq9ZgHswLY+RqR9dY5vKyGC0dUT9aS0ZmYefEu0bEyps4ZGZIbRA
tP0CAJWw3KgmGdB1Unfhwy8bKxy7iB4tHZWJhPbcrehqCrFjzHLcJiOHl4AZRKW5
A+Oj20DIfZsFuHtaNEu0pc62XbN77SzV6xE5ALhydmZTu/JxGaryaPc6DV4/8MuS
SVYYTeIeKjJMhHMLMuWolxr078WjDlCMishgpXt8risin6PVZfdo4tSgeBMeRQUR
sUvr6vHrsIEDHt661R6rY0WlRhKuMzngKEhzKqepzbfB4NV5BEG5+t49BQ75RGBn
+CjzWFxx0dU1JfFU8kZdEd55qLvj9in304VI3F87VfozPcThtFskL/kyiKIFdzh2
XtTyCxi2Rw70FKWgBVT8yEVSF9p7OrBkQ7WVG3INAuZUMbpCuqQ7MJguY9L5Pten
T9igxA2X8iV6Q90l69g+qYr1Mh904Nl2dzrikfszqVR4MqfJgPD/OgIB+u38QmO1
3OMcLzMJUAzLSYo8vVP2F54ch9pAQf1nK+kbP1Yz7cI0NcVtVpp+/TTw7vDPmzfc
9TGVLrmga0FQhlmceC1Reo254g/3u36xlpuA5m7s9c3vgTp6DD+pl+yBJK5kOklk
buzzFJreLaWbGjQVDth3jMC1TxptH8UDCDw91uEJgZzu6HKcpnfar2zpZi2QfBlx
M8SK4nwmd69/fVULAmJNnDTQ2WdLv/MdXXM/h9/5ugTv8T0hm/yiT/y/HiaodqQP
nSb6VTvDE+eR5igS8VHqJ+c6i6Y62TnqPTdrFasStJYbma4OZbs6qkbv+JrOdMmP
/4qukUWL1QCOqUPJQmMCtWBGqWBap9Ji57IdXel85qCPhLhToFP9OVrzIi74nRcC
NBIF+aUy1dditlAPOs9xUR3nEhrg9uYZ/iDcVcm6do2SgOUZGaAtNPUzwN5wcx0e
ioryoZ1no/+idka/4UZvIKLpx3AZfoB47ZpdCeWCP8+TmACpboHsr1Sk24FMA9ka
lQhlDSCU4RVjZCfRc8Qvbo4eDOd752zdwUliQe5GOZu2IXaPBTi+BAFM9KMkF5L6
TnJlDVeap9fNvKEoqzAryZK0f9a7nxZPrS/p8aketnBuRMReZaDBLg1XScgPLSeQ
X/t28g4KbuMPhxLb5xUo3iIm6HFZ22KDReMSVceh8J0wyUm5VHeuDb59Rl3AGO54
N0QfbfLNniHOWltbJaGGmJHTZDmWKjfmbWEnvh8zosxxq3kYrX3BxA+ZXVyEMCgD
U08f28kvMbqEREz10n9O3+tZy817+MrXXzWV0ln28GgTOtvfPHG26ZroEP8o66V0
Bf2iKdD+2Z15Tpng4a9vV2EFI7gBDEP0iWzvzNmfX90FVQy33CrymD1ZQCW9H/HU
kkByZ2kGlXlglO+5Pg7uVHClPxYLuRysPJ1sRkYTMLMqQpZShy/qX3Kbl1edqr71
LXWwPWse4WOXulZN/WhharFAyxvj5Qs/0qCn0ZTSFpu+jTeS1m3jPcwJ0A5KPRTd
l5mdFf/fKfNif+NR7KqT5lh5mGYjYAzIFgv4TzNx/kOJpG+ZLw3hzG6LJ1LI0RJJ
SlgvSprs9ceZ8CgkeZQpFlcGsdE5fhzgj+n7H+H+JUYo11fDwntp96F3q7tzt7zi
u3u9zaNdF2P5AsaHnYdgkeds18slWzRWycaAiHWca9cg3bGvH9numEs2KKJtsjBK
rIT3rZG+oP6MZU2EPNiVPy9Bgr9R8+iuWxyQ9NF/xSTs5PDm08+Pzs0gEIWCHGZC
LTk+pDVle3eLIJKpwQwjrdL6u5suPszpBOC2WJS8rGCGZKTun7SHNYCaqfLj3OGL
Uq61BethDD13mAzGAdZtLPDHzUO4UXqy7GSY5KrSubZlIvr29UVuimwnSLL3/wHM
UuP/Y6F35P7pped9dtBRYS+1Omkhc1/YHhdJhppvbwgtoIM8+jSu5m4v+lwRD397
UqZNWaWsuE5XBX4hU0eJICOJf901lD5ac0FPqRG2ByMTvPiGBuq8t6PLLWTw57xP
1IrLFQxm7JUQ97jLxHnP4JRh++obEvaBi8dok/TpAWK//meubIDZbkLYytIc9p/G
UDq0k50ZJvp4yMGq6IG4iHw4U3wVCPylxB02PQ2aREdZ37sg6foATHc4RCLejXz1
3nSIpPs1MWfgltR5NDPk+z88iiDYakIqWMQHu3IotijMpBFrnfsrDNPCveZFwTUT
1yyFrTOU3KnnbdsabQJ0jc3SVkTtX/4rudJ5diJy07+yn0U4H9Ybu26zfB1DyS3Z
1BaB19Hek4NVU21le9UcEYtf/WqTayte6EDnKReQVlMKjD2vJhnnZarlJXTQVi26
viXutqbT0Crw/L1Zo7lG0HXGIRlbtx2sExYW5UU+HXAFnjkIVPZwPrOALx88Ycur
9WYJeeYYzioo4nM/9AahcRK8J/HsaDCuueUGgrz+Rhny8WcJlmy7vJoV4a+KIQvG
gn9GM6vEjnu5QnKD4bp/4wKa4DwwpZgdzTCa3BazqY2p5bvR4P/Vy9snklWnWl+O
/CJOp3Zz7xqcqIHZvi3qEcL3B0L2h5vMkaDscRqkGHl7fmRZXazz6RAsYKdmSji1
wn+EyO4IFWkB6lxsXzMSyE2zfDGj+ATPtWVJyf7McuqRS5vuyYX2AnRZXfBDiMb8
LMdSjYWtSJzBM2TlxuOIG26OReH9mF9VVt2kCCnZjAAlBekBQtUZy6aB9o0/qqk3
bfwqCA5YEm71U1X/0KIMq/fEUhHNV5fRHub6HEYL2ePASStKbynXhqJ4sQt2ZjWS
bVDJzcxfDybL2RZLIwGiVOqGUXiPZQjn6wVsk/J1IWvQ2FwMT910lES1Z6ir44LK
HwiFa8kvo7mZgjcGel3i1BwY4em+PJg6JRWd0gl/Mr/GndVa4yCK2kUWX8pCj8zY
0SddI8+zaVxJwyH5heT9qnDEvITwoG9eahL1Vx7x8endY57mshxyPnhsOkHbWLzE
urAbzBxkU6eDv1elP+T7lb51cOFK+ZjhRaHOIO1Bko7+psHlwmzU2O2lvaCKqPXl
vn3CZ+QC355a3A4TEiEM1x/FqVxN7Rtwmev757HhvpM4E4BXC0FiMD4zFgjGZrN2
L0axy3KebjwuPPC0Oc7DKtBNPAq4qI2+mhNmXixHRLoB7ySJfxQbQ1KQq1E0OMrt
fK0dxC5xb/5QyfBX4IlVsqSCWQkOjmpDidlYXwyMUpMLu0GOztBpI9t/LEdkAAkk
49buAJldP58qeKxDpH8NEGtUVuphbrLxjgNZD1KyRSZSGKC+VDvtvcFHQQjNGsCC
zs8K5hFVd3E6wtWoG7gsk5tbg80pTPLvl92p971vo7wrrGGEN1XKIFdxLbWn0nTy
yBu6U0ETCZFDntqnTdA/50eDSS8ane4lmXUSS4hMwwUNlA8lvqPxptrgapGluxIs
9VnaRbQ6JzcLi0DmxTF85IOMp2nHfiYAcOW33Y7ufHjvsW+bFMP3Jaf62R7NU0OG
FovMcJlo5m8YkiUUrQpbIjrW86v6m2yPCgm9TmKW0ibyduB4+JW9q0/ntJkBtQpX
ZmCrJCdosWvmSHTWi6KbSJZxWZes7nXwzAHMDUEnhm9+rwUZwbMGJHj391K5KfrZ
L/P0UtWQPL4mLe9sbM5l1wSvAvQlPGrW/ZRPK0VLy7JJXU2dZBn0DyX3imUxIvnJ
uLGddsDK89Abwmt3kcMXGyqRe0Df+ou4aHsI4SlIQUD4EGG+Bn9wjAPpnrpKIws1
Prk7xm8Yl8IXQe1GYUwep/3Y74n4bIv94EFgFw8c434vPFqyAjQ3hUx2FABnNsNg
eGzLAlG5LnBKw3KQhbQ9yNuvmm+WmEimsBE/q10T2NqF3CVKdiD6iHdrHJ3jhFop
yvuaLDjpcryBKU4A2P7qpZxflE7f3042jCIqf9r90+XTXQHUI5BM0B1a5kiJWY+K
7TSwUdsn+1KCksjdoCdVvafMNtEh1hYUhx2xKh5VipUiCl1vjXZpX96X4kWguQZ9
PnrMjQMqgZgCscflpItJehZdzHCrEWJWYEbwdSIqLRDaPJYBpM0BSzKR3DIa2oZp
bgD9t7kFR3YjYQDA1MolkVHzHFkjXdeyEGG1lubNENLCuR0dRgDTbS+VTu/yfFTY
rMgZM+B/CEBseXwsXHcEDw1QtnUPEc+udpFqtGbQLFjyEuACOb/ObLIZxybKGZ1t
dJl+6KOJKpgKtTo3NVaz7XWlHA8RwKqBH+zdkgI7JyPg6QT7Yy1NFmC9JUS/qEAT
igsEXdqnnUZ/y/kr1hgtqxzsss2MK1xtPmuBA+UBy56Pj5H3Dz1YHCbeYGI5FmNO
M+do8zgCmIoVquNP3U7mJW5A3YQO7WfQujgk74mQFt+kpmrUYlRFDZDkp+lK+Zi0
llnzYTx535b/8uKIh7Rp9fEJvTWXsAFXfKmGSoWbsWx6YtSd40NpSY5BoImKcbBp
6L0w+fhZKJKHMwJYaAi+K/JgkSF3wlp06siCwt9n1O3BxezT1cpeMtf7O6z1ZwQ0
3bLi1HSy6eRRWyJu2harREjqmvP6MlBoSyKWQLpZjezLYY024yGHb7ZynJ2Enfl9
zJbIfK3rgXDsXFmvDtAW+ZshffDLug5BNOW91VOaWTtr73HtVCpwuFUFxHNFvKfF
1+QCXR0xR/JIEPq46i6vLfR0YabMHjl+0InnW3nfF/r/efEPIZb8Y62hSC4MTAuj
0P4yIVh+Z8OjjNEQAZLVZfbW1eJoO5NEwIEliLKjsNKX96jboilgwvKJjDgZGZhA
fhcb7XXsKbfx/jg3iUlm592PB1cdGNkO6X6rZDoYF491f1H0Wv9PLBoJihaBl+Ie
1EjpzeYcGWa12RjrKMqHHaTsp72DEeXU/gBetU0Orbe0SLqSsOmw6ZIwIJG8xvKS
r2iBpngfo12cyGcH8oiuv8GMgZSywhKN3f8ErH8ldlaKlWkpQqUfM3GPkXqNrLB7
fnDUlxMFwue2TXrkc6F8OMfv43pFXFWxcBswo9Z7D6xonlZJBAnP3/bGBQtthgWd
yW6p0vISb0KSH3JppllGpJRXCPO00kHxJDZ8dVMI4+C6t22Xy/0WXwXNbGNIAR69
REramNZxPlyvaCtYyWBls2HlKUST3rUnrvuKSZV4iCQ52Wux6n5nNNHCpss+2pNa
WgWNpEW2s2fIb1D/7DMEUVmeAj24q98fYgY7SNKTu53ikfBo6/C9A2IB9YD3K+Qa
hjnTiWsAcp9sBFaXV9EkRK7luhsD8RuOB606lk4NE9v2+DqrC6e6S0eAve06/a5/
FvEuL+RTkc3mhabgSMk7Giuis6WoG0uWDJGqy5pP3e+HKDRmDc1sLV37H4YDCrHM
F7yMFvXR0aISoa61AjPYtsR1yfgqRna4U40E0ECHiTMMzWrRP2CXzm2I9vc5E4pp
Ss0UuQZH2p6NEq7cmhAZ1XEzsbybnFmt4gm1UmmoiBmXZyQJSnDgxcqTdtDhWMiE
t5mNAlADI+62MUowv6ixSP7N1IKkPbs5BpYFOGvIWkmHrWkdDVVA6sojUAxMxmZg
7YWB4t3XFjcWHranmnK8nhGoNNfYksmiZ398rbiX+wuOtYpQhyzhsPGXRN2LqGG8
37/pEvMLlRLPE1qP8fn4cL1gNxKrPiCNKkvDJ25DYABZdKge4S5TPixHa4sY0Nwr
bXchtoWItCmhbeHZgHsX62jqi/DPSQuyLMgCMNmKmf7koPzXbwyrgBULPiswup4m
G+4QsqZmihfZlklhIpSvLC+t7lPxfolLW0sl/rIO7IVorRe0IoOYP3T1tOt5CH8D
sNAOvL9halRbjQh+Yi28bgA57frjVt5X6rzBqmKSi7JIRAAy7LmXyR/39LK1TM1X
7IrR09HKB4F7Imsghwe6TzJY64H8jXkcZf2QGEM2t54/Nt4sD0zrjhRbt61ZcGgT
HnF/FBt2dtG4GCHo5cE9dlAcxXh+WSK6RJhFp6iLJYZZm34JrgxAaWz6jofRh9P/
8kkGtxIuYscKiweosrlHAQarKvKHYIB7ITNGh4YjOGn7YR3v0j/WWw8R3CrSgIJI
awcgFPAznmT50kdKHqevrpVX82PWQ1kFNlRyd9H60+CUI//ieprBiTS4s1+DJeSd
LQ8aJbVQO03Mo2h2fCY8fV5AiC3vdKbWdHBGj65cGbr9oXuQg+S3pONop8/ePxJ4
S0t3+aYe0vrpD/P4IuZztestuxGYVhTWeS7B/7iinEEBti4sN7EjBASlz7H0pWl6
Aswn9CN5/qW0Pdnyva6Va+nJ2QDfCCY4OXXqfTv0kyDT1Yw5cNgT+Iwtp9O6UpU9
RYP5eBspFon58LTrdpxAKN3DUPgw9iIE60K9tWH8frKX1+altQgthm/jlWydb7+Z
Bh3mho5skEb83G1lr4SPxRCV0fpBiB6R7d2xis+O1QkYQE/f3SxUXKH/Mvu8kTBf
HeoAOslsRUyX8/o1plDbdYW/6L49IE2Tw328PLcOkU1xRuNIvYFsXnQ3lb52ugUr
ZkuFZ8ZMWobpcXFZY76HDgoylHLUlzylAwMEdBhXunPDeuBDoqqNwaCa5/Eo7Ktd
qIVVuJFuVirErdI12xX5L52bVASYD5UC0T7MPK4lcF9f+YwiiQziWBZmKCQpGaeX
2gS1b72ylzkmrvsY9JB8mU5P3RSmf/CAp4cnERvWu1akbY2lbHJzOyn9n3wu9j37
uB+ZLfEHXXh3LmIcF7s0OlpocoRTKEF5etskzoVaraEBOSv0F9x7Y1fbyjRigjOJ
lShMihyYoK65yOoBlnxrZ0CRoDpM8VQCNfPYKO3pptgQPZyMTEZ2PDrprbeoIa0O
CKPamtiLN2G9u3Wg+rQNpfcULCK6HusXugjEEnI7+8y0wakZV5+uoZKztdyPrKnX
IpZN/KWggC8uqtUAUSP4Ya+t/2YeMBLIOYHrkbNC3c5yAYauFlIiRBDdDIN3jsM8
Y/+hbuWB1guICdpcJzyrcvVroQlY129zPS0kkDl/GTrBz7C6Ay487RYyMkNbTvOs
ovCQ7vwY4/I7P7bDotF3J+ubXSPH6BwsTAFutIMOCPQh7j2T3vW9smKFs2GnB0eh
QtSIR47t2uTaIszLbWSR/iJssKcYMyLeHKuFIp7rXudV/kK3BBnkrOkSXd7uQf5y
LCNgzohNpHVHlRsjpFvA4wo9vrocZkYy4Fm3sjAjSFu8F+x3honQxjd01qUKqEHD
IeES62wz7kG4Oeml6S/UjweFn2ZjWoT9j7yT7OH/ct/Nf2opw7YXUL28I6IzpeqC
3M3UQLfwjKjNtDsw/lkBYXWVN1tUtHeWmZXEicA/vfypzle2CIYjxf3YXEWrnjJT
UpAGMveSB6ybr5uItsbzt0NXNdJ9cKgnJtseWie6H2KGe0sm9KddQq4TVKs0NUdu
JONZ8XyNbnhDqiVtsPkDXA/foiSWwuWrifFGUs2wB1DQU/2q12UIYSPqI7EVXCyQ
n802/35fM+F9SYjM7GkWsTmt8LqbRzFQTYUS9FO+4JhCL+QfW9MUjl9E1lxHAIqM
tH7GCPJdCxLc79kH/H2fdMo1VTls3LSsquUT7Lf4vqh+pmlXJqzCQi2QR4s6eRUD
MMrBf1xjmg4rvgWYZRDdBnGzPk0ChTVoEw32nP0pU8gB7jGr9RPAsIL/S6eHWHxl
CwtMkXvPhLEpdPdeaAY18mYIfGrOeI/v6Ln2mgiI+K2PAtem9iKiv1hL3lT+e9U7
Vwe3sFZhiVGhdG7760VIASk1FNp+QI9/WKxbEfbrWGepSpRnn6W8bQIox4BT/dtG
504KxlCb6QEicJC7b5VyCfvSTaxaLpptQKaxcD0sPI8OqrkHWZP5XdwH9JtH3Ucz
cPpA32xdtOwptWgZxddDbPUVedmXoy4D3vGaFQeOPPFK+Fjq1Nmq7VZvPVTC4/O/
t0OeFNOKNN5NTjU120H4LeKLiOYsscMI06Ax7o5/0YG/qjuOSBFUDkJQOXB6I19I
kZW5HITNUUFvDQxtEEToWTiLC0tsQ1j3Fr3nW0kTVPccG82jGHlVaeFGiVuwvW0F
Lrmopbz2dZAej/xI+8Ey6TK0IQ9VC7F/24F4QmCioCbRvabdvhqdMs9WiXpcVyo3
y5M9814HoVIdM20dsRDQb0IkhhehbmN9MfX3QCQ3P+IZ2e27vgmCiMylzTj5sKOn
+GZ0hSqdcq0Lss1QIVvYwNFsW4AIwIt+QjHgQUxPD3oDG04ZdVdhEqvBg8sOgsF0
NggfSkwtdFY1zR8jOmvb/izcXCbtIrvdzt7ha05/bMaCQNPajLzjxW1cvWf7h6v7
Lc3QHhhhvVt/VJySfEim7DW9KJs6r23CzNjamnlRi+g8UmWlIzuvj1vLLI7PRgry
1GFpzfIBcCgzTQva57FFeUVv9XXvtWsibt1SHiBdnRKjwS5MoOkxC2fMXTIXODRu
jlZOlmQMhCbm9qBWtZ0DRMkKywA5Hrh1XrhgVY/l5NNuJrw7EG4+tVIKWlcLm3uf
y6I7u/rUBt+6s35PTDY6OLOgUs4kDyzwDVtHA44zJsfzP0aDfg/We5fPVX6B6gw5
VvpQos48j/sExi2MsAb3o/H9oHyQcIVG9UO2lERflB2Fm2R51367dxL9gw+SEs27
YaNlVqLQlQUNY4QFJtiosy+5LfZxnShFZW7WwxJUS0VQ0SnqtP+rQbK3yMkTSKmg
xClM+oR6YQrK/8cQ48vMDMv/eaeqjE/QZQEK9id1JN6obRTkgyzfw++mqG4zn/cI
PJniYprMMDs17/GN6raymaLzn2767Nall2CJY2noYMuTTPu4EbafzTaAWCtwOcUB
dVNr4Pqy9x4J8apqaLigofPreKhOdlOoly+gz566nCppoUtxmg559uixKy8qV2sj
w2JXT4pIKH87WvnWNTEgViemDkGsLs+NoK2f1P8iDTS9Eaf7AVqeg5tlxbcQa1Qt
fwDztOS1c5FVoP8Pn+hjGob4pyR9k7zjZ8cfdHTNEgX2ZUJ2IAab5/JDhb/kw/RL
QoS3zTfDZuzgRUdr6XIRDSCKn7pZTv9sk8JxnqTHmJC1JrC5eljp/aM4DaLL/B23
VLoMpfgPGobNOceD41LC3WC8MtV/p/GYBOwvz0HOY28bc3ePI1nR3/nn2aqTC18z
igV/7xJ+D5hpdIRlTN4Qa8p3UGcDubX31YJ4aUMbHUWfmkzOdNj4e6HSmu/XDYYQ
9WhChRqawPTWVd+I9ZAxQjDEDWIO9udTSa7L8SiZzmxNn5krasIqv00rwOQcFJwX
RyDn+3zYcMba38agUszMuLnpzQ1hOiJgKP6sVi5IxOK958McJUSyhCa6LMqz8mwj
4XrqxAyRqRB3/o+wm6FrnAlXlC4Ml0KaX5BYV3nMFjOJk9lKuiA13uI0o7ojO7ru
5EOLApmycdwc2+56I+1hYJaaS1hQXHLlotH9OHS5wtOLrSU9WK6xv0mKQC7mGJDn
Al4g/m1WLaKktI1K8x/FJA2MotJ8gsudxATR7sOyLfc/ODmyy9kjnRAZlj53YaMe
E7/yHyOphPbyp0O9ACwRSMSFY/pV0uVI+rThN54kkcWKoWykpmBPKvuqaElkuxQo
N0VXgQcyoYsDdbOz/7MHCVtu47hIowiRT6X3NoXLGEHCiZX1Aza79ICRncZ8IlSj
gkG5stLHu0++ykwggTOWOxtuf/EuvjL2VtSUKx6JRtA0gQ+dxiJi6FMdoO6k8PqR
o05efaXNUR8iAToLIVAsZE3tV8phCqakaHtr7diUlBzUVbZ4qUhG5jtdfS4KgK0m
DKRupq9z2UKi3Q46vqtBnbr/TbYiX9MaC9Ml8f5smXbLBe0xlZ0v5dbDKNtzsld9
sIKxsUj73MV89B0a2EHeQL53ukPrU5oLBcXmgGC6TvFO80aJ2bQJgudQwJkI30jB
diK7RqCQI6TTLawVR1piI3x9gekmvnVsTKHbAHEqastkmoqG+u13WdPjbfvUjwiI
45SL4oS4cMFhtCEtqN0D6RnQru3CcnNXVmIKMv80Sy8W9Aswp3AEXx5heuKBuY7+
uDYvseK3Old9Z9TKP9bj/bgIwfsGDP0iEcnSTXWV6Lnpp8xQ7wT1hoxuh+Rc1mVJ
kZe9obQDVn5WOzj1kjm3eTzw2Qx5IMH/UFr0OX1pNOt09/GFL7/LKSxDJlv1G8SI
LjjJyZnZpCJmZoec/QrR83xBXKWNsGdcBUuVyTXZ0zAYnwV3ZzMhyVlEEN+GK3dj
xDwkAoMIAs4NsX1h8SJCGT6he4e3ITKEbVZxwmciD2/MGnVvL35kye9WZLRpPvGk
qqOg23U3REDVgGi6OdAIrxIwvB+MWl+UXg0hhDW0LO9z5YFAV9epIhMu5NHej3Ae
RqD9b9KMsmr6NYKD72wxgYq3x1rJ7OMO02JkY3xiCWs6ebF2/XKg1eKZrdjGIC64
BqqF9Q0eQbA3XrSev6AMSlyYMtMGaq3sPwU29qUMMAG3218q8sUkp18Fz3Zb1OpK
OejanIFNJl/TINUKDb6d8V9MMQVd5TrTnnOaEXirCxPDF9luX27QnuzXwFxUKfkE
/Y9yyBpclH35NcS6via58B/mpuWW+twQYGtvsuESmPxYqS3WRdVq11qKQgRoD4HA
7j8QZEdhF6yNPYrRygGLLkcy/+VsWJhB9ymcxVIX3xpIHt6pTC4RzJ+qS7Bty0fC
IiiLrU4otpPNSLVmaAaFh+b236lkLcTOPzuWoJ+7YMgKSwhvjlGUWX82Wszjc89L
2wCeR+6pEqO3vLaavppVlVTzRFqx45flv9F6pUg12eQqnZE+mdilgqGZPOCp7gqt
474Axpr+wWd+W+7DWtLQYBqCaTrbYHEBVPc2HvWyPouuXvqPpQKREZO8EPvLZmCc
JQTg+2waIWx5Seu+wE8ljbx5fZrXyHgokxH3hTPgJLd5FMjopm16MSOf5InrLwAN
5R0T0zHh8ZMHpnPfCJXKsy+LL+AEkRY2vCqpwrXZc6vhn9FEDtQFRjM4PC27UWUS
JMi5S4NpErgwbKKRebhoHGBdCWzKGEOZGk3sZUpjBP7tV/5UhR0g/NW4FabBzD7w
t7uOvOG8SYliSmHpvRXMoFJxARpXdCvzZPBVhmhaYrCXRZP9EoTMLwNbsTXpqh+r
/F4eKnhdsFnyFiQQbw6VqJrC50/+MgOtxu4lMtkBf/QjUH6ZZCP/Fd+W2WPtKVvo
pDLJC0q3s/lQurZX2LtnLyGPzXj5BDemDsF+brwrvDogENIOKiKa0vOY5hcGswl9
7ULvg1hbSMttzwiT/XOcUt31cG1rukiuSGfSgtzG/MagKqknPZt2Qm/OLwuJx6Vf
3v0PGYfv/ItK97mcTEi54551VhYoPLZstyC8kzGtAclSXJtT9lUNvt7XOQKTN/au
5i9yScvgSP2/hMpjDA0Ox6XTndj4MehsJc7X4E1i6g6yNlI7x2pjozjSsrJeA0JX
BUltVIFw0MlZO9ngvUPExKwHdFNv0mikJU2e3Vw9T3efh0a9t4Bwd901/Sl/mPkW
vsxO3Br5dEIN5jdy51IpyWJyQiyWdAfTG5j5s+nihAcfCdHuxIUobboYHDQgT0X7
L+nn1oHSaT0IKfmimrUyLjEYqs+EHo4jgc6dRN3kA4k2MSzhWxYdXbhoIiRurtdk
XAWt2DjQc4/KLZY2YHl+t7s1d4iF3yrtBT98TJrdYMsNphM97AuP4F23TH1nWQGz
RPgAcJzZ1dlznwffn83c2Ois0lYlYAbYiC7s3GKg+TG3cpCt51MNNTNRwHqaDmiI
0Y7WDEwa6pRbRjgGq/oYfwnZNw9BTL3hNgvF3e3bzRBiiyOmH2Ay1SAWL4Mz7AyF
VFhsO5LTw6szXrYqc5XG1/hyh/5+8xsuYCnqvJ8ef3/5/UqrcTg5pwM99U6pybTs
PXQ3EbuKRUiteZU1ocgyEKOWsTELolLUUjntnKBOYrsYrk2hfhCh0k8RDuQ3sXzv
2+5fLmxICWqa48pMrjf4ZeWy+XxJzrmSY+HOWHP3gk3JSIkQcE6jHZPX2vKeGUYH
DilkkLB/uKwNPXIOeJqAbfnJfvVCwzwhFIoq6Lr/UlgU25c8conVxpZX2s/n8OgW
HvCeR01EXuhiNCUcr9zM9pxgEflAy11fjIsaI3sQC/irLCfHiyWYGDz3YHm7Q3Y3
09WO7uUM1W8/Qk1yjXoDT4tBW5hLfi2ah0148YhgfO3IBx6gAX+Pg4YrS+R1ftJu
ke6JS8A8QvhZTqkyVteB17eqpFEivSX/Mvo1x4d2pAmzVZTN+DTkqyMc8qYGA329
cO1O+s4ENTAO7e4iGYF7esoi6jo4h962iCxTvakNrEP/8lxGG2fStoKC2J7ztclR
kk/sHN25Q3bSF+fhQGtqbqYx6TPwtLfHZcW1/BaPLPgtdzqfzQC7Sy84+l5HHbGW
LSl7TCwdUnu38M0FP0SONx9VK0szsCH4bpHnYZC2RT4zxzVylCBFRdsttr9XyQla
5ovEgJjTcz1ek8tOim24hfRa1dUuArFu0zPq/EraEKLXZcVfjMftejOFfRFMkH3/
PkpTwqHe8RW/BXp73EgKa2/UEQ+R77i7ieFUvyy/nLIsF7iZG0klr/27lSlaza+F
3ZCusUR8msWhOOvWQ+xvObGRkCC59M76UTDjox/jEOvcBngyu9SDAi5vPFArK8xF
6DHT2RlngcKD2JsBKLSnQ7/nauaJytU+gziM1+jjeuPbgZbH4KTfFRIwDwQKQS0v
x3jj6+IgTc7+2S9/iyyJw47YyQDgvX4W/e7G6+xAF8I8T/NyzFPaU38aIDSORwki
9QlDCYNsKFvoAzaPEoCdS+XbH7C+pys12oA2l2OPevBxHJM28OLTLcNj6pLgl9tT
nJ81jVPI10h9SUzJCICVCHph9YHiLmz/KnUID0axWZvDBAwHwrh/9jLJ4rUvPcjS
2xunXZ3e/+MShXFMeIw7l0+qXXYzfGKCn/X3Wv59Ucue/VLOYNuPIrAuNcdjr6im
YagI5OxviUNu4l/AKtPvm9O/kg4dug/3Pgq9Qra7JJT2wiCtcp/b4WJ8ebBgzdaT
JPtdAB+pjDeADWPQCoW3V1wgD6sZc8R2vVc/ZUV6YeiCmUk+dld1//v+qwQdQpNh
Qwv03dw7iyTQN5Y5j+xrXWqrmFEmLyH2H+3bQwJ+u8ErR5P8oTeGJU8ahO7M7fQQ
xPoJN5FiSCEdeai9QAArLkP8DG6PvhDDWjn+xGbtZCbfU0arC5V6z/rdKUwWNUq3
Z02fbfZn2LOUGzbvyZYVUWqFJp8VKZBqGVPmy0CxzPm5yt0n81kAofum7TZ1zUF4
Hfv4khUbotaLN2mmEX5KI6lqBVkmPC23wyaBa5dkep7O1AqJsJeyrYHuFpMknsd3
W6S6kKAAe1qhV/H9McwXsPygC/s6wxrjS+J0FdMrZ3wtcrMDrYaj0s8w4bJJdIkN
/SwsjpRItSp0JlaE8J68l+vshj8jb/yMiyOGkLiqmhNP990lXlcB6SCcHQSgx6lu
0uhm3Hviu2UXp+N3oaPoNSaFaxiEamvb03P1dHlrYxXKUovxbuAU1dABk50PJ7bn
cgygyF2P8M7bfVpiFB59mxaWZO4JC4PB8Z3cAbIj1bioWA3hvix0P6/4YmOZeO/O
nC3wmBLn2R5ECglAtvZsZYxcapNrIdzHQC5LKv27RKbDr452xjlLqXzQrEltzDNd
VF2WTEYk87EXJoyGzrA5eCjSHq9lYJ3pwmhL/HXc4DUuNe0uNNUQ9AiLzFwGy47+
u3f4qYPjCVc29RvZKMgR72ugg6w9HRcOf7lRj6SlolVQC7g+DkxxYbuUvMTMyQGV
YyxMMaQIhWNpIoAMW67c/QSqXb0nRS4hxt4eCU7wWRjWc+LeNsJQEo9jS73aGYkY
GN2aQtUqUbOZzxPR5bTVec/UcIQIWiBacXnOMdmAKjnLorz465rjH4jHka3AHzMK
YBA0GriMvDy0Va4yQHKukgy56nN73cn5P6hHjMxZJOcNPouyHa7+bygdg9Pr+IjQ
N6XpjwYq1CgWI/36v5qADwS2/oum7mE0yk5PXOaZPu3+D5jFaeqpE9WtwR2ls14O
ODydSbZFWJlGS+Y09NLGHfuilk5Z9VryKhziAApkNgcxL7p6E/5yNHUn1wCqL/jj
XuIR3RpEn6W47OFNo9vkenHRUhSGnPzMBgmdwmkWJU0+Zu7d1P2qHU+oAuDLN5n5
2XDl3u3KXVJJpeEks56mxpV+yAeRJKYp7xexPmujq6Qs1XXKzUk9xfjjsNevdQar
Q0geqdJtd46KJ+G49D9Fu13UYRofSaCKt2ramXF3RMpdJ/SQL1DVM9ouwdICUT0i
RB/y1S3LRom3HZDo8z+Oi9g3Wds9hGVGgNq3l8PLkZ1eKxvZuJow4+RgpI3PXpfU
DFNpwKDYYhpRb79St7dFoenehOkyjaI0jn0iE3j6PiPHP0hfHXqlhnO0U/V9BeZE
c+Mq240ozCmUVMTCdoGC4hPBxgy7oJvEmtIBeP2xrwFWLgv9SG+98fM0BT15tlzL
YUI78BDnxy8nJdM5nrHZr3sEgkYc2mEDHh3g34iZ/fuEefF6S/OOW4JHih29EvzR
dWNJYi1TEULne3eTugc+O4ioz8KqaJqzY7PkA3RIl68H3T8w1LaSwOT8so/ktS8I
BBy1Yn46cn5N8yGuivigWq2QycK/l4fjW0dtptX/DjIKpOrXXlNhwP7jRHkxOLNF
3Kouwd++62OKCq7n/tZSa98nMjYvJ4cR/OmVMqD0jDv3N/Ff0j6IkONaKSkJZbEJ
r8ow+/9n0qto9OYcQOaN4gAP4DiEE2Ih34sXGaC6wvjiH/s9v6j41iCtRbf6lD4o
AuHlak14LjzH1o0DlQMNu6AtpWOs9FhHZiFAJYofKCGveZOrOGzF25AGUbN+BIS9
1GDD/CJ4F5WMoBvoyeblACsEm7ZRAJC7VsBDCwhWPj3ZSDJ5Gz+taIqHtkt7PfUc
Eu/2YV1gkPPCxb6STFg6FTvdkeBFsYCIA38Z6ymmoSLTWHWLi3YJWfqll1KsulHQ
Jx0P5/Dcfr5tkYTIwbyJskuPwT96sE9qdS/cOJPqv+mhgcyWlxUrX60vYkoC+l8s
orOSTTIlQpMEh448rE/0xQGR4krCX5eXdqWBdabpbwV8OoqALOiFaZzwZ3rweFxI
PJ3myM+UvgJJmX4/u3N5Aleef7qMJ9VWkE2ZwsjfcnSlYXta5SVF3s4wVw1wPnVP
i07vZvrS0g35nYQDwnZM3GZLb86D4zbgL8SVuSfpA2fvVxbmhGDwzS36n2+TDYvD
FxJdbCtzFZhKg8eBzN1mQHQg5l84+lyY7+rnzYzZWgdyZ+MP3vrYlh49JhOnveo9
KuS2/NlwbbfdrUB7xfHzabhrZzqO55lYQdaz3R697T1FtyASlfNb7B4V2Y2EMmoS
ovAkMY5sr+2l45W9rH+ZbP91OFuPK+/tsXljsp5qE4CMHv18bz/qNZpM0w6Ov4i0
KLzPCs+SzfC/wKozvqg8LCpznUNNojmTP211tTE493lAEIRS7XYTROUeJvN8xWy9
t5lfkt34jEeeJpj8xdZsqxXItESWJr6PQMFUM+6coLRlZQ/EUCjDz0JaHc+BvPsG
g7WCoR78B30U+nHcaNNloJvLBhf8a9PKLQwFULazxO2ox9wpMqbsfdyiLCpdwZqF
iu+OeT/vAC2xSRGMdvqSogvWna0MFvScZVBPk6cYnc+1+g5sRTQHSPrA1Hg/86EM
HVJkl02oq2I+aYSMQgUsD6gxc9plB3V4t9FSGlWc0mXS9OGW8lTr3J9CWV7Coao/
x1rPmoG8GeV+7n3dmUxq6595C3t4dcBR9egnDdJa+SmAh5wNFmhtQqRZkQ6sfqvU
ROYwtOrXvbAkX553N9uwn/m826KTb84TuPnrDLOa9s0R34ZqVSXmr862hlZKEILp
nMM5waWtbXcKiQVLZF3hfX4H5Ch7UeELVzkfVEQbJufMNVrcZfEprsVFCUPTtw1D
ItfuPL86pm4AOMgrfri1h/2sDxEWaB8kkYC72WYitUJ2c7CsdkE3E5F+RKPO0tPX
RsJ2Klh/BDb8bxle+PZRxA3xXNQUE7Ic0esGucRmcUjMsbZ5lUVOA9ptXuDJjWLx
34cGcKdoklYUuZRGtuefx1JsMEezMdFuF6srvsQufk5hbOXgV4hP0eh/bMhbxMEU
ijVCiYCkZd8K7xW/unjGdmbAKXyQgM9ynAgLV19DLHg3BYs84saOLBwhjr16ZNA3
9o5PYso/cUpEK64E5y0QsLMFnt05A1a2K4DMwEJD/5aSNs1uwelvVzEjxJDHG/FW
Sz3W9QUvc2j/YY3w0lK+Xs/E0k2O0NbU9Lla2/QFV1CCNgJdOxdwTOrnluzxGLoO
qEdxyX8AL4OCrHk/cKqD7BLlSFJelLeNe1K66NUvDT+apjKEvfdJEpTGpARUeGLx
WIFuzKcqbbtr0XAzUNFnaKzoH2VJ2OXBuVX88Iz+eA394UomblZkQc17zmrpdDy2
HUV4VHK0ppN8ZK5WGWyRtQikE0FT8JitYQ29RSqHVdXCEyFDgI3T9GskYiLcUFM6
eS//1AzXIxANzKBi99d2G4Q3LtQfNPaLNDIMSHL5li2l3kOQvpAbZ3ljEyRMKD/o
2gJYhKgCMo6p6tfFKmMcjaMw3ifY+cWBotipjcUAHJXHkDqBtskQevADsWbjl2L8
/Q0V1MAcMef3D2zf0u8FFcwxN0/Hy2chPwiETC0NGIdNvAzx+Km/5K6FVA0x98jx
fERn+20eS70nJqiygXYSYpFHK2+qKbK+mSFTM2dmhmel/cglKqvM6amic2uOmyH4
zq/8ceqYKvnUiLwLCf9Q71UH47AcZTBtYftZC+47/mqU27MtwWgB+vwA4L4eh5le
a+JmBR43ca3H1JMs6xGNSgkPkaPWbnp58QzhQASVr/RDtjjn01EsVbPtONO9k256
UnUsStL0bcXp8HRLtZQrvvzDMu5skMkd0ioFQvBqr1gNlIvrP3Jox6GO39gf6Jqy
WEzwJ/bJN9Xc9bx6sh9C0zwLZyiJbER6PAi8Pwpf7ljBaYLh5JypLWpcE8Ln88Nb
0fZmEyS8Nok4HK088kLArZrP7+IIAc4l9DwV09DqQpvUFge1+EnqCyo9utqDkTvt
jyJRJXb9jyQNsaTtK4u2n9Nx+yPBB1QrAc2xFvH40wafaTayJBWew8wfn8faR0Ri
jATkfwA9FqYHlvWp9kPeb8sBKC/HItkaiL9d7GO9DdH1J1AztN0sosOrK1kt+deq
Owxcr6tDoTP1jzzYUmiMJLh8LSOgjoeeVFWWzV3bCjS6AUEa+S641bUdw87LW2N/
zp406c//ZL5OCbX9KJA0GBz1oZCdrJ4/CsFfBTJB/SQca58VRn777vR4Lpn+oUmH
JdGFOz1naBwQ1xEqf6oU93Ic8VUxwts5xogGkYfXuuZ2ts9bf5dr5qlGNBAYGo0f
GEYuhke/L9n0uQmbv3GsgzCDoSyfWk6QWK1/aUQBXWmmp9lbZx0NCybfAjhQoftJ
ZtaUxjt8ITTw2lYEIb9YoUmRIOX5f41nhqgDJe2WlqSmNuUaqFT3d/sPQSpLhFHU
KTY0Dn1pmx5MpmA65WNsIgcCiRVYjw9QAtq+SiqT/m1kci3yDRX5BpNdrQOxu6T9
KU/A18PQAi2EuDskRgwpGhmSAaDNc+2YUlhXtKH+QNa/SW0Mp1v3mfHbUVCEmYnR
tXvzGZ5a7GarrjhRC6/dDLdjNLGZPxXFRWgnG2fZSHXriZ5FFuTLbvSHuoCvUVUe
pM/dKXCxains+HGAh6ruM84IpSvIgz/lmbKu8ZZIJrhP0/PMFaucj3yGztDB5Jq5
KApw3b64x4nUUWNkEQsO2xDzQGjm0F1h2qCJKmtp+5oQPDTiOj+kthnwZ24q3XFa
wIsDoBxhi4gOreorbOJDHvgEW54C1L2rPzg/j8bSV5upIqgD7AXdjMlTX4U2jiDH
dpS8fZLjpLcNh2jF7AFREuRnjHtbRFNo2ANO0SyUEq4spMfdXkWTy3HDi2BsmZ2C
PTqigk0k+uaQhl3U3im+AWlzViz/1c05v4HdYaAr3tUuOs/u+QMENRDGcLLBEDK3
zNk1CPsSe6Rq92zP9goT3iAFeIPwlvg7NFH9mqNPVegtXzdwcVsmwz8J0If7MWfs
huLkS57gmejIxFJiCPuOEYMsMWg8a+hIAWLQ71BAdlAzgi+JcT2WUnadRVygwxq8
EC65XBNKiQGWk2yQgZb+WGEQZyfWVapHg2QJ1tcQ5T1nSrMs+6Y5/l5pppufPIEf
h5nE2rBCbBD18Qzvc8FCiY13K9YJhFPT9JI9ZpaWPGH5Ab/kcnn7DWuLqBjJB8FU
vOciyCbCbLMkT9t43YNKivANfEQilQvDKMnX4GPq8JfiXw/Ov3v1qQ0NpAbpk6yW
brmXyHghU1Ci/BQnqeo6JULtmg/RMuIDjOyuGhqyWreraEaWj8L62nED7V4nYoG0
Qt/Y6WO0T7PDeA2KOXEkj8v7WDNYeRk1+iGgi9QW4DYELzy3sJCeGwok1UP9nlj1
/HsY4mAUGLC8LPBmPaDIX9HXtKeIAdRD9S3VT9ikFuouq+ygXA5dueqG2wqwY2ps
KoOjsENmKzdGBvTkY6f9V3ZS2VIfkG7Jn5l/YqPNc2tInGg4giIIjo1026FT7GpB
CEWZyWcqeOqmmqZzmnM6Knq9f/XnBMCkzpg8b58DmMfGwZ4WHzdbwJxSEOInkynE
FuKe1glUNcpb32LkTWrs0O2K8RTwAxtjPi/4hMVllrfn47frbeoEuCEhbtNm4HLP
VCmkiaU6d5WvmBQORhs+qKFbwHcrpukoVDBALi9EELSocbwzg9hJEjznr9c6lPYP
5TY2YOP4hO5WhgntT5Bhiipe/4am2gWXtCk7cj+DE9M19YMGhXObk6lUFcSyFvxT
ncsk3M+HVkFgfaC4ehupaNgIcYbcKDjRMiB584PttgkdwrRHdRmBx6sjcn0VVOHF
c9ZQ6rc6IInavCSqnjKORZ/6wo/SNCYNY6F2Y1ioTRfkkwW2gp4XkWimgGLN0BEK
h9sOWLgHq7KUSEqN3A3n05Vdrcgd9Lq5S6uRFVTT4wS48+1sIcpBoN9x0Xx6gVCU
x5GVHQdD5ix+iB+d02D90R2WPaZ/Ahz6RQy1YwxejQ94a9FIhyJ3gqUudUL5w4ze
HMcHNF6fvh80NcQ//StCi1gLw6EluTSYIFp7VqhJICK7vlPO5kpXJQfpSUCuL7KR
fXDTIUvEXuF3fqkstUZDNb0LSWOCSBBs8wtWm7Fdds1HuWn/EaoAAWcaIcs+nMHc
LplSWXaKK1iEMeTxB8n27Hz3R45b9URVVzE1caV35aSZN+WI6ZRHt4rOIL40m/6l
p0xAbJ25KqdLuBsCUdU/wOYgcrMGqXbUf5t8oy2kgRAV0x967+WsvtFoiVXl1Z8N
7Jced3wKi1zdaO/IQiJWtuRncpHqyOsgSN5nH2Ocx/VTNqVfQewNp1W3PjCC7JZq
Tpstt9z7z9at4mSEfrGMkZfSfwtzBrvCFkthwABM5rfxk/yc5giI3rN5Oy35RFIH
/M6uyR2ss5lnLQoSRdJq++STKxpsPrmvH8yLqVgrEaQ69yFDhyTn3+pafgeH59s1
CVbaUgcIQjqpOJMfaDi44DKQSeU7taaXdwXZInNONHljgiQaoSnhNr+wJaK1PKR8
UET3m6KVAaiV5xU5uq91MaTH+Uv6BecmDxhfg+SDMC7pLI5ejXY1gpEhUSmu34k0
y40SxtIkUHa9iLnEnpJIdVcjG1QDKAEmvw1IVt7xIYCsSSZ+S/9lp/tqZPEnTGJK
Mgh5cugT8gbCv15dguSdE1etf6t7TORCLzeSR0MYgZw482v88GTHEincrL381g4T
gdgl77e6ACyvbKlJtaqfU5qDvNI1v2EctrKttaCT1s1vNytYCKawoCG4Oorn5s/6
fyP/ppVcpPtjYNKXzOT6IWRSfiQu4loU1+YWlaN25qdm/44KL5UGfBdU1pv4NmwG
mwU85EqMPp9KBAdPVi8ngqL9olkldnfMR7fQKN28ZGp/cQoTP4NqkH8ikl1Lsf7l
UnPSZgRkghp9AmQPSeoGpiGs8Ud/Qi62tN2ykl8Lwjw2YhrVdWlU/3NG0DRw7BYL
mqQweJG0uUSb1YWc+O0CJWqIFOvYRCW4hftM9Cn/8zvWqm1w4SKgXtw8B/pb8PtU
iQh58LiVG461UJDyWaLgPELpsraHw2tNM/7Byyg24APenqIyRgHO9zPNFBLDXJYw
pu+5dPOh5fzeJHwmWUXDOKdEqzjPq8Roo6/bRABGhQK+WVLjyGqS9mqqgl6b7RG1
QBidj+0lrmhdJwu+LYLOJHAeHrmRwzte9z4xyu4D7HDO7sBfAD6VLntUzPA6/xEt
SCJkyHkPgQKflztX9Skx06abp1oQGhlz5OVMmR5hlbGzVW89e9fBNlRG6AOwnTh0
9LbwO1HMikfLU4fDUfnpHnoyhZZCdV8WyvmkNM6acOWVX2FoFg3D0vtADNdfO3hD
Ud/V2T6rVfu8ohce00O08K2mKsbHh0bZAhrv6qMeXBKjDoJdKhaipwmMD5LHNkrA
RBMFa+JQR21k6oH0an/pbOm0/csRVBG8YQq1ekq/5S1woz+A78PshIPYyOhhIypw
LaBnFTbspbxrK9y+LOCbkBtOpOZ95rA0oZAasl5n7O2q6xqUknluHpzDnkqKy5hQ
yb4A8GoiQxy40IL0yY78icw42qbXR8e0+WYu8Xxknuuqm/ooM0XIJW6w2/8AnPNw
bAsMSQRb2E6Qcd2kn48LZH6KHEYNA/tXL1YVx1KU/yLxHlqR7Sj6GFLoX1uD8Nbn
V92Iji0D4IVs55kPwu8rX0YKcys4kBtWNq2F5WvGaMGmRnUc1uhgJsccRFwu8cK2
PolUkXoeg6Wt7IEZXnSXSmDSeM2QBorSkhlMkw9tYH7cgS722BSmqm0fDj9aca1B
obU8CJPXsbr2t5OjnIxOd+ulYGoFuiH7pO5U0EBBWQ645nw4nR6F2e/ajPqqzR0I
CgMy+FIbxnxFlY9PDx2INhSr5BH9dtTiUtTUzySrm6C+lD+hm8GWuqwGns1qGQSV
F6YrLrXAZryeExbl950Wbxc6wbJdPiNMDM7kVyji1UAYzjlRyNlRra55w16tNT9O
Wf5vpNxt+RPH9bkzbJyBpJju9Yd26by1TZW7D7bswK4Lc6VKr9Dhh2CG2nayMMGN
B7HlhzBuhOV+heWiZPMXPIMacE11vl5rcTO5WYsH5d6NyUPc+9bf55lfj1UOlX07
+OSx4kvBpDyERXuGCHqeHqsmmpTrOVtlHeq4UpGETgrNuAwqshcANE9dhTiXsGr3
pN7M7PAgM4BsS7nzPZ1YI1FvhFBwogAFGWNeBr28hc4b39dO7mRQQD6c1NUq+oKS
UPMSHS26TcDx5I8SN2FQVFv1aM6Q0BufpzMcUQVlZz6eHJEV98aRojnJzzIuB32N
gjtj7S7Ew7OiUFW2DopYOndhAvN39rTpJM0hEShsDLqKHveEMCHQ1WAX2BTaS4mj
2lSKcDPVkd4uh73JD2vhOb+ahpct40a92EIZQJdxyUaCposFSKT6BieK6rSUQ67m
4Z6Q8CP+ANo10J39YZ/S6vKkDTMQLlTPMWHZJmdP487jrmjed69QszKg9b3LU+4u
6HU6yMp/XgwspBsHS7kGvsVWSrBodmhzR9BJ+wcjTkVFgejdCpbeuT58znDLaR1W
tV/jjEpIBpop+SV5j3D4kpT0tzUOJwDbKBZzpsE+kjg39kO3A+AkN1UVTWR7mxSS
h+m7nwKKe8eRMxEF8xlzK+amU4nGLuQamm9P2ywVbe3QHV8XrMj74lwu7EUn7xKz
9i3y1i5TCjdzNYgRyOf1SMbifsyBINUlmyubDFshrCmj1jkrU9SFDpQdOVCifHMW
7EDSiz+Zpm2bAEbkv9HjuZR+nhDepCw2YhH1JGTxNuKn55tXfN1pev/VOBIKHcV4
NNji7Kkf/MpGzGWD/sfbRYCrAxuOz/r2NPqVp8E7ll5Jpn5DHBHFYE9MavTsBNuJ
s/4Xlezbb/Y0gir5qHGB0VJwJyNXV9C8NA9tgFYtp+ZoojyGPdl6gwoU+pPN1977
liN0WwJOJBH6mFvjd8Hf8YPXOpTYqnYpEz1FrYM6AqUfs6XX5Fcreqh+3DcEiYwS
UKA0XOlAuVbwi4Nn19foMvQ4K0ZBd61N9cBh443p4d4zPEyteQ9j1rycXr4ooykq
rNWC/L4Bw2ZhkP7O4g+rKecx6LnIyNN31xxPHCUBp2d5SgfPIqYjXfLdVYxaG48M
GO9g0zvrLwGo180Y+lDmnJo+PaAEbP1qUSaJzQn17SdQOW/Rkne6a4YGeere7xkR
FSjeQxa8n3NocB9uP0oqal8XnitUi9ogYktE8fysj6PXS5coRUa3Qvi1E8ZDEnvB
xnAv+Z051l4S60JiG97pMA7HkBOig9Hl2b779zjeGQkPBI4bLJLcd6Yz62jJfREu
hSEJj2hq/SQJ7NInCreptcBPlo4LvNCtUzhrc/9IKMfJEHwZXFme9Ig5uW9Dy89Y
8tzFBd8rtaYMTaeq6larSSoNDIhJc9pnEgPtjnb6FhKUkDZAlyL+nGh3QJm+bcFD
ILLNuaPJ3spKhisDAmw0bVJY84j9/9F3bAsnwCIjAOy8VhpVyO8BeTjY6BIJNngR
FM8kgUH6uMN0FJ+8ZSfeJYthY9xbF83YNICvc3ChDrLrzDMj/Y/4UROrGbijJ9Rc
i1Hbi1x8PVuYQ4Uk9stQu5gYz7GNYAhpYKXyROlFbpvkOz9Y4xjyuX2Yi9CpfAJB
PI/BZsUXDkBD3t5r9tuhouzmAcvCz1Z1mUbV9rpNU+ouXcVN6hIixaSJQrlz9z6f
CGiBasT/5TvLC2S8JL55rUhJHQBbTTljhErpsxJnXCkw5dZy56IYP6VHrr/VL0Oi
XyRqGI4H7LjpMZfbt2lTJEOi8UaLZOKdegTHlw6k66j85VLnzpvNW9cCsePeLb0M
ytRE1buCUV/H1fzyzjl26qWecib4zVkWMvCqjDk0Y6ACoba5h4nOh3WhknguCTDZ
uV+5ipt/9TPnEv5anHBhjjgDmbi18favmQMrjX4Epc2BciNpnhYz5RE2xvzZj3xU
UvgtNOwEjtOeva0UlSuyUDtJAF0U9G6eUxk31eufSSN6fDtEgKEdwgxoInjyAbhP
NdIwql20CMZaJgYlearI58V7Y/v6kEL3NgztUXp/YL9e+qA5G6Tvq9z+PMD8Zonr
rQ7XLDKMR2kCWcQEK3FKTsohqo0qLqOu2WtBpK6/kKqNCB1olwMq3QsZeDwCCz60
+J6+EEkfYNjZlQ0z55F1s4Qm3fUNmu1lj5kbDHlyMf47o1fncaoenlcBuFXJkbBH
HAgLMpQIdD3k8c1P+AfmT+OohCjrNFEY+KzYNWtVgumDVUyNm2EEDX0yIlFPfcJu
zstQHuSuyRYtCN/jdRJJhJUV/ruuU+h4ukhuSIQAcQp4GDoPugijmN7YKSc739bB
sfS3VeHtNTXbY+pthTnWhMmBnFova3/SiYbqFaJusCojVvHoGp0RqsBSJchEf6jK
6/y4Tls7oQ1AAuZnBA17c9ixpueDif132lKPZoWk31bqi5H95wc0swXMmlM5RhDr
AOKFd9pOiR5PsNugioukZFBS+hp91oUL79S/s6ZyBYF3wM8zKh87jDl0u0CgVYtn
TiFJgaLy/YVdtmDro2rL0VYNK2/92mLx6E1SiXzSdAVJ97yYy8P0kc5YWXf+w+pO
Cs1Yqp1QkKZy8gtOiOzEsngJFFVTzgia6k8yuq5eZAHif3alVqUqyto/a9T+IZRO
yJjKZJnjzgsHj27VHmPtyLAEbPnI25DtSymbqRIPIWlnZ2DW90a9mzqppxOjST3S
RDUP36IarIVLLKkW9jFr3G/HIj5lkCwznQ/MgM4GePHPa31buysA9ZoOWbHTiX/z
txLiu1SDEwIV6c4LMwo9D4QbORJ+94MePO4jOOCJYYpNS8tU6BbyjIkF2AOStDRO
vRXlVMWwCoFQ3RVLJJVeEbNDTlq/adFipbXLaL7ZOKmQUdJvp8R2rcl0cQOtXGEC
zf2DIF/gavek4+B5zQtJNSvH5398QU9PERxG6FxHF4nqDGHKy2CD6KaP3EbuJFnZ
akoTHDwYvb9isUxfYzfvGraacYRboRlIz/zlmSuiqlTvksRuqwTnTBrn1g4AUeWR
iKWqyMoThv6bPYD0QtQ2yLuySYPL/qLBAzjS2NNbFDSbXWMu/EpVea3JYBwNac+j
LMB4JomJF6NLSxBX29SdgYyjupd6j4YDBopdDPRm9r3abuqMwIwJbjAnX69/+0ky
cJo97zgwFzD4uPN3x5EelvRHkrgLFLEbgeGXd1Tw6bvUGfuyjynlhJKE7bSfGGOr
RCyJWzf6lz5SMlpb2U/jzxSNMmew/3eN03GDj0Ovc1zpvGXfRQLl+kFZp9ToMkil
r0gdmpMM7q4qKMovzV0lYEnPryqjlfCzihWnbXqkUbs+7djJhPhTtMfDwRZNrIBj
ggoVJcmBWCmAANzxcb6ECkdYWxCXewBxp+iT3KvemuxYNgaM4cag08gx1JDVxYcR
TyHTK1SORGwTJVWm8Z8M6ZDItZwncO8onxbAA9zqy4FLfiVEVisYMJDfYOLZwR7o
odD35TgYwMq34bEeZ84l8DEe9s4O7oaaTDSn/YUz3bpj9wJQfq+gUprg/2wMqK8N
dOnWy5x3Nn4yiulp8ii5rpe3eOrmLVTntGU47cctUahTZScFFvqZEJw6quj/yD38
Ww7nTCl4IhaETdC+4rXMiAZvT1dTRM5aitdIUCBLMxsEusir7oj1AnvooV1BH1QI
13ulh4pAFD0y8IetPXkQhAL/I1YT7yKU6/lsPhVQqwSjUQBwOj6oG3LdEgrhl4Sp
zN2xkU99E5ydat1AQYQVJCSskNRMv1YJbu+J5q2GZEnVTPuJiFl6sM8cLWbfRcTS
BaXNRkgWkgW7wqxgFqGhaGWeaQZPuQ01BUt94A+KzfubTvl43WJr0jh6cAJGaoQ9
rfWn1MCoY4IjbPe6berGgBnOu3mnuvtt/1+C8V+VL7O0y0+Fk7hQ6HYN+aRkyVz2
1pJ5qE/lM4d/cnW1/0fAAAFkEwy5O/d50BEeBmKrHi2vsl/hZlvldrXOIBCj7pzA
lt4A3yEn4NJmLWeeyFLeuK3RGa6xVq/vAopMktaHFOGjQ9zyDgah2GTJkxy0ETPk
JrGqK8LiguFofOdSZLIJtI568eXG3A3yAKsKBRkom8CBAgqXb5U/WTca16gDhm5J
cBT9jc64oXDHpgOlsXO5Zb+K4uISiM5+uUV/5W3bMjjaLiT9/DqqmiBIxLA0nz40
vSI/iGgqMIcrpIG9hwy0TfNn8XpSwaqM9fb7OyplomdLkYX99+QpvzA9xwpTpb0V
oLH6qqsJ8m3up4XSjNyOa8UROJXmuylyiwegMx/gqSvs4LjVbWlB5i0KOcO7GPbd
5+n00Eqq4bjUfBPxPbnSTYMLk2H6jA8uUiaDib8dVtTeaJ5VsXCAybYegtsk5gHK
JDVG2pxrlBLdykUkz4p+Sgzlkth9WZrbS9GefBk93muWCBn4GpMdOHAFj20Cq7bq
8hn6q7NBh3xWzFF4C8kUWa4FR/r6M5S2EqsBxlRsUJ9v+mZx8RgS1twXGetWMPgl
IYqGZfnnjeH88cNHhXx1QBedXFUePv5LImPXyN5feFSwzENFEturlbt5j7UqHgmf
XTXM+LR296tpI5WGlSlDd5fKF9bduqGRJd8vIKlcpwFlAcnNotrws/THKSKMcLU/
tm09dfTD90kZhnXGyoinnYiJA2IS3gbA5JCsN8ybXbTAABS/oHo7+9ixxgoULA1r
DEUwe2mDx2kh7H1SITe8kKq8KNRmpP081YDE1M+B96tb2HAWWC/WVIuxMRQ7aLez
LevDRFitq/vFWOpg++UAVPbC0Cqk9SUiCoo71zoiLZwYtgiF7qX8fwVoBxHCmoAw
WiqFCvl8DDD59n80pwYFP1Okauuf5z4dGyWJgu7S+CgF8GqqrQoQ0aslEKmyYUEf
2CB47PuUl0rhw12uTGy4YGtrorcJdbJ6gUgQcpj1MxWKiyag8XtFYODj8ulznNnP
0uqbI1EpN3HuSAL9vB3VsN75CFO1sbnMv9rdBo7r7+VOx3cGLjaJDuG1hR6+8o/O
X0MzzEj+VvXRO7nsegSEzkE3+WVlTYLKJrx4JCRwqVNaGcajDar4DvoQrgFrgFhL
aFEsjTEe6aFBwkFHy3EQUPQEWKFrOs0QyaEO1ZTNTANB+NY7DKsn33Yk4KmzttDx
fuNfgvbsaW0w679GN1hjkQ7i4IPUEyIvYzh6uaneks4imGX4gy7NGuUyCH9bxM2A
UEiW34tWFIMFzIr4/VYsQ+U7bqnKV6WaPzWusvWPAPNw9oR+Zmx+5HiPSD9f1N3N
3UVU9xCOEEI1ZLU3mgFWG5VaF9habHQOVIvgCZOjDgrS2JtdtUZl9zW60sE1B7DA
QgSMcdLDV6SumX2qQUVdi3akWAwqWUM4Xg0wtMDo4oO4C2dPFEu4+AW5ticxogyb
0fjka4BLhKjnRW9bnzX1H5FrYHbma00JAyQJ+ofX8YPEqxfSlAExfX0Spn0pJVHu
ZCF6CQBrmHXJJK7aFhW9XhaTw5Nelh3oX2JWQn8P6kfwxJo/No+eGjKuWNiD4ZHk
Sr6bwbM1+/eZK2kYT2IBfZgfl4AY4665wfSa3XHYbbudfeeU3/JazrjyQuTbBLyR
LJkb2yC6kym9/sWh/0h7hcjv5VMZ2pPhEMGjKDHjjU5ttagu4pB8nVnbvlTANrH/
NuACU0b4HF69uvWMNAfNn1at/zxPTKmQRyN1wWF5Xib9eCasD3BHG4hRrQar1hwY
J0Uw0xiN/pryze1msoXbxAiwxuyCElBtiSpR0kviO146+VYT/JS3LmgZK/aK9xpm
9bsRlJvQXqtU1Xav79je75Ul5m41PayO5wkEWXVzreyy83ROH95Tpo+hFMSWOSAq
JCQLZCrdkthL2W/cQ3UVKlGaq65/+fLnOhl33J2e6PrEMGZEEaF3d73cwCA3fAED
IvLD8/BU0PXKu19XS4+grzL65/O2qD5FI06Y1HdNlBk4i8tw3MY1SrDmjQeDnSJ5
ykjWm640imbWmaIYfp0T79hWX7tlO4rywKBFCmgXuskwG8LMbRLPy93d5XxldORa
Jd3fLm+YIvtIx9fDLYw/wh+c47NOtefv7Agu/u2p76t//CP8PU9xYQyvH5otuzL2
7Gq7Gy5WGxm8jFeKSqtpwpI2zIAR9EetY62AmPOiZ45eUBxRkoV0yUZPNh20LJt/
F2xgcNtfJmyjxOacVaCw1+cdlwMfXos9XkFbFOve+3zkKLKx7YL84lB3mRw2xH8z
twkhyg+r88zuGAnmlSZSESlbgm3FVyzlxPzlmgB1WM8ao/sVpy/usEFVke3pwnU9
uxyQzIfEKwcdL8dQ8wovCetaGQjejt9wUTc2cuYms5LjVQTYNshD28GZMkPmOQLz
GKNkVwRUBLI0Vc9B3vV87MmDwpJaMxsV8ZGIYh8wUPyIUTcpP2eLIE1QUlE4o97y
/6CrAgvoXmsw8bOWi7vsSFjai9RDUGtaUuqsK9CSD0ph8JoU6o01GhYZVMxM97HE
L78hlevdGHlPEskf7oTyEh0EKEFOOkJNfromyAUaKdrO4TCCMPDo7x8EJB5uev2L
xQjwBEiTc13KQ2gj1KgWHER9ZMJJtmQ3edYpwsnNXf7JiOP0PtD/SzqRVTY8VuL0
ddb7JB6poDy3iHhZwvKQQPjQUCCVkrtO3+Y1q2JnuJfNAIEHcAOeFF4bqlgC+zmQ
T4UBVKSDoIXNCp/Ao6CuM7eiKQ+CAZ2oC6MJkE+W1tMEP0Z8bu8wpzvH2L0fs0JG
gCJtpWJMknuYwKD77ad4HJ+NfwWIxqMHSNTdpTROKxfbGIlKvoxcFUWNmvBs4OJ6
QTFA7z5ztTN2O1qrcelGxTQFU3vaA6YCRX5CYFvwv9BVn1pQCy0/9XrM7RMTGS9o
jpqOmIaZI9oTz5MwV1YhmjPg4Frb1ycx+aGcDDcnPuoR9iyrRsvUfcVOeZwedJAu
x33HO4i7Jr7DG9F7Cc52XWYtM9Xk9URj+GR1czD05ri9ZU3VdL/k5clvDffiFtAk
IznGJMkz26jei7MR+GYnTTRHfcGfYWVIRh1C5trjf/UqWOzl/L0HWHQtX4YeD/9O
IJUKBco5y8qxwa78mNsFf+VAR+A1YC3UNyXkAV4Kwc+JwgYSlRM66TYwZaT9d/Hx
YbNBv2m66NZkdcQXyKHwggBZkvB+SlOEBjGGQyghnN6X/dVk6BRUwx4ebOv7V2jv
m1ajiCYhZmtzzXU510vVvhhit7LhCe/6VWT9UzWrD/Ywzwpl8csoYl8fLJ041hjZ
aLMymMcvjTGmd6CKUd6kVF8Za1TXuYdp3MwzHFfwS3E4kZkfaZtcng1v1PtSDVES
eVGK5OUB7GQKZ8kpIaTWVPslihmbOMMRGqzcmZfrVOy4Cz3S8NwLK5zL+qCEPceB
Ix9ZEmnKcIqUxHygQ33GvydONmYqDnkxerNuPoSyG0dRrhUAdBCC9mb/TT2QF1RQ
AYWyPFvFtECGwvUCOxPs1UxX6j8BGIUrhk1AikPJ2ONSr8vreYAudXU9qWk0sbks
1qqwHRE39a6pbQPgKvYMyFcgx/B2KZ//8GqMHlNYGDD+KuBOFlDrw7RHzZzq0srl
Br4okscG7J02Fg4637DbQxaO6GQf47IDRSEnNE5oEv3rFrrNoib//IJrp3LyWUFS
MkT3RVqK8Qa+lMHlFNncCs0cBZnxBD8NFCsYGP1GLg9bLxYFJAX+EWRfCBUZ3LSm
tEQR8KDJVeGrAOGq+ySNW8eiTNATHLt3ayawb4ndOfl2Obfn91wEbYsX2vTLSLsD
dzNbWjYbZEG7bQBbdvOx/qkZ1aLg9H6nWxz7U7uaRlaX68tiSNu1rEiBF0FhJpQ9
sz9w5tGOl88T0Uf9o/S0YfDl6G4bmK7X780bOI9Z30ZPev4wVa4eDs9cAVHPw3uk
ZkHnHp8d+TMsixQUxWMkZbiDP07n6UhGMOH7TPb/WkIARS3j65weZQlEVhIycMVc
4E80zlKUeKlDHBeaoSIQLHzNSqrtS9Ptckm3HwgDlgjk98vB2gWYiOSJu94HTdnF
Qb7MmAtQTPd8UwHExUjy0d1FgIzFAFnRaKwbKUBDRwWhQSE5xXmlIvl4oFLOHlYd
7Qb6tvxOoPvZZT8MpaxrR51ckqv+Ahz8hG94M1PRPndE0rALKyT73f65CJu3xt1N
meklgUKjwPv1EsC5A6ULZSkxcPAJRunKcAZN6gjL/Yj1vSsYTPtZRCHOOkk3FJTx
WGP4tgbhDifS3dH25ARifrbtjBjXez9lBO+gZY6foB+DReltS4nkWtc3532anVwr
zfL2E+Ozll43mve+WfBu4NMhHrUgcp9ATvE8CL7IgWXnpjCGbJAy2I9ZTtWhJnk4
C0APVLn7xR9ruaYHamU0bkVpFowHLEX7HO4TSkuHTunUTVC90iubvUVsX3GQrY93
3fPZKjMTLOjxPAOLinQUgC8q3Fb07Dkx3eMWfwWcEGf1HM2bJwJJcs0daTldMuGl
ooYJEVjJBNB+WbTXSDTi8qu5TMFnGcBYrYpIHqvZ4u6n+BNX8Tu5m1JP4BV0oJcI
eqZnUhoroycjL/oA7jhpUsR8QnGvj3zrAjVpX4kpvl6GjRsFPLPuRGU/CQDbIbWy
NWqQOTWxaXkHdBRXc1MzxA6SK2AkPdRYP9aP2gJlwXWXH8DoejnnCHKLAweWsXmy
b78NEhN2C0JwrfNMekxCqQWQq8V4xEIwtf1wJlWswCI/ftY2LblT/PUsYsfIx3cm
YqQxXuSCzeYs1OyyivAKtyf8H85u+h3D6tTxdNydKiWbAwj24yP2Z+HwCjH1zQas
yBtS2arUSbtFSntARzMyWVaruieTJGEC4VYBA88vDoBdEU7kOKBl8M/Vqo4rJur1
1Vl8QMtQo5GAgPF+31j24bv/9+pP9UPoXaJB0YfdVgEmHnvcM905TT0g1sgQhrko
QmwqLzz2om6k+irq/iUXdnb3PJGymvjhCK1I+QCJh1CVNCIouyYvhZZrWWnLXwb/
IJJVLnfJ4uuAb7fKaKXNHXChrGBlJm/K0RpTCibXCigd1W8tj/IFngOxFQgGbHWW
cEqC2umden557Ej2YOqFFBeZVe0S1N+WU10eo9UpiFOVHOFLuGNxFN9zZn2jwfjO
RmqpPqThg96bJvoAniHuQr5jKmDkd0UMHsNnCwZHfSwdNTSOeB4Ar9kJYG1vcovq
O38gvke8DV4zPgIYl2/zysbQHygXELrkozWHqnqfGXqRoYGNmfdZDt0MWQKkhMGS
oB9vOOi7w3x3ocqkvJJBjSOPW1KWkrEJoXr2Mos6F/9JY1Q1grvAyYvxsJMrUC5D
9ZcXq8rAz9S2LpCizTzVaRqtHq5yzQ4CP3RDR/W2cFQr7yL6Ihs57ZuijwW/CDCg
GE1a865dnLTkG7XFbiiL6oTUdJAENZ4Hxn9kcxJ1Em+1wn2rgzrVGGiL5AMbaTpX
zghbpuNyEWzNgh8/3BpS3ZPaqoSVXJHxx5f0451TJvln6u8v788d/YmdQGMkfhGp
fvWftlt35UzwMuTyHGSH2VmstZ+ulDrBwOnQpnxRJAd4IarpOLwscXmqDhjrL+Zz
QMe2lwGRf9WAqEx5She99gCJjzeIhlbz6nKaFml6YRBYP0osgxmRcZE2ajqLXFKi
RMEvt6AjQhbnY592DLkU1mhoIWbZp2RO1lqDZfoLYOXgaj0wSx81AxssOiVYdSx1
FnCd5xTdTPsc7ioLf9YZk1LVWP8Bub0tzGgdnzuevfX0Wf5fZr3uiewjg7fiObJd
3BRU2hcP30J7ZJcS3YNU0E5CGRn1gFlYPhhCwF3leMLlBtxaEr8m9nusPb2bGJ3f
bLuMtjeu1n5bQ39h3BR8XifidmVSnpNF6H/lHi9yveWAtd5Fz+1347bAOaqjIZy0
to4ENkPuhDD+DJubIovvP1bnxN/DGf6qaAj2HBEqSWbk23iYzPdA0PEBtVjb0Fb6
pnNxPEsxUZOAHCYeuHJBNyKGRYHUMgW6/EkWweSuECNfqQvs0B2HkVoeh4Jo78t6
Ajxj4hX4K2gmyXVezy9jN0Aoxz/HnT0qT+IKZE1NJQmGjBKsS2kgpPIlFzjKaMv0
uZ8UE8mo5wdZ65bE3gdTouZpJy6tFWB/7Qefx4tLQpjNSYzywq2KmPwAMvobp457
kP4tdDkXZ9N6RA9LsTK+w92wJrveY2sZWAiA6yccL8M+Fa5InX8r14a6jkNMOxTr
quFQnQHr+EocA5yE9CGvKi0BMd+lp6pHOhBawijlz7JTIJp+p2Agnkde5EBsz925
rJNWerez6S3Ox371Hx8HVRA83TSa9GXm4dzhWNi3a6LMyWgOHtNCvpUqnN+I3lIR
5c3/HnZU7DcCAl2Pq/ht8eERPiuxoa0KVwjI12dYzVzfDKqWeJ+N41kZ/DgERcb/
j5K2UWFcWI61V9Q1JNhRiVlXcq75LwE4X5ztxIfzwcHhUr9hhPRiazSlcYX3rzlu
c2RN28qwEkPwMHDcghO9nrwrxrSGiAwXCmbTaijBnUq6607ai60rc5h714W70thQ
NTXwDbfW0M6AQYLJid3iZ49zJHkQhHzhI+EVOdka+jm9wG5dLTbqdCnmCFpOUZNg
veXcnrRAFTDRrGbqaBl63BsX4BXO536KnQqhOP4kV0EiGjam0SAvvjVuoIxbIG74
NuZwhrgOH+ymeNbTjR4Gf535dBw6zrtwVlrOo0f9dWxLeDwOYr4uuA9ZbNSY03Pu
wuCmaZAYRMnEI9QhdGYfj44PljKYOsQTgk2YQuRjGhTeZIc0jEgwcrsqO5UWpj7E
MIl98Z69lS5uKT/0NdXFUWDMtHG8spc9ODfDGC65aTgmax4DtDRIESPHDICRuDkK
2nLHzlWB8x83LemWV0dw/Uo4UTyrODp/PUNCeVU6Fotq3VqAEEVWrPrWHF3FrIVQ
VfsMIrJSnj6L8cOysJfz+GqR1QUDrXMvBGKMpMB1NrawOQQeyih1WCp4pGmmxHrf
LCxIhFe87+J/0PGyHNesVREK5ZIEWv56dw3GVoY8+BWA/VOGHYYhUWfZwRh2bP7T
SdX4pCrr/QLXrlJo0IZ4+Mfgjmt2H7BIQvNIaIhy0S5m/ew7Dhvfmi1WNAV/X5Wo
T4cCfMlo97WDV1gPnKXRm/3Qy1d804jW5YVCJ2vqJGzloCksu8G0KTjpZzshA/Xo
aqQ/CRxDcaLvY3ocwIgrcU8ntNoChPOHtmq6Eb4IWgTkc3udtK1R2JxVQHyH3zNF
Q22KQuLwlw+E58nNP+pm81pEUbECcPRML2qExYw269DjC4TzxS8m8Oy5qOV3M12g
g/Um8yqZTbxxl6C2CBrkLtevZhGxH7ZuDLrRb3OUfjXaqkmFePkFdcKaO1rR0pWH
3EqU8zDnKH5Rj92nEhEMPdflEBXgNOUOHnjdFq1PilHBn7fTLNjDs2kCOkx/wXcF
Tdz00MjbWFzNs3wfUSVCvKVo+tEQ08VG8RFcFuUR7jzZJnCsWIQFDCDE6PuESGzi
xUzOg2wq4p6oHat0Hi37kTCH6RrBcQgzfqk5Oz99C+NITZqhAMSybH5smtaC9IE0
e3n8wZTTV5h4yq10guGcddaO0OUakZrwRpbIP+djF8nTWCrZ1QDJDZAWJP2dy+al
4up8OAoexc8gXgtkma/W2hN+vYQY3ZMtDVfV9mb0ab7wsetzC5vV7vp20raahdZb
BnuN5+0Xtv8bxRYOPUZQVHa+2LOWzqOVsbmtgrIB0Pc9YZpQPwSQPMuItNoPTTNN
9J5jS4QdjIf0j8adPHqr4isnwTcgQRiDHOFinHbRQsIN8ylXbP8LwmmiF40rpONF
NzxxCck1C8aRNvDsSGXdAgo/mhLOFZP/tjWRgJEb3mGjIGnX5hRAmIlpP6NdQkYw
42Fu7ofYoEnizgkHbVKVdyk5KtdiAlQg+6tbxzrCIatjwuRG4S3zI/QiFxPlU2gl
JWBOUCshJgQM3X2fUS+xSZBbD6rhBkyrPCf+3YJNiLmK28haOp25cu0eKqO8T4lA
+XhAZJtNsZLSfz/hnvboeufGQXmJ7F+h3KZ9ae5EQ9tIibFVnaaK4DxCl18cuUvq
fjq6rgcMQeEPhX+twyHjTwgF7Hm3SMx24FVYdXWXvd0ZiUqTm3/WphYG3uuvHlDb
Mul/adCXh5vKJFneSG+LkSahQ3P5/HtPh2AyFhNIpyJ+x24J7HjbNVBeodgzUcID
DmIfdlolzm23+cuBxpEqx2PCB0noHjRTCWGja/38Acel8qhI6lhEdjNo3janPs86
V6S4ZMJL85l4KpC827tj3/95WZKD1t3S+cT5cvN9KQh94g4vTpA6HT/1P8FxaXZM
hXHtUC/Wdq6upkCA49rw27JrmWqxsOvcGYb6kksDiFcQkXQlql5phyqsVgE6oDmr
rlB4FRPEBEJpjvxxX1hvGEAKOtUvmpbWjM6DkBMR/+AyTomCjVPO3Ez6gaU2LL9J
x7BhPG7V20Zr4SXBIcBZ/sNAeQPzZVZjHcgGJHBsJ3jRH1gmZBEUR6/LRi+fHSS+
f2tn/CONF4MLbg9Pv63lkvtcu5BR0ANtO4nFfrNCsyWtEHQwGAOEwQmTF+ynOJIT
FPyk9IbKlcf7ZNURIjDQ3l34A5wumeoHMDrWRXg6iJxFbEyTtmiFauj41ygxO3mn
zYXIyzn0w7rL7mUsKb4NFan7+L6q6arxj99yqIWq6EBc4+hZwuXlcxUan6A1m9eF
40PUOjkYs9a+I6w0WbzElzPVQLd7duxjwAgAz3xO4NR4UOUuV07dnN32zAGdl3jB
X0B1F8bjnwLN0TW17gsr3dsSrHoXAE9C8TOEIxINSCj2nbhKYofivnwoRWfnTpd2
LG9U/b7hyLSobdH8LVlgdoqtE22Fxo1Ozzq4bSQGsCuT3EZtylacv+EYp3dAsdKn
7qg1HfZ8K1fzxrp9/7J8HkMFBvNLPQg3T2MSmvzjeNtQ37w7jLedM3cbDTEH1Pdh
kmzunoVIHHAb2N/pxtYvlypZMwtjJtRghx+GBK4n8QcuQ5WiBP2su6nzmQPfNobx
ee9qDDY3ydy4qym9KfMhc+u9uOTazEyYU/NadVtxEzd9LgsleqrVvBq+AK0vLQGz
qdh+gByM8BBucdl8eSLgCnNKsam8ZFdfCgaDUDAyB1XY3gKs/bm29xuPFlXhQRwT
nYwYd3Z9t1okUtrOIS46Svjtibw/9c7m/WfYPtioHROhRKAGyk9u57e1zmBnUc/M
wyj1sa9iFqrbuLXFMqKQOvl6JJUs4FknqoPbVf6qff4=
`protect end_protected