`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
ddtXksX2+yylW5zu6QL2Lhnb2d1sD00763mmSITNX595NcHTEkwn0zB1Dry37fOW
FufOhVzEJp80NC5qZ/+F0Vk7Ik02dIR0elf3clrjeJRK85K4e3Hoo4xn7YbFUIms
l/8VZSb14+JVGURjfswrIyCUotIzlzVYZ6gzoZwDXIi5gQIBf/gI+KxNXPaKV+PQ
Ufys/12rjO6aI/pPlqSm0hCvftmBcnezN2hk1UeXgOIuKZnogjOsf0iJVX2aOOWE
6pD/psybjbnsNB6kH5uFTA5frkzIzkzl5d9+YDm9OyC+k84E83I/7/j+rk4L2dah
QJOvksSIzN867/4Qt8qYTQ==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="MvBXkzurAa5VTw+1JJ70nePUfoQXBvZOku/SMmg4TwQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
oRtzZL4VJ4iwysPsC8SXYCzXS8Fw2gtZTOskLcDV+1B9Nzn1zTyNtlo6lNICRmmK
ZRVu2BmCc2G+fmzynYlNTnSa7C0Cuel6FYpxCBlOuk3OF2tzAmLAuDyOH3Z1Yjzk
a0aHuoCdIRKv7BrZCdALt03JeUmXKPdOmIlkVGFl8yw=
`protect rights_digest_method = "sha256"
`protect end_toolblock="Jn9CQpRhJt4rnzZPRk+dOpzAubz7omckX1MrFd4p81o="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 3872 )
`protect data_block
gD6l00tciPUa6pDNTk/+t0OO0nC/UTtBwLB41d4inuAUA3i/ALrNyoJVcBnAmEQW
ptbcNp5fxEUJjnOxnedyZEuEBxWRieZFQnkRdF269oPZbWQ4F1RHe3ZVGRa3O+DL
rJjjIdeV8UbZE7a/8K0zyhgSHc+hCUezH1ARo4yaWeDP3TYERMtqE08g7d5nWt/p
id88/GFP7CoKtF4jAozkfaC9RGzKQGXn8z/l27zc/bQ3Hfp6z6D0M8yPvp0BE84m
5B5Sh5+s+EXmGMBcY5TH+5wefZrL7ExQCm07dJf0RS1TA4/k8wh1Km3KkzAIHslI
u0whKwQdXAiV55wjVF24tL7y6qUbmAc9JiCm71MFLR6dLONvRfUCAF7EzfgKla6F
tYmy9dl5BIvnC9+XJEl2iBaykwPbLa+ONlS3JGzESDYndXEpAw+xz0Uqv8gckBG2
pfoR4EgCT8JF66ZfO+3a+Ym9lFMGippBEAGHWc2CXHsfUXXc1P9fC7DYW4n5zN8y
feCWnK/XI3F1y8BVC1RHqEboLqY+/CxMraO6702nrdyILUUxox0tDgBgmoPLfICo
9/L/UebCKf57c/QDR5mx6iookQYmmO7hmEXJFnJ6yGsB0OJLz8lPunj2CUbx8Q/Z
zIspkhf23Qb2Mml3SBXa6CW0+gNjOVV6rPzllzI1eGkcMXv/tG3+amEc6PVKxGPW
bX8WYiHyf2kCht8QSauc0mftksr2FzK4DxHiScUJF7IYjUWVTtexkqnKsF8wvBGj
kjYzDAbgb9rRwD0yUfkITt6XigL5W0W3VPrDarUgSj+M+3jZuPReUKs1DM99TQnI
ZNnjE03EZB6NfliqqBXt4qMm6Q+ja1YP1EPyi4ZX4kT6OuGriVg2gsph39mpfKca
Jxsx4ogfE8CLp+il5ypwwVbVr09rELNIxEHm3D0TVCc+rRNgd94+gd2fCRykb5GC
jEgbefEQtCRTIW4MLLVCfVgzFSC5qUNpRVawcfNNOqSS2QptuwrgnddfOeu4eIM1
m+BhqLL+QjFYGT4HEVt6kQxBhAUzOR1nNz1lqOS46xbB4xsMuE/CKOkB0hTa8YtE
ePeZR8MwwOCNlgaXBSMtYJx26VZkox7DuRyR8hAu4CtmaQjVUWaQpJUYtdywmidK
Q912k04BNFXM6ucXk4owf9u/kmDGErcHNaxaLmfQqfNhHft9+PsVxCjBT0ycBSfv
SOERxG2RHbYMEwAg9gTgchfPx5zRU2Yyf28m7cOx3l1NBs0SNYfOPrLo2KiPZ/JZ
+70kJ6imPVkJcByFZAxuxOzDfWVHNFx0zCbcy2CI5Ub/6riXS3JlzIBJ6Doq4wYD
yZPE9qMKfeYIfVfk05srzO1InfpKFMP+26cVUgUKxcy2I/EC4te+vpP9p/8M/6aO
hd+RyvSHP4cVQtKj7q1aCROBQpWg7VwcjNzvgGHacVvq7OiV47ULvIplgyO18pQB
reGeCUdhv3zzBRR6MACq4NBzZ+NwcyAURPytbflvXlOZPNxQPmYT2WoW1rmPM10O
7MGx997YnaWWdTxVHxZkEdtcFOdMTjPYR28nIKSkZr6FNkFt533vvYB62gPmHqFo
4cfzvy748IdFVoM6kyJg1U9KW3PWjuhtuzHAYNTuKfhiqnuXfTxdzgnvWHUYQkch
RCKT7UQUP5spWrAgCQl7FXN3QEDxS0LvgiDOvXYBRCUyV6aiAsp8PgcGJ4vPyVAU
ZPh4EgotO5bakf5AXVkRTrkkgJ+m1/qIcUVCrIra6pRshq6rDmqH9K2f6w/Qbzbo
pKll7FAy7mL8vPO1OwAjx5/oBLHgT7R0hMImkJ1khjCkq+bg2IZF9ealY0xHXBxV
XH7437DMmSU8ncT5qrjvJtRdPdj5FVy1SXSAYosJgU8Ww7FWgOq/ZX6eHZcP75EE
QSQw8ImGGdIK9ECRXSliQfDI4j2rWS35HzOSuZGEkg6ZN2izC2pAuxbLIqLrw/3l
9dGUtA6PJRgErLSW4w8rGoZk+m6WQwk/jkNX/2v1KP5q3sijI+FIT8S1rGgyZPWT
d6qZ2M3yejAr90MKcUxvrLczj1POZOKSSRsFV5pJf4t1hQhQNbVTYidqvSfwUpiv
wJETBbI0dB+uB3Wu6rQtYnOcj9QS5hhYysRPJtmi224sF+14bg4MFkRKcI2tUE6j
dtS1HL+CtzNRNJ7H0Em7M+4kHkfDamQNanmryEGlkToEPLg1oDi4hLScrzaJwSGG
N0pHEozLEYdx2mWmXIMXkLjCZ20YcYavTxZHnHaHeKUo7n1edInplR9WEcRvMO4K
D8HVbNY65Di0zi2LRyyJOsKYwijibMkCHtc3iCXlGjTAlsH5hI6mSLkYlxKyvml3
AX6Jm6mvT16jzQJ5gJoaokHXINv+pWfGQmcBbKZrhALf0rtYv+cWPMr816g67f5P
mq+efM0U3KDlK68oXNPsg79+NppQ38GvsfJYeYzvuAl+J41rV3B7JZxMWQekRW4W
krZe2axCYXUOahd0e/g7WJCDwPVlJrYqJvZId/kwHS+Gqtd6A4laK+BeRNy8ds6q
VrTTSXfy1sMKM6bKefYcejPtY9RiV93cDuZ6vSi6OgvP8Iq7fGGUV704R/KFTaAZ
PX92z3C3fDH5M60ZT7fng1U8BSBRVm7Vw5j+zyQguwFxagQ6/RTqmNiIlrMQLxjg
GY7a3XvbX3CdeXdkL+0DeE25cXmsyjQd51A0R/BgeApwbbqSxxJpdC4ADli1aWou
ZZ+AYQedgPMlebcsEjpGL3UeQPwgOciGUjkILYQYEamtJ0v6kM25BvB6E24nuN4C
7Xjk7igNk9T0FlRl07DeaHgGWXqLipauCM0n64masoSFmfNTYHhNAc/V7mRnkrNB
2+iRlUFYsUES7e3DVwW0VxXGZGDPc0+pnCZyu4RSPGmFPjSPEdwEUxCFp2HFr6+e
QaxQXd7U3PvEDZ0e3iLeqb1RYat4ZsmPPuBxl/cPotSIhILyim8cv3JRUpNgVGvn
4d+UTy4s+o+jMXxK6zXvjMed4IRQu78CMUGzYReT3HTQnNxYi4k0erQqinkH3z2s
wjqa+KzkrNDO0WcVVyIcTWchjEV4UU+/1oR4Es0MyOkn1iF3QifxbiXTmPJp8GJE
f+UGPToCL0plQ8jICDrqqeLhn0CQDyTVlZsoHM8QI/s31T84IFe3m2u42AGaZUEW
/qpuV6C3xuLaoZmodU3/ECPhBYZVUDKI22fCR6UQT3nGC5pThhP0dXZulhJCuVpA
KC/JlOAQcx9CgrcH5kDYGpOufGs4puX9BssSxqpAI1qFlnqiXW8vgr1SE6TF8ucU
yBLKwu7LcfiqxHbYMPHqA2/xJ5u8TVLp67NPl+k+X+IrziYZdGp0N/+GJ4nx62Ch
fRSY3xAFjYGhWFad+kWOaVSEBefHK6sVU2hBCAHyoHAJbInez4yiD8U7w6AqSS4C
tRl99XI2i/TybnUfh/XbFPxPzYWYOieK6DbuJHzeerZ/5CayeauJkc+vG3pROPA5
ciT8573KBbnC3tTOWM5I9+qQVUYjJZbmwB877HoUvB3eYtw/s+nJxTJmh7rJHpdU
FzEVMrSxS0vvJyu62ihQyzQ4nJsTzLitAzAr9n7y1O5auhtRZBMSYfJ7A0pPh/m+
gRGrsV7C4j2eTOiQO34jvGCr84MgpxMsoH3Ghpa0bZ4NAI7YI7qrI4TGJfDRF8Et
OVX0+GsNRoPsmHwNbVmXLJd2H6j2awsLjTeyPpbBp8ZDHVFU2MsiRGXl6toBmX2Q
uyBHecI03OzyGuncbjtO/8gXeHFFG9U313RWE/hfDTlbTgLa7EJI/WPdyYJgv5Kq
kI4jhcKH0ShByeWXKLsFVk95A/FBJN8b1rMcwrJLNJUTH07IhB6CoEqW/h/9cC2x
aN0vqcFrF2oOtDXc3377Ol+3yYI4Ny1Gayx1YRdTbWX43TULUpTgelYHpqKkX0LE
Ao/x6hoiOB5UsCaxpn+K3KOL6EvvORK306ICnOijFvR0ST08Ve9cA5OEqVDelRzV
fTb3WPq5mTwJS42dX9CNTgwbiLKOQb0+f6KkD4Xd0/gLmrCUkIx+QKaFkgQ9Kidh
Bu1VQXKwFoupZzJEsa0ORYLL20o1Sjp/Igypou/iySu/hKPsJgG/mK6Q7ryTFrRQ
8aoH/4rBMuBlof6bAaJocDWBe9QC74CziLboU5e/Jqf4O2W/jFHenVwwX9ujLGkb
OywuAUwcbcn24SZh9tRlRSAhw4qoHKJUTK8Z8DF+75VP7szyE0RcNxsyS4OL2y/n
BoP1ItLCRJf0zNsdDuWRDTlPmo1wEnP8K+EcRkUUvs8Yx9XpVAx9rKqhGfyCy9DU
blv6FRH2qRbe+47zNkAaf7WKjSTPZFGEdjY8vNOs3vRhFty2F68JeY+GagCYRZ1B
/aJRfalD/90zWc9ZtZUmL9Jf/Ef9ngm73u2p0Zit0Z6WIrp+vt2cqlpPPjQG50CR
eYwxj4OOAsQd04Z9td2I6KXRkpJWHKvoXqzVkzxHFhP2PVdw5JkK9K4iEztJXbb+
YLqPa0XFHlK3B/j0hlGwsHHeKC4eIHnQ8Gif/IGQDWDmAzjkngjd4GnZ36E7LCME
SEzxiz4bqLEf3oz9gsmwdp0gClNTZMDM0Yal3loSP3gIgUO2xZBjdAG5Dww9o6LA
jhiTngeOBzYBzFnWYCliNp/W3r8spTDtvxiN4XP8O3NFvCXQK2s/fUL5aMitZFpi
7lqXS4ueARND5tJuotv/F2K7sORDFmeWOrAgLdOHkQCAuSj45vAaqpWdAkWxFw2l
uKQGBLvKe2WGkQ5GkbyR7e8w7lAF+STsWY5HbyuBEUOGjP6AuEHA5vqi2dNDIeyl
ys5eF7rCqELep7OZUjHO5hfGvTYFqqLBPMHpOflFacHip4ksZ7pUQn0WxrTUOtTn
SvqokBVlKriAHbXzMbO7czUcx/tTSTmoFfwNWaGRVB2mB+0EVmflGJUJMvqYhXQ2
aQEwlPgG4FsD1fqqUIiTJ8Xq9DIEV5Q5CFum94+1PNaqL+l5wx6n1QD3KWRm6QkD
50bKqV3gVzwsVeuZJ4M5H5SEZ2Bi0XrSlNIzYK4CdeHxA8fEit0VX0ziq4O0SKN8
acQHqbgLaJqWEUv9jDu5pXDbL1Q8L6x6K1jTRe9GRq4=
`protect end_protected