`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
ddtXksX2+yylW5zu6QL2Lhnb2d1sD00763mmSITNX595NcHTEkwn0zB1Dry37fOW
FufOhVzEJp80NC5qZ/+F0Vk7Ik02dIR0elf3clrjeJRK85K4e3Hoo4xn7YbFUIms
l/8VZSb14+JVGURjfswrIyCUotIzlzVYZ6gzoZwDXIi5gQIBf/gI+KxNXPaKV+PQ
Ufys/12rjO6aI/pPlqSm0hCvftmBcnezN2hk1UeXgOIuKZnogjOsf0iJVX2aOOWE
6pD/psybjbnsNB6kH5uFTA5frkzIzkzl5d9+YDm9OyC+k84E83I/7/j+rk4L2dah
QJOvksSIzN867/4Qt8qYTQ==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="MvBXkzurAa5VTw+1JJ70nePUfoQXBvZOku/SMmg4TwQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
oRtzZL4VJ4iwysPsC8SXYCzXS8Fw2gtZTOskLcDV+1B9Nzn1zTyNtlo6lNICRmmK
ZRVu2BmCc2G+fmzynYlNTnSa7C0Cuel6FYpxCBlOuk3OF2tzAmLAuDyOH3Z1Yjzk
a0aHuoCdIRKv7BrZCdALt03JeUmXKPdOmIlkVGFl8yw=
`protect rights_digest_method = "sha256"
`protect end_toolblock="Jn9CQpRhJt4rnzZPRk+dOpzAubz7omckX1MrFd4p81o="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 18336 )
`protect data_block
gD6l00tciPUa6pDNTk/+t0OO0nC/UTtBwLB41d4inuAUA3i/ALrNyoJVcBnAmEQW
ptbcNp5fxEUJjnOxnedyZEuEBxWRieZFQnkRdF269oPCkk0yDV9pvM7etfJwkFBW
KkzQarwZWGsz6BPDGoo3ld/vFyaO/9m5K3GGPqsR8X6UT2DFpd+UReyuSb99C746
g1PYBOx6ShX50ZppEm9EYLz3cjN/auXxFgZnIEvAEXuA1/KGky7gmxhw7XF8rhIc
4861PuNz8EX8RxsfMCAY0GpwWgP93659NX/+zOY6EQrnS+uDmMOFVTkcFxcXiOVp
wkY8e+95EcmTgoDJwKuSzKjP3hHUdpO8ICNsPYVa9UKi1bAndLII9j2ldVqPZYSx
ilBtPcyCydLhLccf3anKKZ9fajrRf6QgDyCL2/Ph/8aBKFMBWG0dmUNBPdkeBidY
FcowcYo1rSdDWvIuHbQeeFBYmVLN35TU9ikyegmgvZYJsZOx88je2tT3SIwWrA0a
DR0HfPw7XYgqA+fMwoCj/4kYMMj6t9c/6NU5Mi8ohJVz0l+/XlwMLT4IhByOyfLw
1w4FV24ofgEJjUi/a23QpetJGusBoQqnk0+djGl/miFoUXTt71ZW1Y8DZ2l68nwO
VdaEK1KtBYkgb+62GImr5wp8J4XJ6jxvxZ8e49nBqdboIVhPooGRyxjBFPrG1OH5
qRB21VmdffEF76njHVXctiBKFWboQSnpRbs8Fqy8cVOLCWWge6JmZWLbCZX+hh6I
9FH5ft4lJbRDbk5PoDc2JzTiarPcayn33FhoaItFfxuDbtgWxaBK5lWtflmtxnuw
0yyhO7OWUPAiQM7cKjbVWbW+FJ/fkdkLHO+YP1weHbIVGgNmuji92un2/5qlMMDG
LLAdPmTb+/B5yojTnZibleR02jcNbKHh7Gnv5DSEEu9XS4i/Drjs1wJFj1/5jQHz
90MEAN7jgfac1u3obAD1wxr6Qs+JWyt3ZIWuWLspSPWV0zgW6AkPKQ5J42dTuibd
KGLkLyYzjLRJNZQVvO3VLphn4rCNpS+y4DjjSw+/N/+bRvJb4b+Rdkb05vrRYYGz
pkcJC1YHA8WJqFmXKT39EpMwP4C64xG1JhPcmCVAsZ43OHT/boYPp6kaUa6AWbuj
J5JPGqmwDAzb2gqO34gxAi7KXRFAJxL7NNdUlURxlvZl3Ei0/IXfXeYwtrRSzvCT
rTMs5O54dVRZ6HRP/LSUsp+KX6qdiypKDnWPxcU4kp5nGbEj5siC6OgJQbC7Unhu
ztsCrR6tq/5od3nsul02SE+f/cxByHeMH7gv7fYS1S7ZWpEyftzkLKhOnVSkQANB
fmdPP+RAKA1IaqgVqbfCyior3CZBNlRQCnxCw7HRYyRHVW58PyDlOXDVLkvreCN8
pDTFjZie5zadeVrZKNSZBDobf5surq5630BtZrEf3j/oZms58RrHnmME8s4JxLle
vjkUfotl5jkoRdhsNhp9i918viIgpwMQ0pUAt3Q/gePnmWfSghk2nb+ssUf3tgX3
KuRRtp3Juz9Tc5ui1/8uNHcYLLZ+x8ta2w2ijzagyNXMxEHDXKIXB11ruga1497e
GLnW7LkH1Q4S2oCjqUe6aFT+Ow9AOfM9icv0FpJrkNZo80rfFOgcoXX+791VZly6
3lSIJW/Jfwh6u0tRl3o+Hpv76DZDeAroSblnMJBPatFNGiE9iFcHsvWdyScxrsPi
lbwOwhBvo83Ude4ZB8T+1gNosISM6aecpDUccfpPO0vi2P8iPK+5p/WTwtMXmk0J
Clu1zOmW+e2wZKXhGHjRCZ3GKOrnHp1kTdgrdEpNIWRHjtQYCtH8dwUeAtR4iHTG
2gzJ+CJ2HWPbDiuxM8H1uQORjcrXRvRHw+SEFEeIo9izvE5sZbp18oHf+94eWLDr
n4KOmtKZDVhXFsYQEH+lKz+CPatxYtxoGPROTg7/LzIzVYxxFQIItUCTMBxJ5SDj
Bixs84AtaR6jicCLoD9I1IDopjptI1JLl8b7Kvx8aFUccjZqh/dqKlawUOJBJ5RN
aJ8ValVeEAmUWFba4QzG3ZUlK9O6Uef1Pt5j72zIar3yn7UFKjiyvb2bgEUSpEWE
cpqR7UvTcvCvd+wGKgxQ82K2VP7ulFbWLHXQNBSAwMNY3UQgbDzR7Ui08fV+IcGl
Bk/ymjWj7t1YPAk/R5L7nJkp+anEFdV9th3wfSOeeqE3utqehtBhbWQ2e9i4LaUN
FkDkVsxaz9PrwwZVF+eJ5so83Gm85GViLNu5ermI64ZaAmVQ2xjKtv5OM3XE1v/d
GuLk3+zKYYbe29vUa0EgB9QgxSMWicu9BkXku42Fh/2P6WnkNb2gvHspk/N3sJ1p
JEAx5huLA60FHY+HQG4wP1N199qmXOOa3jvc4ssE/GioQyP7koOu4qJkUj1j9ZH/
PmUqISwb80c9OV9kuSAdHyJ17mPnIoF7SINrtAmgS3XDgzTa6rx1aRJMt2pkZGzU
bvphFCC/iADZy+Iecab7VYszNNCPLn7+389o4dTjJ1/dzVttvbBqnQe5LDwDW9DY
9PV2nEjEH4ySxC6/F4EToJIKOXw6oxWVAPxmINQKvgI4AIW3VffGL2sVIm+/TJTa
QDjnEsLNkJsVrx46V/kYJY95sUofa8wbpYwLXWhNg/fbnC1j1q3pc5Bn9VY93aqg
vqw5mHpbLtzg2D+KmA4sNq66JvILw+XC6rUclFvTA+yzAB0wr2HyBtY0fNBSKSi0
Xjf7o//4I78BbZzHbqZaMVIdLSBeOVWLkUnQMLLd0inNn8QJuM0U6Ki8F8HGCrrJ
EydSEqLZdtlF8SaERm6jjF/9+vlVOIMtCa28D8zurg6KLLr8qHWwJ2mppP3csygo
4ELucUNW/BtTPLkKFyBdGP8Sf/wsJcZE6YpH2hfXDBD4ePxPNTyJYgbam8tP6lnr
b+BzkDOYyineuBPg80jMcI81aeAymRH+MnQur+ef6h3EKYne3KMlzFfRpAnZrgf+
0hjrVCyC6w/SpXr3iXJxRR/vkfNvpuO9guyCwtb4ZVxikQx9b5/NOWFsG/1pWTWr
G0zo29FBAGQKEOja3D7H8lvXxu0WkPZIGKcLpVKmGSAWJRDDYbbmOqEp3eOjbL9j
7ykCOGjwTCa026LSyfAr+u8D6EPfIWIpRLWmq65bEE1B88FT1wexrl+EGGHP9z46
bcWL/HJe2xk5uOvegjPBX2sO/MU3DeUfEEGN+IpCr3A98ZQjirPnTie/HQ5J8pU3
4Tb3mTI7v5lRLDdGDkczmqxin8tcQemnhkL0dK2V7fJ2AxEt4KKExDQLWfealXNB
AFzGgx5TiKN8dGiscuPJaF8fV0kJ0Q4I16NCd3EeZ+V4u3+2k283zJJ07ffHe2Cl
yWkGYR8749uhnqv5LRQTGVt3mI556Q7liuHpTALJYp0FwuvisnoGXEM4NB9w+66I
PObpD0uOajezfTMosqQk0XscRf+tfkxHO0SNWnzkF3HzTtGL/wr3kqzrRmRWtj4m
JqS+K151+l09hQZWyf7FF9+h1lYHUgz52QPr0goWYuiCbF504l1XQuPbtOf4f0U5
OUl0sEcJBECDXZTYYb/wdNmvD9anH9Uhhee/ksrqRxrOg+8nu1RWDYMqItOQVIv4
qgDAnGam7TYnWaH0K6AJuLj6yAM3Ydf6+bh94A44xpkIlH357yfVt0+91NGvE76T
4i94VDrTwovi9ZAbrELiBL1ECdN/iw+UeC4u6fl7AxmksBJc3q+zsBBpiUk5ubkr
HUpB9EpeRH/FUyDXaioKjIAJrrXk3XrHfM9KPGyhGHA/Rk82fMu2ojMzSqlyecrw
StbYJrfT3B7wVyAjGb+tyP34mqIbmEwsAhXD4ajF6tFABv+OrTIE2qynZ9yU2Sst
bYMgrcs3QmhjE/ILQ1kNrZPvqUDBEuy06maTWu9mcl8KpUFRBQXqy0dCfdQPE199
zUQNKtI0A3N6IyKbKM4BSkYdvS5u4fOlWFJk2tsfQvKEeh/hjcmF+2TC5MW7gRPA
b7YP/MU3oUz1/FP045ELItWX+zrVC9i2/FmQDSewryniWUGxnTHbnED6NyLvibSp
UE4WVybomMIPbmrwfAl8U6F7RU1OByGUAUFO7OXiWuqArcYmVjlXovY2Jta7+God
uYJaJtNxGHiIpCZ73yqDylI8uBsszlwaoRIOYxGsx1tmYfvwcpmpBCtumb42pVUo
pvEobyXJdBRYspRGFzdSETFUgoyitHU3M2mOrMwUICW1AkneR50av+iJpyMTSkCE
lnloOxIR6///UFUJktYCtqs07IZPscBta2F/kaGYfiYiIEja/dmRaZz+8cwsVQ7t
RRBKoc+7NH5TKgVuY9ry9z5CaUdixhdLJqjZsnT/z20ESPcRsG5972ujyfpmKvmV
N8K0aCDREHrblOH3PS5dWgbWsh0a8rr65veIRmEngJ8AXG189VJTjkzxcCftwb4c
1+HC23SFBgY9TG7tzhupuKS7DZ3KT2tJGFc1MHk0tG3ivNJR16ovXDZGR//elmL4
FWfIM7FPPr2te3H3MRICDI2ohYNrldYLkvxBAV6IUGvMxZy4pigC+fmbpY8OPwxw
n4uEOaWS5DQNfWMP+5nnIzRjhCIRVOaZo7r+Ylup8GB/NxRoi/QDbh4dqJ5h6fFA
dc7EQUvK5CxrE73gfaOylwiVA3/HYdryDNMyeeAeWwDp0262qabnQ/nU0Em/bm+a
qAe4xpCMZiq9XcnKyhUT5V5vTiyf2xmKmR9+1PjZ0E41ktUPADsBrFi8xv9MBOV8
pVWfkkwYois4y3SRT/B/FBNHX3yuuOCemXNLRji6dxOMZ5Kcpwpy2Im8Fp/7Qm6z
Gz2C+SudjilCa3McWda9H3fpLTdVkbTNtDj73f+HkEwIlq80OUC7/6iMEgcqe6ZL
ZmOyhh0gxbQkvBEg+kzBmimcAi6pTj08RHHG+T0hkTVVAYmoIXltb9NNr2AglRCD
XVDvSoe5Ugz7Tat79fl9zPVhK6U/ctI8p92bge3q4BrXwH7vjLjzsypDQMNOSKaD
CkI7Xe/tRuR/jxQu+nqwzalnFJ7lfFLShbn/Vnjz9j6J0PmO6lLjPKXbHY34/Df8
R/lCOQsqNRUIjPiBHMeuYi+S+a7ZRMc0wqpAhPR783PLRjE8s61crkVxdyyo99zw
lSoidy+HqYkitgDVjOc5iSQTkJypAGB9L2i7I0tQx3OxhUYo4xX4n5Bm3yn3UyLA
RUKZXvuuuDdLF5LStb53lIhGgBmAp3iBBTFjrFoNi9ALtXw5OEhWLvGbrHCcfgZ9
stvKUycGo4D0w6IsYIwuvGGAWG4eefr7Ux5yd6PJkA1jT242jTUJ1Q6hpqcyMPb8
NFa/FtNR0sSqn4e+SiSj7LmkPFz0aivDiS7I2oqiEGPMz/ZcKu3/n2g7uFDs6U/U
K+mpjRn4+9Dlmf1gYCL9Xl5v6+iz+DNW5TlqNPrpLL+gBecMXvvUs5MUBJG6DP8U
4h30yrVZLzwJNXhddNcK5R61Ra18wHG3CrPemerJnB7yYyD24kaf1ZJNvT3JCx6V
ib/d2xVfFkkixSXiigKYagIK91xChwpz7Tg8PUBK3iqmpCXuBgPIaYWecegXR18B
IaPTXTD5AzZG/C7Cb0AmBzZPQOo4SisNCxwawqA/VYphUszJT+vwkkIW93QGiuZA
08TqAqnPwbDNxaZfEX3sMpiOIILLeFqbuPlz9S8fLXDnCgsFUji0lDHBPstgZr7G
O9XgdcZeKc6v3WF01vOc8vdyiqGIJzJzxIuG226zC/tGty435RT0NrSMH+ukcsRU
Nh4wQbVjpuXHxmGkEnZs7XraZld+ojDDKXxDh0iBXpGp5BkQ48EwaJqGR24cHh3P
PCc3Sq+Tub+g+maFB+Pl2QwtpoepPKLNj6uC2sgwuyqvjnYhkAXen4dlI+ZYc8JT
JknwIKOBKPsyMlukP8qc1+lrpwpYB1k7FckMhniTBJEKctrC5UL2IOWfWwXaRd5T
E/DdXvbK/iWVqkywNUHiD0greC3rAVva+kjzqx45w2QBiqNHNyCGX8B2ftTUsHcG
yFaUeU35Y+umMMIvl84oMN8KYcqYvvSoqn9XeXiTsdxdQQkWjAVif9AdyFF8l/v9
PwbHYmKhArC8M9iITGJyrA79sG1EmXvXa+Tvdw7FXWkizuaeN2Nje8m0YxNJWxks
WhW8QvTvyOeToT53RNIWGXSVHLHuQFzUkKFC8ycr6ga8nSdnXRCoXtyBo+TN1fhQ
AUEqEfApyQJJ0oswI5cQvN4UfYuGPfEtWeTdmyASJY0ay1Y61muaVkSEbVcWlB46
3fnJ2CPtNS7aZHJ7qG9eojmAbSrjDNHf229UR2Fl0BwavUsrs0bQOHCLBmR2im4z
zCYjq0FRGR+4y4itr0oSGwDsAxMy+cSX1AJEZBhOiHTgsy9AGLaJkF+Sw8J0PE7A
gF0QVdTPV0khaxDDgSWk+ZfCU9i0TGcfyYpV0OmhlUAHPwMJhrg86GPDa+kdeo4w
sAqP+laEmtB8JTW4DyBFgjm/09IWz9GtULpF4Vq/3kBWSylrBHM8Q7qXkRO76G6t
sslHm05pbxquJr7XR+u5ovdIppxolyzPq4ZtBXcjQVAZiEDxCdqkOZeqF+DT8WAe
MApOBzeqAXX4sycsOjqNLj5dCIflQu2oLaNiXMQ5AwMpiC/Yqae3xe8d0PFisGaC
RhDvA2yzKnlvLy5ranZExr7sJRMoXC44oWIQsiUn44DdpuyK4/gr4V2/lgsP6o+2
PqnSoYM2T/bxhidkhGOOzywB4CjkobU6krfYg0i3RBX7RJ4rfaBpzl7ZqV1wp7aD
Ftq8jW5tuseetLPpWGfA1vk+SQ3JrEEVGYYVUDkxhyjvd63cK8B2+JvMI4sOyuru
0VYZ0yMB9OgZZcz1iC5L/O0ylujWvpjO8hzfX5VzISfFXXZml/7JP00DYSGfDeaO
YjyzCeLffOT7Fcw19BMmLalbOVu+muwtHx+jUDwBp6QnZAbWOhGKR/3Ao0gYkDRq
kocyGgv6U+uXO6jJIVYz3wQ5qkIFCYPLswln0SjFdK3Ozxw4ofpFI7Ye7m9x3YcJ
c2AtKhCZ7Wh+ZGrjvJH6YJLy8z8WpOlgRmQq/sNlpXp3HkSZh7IUdBqUv0F9hK2r
qcpBblklOrnBNN/R/dZu1hYdVn6WobNZ5AEFrXP1x28uPAQe9oth+YcilKAciH0w
bFTZI3OAc9xjeK5ArRAGNDQJfqeXt6ATfgz3+h2qROiu37V3483ZnfOsTzCE8VVQ
t2vDF+Rfm9Egj8lK7kVXsmJwnOu37dfr8WSFViMUp19B/tY5pQWGRVHf6o7d9Vge
INeQiwvRw67XhWaRBDZ6ujzfh4rjApDLr+KoupEnxBpREqm5BhHCwocxTwEMZQm+
1qYJYJcueb9JRBA5VQK/wa+E6O+ZNM4g1LC6yfrdXaaWgrfWY7Yx5QPkV9fxleyr
fhw+pn8fGOmQaYKDhy5ByHrRAaELPMihtWKiqOQlrXjtnKZG9iTlo3fOASU29ujH
22COHOI0S/BbKrk1SUP9W+jVRmW29kqTWKep2NTn+Ww79vUdrKjg7M8oZDvC/J/v
VMrMmCaWMHVuByZyqFN5gRlImNONQf12RVoLcyzn0f/Wvq2/bWq25yhu87SykXqb
1EuO8QeAng6zzgRE3KFu+ptd614guNqty51uCBOeLqqAfhMHmuMsmnF3YzIiyLxK
oxmtCPcY+V0nwHVPslN8W8aNwnP+yBuhASWmRfIA5XyUwZ/LCL26cIqqQUjCP9rK
WTBlh1URv4G4SgM3fMMQjBtH3OzX9YveiixjwjuhfeE+f1dbbzGZ6iLfIcwsZ2Qw
ulmGtgExZXmhnqQ+oOhzFLHLnFrnE8dDKP5N9+DXEpW9exw+eMvx5Z1CZ7JWadNZ
ZgIIq2Eo7UuFyGlIhhymtMt+yQZPut3OlODgSlD6GLaxpxPwFye9aAAJuYZ5aw8h
rcPvlzo21fIEsrBOGtO+i70ZsoIHxp87F/4vXJhlQSkIxoJ84d1EtWfGo4GPvpQP
b05D9nsJFD4rbGD4A/8x0ONzyykXT6l9E3eUbUVPbUzuZgJpfS//ZulCFbCThH5v
jk3Av9Q7rFBirOjmmw9P2+DsnElZ7h4IpCY2Q2vuK4jAGgKPqIRuOawMppdQnSpM
3F1rwPFzEq2/Uphs7JJmPFhtzeb45HOFkjyr8IB7Htmg0k8sQvOFNd/oGfByIhOn
wKun9qWRoy71dLmfsDQEAIQqHuij1f7an9v+okgkYQ04PQJTxX9vZYdueA50NCEf
V6CY/pzgMhfECedESTRQtln5vRYyCOznHqe6w1oI47bDQTcSHYHSbf+enHgf4RGW
SCbQPc5kwNj4SGdP0nM9tnkPmsHrbhFTHJjXdIDr7naX0Az311zd173zbXTb9TqQ
9LblO90T5Zm3sTpLlk9YXn8KIi1UQCa7CKVgbt1grt/BxUCxB2x4YPbRyu9OymVU
oiNczJEcUVwkCSVLdDlBMlJIQ6B64N/UXgv3/gTToTJsQQifv7p8oP08+B4bYExc
12Co5BuD5wW5PI6rGe2GvfgsnMDKt1+PQlwF7zk/6t9wNIUKhDQtgT9IR80j3Rsa
KM3HouPvppB4P6u4TnwsNzQXGhwlhzzPbYTU6Xqdk6QwoUC3r7pnBNcLxAxmstEf
eHJv++Oj4dkZ9jsWg8KGx0r7axM+GSgTP/+ZSfgRnFv3phd/WXg+oax8vrybZUQj
kO2zmhXY6jido3+5beg7E5s8HIK94J2JBNQP9cXM7KGVapbciyLZoBcmXPA+cJ0Q
Y4RV0F3MDsy+JDEKgMNwqI0ej00bWVOG3UMcOIcRKDUx3/cw7e8Yzy3Z0Id1XQyW
+FuAWyt04h+MUY3EdaH9HAr6uR0sLzbXMPO7GGdxuzUGDtf1mb1EUcUHXTwfiQ/U
l/z9I7hfD/Q3i211e03CUDuJ5Y/y2ydfd9E0Meflp2YqKS6MoRsurLFumS1Okp4z
rPZuLUbbhsq+Y8d1jV5wrG/9L0PjYjVO8mxOGLrAR0D/7vUSGqvrfMVw2aX3bdGi
2u2JTQGPgcLGMTBnFyJcvS9CP3aKVaPTf0TChcbspR4hebjKxP8Rt6gpTv2BMZ+g
4l3kR+KC0UVjbTMRyO6r1l9zO+6HX3FKUshKoUp9JnGuHZKY0SY2FBn3S4OtkRJt
eZ3rKnBsJmMkO9S8eYy4Mr1jOIOVQgyIBY5Pahj16YZv76EtG2IOS6HLK4J03hsy
5wbtWKTAa1e4oZvvi2gCmB1QqRYXZ2Xxl0zMwxciBuEcj/+YjOHjT3a9EaFYcnPa
EPxjy4j+cRFWGzSH2XnhvpnZGhWnEEsgdDT3CoJZdhTwYPosmtlo31xBMtuqZQ8t
D78P0BQcd/WsedYl9sC4Ky0lO2VkpUNIU1SgalpbT4IJwXdhftkrNjGHU1g6l9dp
My7pWJXq4EEtuB6D+0jC0qAWo/eO/Tb7ChptXO36GYiwY3mfMOhvTZ35/oQtGVj6
3aX00NatDaookQONkVgHGWrMHhDdQxtuviswbjM7OTdbv0T+jhIQtM7qn4yVYPkm
Z1jvLCntnCYY/Q1G7vZlNGh+6WMVAtOsxXxNnMHL/AajOuNzdYT511CpZmhTZLlW
8/Pl6O88IHqVsbbGe/QNjJ3QdBBXekLtBfepZz1hC0kgrXbjfCtb85Md64d0+djL
ZW2nMQCUb7MpQj/N+wElzvpq2HXb8rGrvvf1nPv6DnCM5D7wLPKbueCpHidh4hOf
+hL+Qi0vRM0I5pKtLIQau0vWPD52v1mTkpXua59hROlH8YyGB9hs1QPvCFj/sqjr
9NCbyvatOb5hTeqoUnpGlrp1UitGQ88AsYWvJDILUJBaj7e4tTpmEgNUo85Aidkv
2Aq5wucQFKRIYFsTK4q+6z0PENoOZyN4nfvM0KqTZCLOU+hleYYDaQ8C5fvWq+AD
V4+4xPxGi3UlkUh1OXv0aO0b816SBvGEd7lAQqxjKp051FKNEs2jAtl02z11DMpx
GnSi9VwEDbZHj3U10ZU6ZIcBeSpOFLOj1zO4R6T2Cpdyh0Vq6iNdpdEAsL+dhgVx
GdxC3cBpYyE6ks4HDe1pbevIBQeomlxhqYF+DufEa608iScMFU4x6zURv/2TZJ5X
Oj8qz6HU25iRipdvYPIGtUWJi3Mq6xbPiMmCCfk1D2DL89dE7gKvYjmX6pfDG18T
X1ZcNvlP1feN5x7Xhp3v8jBl5dtYVK3YPSXgu/tq7uswluahjttP5DNhrAnsh2sf
YPToGfV4sHzjgcNcG5/5RG1ppjM9pwt6z/PxiyMrMp5jCpq8znyLaCJ1xZ7ynnDc
zWmwgJM6dXvCC77ZU2W1S1/vutJtnq+DHksa94IPLsPF+pBCY3dKUxM/+HoK5F9q
TnFWDCn6DIbTbHVbJG2Laan06IADzVGTbhTyvfMP0bguDzDaJ5ngJTU0kH6Ao9jW
Itd2hUZKI83LhPbqqNaCoCdZPNacCldUygaflKLYKb6VbmUdsYllGGZ3RBjp7SyK
frrAbtwj4XZzG5HNaRqowQHIaJDIcf57XMeZ15pVF9fXJ3+dq5tevaZUDlwpMnaP
LvlGZUTpOhT+Il2xy+ByenAVINOSzlrsTBZNQU5ZiveTauADuCun8gSPwG2JrpZx
euM+zZddMxhUGsXdLcenUNXVlDuoBO0DHd1zrK6HJWGKoantsvLq55fLFIGTdibt
WA9xBmTfZlCgcuXNZ8jHtsoC7Z98wGKpAWzEqF64UWQbweZvsKLjZxbnrCakZc8I
olicLd/AhHYU9tHZWkUZiU7HUm3JYN1SWSnqN3yyBdFCc5OT/tdhJDpBI4iPPrN1
Yb8vtcaNpd9BG0wI2I4hwcklOWe0RgIXrvYZk3oHrN7El7851nwitc1mxmJDiqZD
az4+Fmt3R07EueKoSFqj5PGFTmztZbbIlHG2gxPCzdw9YA/JSk/HnAZ93JZchDuj
zx9upO4oSIiFD4/OVfzI/qbCo/WfXBOIpnwYYuG/y05m4oafvtIS01LM4mhY4CPs
+2htEewz1+GLLNHD1k1z3Nc6FROSNNJzI5Mq26wQ90ntMVr5xHkK/P/427n/Mc9Z
Fq5eXzoMI2Kuuw/CgaSFeqUDv0mHvAEIqS7tzc2c6cMSd/sXJxtOZX+YfWU6csxH
1pUmMg3QUKuuwfSf3gocUJKIDfRmniniFu5y3jA1iqHRqqMKJAsskCioogEEl+ni
fN/5r3d0+LTAmAvPFlnydZ1EGdFfPibvHNiIc1800ltwMyYmF4j6IoBtvales5Qw
3ti1wwCuaXaXqoTDHtH2iqU1ddkgmk0TjHa1ah4l0p4gIa7L34tRkv5KBuqTJYju
RjFZwOp9M+oORQJH844NscotkssxX3YBKsA7uxxV8GLr6O3y6hUoQTvsc2UtgWk2
Qmz8rSnZhqnAx3ZgE3fP5zMMz+7eyzwOLDtk4iEOzQTeZ20T/5Y6nQZRI2oYF4gy
rrgaoVAfP35/5UL3jB3w/z5IhU1yG0Fa8fKB2hUQcU1sdUMowfYKz3W4nq4t8tXH
5VttzIfJON8hAkuUpfabsI87Zb5O0SMWs2io6B4MjBY+zQ3jsPHIGqsf0li0HTUx
7uzCJBhehFI4AxB9Y6vWgrJiF+X4bu9jh2okR62/KZHR5YwAyEglOYL6sZaGWwho
CQqBR7gWzf42/lt7YWDR9QpKGIDc/VBw0LMhalsN+hEamZHLsaI6OHAIdp1rnKlm
xB+zENQkmla/5MiarP7g3hLceJFIPN2eVmHfcFIJo32tnkB5xQGo/2Ks3m8yrzCf
7UaBmp0Ct7bIAnvpiBQmjIAUrUsxFd5IimDsTLzEUNv22WIA7S6atYfZ/SAwvz2Q
VYtWD4iYEYQHfHxvZggogpky9Hl6UkH9Y5916SqBCBH6FWCw/pbl/TlByvpATkKC
GbMmOMkY5qoC6ha1mPkzeQ6pAZmhntMeVMwBjkIloljnScjMu0MM4DV68EWHwzI6
uYzyp93kSapJu765mmwh3vxw44hs8bu6Pc45PGhVQCSIekhnFBFMfXYZP2iAbKrm
TwViPr1xoq0WrEic2vuLMx9UiSjPtsCJg+nmJyuKb9pXvr/FgcixOZpCVjfD/+AD
OByip4CCkp6J9/XoS7cKq/o0wmJmAX4V/QO2/BGV3VCbMgk/IYi4QK0Ny88I/KBW
72QQCJBIw8MprSO1q3fckkoenPC0/rB+iJixDlTs4T4BCjv23hxeJjYPYHCb+G2T
Pdu1tTEW3mnR1LAf3AnQOrZ2a8A8X52M1QxTY6imVs4HernYIbTAV1I8VRwhZrXB
v4y90JrtjBrYQeY76sYxW6yr0eKLP7W1bzveVv7gqEAlXVmwMUg2UeMwuEqwDVeW
1sxhb8d12ZPnZQQTttv7bFMgY2yZHxy+dMquHrq4IIAfIkoJJHd3u0batR1rTJQf
Ew/L1eAmZeyEp/OY/sS6oof97g2z2yyZ1fIvTJNoXPXDtGDqdy0E8Pnl2wOOqMZE
6XkTDqDC4QuMXTZT658b+cGokzOYrf9BanHl09AmryD2V+8jC0bqS/vuJbV7XlZM
fo/2rcA9UdI1aK2A2u0DxQffoLuNFyJiZpJzNzL6f+kMwnU+OAM/1v8EU+s8vvM0
bkk4BNGXOtNgECS1qqFvjVll0k43q+hwBbkMiUXFlZYZnP6iGyR3D7YN0337EKeF
OzVbhvAOKqSCJbuk6/34MsQbOYEUoPb2TQykp4GCorFU9L8iHONA0Tln0lV7Au03
kkw6Tx2JPnWjjtLu1F5/aBlnPb6sIBPu/8E1Ts1zeVz+ke6wBg/QhQAx+XkbMv3g
j7JWkQXZFW1RAEL385Z7ydDlJPBWC+AGJ+Pf8S2sVQpZJ3+WpZt8OhJAfyH7Twn8
QP0S/hvO5Yyyn/7+Tvpu+0xohi+iGhsx7WFFaYuCzqkZGDrOVdQ3XuWrrBZwuGwa
+xcNfT9gwQQW+SvFALgnwhklSRafvE6NVJCn1+EXXtY9ekyjKt8Ka80g17nJlhSk
mcfB21Vc/b/MYnADhw8r3RLg+EX50JT4kPaDkIipWeV7xfIFrRBk6YKNwJ2xUfK8
jg8NfF+lduwVgKxQx4aHGm05jIbOQlj/cJ0xUR+nPatw/vwZiZ8ZhvEYCa9nOYh7
zT885z2FvCcbCtciHmyleyZTh6cksxovsdPfl7UbGNm49XLf3hx41bphxIOWtR+t
eE5+UNvsXyWrcmSQ5PRRtTipVAI1DT700MPgPdwcYPtSiawu+jlb3yAdH82EyxEX
A8bamG4empt/f7/dVxnK6pD30sFiIM7arz2bQhCjDliW4l0dDBD6Zt3avLr37ahu
YRgAgxccAeQ7DLcHDfv1/aIdfxHMGpqRv3DHGaRSQx76hArEjw1M7pGcWdgb7W2J
DqR0WbZN4FfB1x+rByE5DDz/RO4EPMZ2h4o9BhjsUJX190gc3YzO9ZMWkoStji1X
n8oPkD+NekdQyZifjG7wQeLlWpXa0ca+9T759IehMWwe+frlReQSD8w+PmuLjyOJ
46hdie/zpSuOtQ+BeWn3/oWrC+w24ObzRpcGNKJbOoJeFZKMMZDyAfamGxAwUlyI
itcfseHsuO8d6vwIMcEfZuSh2CXu3/oJWteBWP4diwSICWWWhbk8aweSCMfiCAAg
9x/+D0u0CDIY5h9qSzfCpXyBWgq+vCGVz9Gve1el/rWtC+cmgR0iF7rMlmkl9Jtq
lfj5pk3pfXuOk5mlR+JNucgP3crLx4wO5h7jcOomq3poxcP9sfNH+HXrLvKm5xbW
XMXRQdhv0BfGPK1rHrqSNzSBmB00OQOnlKIVML/gScR61eZxiYWP73WAcTUBVUaB
QXFXnmquipnQIM9KOec8WJdpmmNRl79HnTNRXgvthJpIm+D4NRlRPp7w++J7AFfD
AF2I9/EbKXR751zl4yW1pN/0voRYlH7IDvxjhdKg4ubWnAkLdkroZ3rwhgIP4+Gz
x8oKLEiKhGCt5U9vc2o9vv1i/oQ1EOxJretMDDRgGs50swNCfBxLuGFHV4eh6oqd
kxwwybHdXRKtUid3JdmJH0FEy1KhgKx4qvPZw1FYCn30ckrE36+YHr+Jb3TaHJ+H
4EhWRvJP5o1j0N3cqmPonFJsq84pmeJ/ieBTUiOn5JWL26fOLUBPW+0zG4vKOszp
7HguEEmIzkzzPMJFXIWva45y4BlC+usQKxAZ5fP/2WfBXkvdmt1ET2lJunBHVJIH
g7j7GBBuOV27k31q2i9+OUe2lfhf6J0LzEmtIfuzU0F6W/hz+5mvfs1poBkZ0uv1
LMPIlhO92muZeP8XaARr4T6OnlWk2IB/5ZcZoBlTp2mY2zyfDkdeJSKtQsQn7XAs
J+pgfZE5HeEVuXTiZ7oYfA+f8CeJ2x8XvHfpHIt/QclhFeRY3IzJSz+eH8KmIepe
ZGJ9UIs5iJfWPwP69srepwKJEglK3oSbpjvSVwdd0Ofty9Z4B5FjgRqzZFmGU31P
Mr2TN/5MHjDLEPWBznaTrgnTHbkeLjsSh9uerGX+49F/Emwy4EwWrjAnVIFXGUqJ
CB14iCBl76gwFOm2HgVsHODoqGhvmby+vKO0Ho5SHXxucXEOyJa6B26Mccpb5LMJ
6fT6tgAjCXgpRfpHw2AISLUof+FOPM3DEWjKN0Sxjd7VAHezE7vrec30hJsa+6KK
+AF7kwzewcJuX6HnMzrBqCohUVvd58oRkbaco/LhHhToraZg6o/Wkmy+pF4EkofO
QLRytyaP7mj4VLPws0Tv0PesxI6hO9OCGc8VjYUAaI6sVozohe1ziFvI9878q6g5
sbN2YUDl7Ap6OrDDZjTuk9ksEkL9hzXX7wVw9w1qOfWssuFzEX5/VGBgI3pgjrcg
bv7EOqFkQAZeE3JqGJ/JOzMP8myzIvr5kNdipyK3LvJgcPY04HFJog16JQpTcQtr
p8T/65bRozlfUXsxKJ3X1CpjCL376YniryINBPqQ3zBGbdQeqRy/dDlANyFkMDoh
AWCxd+Dt24Fg2zqQZ0+A4BZaeR41ELKraDDO7GW6T3M8pjDe3nKlF7NGXVVyQfiO
MQyCba4r+X1YiBUeCKZYHO78hnel7ZVNw9YvqgO4yMqnPer6f4Z8f67hdQXL1Q+7
S6i2IdZrydYaQnE8WkS/n0goub7aJX+wAHPAoKi7ljv5dYD1vDNCD2CEOvTXaet6
RUraMEBJO9IXhKEppgzPC2rgtO1AIYDglMA6qqfihbz6dhyF2HYLtBbnHZOR0qhD
1cyE78j9oXtYJSmq/VjRpT8Y9JG7lppbJ4rZLmdtgWbaSqy8tv119paFUO1ax0H9
UdlmR/1Rqi062NeLe4OnjNEF4XEgRn6WjCIeBsqVqyDeqYWtg36bXu9F2BaZ7T7E
YCpdk8Q9CktcIw+b4QQirTUc9wr+YSyILzqiH7+pUu3y1bX2qQEQ9mtoWS5Ny4gT
oPqOjvO6TtIIs3Xed2VOqY0rQxAQMC5x+AOzgS7856kRP9VeUxz2g7EdoBy6x1Bl
CJQz6zq7XS7dqBB0P1BpkdS49A4sNswg3U3HzvkNWesAkGivcTACMTzLJ5NhQ17X
T1qHYs8ZuEH2tyC4HZJzlpzsxC8c4SNpnw+tFfIfx+ay8tp19BwIRrV+HfHx+QuY
2l1iAfsEaI1/Le1hNDJeLbBteJBmDWoxYIL4ij0uJp58TV0y0rylfbnSr51r1GM6
K2j3SMpcs2N4usdMu+yJCRxBoJwzHn3NqUVscOjCEy60yNHjJvMvR8dlt6M8MCDC
C9mt8mF70TzpviIv7DefkDoppgFGkt9d4b9LcMAnMvip4mWqGNYv6P7Hb27UDnH/
wd/9xvnyfuoSfZgX/v99cOqAoE7MQ2Fw1P2gN580hhwA+/cBAgphvMUdr1v4RbNS
cBpIjFDewlhyS77/3LsxQD9M5yh1DNMnKggYLW8Zc46zFj8Dk18eFT9CEMwEydP0
TLrjeTHDKFfW9nx87Pw1XeukDftmIpnNHpiiQnzEF0DoBhZsP9tG3B2WuXX80ERy
8+pqb7sJF2HfqlkrWPs1To8oqM+FU/uHOsvC5/a40Bgfn36R8rWoZPfN8rNZIViK
VM1OfGw33+p/XlpmrI4VB0grS3GnIUCZNYbDUO6BzViBpcz7BE+CklLzTk01qaHF
38GFbGVRRPZe2AgtYyMtOEkrAOfyAqdYf7RgYMoYPNAbJmheOCbdR2+VcTv8HwxG
yX+zhWpkAY5oD0BkaigyQeTKbyUauZpeTYrKQjialgEe95ZE5L1PZpRPd6RMHLQe
4J1uXaTxfnE5sCvbbBS25YC/eq06O9l1MDGkJTLaaIX4lw79hYXcgGBF0ihyu/wB
9wuXZ7mZoXVrT9kgutuj8vR8u1c4fo5x+3jb2vWbQBtNfwelBNxDOgQCKnJpzUkN
3544xsjrULDKNQCWESyApfwOqlXG4Hl7cVjGuqh5oIoYolDndCwEGvKgRJNbtLuf
0dh5E7hKFL38cO/ZZUlSz2aNUY+BJ4YEzzIyzwPkFHXdObb+Xpt+xx+mHw7jE6/Q
DDGT5RQPbmCjH5gobOkrGy/4f2B3pWhpRbzfwGMhP7QspLPyVWeTnOrrCg720Q6B
tBLvftHXFcmHlCWxuDIUca9xjXq16qH++VSHggs50k+Z1Ea2bF0LNwtS7tAOW7Ms
xgmnihyonG/YQPhz3tfOotaw/GReGX0M31GcFKiezPvDecsifp2mZUXvEaZImueN
DW3d0hwtBg0vX3crVLRyCiayFcb/W1YDZ52YXCFtcTDGLyIKD7XoLR3Qi+dtd7aa
ZwSFmjM1rja756GXF7IB6gjMo822chHcoIZC+aBkq+VoFE/PytJVOsE+UTM7ZaU5
Qebm8RCAHfrrlUD2E5rq7znZdm1k8vA5Z0+2a0EhwCMgBg21Agd2drbWFejg5h7q
AHxiY3R/iPkv5y3hwefh+h16Zs+7xycUvbI43EIdBh/E+tO8Dpz/95xzx9n/gYtB
RBxsZTBkoAbrvHCWxd3+DCN5ToZhwyu/7kxG8/Ckhxpx7QoX07gsg8DlQ3hO/J2m
5pRFGyQkM71GsZuz77MXIapFNmcAK25vMheWO85BWDoZHncMEY66bVSpFLGLsPn2
IrXeBmvm+fVFLt9qMNJgJqi+w6WwD+6F8AvbZLtoBPaFbeM0+lg0met8AYPq0TFo
eYbUO3GPdZ+VCEhuar4hOWtXHNMz7n60F9IAH+UR1vz2CZgaYY/6BzbuHLV14iTp
7xg2VvnxxxGNNrGO+mmqHEdU1P8OjGxEIAaoyx1QatHleZ7k6yvk/ED3JQBCsgHz
AsuQ/x4K7JnR8HyycEA0gy+HrSYVnPUrUzF6H+E/xAlIAugZCDKyYnI3pGnpkvgh
w3Y3j5AUEzOiG7hKq++Xbq4B78EZqZSODBIlHOD1zsuUER/8HrgdnFimebCYkISs
NWwHmUJ4SV0PN9d3LoBoJ1TAXHdV4mos7QKlnb+V4xyyJo7DuZaXpOgBf6xnXMvq
laJOP19oHDtg+SIIsu9u2mCRuqZXnE3dN9/I79bPWWm4w1nLvvD6v5YDk53TxhAp
2roYZurwvmxuDbG6+iZK7kuQSplmnrfu8Et1Iz4wLlCFf1SIQRm5bYsFhCpVcZO6
6MnzeM3WgCGvPSR3m1CELkp5Zta86pxewbS7gPkZeVObflciIoCoDykb4j6VonEU
hpMNiZa2p/LoRvtTdg+gX2zO5n403Pq+STTAKijNe2WMXVkbhI1HYsiUCOL/NZxl
vLhar1dwE3eRxUZDkRhdIyjKALOPMKHCwqLz/YE09JiFtRFKDf0PgNuO18m66imq
v/nKrIXsNcZhpg4vN+wh4/feO41Jwly2apZzPSOiU1yXcHhZcn2scZVT/OX6Zmpp
0ABtzXonufjaUjn1mFcy7j/mo2VxwmdXRO/Popg98joBCBFxGU2OK7rTdVYtwygs
3h/V/6Z0s4+OLyCYMBe9YFISf+l7kIKAqWizfxYrUnjKZjvAoN57vel3oJ9d41ze
qP09r2GaiUrgsBfO0TUw7qoko4OM4zEJxD4d7J+6lYFmNlyybyRUAkogqJG/QL27
HMzakIqF/XQvPrfmLrgHKdhVcofa3wZwXvic0Es8D/r10is0IBlFkwACBMogQ38t
qwEOF5QN3t4VEH8174nHiSi9pX+jV9SNMBH5dxaF2sBGF2/CjRcKpGroA+Wiwwx/
dbI5zfzLM74IJCjV3GP1p/LrirCXjW+G1w9sycNBaEpdIFYn7d+YA9izOXEBr8hh
hBuvlBFXMPiBEDN/PVxzn1Ibxp/CnfCgMtrybTj1ZeKPJVFsnOcRRZoHW2/UiyU/
1H3q2k9AHne3HSOU9MgoHPbfQ5yINRfZgybpBsLSJIhsmv/1poDhQmBBbtM1oPR6
aXRPFrWEdtsrqs4Bdv4pIcLPg1kYAT6m4ni5fX9dkrwMmAwAKwH19YlZehEDT7Xy
TfEKuh1mEZSE7nrlReflwd85vP9Au/MAs1GH9BJmSsPyHYSMKUi5pvmquoygcded
ICKc8KGSPNsIkIxK5eBvnsj89IguMGEGd4nabyUa7eC84n1YJ5ZXSPYIRTpSjoNv
ol/zgyVUH588h/DSE6uamkqFKVHkhvy3Yj6h+4Q/ZsUVRwlv9V9Y9y+UmLm721pv
HFmLK5PjBJrkdJLTwn2+fFDUToCoUHNAK8q5uVbImfjPPP2d5Z65FixRyiLMB2J7
G/EYqW1RUi99I32AbNehy6x/uowM/ofbmV+Xme8XKP12FaGvaWef5SygKw5meGIP
ZnHaewZMGMzkHtr5gfnmu2Xc4m0WtqBwaMI/aY/b9kp3oqgWfkVMpZ5SVaqG41Dc
gnjXQPySFIyaI1BaAQiw10jnMAJ8XOGCrvilAP5OMpNFC2pw9jsLYz4WjaPYlMlp
qHs+tWdHZbZzqkLqSDz6yX5Ke5dJyiIrpRe5mPHiTTjMZ/pp9lq3q18aD2qQamPM
LhqdA/OVIEkTsjWhWsl8CahlCMv8Ea5uQm+XcOwl7aHNoMEzs92EavJXlXTtJFN7
WaGnaf0u2A8q8NW1FqKG1t4g/t0/YBH1s6elUDjdCPo6Yig3yzeDhwMOP5gjMu0C
g0o4ehXpxKmiQzxnShLIF5yYWzN1NflWSh5yQREqUZZkoF1lUuHKul1kNiCSu10n
Bb+nxHGka0ag58Ixq2sVXSYLFmYlTsWd5ZP2FKZRYSGFh4dKxlxO3gWMDshWvEMc
38zqc8SxuxOeVHQmqrCNXUu8psw+pgdT+srLbt0h+HvUwjkuhm7PTK/3rneUna1f
PQT7Wbo5dEylPZRpnx/fzWCF4oDs7jWgIt6wPiHQc7GOE+0EIQE21kHxfvksadJp
H4RSu3ItWJZLx7MczWTzGE/5dODXpU8oqysfJ1A3QoslIfbfFCT4mr0JWE56uYwy
St6VxglElp4/zYEHIq1LTyRtghJrN1dCiLLgsx1Z9SjiMZjXq1xdZEFz2FueDIRE
PdVxmPvrCGdery1QLkxxF9DAf13QcMlBT+8Wmd8k30fwQThEJcp5EwTf/P+S0bJ/
1Il+zmf647M49VBee2/XJ0+NjOgo200dpjb5hHM7cKMKpGI9zpAwS0KkrBFWrrAy
fQ8TPYYH0juMX6YH/Z3+KUhEXn3dbn/C5huC/YMGiTq4ts6QcSBrgH1ES3la+y9w
a+cY/DnF2cpOV3mEILi6VGp4eW6fBuwlcXIlEwzp4IQGm/fE6eVX3UnP6EcPE558
HvcBP8jBlyX/jMCpbgq9U42MccSyNnlxickgAj8KVQpBd7ZQl8NZXJbJHkPMdm72
BSE+vBaalcnSiTEzlH4EQWY/+18tVXaRbR41vspAQpMbCge9bdcIUhWzugi39Uyh
OU7anFg300VVroyjAbkydbnRQP6GWYt/10NYaDfEaIYrwzCsfjs1pVF9ZlgGyrTg
C+4jp3gwOs0cvZyVwVFGHqhzhq+SI0763AM0CyrJH1MUnCvC+L+CSItyyo1KD3FI
S4vYCoJEGfzG1PA1Jx+1p8HU39gOVVlbTqcGDc46cUnB42MKzW6pdOt1PhytdGRB
aa3nr0zmdZMcz3ZWCYJ+jgCuzJxYJH5jYH0sJHf3JmfGUjxMGxCtYzFJmwPJFLpS
YGMFrHwTMwPx+EaKyV+GSydyusC2nSI/EyFtInZ/VSFx03gFXTr1BFQ3tM5JCRq1
BdI7DcPLql2esrNQpmfH1DxwAJfi1jAXhjSeK+fJEQuDwuPaxFk6BUqxN+h4p6gO
4e2hMPaoyoocmE8OdgrPSCeaTZS2/wPO9Uhm81thzk9sMaC6zaJ7W6pEGo+WMzVI
voreiBBalPezTb0i+jTUsvhIlgsxSSss+5mNl+q1Bok0cmTYJCdgdTHn8EGKcWHs
T93O2+Z1auInrgAkZ0jdaUfAJsIOtpJEwr+LkK0Z8IbRM2ghLNU+Cm3d6OfmyT9V
xqrIkPRiEsehsi3IRt+oZDoyaoAo1TSj0ee3kiTiON2ISzBx6blIFaIX7ZWSsUrL
d5xxa3+VSu/fKj/hJI7h6XzrzxyRvhev3mjJfQNddpVAxHOHSuc3aOFOJyshTWkt
txibd0YUj3SsC2UP0Zdsb4ug4dA+MFtlbcoRapoAPCsBMuc1urDtTcwURp5Okdoe
qhf67uZ/ONIUMnEeFlN5+yddTnXpqGnq5xpa/eXXXDcLElfTl751bioju9tuxF/P
mzFCJcs4KG8pixwdoFZ31VNvrP0ke93mJp5UjLAIB2ldsxnDNMyEDTcAeaKyK/qf
f933U2X6FL0TuHRiKmAnQxfBQy5JCH13ty7cG5z4lflFuZiW1Q4MqnkWg+pW90zq
ElMEhdt2PPLp3iGlXAkLwxByivbTloAnwEPDeQjYMDFJ8H24SPYnkA9nTTX02QQU
x228AN3yiuBgeZ0Mhf0k8ayOJP4YwUTkjTZxfE1D2hyrn4DtsrS8IjgRClVLmgew
198X69/gnv4+QRHr4aCnleGHdhXthzKoSgM6X6VVhkU6YNS6p7fVoI1ocvhn3KPn
BCgA8x8k41Qlof3TfVS4V7OGpmlftVhUUB7+p254WvkEOipgKAZLd/wlgy6SiI49
MBREdqMGi2N9EmJ1m0ZtvN3UyTcls9rsH01+Aj1nE4HnmgBmwT7OKPHEMb+G9kGk
SSXXKtuInMRtPrntp2WYb/z5Sn4AgcKFd43w2GCi0ncMkMvje+5PejbJjFA4rRrB
hnawHzVC/hzrdIrXpDtpKKrs0iWlcR4dcbqZI2mCUxWoLXnHY3vRjnI48FguIM9h
lrdtIXgWUti9ncNY9gHegV1/pl3fTLfMKIV7DX9TWF3t+srfki6S0aVYKciBhjL8
Zhgw4eRAg3wTn0yIcc7cROPccTsVdEUXqewpPEcVwL3hBF6+S9SBh/Tc2QLeRgVA
HXUBmcy7Ms5oWMnREJD3erNWFCnyFui9xuO1Ah09uZJ7Zhj6iKvYNSW4ooQjpvtp
Z1CpRWRJix/pqQIKQgVx8+Kkta9pgVo8f15L94wSu19yR8z1ZB98ClwXseZrYAhi
G3AZvscsdST17ibRBuKvTsRs11cuBsz1HR4a+MV4gZ5FfE6Mpd9vH+0I/gCU30Ev
fObzZ+5yGCln45C1zmRZ0Rk0W8VU/hM/rKVVb5NojuLO297XqjB9eeF40+4vshgQ
R59efwE0wzEebqBuuWqj0JAB911C7ZUNG3rU8HAs9mBXptQUHfac0N77b5JBUq1Q
8FZOC+dN+Fj0CLtB7zOlX398lqBkH8sb5Piwx4dtLmhv2gwgOTweEXa4Dad2z/6I
1jZLBXrtBoqJAl5sZ62cwroQ2uft5g2BbOJm1+B0VL6G9dv+n5LIuIVxxwSDZNBT
wTgLvq3FNAAQq7qiHOwNxNahW3l750UKGGwiz9zpZ9n6rHtrjJqA5bXf26mm7jK5
9YXfO2jprc6dTg9WluTANGK02ZYUEu0LIxg+0+ytFvVhdUAU8WJFwbp1Al6ThX/k
Zb1HWLIqfOtYlBcJGjiMVivv+bjLJAh3W75+eq5k5VRUiNfH2MnoETfcASuxVkAq
uWXazgea+n0PmWaHYgJ+qkVXPYjAx82xVhi7kc9zeIT5pcni7Mui0bIU5CiyRpzF
rDEz7srCIgc2CmNEobqWwaZmeNTbQ96cJbb0aIN0+xFIq1iCjvAkFtSAtvOl/OeW
3uZLG+a97OGP/FKX8duu4ufXo0TGmHch3IaPdGizhaiZTZ/g0OqseOK/OnJNnY5/
kkfM8TyLd6zChYe6SHs5ikWQczTxqBPheBM4ZL+zGcTixdp004qA5UIzX56xArmr
iz2e1bHBaftmTgmx1V343LgyHRSu4xfR8bR+nR1fEbItU7a7Tjk8o0EXeGpqY4wM
KS6zUXjACRvuAs4PwovryAak93Si9yjLbNB0NmJAa1YaIikvla2C+t+qijWz0XG6
iPBz3tdr1UXYutoHDZ/1MkAlcAw6VRk25Iw8WflF+qhXwhaleNH2CGZj3/VUQhj3
4Kh5ViqcIjDQiWY57Qmn/2itWhBJINWt6JP1/7UVIpsor8Omyw5NZ9V5ouAjjfUZ
IKXIjB33+wt6NvlnH6ZHliT3CxrVKHYf9Bo66Nu0D14EQUIi5v7gRIBTBEaiTPzg
kPB205UuShQLaGUMovbIctD4PiEjrCtpHXVbRciQL0rCeHP59YamM28AJGE57aOk
rYokZ12jbDmO55mRUAsOChCA+aDD2k93vecLBG0L4nugS6Ur8L+bYnwPXb9+1//w
xuNeCyNDUZRNxcU7Dtji4e7Ks6P7mytzuZdqxrek112IeHJVbZPW17bVMI5nq29h
ZPkU+FpSRICfGRsZaWNTkgugyK4G+JGUpg4Bj1q8ZxUYDZMmQFMi+MrFeQ7KdYoB
j1fCFFeoT0UOawYzXcpy41zCKSBq+95mo4fewTWVrbg3u3mPCYAYT0NX1puHErI6
wz1LXKGCRMpOzZeFdFK46DpecXunY5m6zVKc/KRmacyw3s69/RmOqeJJ4THr1Mw/
Z3ou12jLJKcWEPriYeIm4ZCbFvtjp6/hF9JbqHGAeJY/eMwUbeKJC/RDvUelUKBP
vOSvKtiopVc0sMXrQBGnzFZEts0ZDsxKt2Ux8v7mH4jiPcFaep7X3bQQfohgbnCC
BwVuQSTMg6OaCoRUvzpuz4Vu6QLveAWq5+GYUuPmpkiEu2uahS7xuHnGMyFHYzN9
i0tP9gR+uzR6rM6A42g/w/pnnASyqIVv7mGGp/XsUZNQhz1CHIrSE0CoH3ng3VTH
6Kg9lZG4kJY0y+hSWBs0qDehln4Ak7mmO4t4cker/76xqr14s489DH7srZKuQ7ma
kVdACZRKHcpZWgealaS/p1YKmw4jwsemIGTW9Nc2eAjNRHCWLCeqVjUx6Ltq3GQE
MLKdMOgseneJzG+WN9KIIWzaohBRGf2Yza6b52cMtFsbEQj72ytNWrDmC/Alm0Jg
ydkusf8Fk2/+aX4bAe13jtmScWqVHHxOBAyFR1la24CRKFhjrGwGrU8GqSkbE/WU
hj6nVB5nwJDQ8hXYhnBqHN5yoK5XWKNE2piDIV2l6H+fV8s0FqCg5m7s3aJSs3GH
Sb2cdM491V9XtYKq54jKcc69fVj6g9Uz3p1bYZDhEiAEZEOw5G7WrBKqF42Yh6va
qOzQqZXyrAz9b0gMtd99eXGlWtBccLh3vIHdeVFAOLwcV9UJZ75OnNodyPUNFPZi
hgQqLYba8BIvfjAHOo92kH9vbVgjNc4FMGGbeCBC77Rh/OCbJGD4NcK4NlGAyAnh
5OIYam9iDEkBOawJvXJ5woNeE+8QivqtaVNohpUNy4eRHaK6KlXY9EeU9tHztsIT
+EXjome3vS3dM97TWlMYCt4FAwHIpkRNzSYIh8EHAYOWdiMbI2+mu2DnPzuObTBo
v1x6eUAWcXB+ryP4IV5a9d2MQGI3nFSKlsD8BeR2zu2KbQ5xnAVZnTzJMMw1WNPz
rfA01CfHEUsfqayOBGHvzHBhR2gNnjHWVQZmdQF0b3mHldKSSQGyRKMTfiqpQcHS
y+YebVxe1CzOTZM08nqr5rLa+CcVrP7AdfGlXJUVN15UOfIMgufGHiC68Ep4u2Y7
106IsoGJTCDLVvnR2J/YtQgUKdn1Pg+j5imuKjRNf4aon6fvAH6vGMQcHshVc4iN
8od4weYVLDHupFi7Ludi2rnrwlw9fJVvXyEUSUDAhXMNrCVfg/jYd7eoctk4RPnC
gdM8Tk8ssRtgyCqeKqk2ARpTr5cpFbk5bPeEcJKiOSosUAetbgs4BbCKAStioyFH
Kz0L3tqxTDshxiPu37YC5TSfdUfaIcjoj1y4sBz9wgX1Pu3uMpBD/QWXMZRBsjM/
tfgFHiWCSB6dNMCXjhGlrJ7i5Z9w8ff32L/Hl9hpqdHAo27Kz5mZiC2ZkQffliTj
`protect end_protected