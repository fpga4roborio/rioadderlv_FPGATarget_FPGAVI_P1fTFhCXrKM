`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
ddtXksX2+yylW5zu6QL2Lhnb2d1sD00763mmSITNX595NcHTEkwn0zB1Dry37fOW
FufOhVzEJp80NC5qZ/+F0Vk7Ik02dIR0elf3clrjeJRK85K4e3Hoo4xn7YbFUIms
l/8VZSb14+JVGURjfswrIyCUotIzlzVYZ6gzoZwDXIi5gQIBf/gI+KxNXPaKV+PQ
Ufys/12rjO6aI/pPlqSm0hCvftmBcnezN2hk1UeXgOIuKZnogjOsf0iJVX2aOOWE
6pD/psybjbnsNB6kH5uFTA5frkzIzkzl5d9+YDm9OyC+k84E83I/7/j+rk4L2dah
QJOvksSIzN867/4Qt8qYTQ==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="MvBXkzurAa5VTw+1JJ70nePUfoQXBvZOku/SMmg4TwQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
oRtzZL4VJ4iwysPsC8SXYCzXS8Fw2gtZTOskLcDV+1B9Nzn1zTyNtlo6lNICRmmK
ZRVu2BmCc2G+fmzynYlNTnSa7C0Cuel6FYpxCBlOuk3OF2tzAmLAuDyOH3Z1Yjzk
a0aHuoCdIRKv7BrZCdALt03JeUmXKPdOmIlkVGFl8yw=
`protect rights_digest_method = "sha256"
`protect end_toolblock="Jn9CQpRhJt4rnzZPRk+dOpzAubz7omckX1MrFd4p81o="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 5808 )
`protect data_block
gD6l00tciPUa6pDNTk/+t0OO0nC/UTtBwLB41d4inuAUA3i/ALrNyoJVcBnAmEQW
ptbcNp5fxEUJjnOxnedyZEuEBxWRieZFQnkRdF269oMQOLG0c3TvSNBVgViBMLp4
+Gp8V7J3/FrovPpuZCZmUW7dFJuRd+bl8E6RNPVaUiqAd6EFglfmVY90lkIFhcRC
i/2om3Na0MDp3hXNOcN08ZVuUgbUPxdLByLvgAp4zZLJVs7PSs2c7Mg/zvY34gfP
WL9H3KJNScs/fjGDQGxLEmZ6M5WxuvPuS1iAV7hKEa+CMxHq6EHFBUy1DOp/fpPH
R2GnSKY1yWftYwGqU5Lr503621/cg8RlaBfVNwqdaQp3LOf6czTCr74UmIMklfRA
oYNNLvdVEGo08o5eOMhNlDnE7Z804KJj3i4SIHds2kyBLbDva3z6UBgtr4JVjASl
ky0FAEcf+gQmRz9EWksSZUXRS+WC0+crJX+EnlDuhJ2HgAcV0pD2MRRrtOJI8yJe
OnHtDp8CdWbKYauVph7G9y5z2KTgg0IAUz6iOSATfAtEiuL7yeLTQ6kqrtRJBr5V
q1u41jjiq73ZabKVaFrtRHPBcmvf/NuWB1f3iPWbfovaWG4CClFv/0ani070rM7j
JLTxj07PwEFmd2tHDpv/W+0Gp/8NjClO/LdbW04pBMFAhtghBpLksPlJR4dTOjx3
DxSHSXwR5ngoVMRjMMbOSmMG7Ws09PFcnpwvdiaAxONK17YVETOKKwzTrIjID8uW
MnwLVvXt9qZlqJ3MTiHv7pVGfznuwVrhW3Cs6h0tKKcv7V5FO2cQ7c5RAIAK/aLd
jDIppMuml0bTs/aLYP6VVIWbrXCXpFxqwjovi9PILQByOaVjv7FhtNk9ajSD1DNf
WbXW0OtVL8uQDYBAB/09Xv/L6qlRUHnmj711uiO06a2jt6h+flq8ra8xCQFvnXoV
8pd94Es/gbE/jQtDUiJB2T8x7iKpjn3au1iUPrUHiVDfE4buwB30JyKRU05WhY4h
gRa1/AiVRTve59HVqvr5KLz/EUif1h1y8x5JEZAj7+08sq85bjPPBslJk1ZL81hI
7dYV4oGBhPrrPZVzBicw6pYv2DOtKQggDLhElos1TLpZOjw6A6jx92Ph8WWGSD3P
9BUbo/GgTXg/mzY8qj/NmNZq65YqI+ebbO49OsFLD57A7gAgH8NbHGQrTBVXLzMf
1SvtwCscoU3JVwTWRfInwRd/XpX151rVALmtsDoS9rMHn4p3wsSgqcP5/MZXKjS1
PNMhSsQSHwNGvW+OOp2f4OihEdoiBB4gvpdEPXPM73CqRfrKO0y+pUDa41rqXf1u
XBL9+QTKJMarTEndP4cDnkiu9NbzTtq1kpMEw/FbNFU1x2Ld86KZLROq/5+ruidU
1PGb33aeUZmFBgLFSp1a/eHc1mf91hhKllnY3Pb27n50RNaGA3GdfQXUf43SPBIb
1EaMLLmzsotvzSpUcn5LceVOXPiR0uQbZy4+4sYYA8VpXqP9WUadQ8ovUQ1nxPEy
WDQGeUcZ/FUBjYJOYEQvG4N6LPc1HrefJ3jkK0v8zz2nxfURrI1PDugI0XcB8PpX
sPn9z3tVVXiOCeh0ZgNrd6Mbi0vnxK6ufcDhwPvt/4a3OVg51MbIdN8txlMifMtK
BD7kzOAsB6DsY8BXcPPdSC5qHqDM6ALOuj6uPxWfwoUV7DdBOJj6Pk/v1+1gOFU8
FHw9NexkO5cLm4Qu0aEy8WbG6CG0tEuqkksW00lZyN3cx40yu+3BRtXg4Oum7E/A
3UmIZRwznQpRtwK/MjFeAQlcAGw1FIvFkEr485lm+1ZlLj0uCtAFM5tS8t97uROF
a6bBTVH8qUPlLpi3iRjhSqNbTxMMVkJrHo3l/pnnSta69Eeeb8UHBifxtLj2srFr
1+LukNngt8UA+Y7ct9L5D6z9USFVAoKUuqyWMWSxNADDgOJ9YulsNmXcVRIa3t9M
P/bkC5W1E3QlSH0Rd4/lZcVXGG4GJqJnBeTTpH8B01MjOT449QubRhdPHB+K1hWF
Nfihzw16XCR+p6VYd1E7uFaef6AaFd1UFPOAvPzxARBQ1R/UYedsFxSXoLz71hNs
fzw9qhkGUOaUsVi4oq64d76Nh9ezoxey5+pi5pP4/WrOq4niSAZR5pIfcQChpg+w
shV8X75QBs19tBYIkZq+wb4aarOqZJL7W2/TrdMDZ6ZBodYzHwKgT/wzr+6wLR6c
AOgrjO9NCu5rHYANKjKX5O4lqnHSmU7s4BEX4oL7SU0Aq6x5LhsGv5dsCT+v0rTz
xsI+wunNppOItFzlYxgG2eq1cvzbgOw9OVTvMJSI9BwQrLEt65fLHq6egRFiHR13
KgasYx0fJJtTmwv2RzXqo3aUwW+m9uwjyw75Aa8q0I18fKwO+vZ/3pV98j6UfHQr
wednRpugen9CVBXFf9h0doI8uN83w3n1QOhXoYUqT8ygg/Qd66ovkjx9BfcjFC7g
y289eqO11/sevcUTCYN4fw4lIBp3ubDBGGrqwMc0ch9rvLUc+rL5TrxOuiDBceD0
czAaDuF7VGEto53o8+gcd7j8N2tDkt7aCKrjcGGfmdEBlJp8Jd5/+BkPJYwMrpaz
F/iEgtCBvuV4B315SI2b/QFXboVuOSOgwx5sRMrArnbnTCLHb9lEtwayMD8iwtdM
HPcGXv97LcK30PxgSQyZfJmC35VqjPYTM61/vVsABQfM/FvwLQ6BuMUaNcPpgz3g
oqgSn+JwgyQpPo2/9DLLVf/DQEkRPNChaUeLPMSOuDwh07c+o8GwX7CifxAvgYKU
mIQUFQISaBsrnrGLdymSh+ja0WsP7lnaLZP5BX1SFp7DGvHuid1dmKbEET1PjvfV
imD3VOrAw9Fy1tCunsz8Z2xdbFIfHXXFkuay3Fmv4Ls1JL+fsQS0m3u64de7O6W8
Vp4A2IFUBjX+eEugblFFFXUF7MvtW4kkHRzlHtuAvdXX5zuqQhD1Hji5BTrZ9wF6
F/iSw+/TlxYbFgMO/UAfZT44bG7wHCg08vEuPCVkE2lGLEtvSIL6WuGasxKWNHJi
i9kwFL+SeUh5RXX882dMqk0mFSNeF+nRqY5WIdOAmgUReoEepZXAWiQftI5nV55o
xP8o81u/0CD0w2epo6KboSRnzSuRk7LhzZS+ZgGJJmap4f2B9WVAWdj7sJ3bnYiV
0m9Gz9IPY/EOnHqQrIeGSKSyRW8nc7pTVWyvTiZMfaOYSJ9IU0aOMdaEACK4+ZgR
ezqUHW8YdflD6Xkg9PnpU7Io5947+8grI9/MhXwwhuDQ1cfECT4bW1phXv43t8vF
MVCZL6S50JgkHBKtrdhomNg8TQKiS9/l2yESSGdMv3kUwzB6mfojhjiOPjlLCb4T
KwKBiFbTNNo72qnwUyDTsqBvWwX9LCmGh5yFRzaA1xhq3FyWdYfqS/qgDM+Fm0+T
IKNAFxlcB/Rv+lhRKdE5C0GwBhbWqFY4EB35kIEYYZAMZUsd/V0AqIwa2aTK3LbL
mVeJHxqlw9Kp+kTQL5PMxtPvphVA3krR70LurZZtI3aBLs8MCzO0TkQWKZrJlFjF
uGEmgEr6nwpO1O0yPsfXCdKBCS2LgyNXjg5yqKTST8hOHwcQ0wHbeSHR3wyhG8Mc
uIvRSm4mSGKzBhmkrgXzkHxbzYO0qHHP5pRZt5LFRRyG91EyTKco/ZhHMJHPgHIl
Iaaptun35UGOWR+SHk7q+ibsFsoLJGhO3v2jXccPoG0UMLqwAU5rPuQK3oJbzfD+
0516i0GXxHVOUccETxiVcoH2ea94TDIE9X2AYkv6P+nE1h44DNqzevZHfNIT961Q
KrbJjU2fWFi0lTiiVMLP0qUnCLAiGlX5GfkcAI57Xp+wL/J0zOqgyF2/X34Bptuw
MvMh6R0mKyPgjHclZVhAbSyL9kbKvVdesk3lKydeEP/jQItz08tPc70GUJ4qyn/9
RvJnj0K4an3aFiKH9BphInp7XTsS32OeF8zhcwFwo/GMcZ2KtZFoMypWiQ9MpKjG
zHR9MKtTy05lv1JJOGQeovBsis9IXTBw2YUsxT5ZMbkfJ14dj9NGhs5gT186M3Wq
x8VRy/XwTwacDupTJsyegZ7+DWm2eSStxQa9UksqV204rlbSRr/2JYvQEewjInPH
H3Zp0Xzv4nG2ixS/voyd5Xp6eJvnSmEHyIEfqDTN8vkxqSPO8Ocmgocy5/cHNw1R
mpOwRqt4b0SKT2rJRYvwPKAcgQhND3SYA1Za3S6z9/iGsS/0vUgDW0VPDrdjETWr
KhOcbl3oN+pHHYbnScULwlKJwddbVp3wrlKWntmNEcDhPTnUDViAVSNbMERRDp0a
6mtx/IKRYIxNCJCUuKVuRL1ZOjvXOeQortOZPuDl1ME/yDeyTiBENrbmDwonV6YB
nVVCXV8d8zRtCGzmTu2GGcuFcrlL+y82f3foyIhSHTyueYiv/2uDSbtmkGewPkzx
b6LiirsCujQ6KdTOsHv/qiuH5mBmYxj9fG113je8i/bAwd6iOH61RXWkCwMn1jhB
Ay584g8ZM2X4OXIHSz4YzHtLtd3bpQnz7u5XBsYVjrHA0hwo7lJ2zZYlfC8L062H
thALuDaRUiGMCl/kQeZ58R1QhvmkRg3aGPJDgpjrBxwHZh+Uiias1p/NFSFnVLl9
t0OBfZSX67gb+y8N1LtID97UWNfRSb/0pWpdLlen7w2klRt7FUNFAndL7ryV8A1A
8keSxLZOUvn2U94dni07/WnOJ5tPjAeUxiZTX/djr+p/hzqtS642Z+AU8M5o1eIg
CQ7l7JxM2uKyOLaT3sEejewhHDP0084grlBk+lwxR4ucf0+t6P4ObdZNE+J4aYSt
ozVRwgBCVCRjt1sHMK525mT63edL8+/3MZfOivSC6g2eE3/i0KuhUWxjcHyVJG8s
V2CIVuioogULhDrE/7FkA4F5OGea+NEb5E6B+kD68/bM1xIUxYHsXLJE04iVhwkS
wDIgBMvsSWcowsHlXoAqrw/yiZDJuAouK1i+Etpe8bAwllYVnegRR8zjcGb/Cv1A
zErjjBswoFOk2NyL07ylvbSA9PSyWC57oeGmMR8CTiOA87+3ADu4cF/qU9zH3XCd
IpcXBU0hGYB+lYjZP+/ovozuhI7yJ2fKNZ+/ojcDIL0ZQP3VlaI8mdwuAFCVPjDM
3kDS87dYT0Y3cDvW7G7yrcfKkTonsWXDVDQgX6IV7bHN7Sbhy/LHdwljCJeLFE8a
bl93IcwDYhRdzBkdhtXzmrGAPQHg15Q+7ZI5E0yYdX8rWkx6aPdpw6uFHn72HOps
Qv5tjWoGd/CcLnYl2IzJYOptKkaHARrWvhTQNCSB1FBsgDo/bdphWwoyYAnmVLJD
TW1ZlRqulodruC7yDTtBpTF+Qe8NGlHqSEF6npQrljuyIZOXWmCJP2CdHpWgUwMw
+Yr+VWcBs0aTVV8+WI0rKXBOx4Na/ha+C+CzFgDtPvyiEasGA71uG5V0ZjtB0acE
R+4j0iCGGelJP2OfrgjirtftpfpaToBe6SMLGMh/L6hhMXf+w8yBY5b7rznTxO2G
FKhQY2K2u6lXL1dCIwfYtetB9bN+aCGTVBMByBIl0/xhNAH6g1MSiXPISR2seqdk
BKkcxHDYdnyx3OBOzpmhhx2Fs5fFr60iLHp2t+p7ZsfmDegRiGkCHb8pR+tMBsJv
6Bck5Y8sCS7xeq7AIRmERH/Qg7WO+zrsPVEOVU/unrwSQKun19TSwQXe0DwIDUCC
5J7DDm6CxLzadahfMtKaMMLps6x2aaPcDP+pp/GbA++mxIcTwRK8irQ1js6NyBDi
tAmkcBMi9cBPu5L1AOG3wt15IidPoZ9L+3R/p+RDd2/ApiBt0RgaW4BGjuSajscc
yqq+7I1pHHD1Quz38L7u5Sgrn1WiyFvvfruRbqVYI4g7NvHboEmS/+ziIKnAntrs
K5rtwckvtpbjIojLQzr3QZZZh3oK7uKVugPLemORmm4b6BgkXbfa1nWR/DEw1b5y
CnO/iS5X7Kxv4KUqJwLay9uvLTxutWtQU7rsPLaCET5zUN3lI3Bz4hI3qd4l+bBS
/NaY0xQZ4AtcBUVMr0EpnYU57KBSTYejB1zJPPCzAodXe21/Bjl7nrEEbJVL+0RK
gKWCvjEcUg56sIqK9XWt5VAc1UIoZdSze5IKFjtA5zU25ID34+N9NVvdsPT4MLEM
bjbTsZjf951DFr4OMqutRkL0PJo9R+p7Xv6EAqGStszuJHI8APUsaVHk8WJjQ/rI
gSC+ZGq+QnFnFIU1kQbLKWj4fQnhk//kcRjK4ROosc+gd+OuyHESJjt2L9/ls9xs
XOqPBPlSSE8UWLnmPQ9oavuGeyOMK1KLUkI6y0n2VwHKITTpGzwfoPxlFHg+clt0
4yubcwJhSHAYImxbotcD1Hb88QRB4tb+UJsnjMkJTFNMdguGnO5l1C8iOgVWX7mz
0EnqfbUUlbCaCrrtB3Y/aw50mSMGT/ZE46n1+QYJWh2e+XiQV+2nxsSnrgcLbMBZ
zgwJrwxYYBiKoFRQvn0M6BcRB+9jqEE/O5iNhw0AaTOMuaXycnC1Z3ue6hOwAE+k
dxX9jRuRIRIgNItDdh/SUGKrdJnU72uDa3E0x2LjONy8kVtSYsWoFzloe+38W551
Mf88ppmzDlQnLMfx30afdaXMUazn2QFHSEGoaP2ydZFrv243DYJggvsvcQPR6iRd
RTKuRtZAKFjmgUqmdN7b0EM6Ydhz3/5To2MvsQaUSaje0Qr/T/YKyv+6bcYdYHWr
dM8/8seR/gvqOlgJsDNScnZ/iH8WZSzgK2tlG3x95G3XxFF9Z6Qp76Nr1st4S/ti
rarIXouf86XKO3k5IhmxjuhX1d565T3iTw30UljpxyraAAQeCMth/NiQIoOoQbYE
1qbFDSY1gxYx/LpWzJpPGe9kMPKTTckS2AAedWW5hxwVRR33k6R6zYjRFFSN4UbO
FEZtR8LWPjanB1e5N4qbPt4kYUH8LlT1AONYtPZxPHKX5RH3NOo5ywSEnoqZL8b8
yPupzqevDXISdi+l4gB6yate99q4H5ZVSvbw9a7qGP5FN+loi3fCD45NWxNmrXYS
GS3gZDSneFBNgSf8hUYynlntGH4mVrWfpEeNAB/4shs2V4wytMqtIU+7SBMKR/PT
UQ5Kpv31nvkM+8Ugic2K2e+S6tAGx5gcxXdtHUKOVYbWnXFAQl/PtVczEEJimthT
pvrQ+O1HOBFtrJqAGN+7P/mLgCnsYvQ9JdwQAjZJTVvaKXafZoqzsgTvghRB0L4u
rMRy8sy8/ZFhtKHL/QL8OuZvTg3wVzGV6HbbMCAtwqTgbRz4WlC3yeoe2naUTT07
y0lsfsI3OYD8FsFOglvZ+70JCs/WA6g1llMc0HCVDT+2x6Hwey35gMDId8BjILyP
pAgVIRZ7vV50DYCivW66awFzCad7Cr4FOOFXXgDWzgtD4WECuo9gN8tlR6+SYKYm
PSN4qi8txgul4uX9OQAZiLGIJPxx68P7Ya4SCkF97551jYdrNQcDqU5oFQ/7+xXK
DGKT60xA5UK3R7NU+zLTPHK6Z1ZcDHomaOXVzi74uQ/VD2RCi17wG8iuVTjgF2rC
d6wxpQJzDziQG0Il3AO7z3zPkIXwShYmLsQr0olKGXajt3B4JHE/8POW74QyARKN
Ixvn5Mw3k+WEwm20Nd0vXEsOP1JHPmD3s7oYfbo5q9uvtHv2X45NJ/pB0z/GYmAX
`protect end_protected