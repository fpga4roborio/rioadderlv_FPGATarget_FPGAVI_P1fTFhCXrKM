`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
ddtXksX2+yylW5zu6QL2Lhnb2d1sD00763mmSITNX595NcHTEkwn0zB1Dry37fOW
FufOhVzEJp80NC5qZ/+F0Vk7Ik02dIR0elf3clrjeJRK85K4e3Hoo4xn7YbFUIms
l/8VZSb14+JVGURjfswrIyCUotIzlzVYZ6gzoZwDXIi5gQIBf/gI+KxNXPaKV+PQ
Ufys/12rjO6aI/pPlqSm0hCvftmBcnezN2hk1UeXgOIuKZnogjOsf0iJVX2aOOWE
6pD/psybjbnsNB6kH5uFTA5frkzIzkzl5d9+YDm9OyC+k84E83I/7/j+rk4L2dah
QJOvksSIzN867/4Qt8qYTQ==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="MvBXkzurAa5VTw+1JJ70nePUfoQXBvZOku/SMmg4TwQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
oRtzZL4VJ4iwysPsC8SXYCzXS8Fw2gtZTOskLcDV+1B9Nzn1zTyNtlo6lNICRmmK
ZRVu2BmCc2G+fmzynYlNTnSa7C0Cuel6FYpxCBlOuk3OF2tzAmLAuDyOH3Z1Yjzk
a0aHuoCdIRKv7BrZCdALt03JeUmXKPdOmIlkVGFl8yw=
`protect rights_digest_method = "sha256"
`protect end_toolblock="Jn9CQpRhJt4rnzZPRk+dOpzAubz7omckX1MrFd4p81o="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 16512 )
`protect data_block
gD6l00tciPUa6pDNTk/+t0OO0nC/UTtBwLB41d4inuAUA3i/ALrNyoJVcBnAmEQW
ptbcNp5fxEUJjnOxnedyZEuEBxWRieZFQnkRdF269oNLhYHlyp7RoaKwZ2iz7cC1
rOPIQORbL9OPDjr6kPO7NmlAZeKplw+w1zLsVP9r/nCBwvPO1jH9YPjYWwRby2+s
VawPF8HyjVrlntW85lGf9jQYUpwbzKhjF982Etzl4R2sPPQ4HGJzlLeeATaw+zkP
WLBSczvlGAbLO1rDdh/kecTjaJdS+HpWhDXDoi75/Q/f3gSdciAUtRKYIcJwsxSL
Q5HDFPbYEgcLLPyJQGH33kU3pFZBfEXzGXh8p3F/ke/FfrqG01cdu+m569opyJ+L
ys3KzBz5jn6c5re+DgCjeWkWT2+lbVyMbaYBHuM/ccXvN1o3jpU+Dhrnc/Cn7Q70
Kne0OWpDWZLohsqfU+44YlyU9UM+ZuVDG7iIh+Rsyt11KneCrzC4m8LUOiUoLHYn
OGNK+ciTK6XypvLGntpp6hn2SfAoQ9PUzSJtrBlcEmg5QOdahVrDysS0jcoLKmDl
jfI5HSf1aiz6lvHT3eeRTULRdtpaSe4tGYSLxrl5RlxwUntDh6L5N8ShXnnlQ4lD
2v3iLKITJKCZBIvjBMVRQ0+yyNhVZyqa/j18LSSg57zbNvbkb/AaYhLp8Y01U6DP
J30L4437GCuV+l8dL2wZ9BN6iMYT3SBju3tlVbrLEcvZrhLiSihp+SdLSv9rQs43
24XpkN+9GUveQh4MVw92O4wmIW1avxBK9Olfb9Lo0lN1AHVku64YOu66UqYr6O5i
RRBq2lWWnM4dJjva0LJZUc+1jpHezLLDETwa886ey/FuZnpqMmJ2t5gX2yOLDbR3
vHY20PUN9YtfBjE1NnNA6QIzDOIqkgWL0m3SOMMWH1gh4MtNkr1cVDpJS0nS2N/r
3zq/Gduft+UOt9QF53zDUuv/Rv1ZXqQygC8K+Y1pyK8HKbWjQdi/ZOfnEVs43v5T
Txg65xiH/NKvcUdvSXrf0baQ0HNmoypQYGBNqB+eDN2MNMgNXOlJdsAlIEA84wTn
D5m+m1ZspCUShApnYcs0fWaBP0CAy1AqBEk4j3FSYG+5jOj141s0+FXSWDt1JfFH
kN+H8dcFcOQf7PtcThidSzk7Gsm/PeFc6xZZmG0bKQqY8RPi64j3KQvbkrM+UDql
FuzvH7+0dxXYz5/0nsyVqIzl3bnIrslpVQpzZ6pZ4+ADkGPENvxe1f9J7qvNJrO5
SJMkmsjg3tYL6Kd8HKheSBp7bMNyCM9PAajRKkEDwFwuxYRx7y6hOhl1vZHRXvcB
od3yCk8cTU6oIHXYxNIZeX6rt72U9IUU4S6MeX/aT5p/Lv/h3EX7tIuy3J+6r9QX
w6JPKaAvGCijYtVOBYHMj2wzM3+QS8A4eeB+lWo2hd9oKsPLnLo7qgUPPm1Myf6l
6llo0U6kQe815MUJnPwbl2HLMRQJaOXeJMvoYVBH8fUF3mgA1w1jOL0sZrobUnHO
IXtW7nNH1oO3nbJonb+cuBKaGAySeVRw7AvSv82ubNq7lFRaW7kNDcF1DjCqRRd0
dMKbI1cgFhqMqDr20yt2C5R6TRVEJVK9fGAA6g0Er+IKcv+UnAB0+ZCLO66H1v+H
vetzxFLAbJLQKOMBGWdT+OR50ANbd6AzLCNdcZKlHT7LqpIS1Em0HkCeucHpB663
vqDlIxhmmF0fkGGzdAR/9apoeYKWuQgU0GErgQsrEs3WUl9P8xK3RlMKwgsWjH6K
yys4w3XJXv6zYB2BR7KUy9uI5yVB14EvaC0dj4ZBpWvvKvX4txbHdRreyWOQJpdF
s9QGKX5Y8JVL7JQYiaBd+1tpox8CxcrfNpXRN1PB/chj83XBP9cizetLo84gUlY8
dZTO+4Rh3eEWIatjLDJzkOXykxyyf2KF7zwz06P6OwZ7hfriKW7QqWIXoPmUBnGu
k6eK3M1ZoMiHevgBe97lPn0OG6YccyxIcEi39wypvZCNQRPBDz+EoNXuUSd3D7Q5
N8EWQ14d5ef6YEyS7zOYGV2FYAr2NXYxds/6hO2dDPsCYJmLcwjobovZFwweEieW
96n/t+80XID4LPsoy/EN7Hfh4CmeaV3OBbBFFm8hhI4LK6GPqoU8QncaVqq+80Tu
ojxr8BYRARZrZVZvRUDrMEg9wM/NrFrbXU+3nOXWDVynZb4pHc8dXiMTwPvu4D7q
MwpIllsrfvd0boVRgt58j7EM9WKaTQRDfrnTxIqkl96nwWNL5tUcBEn9lzudQD3g
HN75G7pcIcbIpuc75d2yJc+lxcNilDO1NgOD8FzyfiJqRqhbfAr+ixVHaQBc5qbn
QoAAX/C5t7uEQd/5zQe+BpYeE0FJOZmuTvNix3kuUfcg1O6Q1epgp3EPzbZmUpSS
JVGVGR3wC2MHIEm2IcebP40xQ1cMYQY9+9JXmdDeayCXcnENnzqPYU1FZhmXoLfJ
iI+pU6OAhFHjyVu6IHVI46X6Sh6nRmGLIOrhIQdm1ponVt1l/FIf/FFUiyV9bkuV
ojj+6xddMz00l3AuCUFj0WxrUuFxupQ/mmXgc3+2Mmj5HO8eQ+aIAIj1/gG2OyAu
ljXXNQujDFTeQiwpkYG7NtRsYcwx//Oesn3NEbIn0Efmj0Bm1Rs/45TQ3MqQwdAq
JDlQ/CUDX1RQ+ZRLiPrx1V9196YbhkQc49kl9+BBHlwlFyLX7o9XHX9MkXHDpW/l
io5yQ2ACswDuhdyx/ajLttm1qdiLWyKKIgI7B0PYwxokYSBmzNc06pDfI92F+APj
zK7xpV2xFQKDBYFCwRaUfj5wZI1e/poxuhff6JzVskhicAtvDKqa7lUbOqwKeSWa
1zh+1gGypTgJaXRTgag6vq4bNCslC9D5PqcZhs3foYk/ls0jAIRzTvhcV4tqSNta
CwOPc0MF5mLKag324YUzbFm1ET47WoCa/9eUcNfwQtSpOOVvRL9CVCIy10z5PYtp
aIcCHagT0t2hjwdWhloEkIV2uqctFHT18Zk28Q9ej9RXomkzc6CYQbFsgjQ9a3+R
g/kM2EprBYyQTkP7ci5lFRIh17KCZB4hoVObYqNwodcDHJRaemulgy0OSl+gocVS
zUx/kg5pvyqiRULNjbKz5Zu9usk5GY/K1/h2BjUNR9GB3Wsdz9PGTbGHS4PFEux9
FFt286yjgWpwTeAFnwYBDOBS44aTbEqVPSACTLq8d6qWGaq6k/qYMsbe9Y00pOuD
M7o77WvxxpSoPQwFXvvabqN8Qv6pqpyTRTM4Kwuclp9ehuoDX91flCZv0f13d8yH
HavC1L5fACO2kg9ERgwH3gfmnJ4DSVf9STQ0qBGAhfsEJFLL+TCgvJfA2ALG/s1T
j1/QDYbtX5bfoLheUIrTt5b/sQqKF+ppTLn0mxuY7pGbQUjyUg01pPiwi6OEe5mh
eLPMSVEqOP+MIPyPoIJyx8a17bENMkmL8a8pYR+gt5a3G1Fuutsdf1Bn0UcLX2qk
Z+UCxeDcif7UR9OSHID86WNJIPmGVZfNMBoVqDu2nKpEXAb4wZgGn1w9cjEn4xEN
xfwkkYZmVwRoVk+iiRGQjaMrlVGrU/JK+i45YTKN9C2ynFO8PBeWqHVwuwIc3ubs
3HmgfSBZhCBYzijDdvtPAtoxLUC6n9JEh/guEN7tg5G2pXKEWcjNCi1yq52aovYT
UaYgYy4gl7cPMqUGaQUOEhpRvKIgeBs+ucrmz5GXyIGxOVnrEjvjyXZuiPwQ9ph7
tA7eLrYLMdwRFXeaoE1JutCUt8CwU1Y4Yaq1iE4WRt/2R8N2NIxcEI1X6apfGLrt
fTYR3FkmWJjLcs+BDvfEwmTiT+j3C3lOOamVcUEzBn5payCfHtUgWyIk6zZxxsIW
iYbnNOQSCS5t33b+jb/dRS6+QitHvVqADD0Ck2z/QzSP3EwxpgLbZjb2JDjFsxIc
lbs1mpkWPe73DCcQUOIBn2bcLFXDbJ9m7JUURyLNySl4AZKB55jy0h1hkzC0vflO
P6UoBC08UkIC0v55A+CVogg8z71qOWr8oaFVNH41dm4Kql5HCsatH+1J3w8dj4vZ
WDzB618WWlQk3Omn0ud4417tw8snBfLGyMS2cv2H1J1YLaff6mCulDS0L4VDeB+U
17dWm3vuPXD0CJ8J2nWSRdEQvr1KVVnROHmP9v5nMUubW/jln3mV/hiHYraFUjji
G0CF00mTGZr88fo5fRj/wQ0iomMeMGbxLwXLD3hu4/ECbaxPDD5O46wtR37UtjYP
HsUgPG2WooalZhas6PvZDZU09f0QwRjFNQvnopBu8MnHBLXsY2McgPJcvdXhvMa2
8I9PTNcM4tp7W4EYWZAgiJb0yNeRkIgx/xkP8wHXmbNtAzmzilP7wsTS5gQNVYMG
VQ8ZMGgBNFQlCEXxcdp3ASe9XWky8ROHZcx/RSxzEEGiyo7P9EErf18pICu0jUCX
UZ47MoGNN8m3LOlSUC0wcIN7Z70+zsXEq9VKaeiITRtlM7vCTUT4MXEC6YpBt6ua
Rp+Uo0zojJ74iK5q9+WuLR3vaeOF0CCZDq3BmJFBGvZDhF1XviTdAmyhvvn+Fe9S
jIt0kmuNCcPCbDuPWTagsTE/939ebjlFN3qevUkBX6OtaEqVK5s51TJBRU1sK4gI
FuUIR2pec2SiBXs6MeXtWSDhqrIVCJLnOGfH4snDccghLW3II/PyFfyuyXBKwuu1
G/lUPSLWKMw0iCnzy5ZfobkBtIT2OnjyvtW7p9TmoWgpG5rr7RoTwRjEBqPIu/K+
qHlteJj5CSsfxk6Zy+0rh5HOemevscXTlfksV1TBdvkYmy24DsTkiZY+pbrgNk2E
SxPy2/+60UlXr7JiXW6sae3GjsjhcDMUqIAbO/HDWM4azjdDmHZyHhDq1ZRyLR5g
wSWcKE2YJ4FAOkMxadKrhm9+a5xhOnArpUc7qf73jAQVyYH7lkqYQ8nYrnBOfYgI
SKLHF9yjnOoNvp4Bri7N1MeMQ0w4KrKSBxYHc6xI0Pbk5sv0nbE06ps2Xdvbnlxr
bYt0Yf89BlPmSkNftMarZGz5boopZNkWaq4UDbDaBpvQmtR3zQbjLK9f+seI/5Sm
pPqcz4kl/94DZ0ZspAq4YWwz+JYsE+7rNIiwcvSpQ+gXV5ldL70sw/k11kN4BlNt
GAFLyfLmrgVBo1/ZGze+nOKye9yWLpFCV/22GZOUA4oo4z4wS0b9IsvcXYSgPHa5
0QBkdCfMZyjMheeUQ1AW0uWsTsj17n2Iu3MDnCkMRjDD9nPvUPkr5dMpJlVdP24k
jeMQGfmcfv7DdGRRCjCjVNE1N+e57dLuhMX/DwxkyZX4Uoti4Uj8qBJwXWTMug9K
YnNj5Sg4TUQbRWLK/3DiF4UJp2wSrlXloal1FLkggvJwa0S2JLRksdJdlBnOw3MB
CelBWLyQ5NQ6vJAGj/Y5klqgn5EHKysiA+TBzpI/kiyOcphDxQepocdgr6glblx6
f8zlSV1f0pmeRl0uuOKvwMcsZT4a2A1cWQ64Cb3vUmFeESMAQVl2jn7pLsMGxWI4
bG0plwQWVWK+PUYc/4nIH779LoM+lUWyOtjQOZ6U6pzm83NN2NVpWX5ntjNXPfJB
BUEF+fKLgSKkr+oTbjAy7gEOZh00gcX0wfYXzDujcX/3LrgWkzFAtBERtswP3TBK
iV2WnHKHKZeyE8X2GEGvfjbycov+LF2f9wdTCs9E+VcgKvb3BlDTZmSpPYj4ihN+
3GR5XZ1OjQkQaA3sKuHVxhXoq/gfRTOLGjchvDteq4jManmWJ6ipIeWJ9yZ/qrW8
59azlkUfHvxltb+Z7k9bKhBKisd57LBCrUqL1nJfteZV5sNLyDnW3ro14bQ2vLuK
O4p/v/BIFH/ERuzckwy24gpBZhf1y3Pidhl8010NdLgWO/dxIE3798lfTAZ2OxkA
KdrjYctOlevNe38+XFhCH4TP0KeZ4AK/4v9N9kxOtnYxPPge34UEEJlMXbD4rlxJ
C9Y0FjSv3x7Jb44x5f06RuMG/qL1W3UBrMolZ8VOp0Zwkowmk9kCb06tqYX5BI5+
AcdlvjCemAHhk853HRHKdno7M6r6Tl7LHxUcCifjD/HgxZ3CRysr/+/2mqSu4lu6
YIqr6QCWroPUGSEHMEE98ioTrKqXXpzkeTbGgke+K6LrBb8twjpubuKZskwX1PcI
+oosySrnER7wow29mTSXaZPbnlOtCqNgY7J3B9DYJRDMcqxKPROafzaX8m4kmZvl
jQAhPvw6kbbc+UFaeufcXpyJW0X6RHR/4DA1XHbChrY4XyOS+6vDmurwI36stsK9
1fTHzEd0kBQt8XZImSWymJ/iARwTD/2EJkcdY02a5hXlyYv0/TrNbgTSwaur90uj
+XeN8BqMK6jcu9Z4gjOGwXeE5XuEzuSIOpdTrBmIoukIuAuk4771cu/ghQaYL5Hf
JkGVdWU1E3VWNNCj+0oPV2QXzs4nJ+c+bfbGqUn0bbvAVy4DdxwOnldZ6N9tB+k4
1DpJhPBRWg5Bfr94SmAHdGKIkEQAiM+T6Zay8Nh09HgZNVYmQrXt/KDY0FvFkZdE
DQxRJFzFBUuTg8qznaU2rbc2cQ5L+7deBAJ+XnDgXiowH0irgfRFNTcbMHHQ90ot
M8haYzjSdqsDJy2hgOSYiPu+CiyzWNa0JAbWbTEzR+yJdDIlIDEgfxcKD7uSO6GY
X1/1MQdJjCiGRiG6vgO3I5NU51cC8UvYeJdBujXIIZtbmEEya8HxLi0I75twLTrR
aiiwvE6xwX2MEO6kAxn+2aPGSrLWYXfueSHCGKcqfMYe450r8NWgp4gBRnwaA3p/
HoZvXfgShvUO+T3L9M2k+JP4jU9THVGGjBXIsGZRyXKZFGMMfYQ0Jp6iDsOn2PCv
809o35ee+VY9AsABnfxo0lFDTZcLJHrfz2CsFPh7jIbZCw4QmO/qRYTvmBBOY0b3
kbtQIDXBB0Z1jfHXBBh9gzsp3DiyGH1o4gumfDZGFIg74T4lLcB/ZP3AImVWNuN3
7ZPzrc34E7EZwF3X3y+Jbe/IsE7DWGqk+5mwISrrdM9GWienq8KcjOYpYZgdKzkI
Ey/QM75ZH7r74u7d2I7puwNA3q0viwDQ0JFvG+e7F7gecEiGra+IHbaxtJjqbRMV
6fb47JzZl7J3XCchEoA5ezaTkFnMG+z3DxjnHfVsa2Vpz/8beZRIpjMHdGW5GsKP
qXQPa1o6IH2i9i7MwhUV8R7JIJmn3oIjnrBC8QO0N0YgV5vKmFQa9CIvfgPOQyNF
s2dF4uP3hgOpMHkCpFt80Mm+8lHQoxLrd9ts5wsrY9PoDdx5YB2NPkBbkPq+dwLu
RPv1l1jJiDUNAwR+Mve/La4MGe+MywUMduICxx3Z5YFayf3RZ77RGeEtCTnHo6/D
h4Cr68BULqJvFejZNM2xuTxM9+6WwWD2ONZYD9O7IlJiyuIzUwZSxGsVwz67tTEc
eEMmscVRLXclvvzmPVHDvByRuAye4PzLIPYzzJwujhoHcD7UE2P3ve9+IdcnDgmc
QW0Fauiu7HN9jNlH/yihI0VGsOksVYkOF6K2cxRpfagHWH/sDgxzTA2Y2do8ERrJ
Cwb83/lqbpztFeD8M+P71f7pD9CPTIP74mFaco6RI6AG9VEbcmbNB/GMQZG/9uQQ
2KPivwRrcUuNkIESk8+L6oyQmD6Gz5YJzsFA5yt1isjDLFjTGMzHITsuBtRP8Den
bJffUGJFLGGRQTbs79zzwMz2DEbmjNuYPuyF8y2vFjN/L4s7igg+n8PYmf10El2v
hdIEehphRbgkPB0I/dj+PlkWwXuiegPLmxdQutoW3Tgt4n91wMGjuFr93yrnqI0G
wqYaVU/oHesRQC7wzb0q68JE9DhSffyVFUW1OxHaThHs2ZNLKyUUbiaqgWT5sqVP
MqZqTcsuvkxMDROfcb/RvORVy32KTu1aqtRZD3M5hlft5NNU0XSvfj/dmDvBqMCl
4qKwVzM+WaSG0rOIqTTRYYQaz6STTbc0lpDcBM+KhF8msX9w1vaFayPYZ7VqraNc
8vnecLEZFl1OXKI5vmEC8toPur/KJlu1YZIXLXKPQZCx8guvRdWi+oOQgD3Z2HmR
ojM53ahvR/7breBMDYGEQ/JitBTzUwXdngNt9zkXw3qUrBksaZlKBGYuM0x92kvB
vlV6LYkxEimso/ngBLyGYXTKJfNmPcCUixQkMvJ9IWw6ZSdgAwlferk8fUF63Qn3
3Pjnm5RX+xil1n3bWDOTv4aO+MdR76hqq7NQ1HgZpPDcWGbkXMAIskGWNDae6/N3
7fekqRa8bqHsft3U8hapg+Z+AjdvkKCCPwrMYwk+ZhGby5XsONA6tSgOMqYzzjIP
f0/LhiC2jaw53klTCR4mD3vrjr11Cy77bxlZr5BHUf0pNIwmzzrahyfMHn+B9bEY
SlBCUZcKNBYpTn8WgsKvG3TKj815gAwHXq9Q+zmiM5Z1HSgh0eu7Yba5/63ZUG0i
61kjggeRIgWp4civkolJQytViQ+T7cCaQ+kydh3acAVjuQS1MU2bH29Rs/b790gf
/7Nkg4M+MRlFh171G/YqMF6ipEiHjSqyXXM/8PIBN221XejkSf7Qf3O9rhfQqMkW
VNlQX338o5JdJuwSFI6+U2uqIlweHMgJRPe/0KfHcKR0rSZ0feUcD1Tn+/FioaZ+
FtaN7Eo4H9TgO2dlky2JkTmAbyLHTOkaeYFIG9MuUnRpmNlQ4IsLeZ+FpDofzgzN
T/hDbrOxzrsWXbnjkSvn2aXrs3No2oQc3b0l1URfLFNrgZFvlsZ0tw/zaN+ygU/C
pW+lbC1TxTsEmqIEHKRdvMgG+0MojF12m4PuMcSO4XoU3imG1drM5mihmV53Vufw
5nxKmM1HWypQBvkBlEhX6/LkCuQojU+Wf2yRX6FiPDCGx5aDiLnvEwk9K0LHG08b
wV1tCjcbk6RqBmP34Nho3ObjRKdYlYrfmu895lTvXhSxwvkNLWkQNKb4VDrf9AgI
MC0rN9mzzoc2wKgqGALNKgYXNgoeTkz+EQ/vncQIXV273hEhe0T2ynGdCQmDvLyF
7ypG7ka8aYfEeXCO1BdaiI7dcBODJ48jJZpcjmxvMXAdNqCCXggvTfnnkdd4v4lA
2G2Rl27YrxdXy1y941+O6YXflStJAWFokJDt1uYD6pKwT0dRchxmxXjTgh4LbQ+m
1La5ECB1pQCSnXwn0GBNwWYb6BX0v7bHEoLZHE8Q/E7mVNepfHWWv4+LEEPirdS5
xc1UwB8VvfRlqiMp9vE7FXB3rMOLj6WiU5K7zZ0CIR92C5TlY9qz0EwrXBHsXvCR
b8xvAF/wO/ZEReTqaK+Mx/+e80Xd6lTJ4u1MqR5ex/xJ7rzBBHvW0TV9yT1poEyb
nXk2t2/g/7LoiQczvxSMBH8fi1oraqauboACi8dc+cE/U0HImdvqRHQQyjwrQLca
gfe6Jf35nHRwaC/AeJd+lEwRM02sOWv2ppgYCXX/fXc2eOxqzLC0odTBNptQ9j0h
/9okYG9qR2XFquOz+Ic/UlN5MewYfTeKgCfTAVgG4rKUoYVG/56iSK6ZXX7eHWjb
ErSOgNXFp485PxjGhm7wGqClIiwU1pXeBqqTvV3Ct9nh5eMfF1qzyym00l3Bt6AO
pWoWsEqSE1A0KiHNs4DCFCCZGoGA4eBsbcc1nodhpGnpl/6nsGvasrLr8oZcSbZB
zv0t7ONL6hS+pOw+abCBUoCwS8Usz4+eFgYoYcwhp5wFoDnsa2OGw3UrGMlOoyg0
gEGgXe6Lvy7MNHVW9TTkl4l8vUF/DP/Ymy3UhytiJu6DtVkzk26NkYDXRY+jupml
vfSxk/FTrBTvSgJO2Qr3ur1ebLfay8WYRU/Sm4la0M+xqehBpUkfqI4F0g7YCOQ1
TKAewwsU+7v5g1Fhxvl/2PUblWneByym1wJvANFsFt1kAkVpgWNM47lNJbz+nlK/
m5XH2De3Pmk/7bRCpqvKuK9TL7gY+PVVrpIsbyfDo8xVNyzSr8xxzYABip01ad5i
MK1YB5fQvPSFmIRg/oG7qKTBMQi/gjRd7o4kb6bs4Cs3R9uuGild10mLatkHapV+
MCQ2PELzzQN2AzuAR4ERn9maG+xWALGXd58yC30DEGeNlZD5Y+k7Jes4Y5uZ37IN
9WiVo3+9nmEqv6LaAP7kAnZzztZTQqmohGGuEQDCakHKO7voxLmIApMWDR3+UVtw
SU3ZnKkvggKBW2gSpBwI8cRVKT9U/IR6PfO4GQpgQH6O4cbrONTSr2RGU4vrlsqN
oHCZIoHRpuCwFsaKwYQTtbaI0P6k0n1XSmmzkax2vRpgAFw1UPRgkxLS5tFuMHOh
WUEdwdO72LECJoR9JESRg1ncgPeWEtIeHe+AsLWJCK9+K6sAIP2p1+g7zju8XZ//
XibAlzCEUtBcJyNtGtwN+vJGt/6OvAA4cFO49SrXZnKwrpccARFP5aCNWA2rMvff
+Rzqhpe/mCDh2cmaPAHzzL+vN3hA7fi+R7BMnh+MfsD3irM7ZONltXg7RPYDqXck
eLXb8cU+xAFtjug/as5d5vGPj7Msh7SNSKMEFwEkI/wqPwV37KrgDo0+Vona8Evn
md8SC9dkltAPtr6UJRjDDPDcMh2JS27HH2yvd7r+dS2FK8vmdmgd9PZ9Ju00qt5+
qbLauvHqGKoFRKdkXMfzZZwwsvDEL8sSaHiv5Ow822qw7gym1uk5eRUMQpBKBgbP
ZeMISe1fTCvYagdak9QMG6u1w0y7pJ3nvD04HIMQZitdw1NFF6oWC4e7pm8R0bKK
kWKxBvAWSS7aJwf7TV7Hmd/FWnCQDq/Ymb6Z8zgVP9k7WbW2a5DIqJHULcwTCt3o
4N6Z6doOPNugpoxXNYVusBkgis6YhRTC5MuWTH/tnJ/Ra2Zab+zw1FvAidLh8CWT
1hKHJ047rxaaxA+WenAx13mIMxrE/GjbYTgLaqFTystpxr6UARoRbqkmXFu+h20/
Doo5yQAn+iRrhuCd/qtlP5uFEtxUW13MjizNKP7tHuAacbX+0wi8bJA1+Z1+E87l
KuU/XNsji+c3CQuJsDpaY55JBBNhPmnIaKivWkzQeA4EPQ78nZY/faYgcuTfybOH
MNVimuF+ozfpyJhtcamT/gMUJXIbE+A/tgAZMmrrYGyUDcClGo+SmCcGOuN6PT8V
jGcu05E7eEDEX/rlFp4ouZZJ8sVJrjnPJl+FEDyrteeK26743OC+vTJDJd6fBzh6
OvlXO2wLnkuXeKC2y0sfcK+d09EzF+CaalaQjB6xDZdwXhmlS3VCMRikMA6Us5Ch
oN18ibTPuGapvL7qhvVesZ64OZ6II5IOMAGKKMyO5q99r9spn5gRky3QrsNtVvPb
VMgFKaFsbJSgazmplO4k0mARaZ0LBoD1UfggPeKrAFHLUp9Qnvb2ou7HnYVbzpRO
KsvYI0YxTR+Dpum4U7yz9kxofKuQORD6l2WoPoPwvrwZlPeQ0/N7BkBrbVTNVQAS
wRpCVwIAWOB9IgWU67E3HZumKfMYxlqMY6qzBnbcBmuz+KBW1jCMz/5rEsbWeIsi
IqjAuobIpIWrQwg0oCjKtUrYafHVf1BuVYERN+xRiyS8T+KzG/j9ISUz8Uf6RmkV
znvcQHq003tQAPurytQa9+mFO35gBuhb0r9sxPgk1I9kFB7MnESV54uI5/ZdpvKm
sqLFVle51HhGM3ST0M4rDlOMlrjRPYSCvuIyHDF3BIryA/kqkb1+Ysjt3zRI2QUN
XNjzMwlrIiRitA20/+v6qNTSYyKbEebn0qZJtMYyLVczGefV/BB4Ks/swCz5KFBE
nPqnWmpbJfCXtBIf6LRjYFBQTaaFVYLcHfWVH3ZG1YHxYLpIzDsrdfn0463BRlGY
CIoXvw0BN1+m2cio+/aYTFZI+zoML136sM5ZbpEyHbnX30wqTuL8NSZiVumtJHdN
JHSkrtUz0Fa/3Dpux7uKpshiZGJqLlPsi3HTcaYKdHpoQ2V2wpcS575xk6edbvs3
etjCUV850FRLsl7+uTBBajU9oqCjE0Iv6aeUXu2FwkblF+6tyOXbMfhBvg+tD5yX
cmwgmFW+0pUVK8rH8n6X0mxoL0X5V1hTxmjjK6b985zJX11a/FdcFWKfR5Pv0O6a
vh91diqowfLzLKHPkyoU+H3ljHafh7Z1SM4w+uY5f/45vg729zPCQT0ReXMMGmNr
9D/ctVOQzhN9pZtcycW/GeGRcMJr5XDB4OCW1npboBW46oOjzlGB5RZooDcWCClg
kRPXuzzqfaqg0zt4IzNKK6D/C1Of33lPh33QczLLuO5O6mfdscfDu8iFXwcDHagT
Be3HxJFp3CT6FbmDD2tOdMFxvWL6cZhZVlg7l+J8FdVp5t8WZrOn1Ap0K3ahGMr0
g/9RKqiCKKYDFKsQnW9LkGe9G1IsO85JmL5b9ME0KC46xA3DPbzZ7arGSLJeKy2h
cOAWRBCljru1KXbpPl9mKazB2pqyV0JjcrsdZHN91wmzwp3uoNQaxtNRtlS5L6Sk
9Y4dMRws5K1iWqmQZ5Z5iyTmbfcLNlkoIF3eh3XvqKtczI9XqySjow7ZynTjiqwm
BBV5CqrGbvKAWgPSFqPspJSm/IFvQviHclN7sIqUyGMZhqvQ2dfo2T+Hpb+eEW5h
K5wh41ZLsM+vc7jnNrWzvGemmZiT1mJbh81hRglSk4/rYHaO0pGTPoAmxlmXcQx6
fqjOzKz2Y/Z/+M3E3tXm1Cp01HdDhLvF8/sR4s6Da6d+ebWUGc/JZ5EO2wx2gJyo
cbc2rbhlNchARwa+IqfkbKBzZ9EtpiTOJBb9wy8lZwBVywi59uBX8aXfbhaAyE+8
UbmhpXm5+fVZTMDxNfXFNunvPk87u5pL+urmHNsM1Ak3cv7T1QcKjt9AQobF4n7C
iRG2OMgXuUpKCS1csgjon6/vI5DxKmlZMda7VhF6knmDCZn6vWHrxqh8jPYjpS1m
T5lNcXM0Dbjc/SDvcZ7a1cFmfCqR33JakvwJfO/Nj2tqgjEi2fwQvx3eQPdvfRL1
ejOxOsdB8JLyXPlF/ERYqGLZzXrAiHRsvy6S5WVoI1gRIGAxN7PlAcMLQ8dv3OPr
Y6gsICcEpp81Q11E1bxO5ehasP5iI3BWUaU1u7JnLGhfP87a9uGT4D2tkl++g1DE
IaVXGQjoChnqc2h3TjV3zb0/Kii57OggpBmd+G2kxV/1lgCROKnnPtmu2V8blxk5
o4rqZ5G5IPspJxEEpgK2DXK7yfDCb3tX3NLRiFhtQE4uv3JlhFzyi2wuQqtO0cXd
C2lROqt7DWjYbAtDVh6eEr/wuZu99nQoeUmZCXUmmw9TfIb3WMipreruk7p+SM+7
RH837IXJSk/Kd28muviRvNhKqZYELllebmAc+Wj2koh1+BIk4fN7f6a5VtIwPyDF
fCh8j+9c9vAJ45J4y/qCNB/Ve8pMJfijsl8HMTo2e0JFOiH6SMPe/04wGbhFZYAK
c9GjtKZMhD0D8u2nJm/X0hbDf+r727i4IBofDcPO3GKe0SekEqMq6hGNjQcy0W7i
4o0zy1kUfD+wehsR/kDbApd0BBpRIJx7PmgQ6qi2arT0tuf0YtpecgQQ6Wt1svuJ
jHHJjnCc9y7M8EtwjLxDUKxjT5VyMx0NTZxeWL/DKXFe/zpFyaYhVz10DW1D3J5n
87JatXc19xfIWmgTqiFk6ZatHJjpOB0z9Diqr325ubzANvHWQZjsp5aDIVyBiLy3
t4KpkpsQ5yT1Umw8uWiyQPDXFFZkm2My8tYbU8KMMRM036ROGN5g7RcXInha3jRg
mhTAvACvh4Rm3cxwc6tAXFkRQq2sz3VQ9j46OVZgzcrIfoLOcFs3F+e5IZAkTJ/D
jTeH2H8phX9E0nnzAE9BKR5hq8f6o6+8EA4RjDRjuvP5cEFHPjYnCy0TMU3x69ik
pY6D5l0bZBL3iJptUrtvb2EIHCl7ZXO0S2ILQfangLorWmOieTEI8smoEi6fsIB/
maCGvMFE9r1JQo2U9InlukASuaptQU0yKc7xksRXlGlg/cqpwYCQYZ4v6RcoDwIe
pQB5xdBQ7HwsCstCYeWVO876OhuE+qzy1UXm4H/lZfIvCK+zxp76nfVmbXpu0iXn
urq4DlFQMYmsOUaHhrEngF0XrChhT317Po8HxX8CHQs+lCS24HDvL72Ef5NP4H3Y
D3Y6GQJwuBCRFF0b9Y034uUsr8V/jxwJgHx63NEkybF1QdOSGfR+evgbCg11eScO
VfVkjHEyNcwo5GlU4ppunhnqvDm5mwaVtylZgCWDrscaFufyee8hVIMrXz/V/Wie
kmDMq2QPSf5yUKtgM2not779wMrW6SpU0qr3LI28hj5QeOcNqqZTEypPHKUYebI7
DgTFXJgcV2j8AAZ3MuslKCwc0NqM7cnq/j+qwN9q/Qzue7LmDC+LYlCZZZn0N47l
uwnKhuNByO9FD7X/oZfhhb3Z41dQ50asEtM7FMPYqp/Xk7GKBODeeHs6vhrCQHLd
Pn16i9VA7KPBUp9lMhFNxYbB0O3tvRc8lA3hlkRPoo2pYtgJie6ArpSij8cp3ki8
lSqAZ9X8PpzBO3hlaLyYSJI1qXzAege/G7+WBQg1QzfXxRkL5wTK8EAt5T8leuWO
5iWjvOPnPoU2/YYi4d/7r3EQC+6mqt/8wJWCs/IJTvssyxKIU9BG+nJQbCATA2wo
T8wDoG0fTcV1j5EDTcdxyeES/tngF3yrghi89Km2yPnum6FknwJvKrxXc4tL4b9+
sZJvxcYOqIrdEe/57wLso08MBR2UkzwibM9Is7wHJuVzK91Rw/686ivQlVqvSGe3
l0BJV34Z8SPHASTL0/rqv7LryyFAyqFNPtyvww+AmCHwy2W9BL1w0ajO74XAsKuS
2n1u4RSp7Q2SgJc+5eRkPPezUH5cmCxiniblOPXINDWot/yANz+7QroH0bmHwFpH
v23q+bd7Lw1b2QMjnolc2ULDOe3o8BvgSXADQQqJwqFhaI9C40R+cSQ3XOg9y1wf
ZjMsEpcjFliomIM4OFp6MSz0SL8e1IIJZMorffxYDOhbjfASiuHPpYCVoI0cAtOt
h6xv5XC3i00gV0/xR9YM0C/H6CM0ah4khGefCemqOu71u5UPf1EiZgisMcmrxaSs
vGCSRgEP1u4AoMydiWeoNQHEvIY+KfXYpENjkE0BVS6wW/uBjusla5C0VchvOnrO
RRXb6jn+Oafbsdbvf+aMXXU9tMVndY0hYBsUUFR81M41bsSQ9OIt0BDGNWx9bLdy
ZJ5cCle1OGlJgMYCDEqMNTDTopn8jZDL3qbUOUjbI7SaIR8xl55wPwnTToLu9LQw
Vw88FSoC5nAbdMZSXmBY2ADkkTQysNljudoI5ZiSZfth9KypBn/ukFVJyfdtQuWd
7t2xBSSdS7c6GwVIE6ccqN7QqE5cCmdCf3+vtFc37P7k176EbdMmzrt55L4Xr8YU
YsFf07OozHdVkIkk/omw24g1yt+DKqrAmBqWHeGwKv56qSlGGdPq9KDuHPqdQCkp
k4PgiOtxReo+3xiLYPOya8fwVhRKd1Q2Alx2RKQ8plWw8Upv6Z080rIDqgcAlYtK
QNVYGmeyKMEwwadS8Uz7h8DfcY5jj8qoFmTsGmV2+Bddy4RC5Cuhrfss0t1lnesJ
bIwa+5lFwhG6JFX7zDWJAuBFWIUPt0T2j4wx71b4URbKrVfFffNs0DkOlL3pKvVS
VM5j7kARpfvYAi39agaa2Nn8rQDiKgAscc/r5tdFNEqZ+ilILgpMQhu6ZHMPGCqw
zXpa6uGjDHalT+MyW9ZMLQW8mvFKsI0KFfTH11K5YSF8SOyOc1fUKyegzzTAbjgJ
uesvqV9V9OyN5OQyCGUy55UNZCvMqwg9Q+cQt61YqrARFHGe5SO8APP4JwhcPqH+
3YDjzHWy8v3q9lcbWXZfzr7SMLOZMIhyUe+gE4BBWSXoAoxsljRmVZ6mhlwLCqU4
bux9obKLLaOomeVq+AYdEYw/pKvmkRo9Xr5oROunJ6cgtWzthaGYqc7CYFKCYj6m
GHpNi3Ith9sXx2g28ojFcYd6FY2GwT4JCCCTpaYv0YfiYdWu67y0Gn3gSvc/t76J
dyYFcXahOXC5NLzG6vHoWdTsvGsavKtwN2/r+Jj9M24Wl6UDEtK3/6TYgqMxvqvo
WRA9V9oxVskJw4JQVk/AzYNAiy2P9txa69aox/RrMHjxlWjA7LKVwdJI5nPEt6RU
ZhajDWVtk0Zm6L4RcD11HNBP1S3oO0hX1bedNHC6TeMHXxs2EFH+YX96TMH6/OQd
DeJiXBiMeCswMNMzFprLxlI8RXiIdJJKqTBieBx3G1AlfyLvRlY5iP/Q+EANTVEH
SohFzxmns3SZwNZudBZ9jzN9ZwWqRDlalrjt0yK/CaftRDP03cQ6a152CO5CVlyz
NWGyZVDNVFkt7J6mv/U+xJMNG3KTY7wO9ZkSWU2OKE5JW462H1ovm+uJMXpVrUeX
EnSF7NBxSypJAhrtFtMKPTKuuMsxPYmKXmBeOzlJ61uDZZ1Hm2hB76ehksRKdcve
VdnEIpX+rv6Ovoyl5uwJlGTLjOHVDV/UuP2FRRBPc2oi3lV7f4jqY/myTF/KgDWn
gwYq4jzStbsmUU12mOWvlNNB3fQX3eWKJJI1rxRU85Edys1dSfAXRggr1cfcsyES
BDvYuGq+E7InyeaIRIMg61F0cUBO00JamTRGLi7/bflQtiPIid310CH4THSVu4rm
mV00L/ZdwC2/uE0Ggp2lMmgcASTGsPVQBmESUlzd0K3YzdFDs68CSAYiJOpNib0M
ltdppcOUshiDfbceoziE8zSmITFEabh/D2uI+X7j84fRxpQsWBhb6CqRfOyxPH+g
5nT2SHr2ufUSl8BzeK8Afsn0gcoAqBIIEDweqG6VMWeIU37XVbGLNnrKJ0F45mWT
docDqC+BoGFYeyM8GiBo9XLi+TcwW5g79Ltc7ZGGXrjVPCThxV6eSkQHbQlSFvAt
5th7X3icH34928PKzgvq/ZaNR80c8Iw5S8TvBp1LY1Hr46YIxIBp3pcLTc5sblir
QvE4vjywU6/QaHdwvvXg9QsiudmrdKTCloslnk9zZivZC2nzTbeB3QL3PSStkmTl
M+R+QRdzYJW+PnDIuvN/+H9j+y9Xbn5thPPBL1K6n/mpqeWkIKSLDVx5wC3Wy1KX
mtDaEJk4/S6fChjbJYlVphF5z6mM5Y/7H0umqUqUTZcmiMGXbiFcEyiLMZnaCCKo
S07hxMlWhKCbEnYkDIFNr3Gkq19wpHq3xOCQdADjj+uvreWofM5r2fv/TMGBW+VW
eTNYoeLRN6IEG8AIof3jWpmX7wP+zMlNXVKbw+Y9mBhXsKJdIE4rRyxPj9YpPIhU
ZX8JUnUEdOrPl74kryoQVc7Mfx+gTyfan5reaHNLgxV2SLM+uqJJ3I9KScbFoVj4
9CR86ndLkXZ84xJihnw57lSpP8TEpaMtheaAn8pwVFSP3IDp7TqFoKu2K0GtG5XR
OaqrU40DQ99WhtGxZoIgT98pHFurXMDevJFqK1mlITKO81AaghhFE9DWXyqyU2cK
rFwBsigz+9v8aJBGpcsDFLMGufqNaKj73SwC2pq667IxTeDYFB4nqfcp6LsBNgYf
/zzqOW8Gi1mA7YQLgkX9wRhgH9zPZG140RG9wkf8O3jSrYlfEreKBPwGCEeusQB5
wZnpmd4569Y0irs2et+3qqHr8lnGvFVe283z0EnWGILaW/XsG4jsEaeCPDjNOL3/
COGY8sfAl/fMcStH5L5IM0Aujq26NYiUoRYZ4ZQWXFO2bueKzdpykPS39mnoriz8
2OCpLuCP2Qnkve/7uqo2UVPT1toO1STuuilQHsM4ubNMaEMeNniTy4MKasJbdkee
LHUNhV1V4+mmiVw1qS8IVsZLDAxJ96uplZUUjbjMSMmDTcWn6wkUr5+iO89MLY51
SJnANS9duCFqiKt1jBXemxtK/0Orewwp8xXLV+duUFtsX/qTetBcNk3BoEZ8Z/gb
eZesu28quEB2YJ72pe7LdQ4BHGSFY14+y3CmBnkSZBOrWyTOStitp7VRqv6geJCe
MTwm0Vhy0fZ1kaGXRYozeHBXedrEY/MLSgmgLXAYum+1IR7CYq61nxAU0Bt0MDvf
TXYqPuNoWvRlSbMI4mF4HetDRv6ObPT7f6qq3YHDXz3xCaXlrJeCty4fzn9jE+nJ
guqW5dQanqQknJu/veQUicyHBQsowTvo1yiX/+52VXn3rLsBgPJfAEGAkqvboPjH
SQUkrl5fHQbd5tnDYZ/949jOH5WsT1xgKKFJAlon3LiSZY8eqaXozoOlHBSFzM+1
jKZ2fIUTPFHutkr1ted89uKOWIzSDuxtEDCYBQCVChHNzP6aoVk30lI1ttupTiDT
Zi7yluJBGkzibeoQyv+JHg/LQ1Is4u7O/RespRrrocv7RUHYizGaCKHiRWowGuEd
RMHvOswdI+zF+SXXoKM/WipGqYIE4WDG0n5NSpMq25hfZnmqaYK0ZgJ4O7zAZ7d6
7B9mfia1gQUi5k5iNJb+NSBgwALn7mUNaNDbNMh0KEyEu5AVD+W8EnX0fVXNP/qc
pi0hlpSDrFlQ0RuTEObhEinsHi5ZQ+bbHkzTwHHSqM5NYWmPWxZQW1AHngCJNE2O
/2Ei1OLc4LXS19Re03dRgsvKEVB1xzRgJlaTv8DOvxz9xkJJKlkIS/KRPModLMFg
WaCTFTS/6cvyyyuW4S870VQBOIg6Se1r8GIt8MK+1W3dmi3DUzMU0+V3udWdSxHr
57Ue2ia6TXmUdK3PCvilqrcXF9LT2nnQ8RO1j1k24XQEePwdr0N2h0LzqzTJvFyf
W1nxNomyusmsWJciJ48ucMdIfWvJfw+izb+cOn/5Pm5jUuS9hmsGmcZDZ/xTrvxs
CtR5m3xDPrNEsc7M3OoOiL79CIZNCJkEriPR2vxphCGu/JEdICQ4P0bAr72tebG1
d+fb1LH5oICOBHEA0NRL9zNkvEjiQnNILkpHyah8+wlM8pPoPmRvsEjnhdn8WAQe
OnUQoDlKhi3TlB/6Bvv9uR1WqPjFjc9FS8Yk73UNNPUgt3eXCpBdAeeMfgT1TZVC
PZjX99ZLHU2NrCYQ3kYaoWJUlus+luG5/qfyddUuIkqkPaMPvw8FZgBN2SfVN6c4
3SZ5u8q+5n7rvujwMl5znytF0M+UlhPPHxh7KBtquaU1CZp6eQ93W0tmjpjaPf8y
iEZ9C5Innl2Yo7QM0Ggs6tTFszS4C+u0VlimCYtOZo2+BedFjDxOO/nW8qHyA1Hn
4VIXxElO2H/Jbxs9g+4QAZ7dBz6yyJXXFgFGOxvwK6mmBmf5UXFxz9sQU9z7AffC
HzFY1U+Fltnz0DoVT+9dIFqYqIIozR9ODUvNyc8P1p/bhurRCO1eWm2M/tDG5gk8
F5UTKGBCI1wp9EcDTL0YJ/AZEtAo74d5kaWvVVTksH9g0BzZr74HPridz3b600eC
3mqi7Iiewhu++A0QpuSMQeNxEQ+OYq1XRCoese0fZNFsz2nyaMa6bo2LFO9037vr
U+gjyJpYxf+mNiofc12mL6fv4Z5agPa5mzq5q76N47NMaKCORVC6I5nj9D/YqhsB
H+LGOckqk1qZrSlyZidLArnWrXL5tHRe0sYWgYSWM4n/hWoZz0mHKmS21VQuKdKH
sAyKGx6JHJwQsgtsQvvhfC/svCl72hcszbeH5T7KjNb88po8+B/NK0Nl14FbZfDB
3wv74/5uH0L1gltNQP9r0zzUYw3vqyR6EckrrDFyIN5kfRY4fRfRxg6TVap5VuAn
sbHzYO7+I0WMQwIY56e7+ALxfsXtLUq1xJk7f1y7FUdxK5lgUahlBRxa3tP9CI8g
OP2rjw13WXxXqgdzLKzdDS/qEBASCo0XyrfU0cU8vndfS8nmq2686EFlAOXSFr3S
NLW60TqNi/bUXVemnzbI3pONI/b9G4cfRV1MAgd9ZosZ0kuzrvR0TNzHf29W6CZg
ppuqiwqbdFdpe9rYyUiERcJ8dh8TUuntRzWX4jnn+C6UbUDNNaDhX9YyP6UVHBXg
grquuISKnFbXhrNYI0hEwXY8L55FAv8aMUnuibPum4XnCwPfjdod1UQADeRbao3d
BpWRlFVmKZ2Yg5j7LbNJEjSfCGjOgFNEnxqiAv21AADC6krxYwyXXJmGvPvK5TuE
cjwql3AcFSNZOuoJ15KtRQNr3XrmCdPsZ3InI5+llWIRigR3tecB6EVn9SBz/RfD
fngNFI+GrLRQ2Eq9zxupOmUnlTT6Hc9ZXzUf/idXNw/Nvdmdmm/bmKSWyIouKlEL
32cl+/XPEZGS/e2UpS27QRXHccE4TAFIPWNMFEQqfXYKFktqicQXrOenH4/KQoFc
SXfee+7VNYwSmNF7QSsiiDXBeakoj+TFswCkkjJG82Hq8Z60WbtS1CpFx2D+sgeC
U/iS5H3vp/IZp9tTWYZ3rUJ2H7mEKK4NjdEskZ93SVO4Mjv3X4x4q1IK62Msgi6p
pUbaRSAYaI6TzGI1o70pJ68lthsy3MGmPKMcN6nh4MTabAbF91Yzr8y0ww7Sod/s
FbXsZlO3dmeXGjGYZAfEW7OxpeOAGre/wTRXZ3eUQYBIWGYd4YcEdyGfwzsbcKoq
Ciln4i3xdKaDASClLdLuXm3ck+Tmt82rPQE4yrHQrx4s6f2i2YJgnO5oMvNskTms
M+JBD7N4BGM2vBPhamx+fFIVtaJFx6L6H3EAqa6JNFHe6ZID5u5N7V9g6anS2HL5
+qOekxAMs6aWBePnSN1M4BqFonyqoOLTkhffFKUy/Zsw9TbzudpSuwspaxM3DoQ3
B6SNLIAGUJ1Dq21jej4PQ0TyDHmazna9lVHg3iNpeuBMhuvY3pW+XbU9cJ0lwebv
5my7s5Hm3IBeo8FwUV/obja0VB8BFFkuAq9p3NANn7nUjBKNY3FUm+O3Co9nSIot
nZWi2E05WWyDGmHc+cRwC6quRBfp5bARXIAkp0K8NC9OEyIw6FTQx+3h1Jp4WMvG
Y+LPYOXtoYM+ph6nqXqadrWKWF5/GoQXo0CQOrHfEaFpJC1EAT+hRGKgn4ioJb56
8CNVNjb31tTHLY/pi8D3oii/+Bg6S9TsOoxYAuGQJdPf8i2NHKu/H2hpinMlhkK8
W5OwVXBp2VcnnnfCKbFkDxabC6HfzZin8YXYkRV395Xn1XRCo6/xu5H+EacmHqPB
aILlPRsBbPbLcYA0njRjosSqqavaw5zoVJYWwnrzx+U4QzXZ8x4WiFZaBsy2SDTJ
8K9SmCLgtvkGtZYgKgCayM2VkQbwK7ehwg67460sRO1JMqORe6SU0sTi4MRPeXKY
bBK99e783cN/AgtPHfUBUCNqeZ7BHkoVhrdT/MrijrikNH/oZhCWz8FwmlSPzmBY
EY868Ezs5/jyNwkyub6H7+gGGetUgHMFjt/yzAOidNlozI3+Qp7r1KHWpf24nAY5
gnFE0fUvYfm2guEk8mxWNLcxXit9vrnA2gBFCkDJhelh048HThFRJXNGrI5YgONw
1VavI1LzWqPVBl7aYu74S/KzrRMPwvikIqtRPViWNiCc3e0+/r93tITUdv+/iZ3i
rwtcAvISKWGRIeMvbgnXYlBw3VAyfO7J6B57QT9bq30J6pcSXJ+gswbVWk/ZTp6M
K3ggsIBAd3Z19zedozcpDPns8DK81GOAGgi52utb10MeS4Z4UxqGZGrRvj0OCZ0D
8TrWEckZym4wssukbQ3XBHloyQgeCVCayGCtDT9l8wjCMtPmIF0QGL0Nl0YGKNQ5
UzqPQQvfggl0z2plibkD/Jtm43wxqfjjRzZj0/c576ya/CuY3524QwFs56Wbt5qB
VGsof0enGaIc+oWvRfoXr4lZ01Zy4BwGx8W+vtaITwllqnL+SNbzgMZafIT6JPtz
40J5XYXYkUvyvYcfj+5OZUhjgcXPv+QQ+rKBSjGpVjz46byYk0u1Y90/EKP9t/w+
`protect end_protected