`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
ddtXksX2+yylW5zu6QL2Lhnb2d1sD00763mmSITNX595NcHTEkwn0zB1Dry37fOW
FufOhVzEJp80NC5qZ/+F0Vk7Ik02dIR0elf3clrjeJRK85K4e3Hoo4xn7YbFUIms
l/8VZSb14+JVGURjfswrIyCUotIzlzVYZ6gzoZwDXIi5gQIBf/gI+KxNXPaKV+PQ
Ufys/12rjO6aI/pPlqSm0hCvftmBcnezN2hk1UeXgOIuKZnogjOsf0iJVX2aOOWE
6pD/psybjbnsNB6kH5uFTA5frkzIzkzl5d9+YDm9OyC+k84E83I/7/j+rk4L2dah
QJOvksSIzN867/4Qt8qYTQ==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="MvBXkzurAa5VTw+1JJ70nePUfoQXBvZOku/SMmg4TwQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
oRtzZL4VJ4iwysPsC8SXYCzXS8Fw2gtZTOskLcDV+1B9Nzn1zTyNtlo6lNICRmmK
ZRVu2BmCc2G+fmzynYlNTnSa7C0Cuel6FYpxCBlOuk3OF2tzAmLAuDyOH3Z1Yjzk
a0aHuoCdIRKv7BrZCdALt03JeUmXKPdOmIlkVGFl8yw=
`protect rights_digest_method = "sha256"
`protect end_toolblock="Jn9CQpRhJt4rnzZPRk+dOpzAubz7omckX1MrFd4p81o="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 20416 )
`protect data_block
gD6l00tciPUa6pDNTk/+t0OO0nC/UTtBwLB41d4inuAUA3i/ALrNyoJVcBnAmEQW
ptbcNp5fxEUJjnOxnedyZEuEBxWRieZFQnkRdF269oN0lnKwzPyL7wDtCUIDMRLB
IaG7tV1ZbGuabQfot3zIsvRbbhJnBIB0Rmms6up9kjawyojpxEoHIq/ROpICPwUT
CSNTtM6k8J6cTxcwWqk3QM9pWZIOmkv3L7CDgiddTFi3uaImA4ZbLSpbuUkyjtZS
gr3Ya0kGUtT7QakHfEOtBpB/ouopISOfx9p+lATF4AHjtWQBAy4LlRuCk9TySsD3
XTOU3bp5TJMFH6Bp14MgXEvx46ns/gcmbWb5rlxVxlLwIOU9cpBkaLZAao2ieeaW
Jbjr8vcvfiadNy0q9f13J/VUjUTSnk8FMNnIO++ZGw0D985rqY5qVX9Q1XUxWgDf
UnaPe+0CCCNZCjobC0g8uFLIacnBN8I6AODXn+GI1/qmvhGPy3BsGDhztulYFN45
HT0OmuJYAbLPfp8oijJKxO+iP4ArXMGXbBoIoBlUvN8R+/RgDtmqxYKlOg89lbjL
cmnA9ljolRD7C9OFzsKtRzUKlX42Ao+NOpdWUsUONVVSrkPaUh/bC7/09M1Q7DUC
eMQeEZ5qNnlFNef+y5Abp9Iqhr4UgO7P2gGhr6B5UTHcN6A2onlBC0vPqdJYgC/K
K89s/tv8ZCCWCnxRKdjjK1WZXVtKd40zBJL8ctr2iZ1LdyP/X3wuWJBzoEJuH56C
Fbi5c63x20nlYjwITcLr/aRCyinzU2GZfleBFcg86/u4Je42Pg77NG1MxesP3muC
skfk/dg8SmWCZfxMIJUvENyLQKxYsuiHiQvAFF7ztq7Wq/vsXCqlXnqrZo+cfgfi
Jxe2R08BJdu4Kkkyoe1vf8+xEPHAQlN4h+9UY1lwflms4S8YqsrPVkQkEyhScJ3Q
gHH9cMUGNXnI+q5F9UD9KwEjyTx+N2TnhQBYU9TuuUpaLc7XU5eP6hJjg/nRGObB
lo5nExPLXSX/0iVGv6209DP0ltrccmL5Bebyo84RWfQLDfrZpHQ0r6xt/iuyYmig
ZolWXsd0uZMflsFp9qcQ7wLST+s06qrr+uOiqKOAqc9IQkBPlJ6IvotTkfdd6LKW
gR4EsoNxeauWmT/uV0YK3U/0n1kHL7nMNE3HL0Ck2iVHcfFvW1SNEyf5OSo5ijIM
509N1fDJumHRDqEYIEa/6ghi4W+fAQ+l+cZz51RBXnbx4ePFwYFjP1d3R+nL2SYB
hjleEIVhzOekXMTV0rA+EaM/3iE1oejidmzntky/F3ksl1o5894WVYvVnNSNMyk8
x78Vn0qi1oYlRVYkB2OzBCqRxwjKIjeo1eFNkst5USVV+NWTTvgsxeJ8ymOA/TS9
4MJ0xwamuBEOjiagDq2UBrcB0Y7iCCoKBeu1mO1pNTblIf5K/kNyJYJF+aqTnAM9
j2mxecoflJBg1DLmVA9+N0HSRFxYssrq8wViLomFEdIlvF+t8fXZ0zKyEPDI+fIl
gGyHL5VvV6di2kK3w7Fya366FYEUWeIRRZ3R0ZHkQs9inslLfRM4LQ+qiWGaii4r
IhXgWVDiNGBKJnJrkV+hy2U/FSO3sh/glSlF7Y95PriNa0/5JK1aPg0EJ76PJX0j
i/yhBXFCl22ciltu5HpMuzitjChb5Onv9AQi5TJaexovb2CZoN5Xnyuo83Qjnrom
CZHymwjbvnKyNIiF4M0qBteFSxBRa/0nCbugv/wB+ToVpCFM7D8MohldLdnvEQXe
2kiWka9bv7TqtYRakK7cdfiq8fq0lN8qzlOXp5ffHYVNhct+fgL0mPb8CsWacHxU
hcocQ1d6yT+a+oFf2OZG9B4t7raH5ma09obu2a+5ZfrC3MVEQhtJlfulkngOjsWx
jUrpLq0py0CPuDPp44VXgNK42UbZpQ3Dpsifl36b40/MtNOaFm+fvDRDrONQuW87
YOo+QBAK5trDXK9o8rDX/ZC0yYQ50KXiLrQXl5R2mU/A2LUJCBM5vnVyuJg0nC1S
AMqZ96t7cIJFGe7s8SNwtMLLbKEinw6Wz/L8pM7Vf9NLfm8iTAH6C/NQHJSzMpY9
CBkT7WyyHTljLdCcehdTU7qUpZX8KeoYiwazGgyylzkiG+LqD9g7Im7cxAIsR5br
3xyF1UN0rUjBy2mLxxqnHvWX49V7zxufOkUMkU5MquIoMZu7vuYAdCPU+BPYi2eD
MTnWhud3WYiGOAmlqDntX8Tc3mNztNPS5Us6cB8SFMK2jncJfSgSKLlNVriTpiUl
NqjFQSzcbuzuk8yLNDygM8JkjWKewbICm3Jq5WEBrOYaeEj2pzhHazaEWmNwMfXP
xwjj5Oxu1DU022fSHyuqBI2fNWaH7Y2b5qJRJcw5P7R3g4Xhg0Z+pN1Ug3Fbdzn/
6WOclMJYLIr5elUB8bMM6fyFv4ZmvNvXXDJNs+ip44qIs8/ndg/diZUeX4yT4IQx
NeSmHu+FPIXtGrIFHKImu4Y5FYAOqjyS+3CQzGxEajpqgwAOjTqXQ8o8lSRLCKgc
Sk/2kqBZzYDlQ21JU/5/O7PSoCTPid5A5WbgzVpGk8fRK05g5zOKcV14DDeH7zze
eBtT+E5ODzUNFk55zSBWUklFnZctwis+mVaRzIAsPd4aMcZuJpgmIvsdqtY6/xx2
8C1UvhHTwRW4fNLPie7lC74ryAGhL+AkCtEiKobF+R+41AkMUbWLPf1s6c1rFGlZ
oytfWPQjVXJueoMcXynSIMP16BIZUSW0BrTHaoK/8W2jb9pmswjbEI4a74jK97MR
CnZMKYYfJ0XF8r3IiwKPk/U2m6dpOkhw0/CV/hdKORBEDG6UglcgTh6eBZxU8F5E
w8PUrxAf/ktRKKGIZR5RUoXeUzLdY6b/1sL4TxQq2rMjO41wkbOYNnXaWxRiZ31d
hfSl2iatKBQj57NJkzyj5MRRCjWcLFWx8LAz9fMef5B5a2m5NrtpotZrGSbNnpsw
SFK84Coh0qZHj2USSfztHnklZ18aOAMAgwHG2tlQbzUb7fbrs8m+Df/GAHI/oDdv
5wqs9Whv2W4ZSPs106+sjAKeiPYSMdvOjw92Qu6hAhPxGFJaiHzYQeiu6ff4T2Ij
gf5gNOGiP1UEfniklgo7irVjxnkp1DOokRtWwzGaRN0ffOGhC7L9zRm8EgjeWojv
qnmC64NpC52/4JvoeAbSKwPvNSdYmc/VYH7PDoTNnemAyhwRL816SaS2VWPqqX7o
48/YEz3LOCINZY7SeueRYH8W5TtK3uhKWXleS3FYLZ3rlKFP/ZKhUJXXXsPdN0O6
nATxB16ghumxJX7z4MJIqHPmQjvLArcHqshYsvJBHLdLo7dTQD0l9Shes3JUr2PC
0+3F6FQWbBP7c+VLF47+9Cb3Uc1hn87V9VyeZQ56lEQdCn+3Gzy9kqUgJd6rYNNR
QukAGzytiWcGe+/WCg/DVfRBOo+EM5CSHd0Z57IYuNAWX1PqGlA3RD2E6azGq9Ko
MJBLeCcSFTUEbCDt2BKBqx49SPHfl20lvZedR21OfKbsWAJNPVRnD0UKQ+efcFbB
Fe+RQ9ErCMV5xCC+azQlr0Xid4YW6HIGB4BY/FdTNTTWK/0poYGoqkpnsP5Xo5ZF
kGI6L+sHx4/qhhm/N4RpNB5cBs43bOQAP8wPJv2tmcEGoDseGqeaQ9tVs7ALGP23
VakGVDpLokXwUBSuSrFsf1wkNG9RBMSbBa2tRiQZp9MQbRe2ryzcDSfJu95AwqDc
utm2IpPnuyKXhaX5qrN3zJh+SHfMU7dj9eUc2ixyzrxL9Mpl1ZslHQsJLAYNX5iL
/XyHiEvDSwylvzEy3nyEJNx1wR4USFUW86EgxAkGKYSKjHH0BEbiCcXbq7S1LvKY
1t+Zbru1F4Q6yvO3KALNViPaTrCQdN0z6H0EOIQGmwIjUxw0L7rRunN3gmGoaqZR
PBbcDyovfLsTnmwNt/sNrAm5DKVyTTOI1DJDQXHYUTVE0H/p3+yBjj8W7qIKQB3C
J2siN3oO5UeGZi/uUlIomRFOx0Td9XvkIjVFK4Wirbsy5K9UwuBTZ7Y6bkOxCaFs
jyh7/GKEIGSpjfIp/0bK8RZDCrcuyfrtytOxiDjenZ/A10ROeuH/NEdVxwy6MRI+
3FfE96BhRNZ4FUkJrfGhTz7vynnnqvlty3ReiC+/O7tnlWrDvYfzpc+pVeqgePdj
XYV7Lhq3bVsgehlWHPSJlMGA9zecyiEtSyjXxcbHci0KhnTXnHlnZpwrCFHjAbx2
5dTdIym3ydcguIEv3nGJJ/VpTw56b1Yz8JfITOuIQgEIpRVwMZnf6Q3qSgXReQFj
OIC0Bu+5C5wFN3MV+hmIs1H9TS2XJCZPT8uCZDHb/BY2PwMGBzbHLA9v1YW/+Iiy
jtawDCxrMPNm1JAjSb6wnXZLxNqn/YSriyZvfFcqrsgKhWbpLLz17Qqe4OZAcAb9
y/nlmQUYO3PWXMIwuFBLcPLvVrHBpFYefspuILa1/yrG9KK4FCfTCjrGbEEMiNSG
u0Csl9RcLjPk5vfLRdNPMZ+DA1gBjhAwpUDEk0iEX7fJkiMvs0dcDgwx0lknmG25
QZBSP/7f31RJf3NVHW5YNSQeBlzJ7xo29N69Ooe3GB/OA9Qm4wJw9n+K4NYTFCIz
Jn4JlfKvYetclTkhCBPcxl2HtsYqGQjqB4S1pPLglBsqzXW//qSUnHOI/OeU3wN7
rk5I9TT8xoJ2Agfxf6N0tx4LjnrAKw1+z8gajHFnBlXefsPT183fKqp09xKZzCgb
a7xYxOc3rgHd4nIZ6yeD+uDicZNzPdAYvnsc2hybwJBN1HNTb4FBy853oYSN7yNO
Pff0yCoIRfRy2aWO84jiGJHhXxqB1zezv9XFhoMG+mi4XnVT2xgt7+vvDvpYnwT1
aKkSKm1z+OvfguPbs+1Tlu3rqsU++L4IFyEmgz+PuhUu7qpX4rLIX/XvMf0Tt+xm
bYpuPA/YQrk0NZ0kp7ymx9f3Z4Qcjndt+57yL4cATp5/3TpSndAJyNa+5yur53dl
KM04yMbEh8eC40c+yx3J9WrL9cOHZvFIrqEQnNe7q1ZdTZ8mXUKQxRj3gYq4g311
+bYgsF/GHeCzY6hLUqCJyqv0285kNa0fc1NtjaqFRjLzyEmw9cXFY2TftIelFL5p
/y898jka9HvA0YoEwRK2uKq9ab/KHPP0d+8THP/et/iMidwUju0wVrZb+Fp4DXJI
TA87Nr/x9cFNEm3LH/nlsdDQk5ocvsu0CBdTAt+zW1IU4MjcDzUCWRjj7oqwARub
qZ+hSSy6Z/w+qP/vwNA8DYmlgL8aUmZfBh1/VzpSH++s3PsszTJbN8DN3r+VIobO
pHlv5MxKPR4CJzgX8ZCX7kd5jsPy2MjMCuqAJcW13gnicl1uomhXSlucGRGtPMCA
VfDFaqqcd5bZ0ZRKgmubvCTwTKlxQA3pbIftRcsZg8hIh0w5cUx2N32UnXe8hhyL
nzd3VH0FPJWlHOA2MOWvQJ6QtYBUA/vI1bojPgHNz3VvxS0U/U/XWASKpzJFop1+
wdH0PEow8Gp6Zo4ooW39pkEAm3TnXoPaqvwJmwQofzds+yjcFniOU6Ll0FDIZzym
AkGnX8L4N2tPN/mN1M13Qwiqb4OX58cxW8axjXf9XE+OC5EMBuodECNOV2/IvSM5
PlnnTHmoZ+Qubcgh7zW3Kc9f0CrQJGr+L9PKIfOa+nwHBZ1AhG31X+CsluIvFnNx
qiQ0BpYVRa/binQIy4qDTYpq0yl05y1uNV10kLw6EiasNNuPFLsQyWqIdiKZ4zuR
eCP/3YdMaxKAsZlEZnCFQpq1wh0E3nrNZL1rddEnnq8NfeQ7hZEzwKtQvM+MYlhT
0HfmMMwdiYMSIpoOLGqhZIxpATFgkBX7z4nZpL1uyEElvVfmjPFpnXrd4DY7HcvA
Hhfv8gvGLVCZsOdwpDlyycPlWLqWGZmDNX9+kGzWWfy3z/2LRIhnYcm2M4HIZlc5
Dhp1GjsYa1v79jbIpEiadIICP1hoNhVDr0hsZ/ixatkEhXrRNfAVSZDg5+6Jv8+2
JcpsKBLi5TDyeXsppIZMEaO6xt43Gal2dCZhTXITlRFK2UOvRqyvzbLPCLoAMYDV
/lWhMjuFjsE1xGY7MpVfPkwbJDJj8lhmU2PDm/ttnzXSMGErtt+06uzB/cU8LnR5
dhE6PUYgLMuIR4Z/NMV6MKTqmzFqLd41C1QDQ1YBVb2/FeyoHuyn58wCQJscefw8
upo2o7WmJmx9L19q53asPczMnzrihO6PEH2pmtZMjmiSwIBdB7W+AKmt3qLlBjYB
m5iEWelbaRcTJHnTrfuSEBI+2a+M11v4fNIcTPSh2CpD89CXVei3LGfIH0fxxMXt
bgIK0xjvnU5uFWrNXY82PiVhAMotu0/jA++eHOjmc1jYSrGRAvryIftQqra9aNhi
fFNnRcFUDRrxkpqS/JO6/mhscRz8SPZF80SV2gOU8gRdgSjPetWDUiBy3sJxf8pX
HjrWPpsxOOcIekYCC1NmyMjCqzOn8Q/CgFzsW9Zd/wScLhIr6VfME66GjyrZqko3
LL0brOddLKX5jbmshVqyiMvZ82rqaJjVB/k/11z62wFgrF/q//vT5yScYPaAr8UP
+puk8a5yaMdoZcNtWQBp7Vdn2hDSPRr8gUQRxR0QZt3F9Z4e5rovknuf8buqogyq
9tae5LM2LY3+JrHO0p0nlaq0uYQJysWZZ7fpwvVnl4KdSABCesPAxkkDHFDQa3bX
o/wNee9pF9QIpe3BQDf6Shni/PwrGVJFinG/nKj54hOmXd1JHVyW2YQJlMN4LLxe
uPX6zZGBn3LavUsulhJgLYg6NGFvZu8+ZGBkqaPun8TT6JytV/63wlN//iGmhTSZ
M6gmtCp2xt0+LfXRZyjueJPlK+H0q2p2aMjiGKdHNjXVJ9j0U3x/jBJddC87CQMP
CqpVXSKZoKTGC/Uir5I+XiZxCeBKOnxFXwzzM9rglZswjPGDORSiAYIAwe+dabba
beXfCWGnyaMeRlB+Q8RRlNARTbfV3OzcRE6SETDvrF4lVOO0SUrkP/lTx26CWIjP
I3cq9diq4d6mGxDWbHWOm4tezWjIAJGIz3qgdteWFOnTQfW6q0wvMPlF9rzLrNAo
VCf/qEeIxblstYqL5uJWQt5Pdp0i8j2Ov42btmmh9Hub+eiE+iKY4UBAl8s4cq/G
52gURIkkx1NMJ8BggIcdc0ILoniBedMCJr0DguwgkLhC004DrC65BhbYMLVjuz5x
D5yztoe62eKZyhU6gv2v1vSuuNU5pT2PD8N9d56XY3PancWf6me8f3qOFQm0Pe56
/8nVhz3/ccQ9f8XuRJiHgsfjOzJJkmi02TPFwYcTFkbwdOt9NGVy5zA/FxxVAOyI
KiRtwW0ItR7SIGZnX7sBHfZz1Zdl0kzCJ6PAsQJJg5pM4GbDWxWgbiJHVpTg0YK4
6FmwIRcnOy9HAURhbFImBWyo/d0p3jjqCVwKKtO6VDoKzum0wATC4/5fOWNS4URW
vyj4GSHBF2aKtXigS2BzfUTnNITOsStnmLYYijCKjwCZtWU05d79KUzGcpeB0pnl
9Nsrupy4FXQ0Wi+YEUXKm9usAnJcEffH0/Tc7jDeAb4QKrqsGuwHWYGKZpp3zkWw
NYfWAsz0wOc+JqhhDyqq288Wom2+IesXLLnSMmV2ka0kUB/7SBIx2DkZPllsNem5
U5O6KykPcPOHt1m54l/rmcHXG51EKEXzVmyVOeiiLez0I5t7goF8AMhFPLXdVaNC
IuYDH54ThdzZb/kPbqpxeipFNgauuUwROy88ennnsOrU4WGecum7gxKFFvLqYy1N
OQhftzyv/Ez5v5yih9Hcmy2j/Dx0gnjmDhNx7lCb8FOILuSwkgBY8Cg83VAhjDJn
WFQIc74TCWf6GadmRhXgW+y/nkbeh+xlQdqayD0zqKBbYXM1dOgfZuRnaNhyt08D
bSoMi8pRl8k3my5TXtfLQx7KVH7frPtTqgEI3CzUG6x7BPq/1EEqWFuBVu9FQrup
EFwJgPL24zj3cKshAqfzCvofM+i6gSeHFeL4Rf8GVImpOVWYhk+Ia66/UrVhBPxP
9fUaAzji5SqumW9rphvmKBDJ13o6rS5IVP0AdciAPr6snEWHYrV+1F/uwQ+SCtKc
AMVs2wuVRTdQG4pzXn9kFro6fY5Yg8OmA6cBEPZ9pBVBbF4dvx9IO381VM59o+Vy
fPhrf8ycl2+I3u21Sp0BEhUCSaUDVNuLrSJZipIVSUUrEEjKK0M3b/3EplIJOQ9c
oUbcwXU4N3Nz+gvsjqghbclpKBtkBpzhf0sv7u/9keeldjrv5N83fC+k/+uwC3ei
DfaOT+kB+sFb2dziG2zV94mT65VMbU8NtgKQD9CEb0ePH2DtBAQBSwdWB+Fcafwu
o2Akzd2Ak4P48P1Q5H08WAlgMZttVh5uQXbFCzmgQakHoWlGzTyJYTojKLPEJKdi
W9V8B7kRLrXhsAUlhWBuOxfYXPWi0GC2dioxe4RIDrUOFcgxMsQiu3MuuaxODEUJ
k8qDrPH5QFttYhDdpRHkPWpWlOVvyJn23u7guYbIGvWck8SjgghtJTRep6XoLzh2
Yryzk9BUSH/V+5f5Pid8yBlnqGT6XB8StNeag+wT49YTymaiVRN7r2NNLlVpjOOh
Z2e0RT2upj0xWjAQzHjObn497hkPUMOcy+6fWTXploMbBMyfs3hw5f4wCeAM7UP5
QXkOO3GnYvvI0WlpHwiYx2Ilw885TcGet5lF9ZgFZKPn8/61B7gV530Wbz00ELAJ
LbKzaelJJALd3yEYNSl0Yt9TtBWy4+mP0ztQTLXnC2rH4CaXoC4EF4gW3E2OhamS
ZwG8d0QSfBvQvLQ/rIdXwByNMnH6D2k802m2anc+0DJ5fPZw42Fze2pUsZ5y8ld0
bvoNYVfOYdzZyLPwN7PCGv+Cbgxiky+1PZHG6g83hKiIjKXtLahEQFpwDdipxE8w
Dk3klOZZywypmqHyS8qIHWqhnZUBybliiYxiO6RC19nfrHVvpQmlWyeVboPQC77J
0OOjU6asFlZ+gxvWwtGSka04UKhyUBbW3JfAybucWZ6rIg9TAuqx6sx0fyr9ndiJ
H+ZGuJE8VJ6t544Wz+kvNL9pe8/RCGm6n3bkKcjSsqS8/y1NtY1eeZjvfflYybfA
OHsEDgmXxx6h2CrTIDX9PGZvtViEqXjNyAKNVylEmzUEERKbSmINuHhKY3KCcDzV
OjzwJkBZKGP4Uwcfox0Ra/PwgIm9MmmNbVORdQhYWAhWEpjF41fuYjNk7nZnr8WF
U1Cd6JVLlg1yDHzG3IXOhghiGlwgQCiimdMMR1ZECCWzEg4mBqula7KIxb3nzhO/
QQu76L18SMdsUD4zpSRKPGENQQ0rsw+45KD5r33a7wIDN7vo7GLmsrFWIIC/fjV0
jF92LGKVTPbXRtLdEOyi5xLewUjNH4r2SjZFH2ZaycJwMaN9QcAf9AbqSSFRC3Mr
cPBSm5Lh28hsaNQABUOdy0ChmtlJRFusO+DUXVEbVhtUa8f/PkZ5duPXW6MQVhJD
VnMEXicFSiwHJbBIX6wzoqbs3gG2ZKQ9MqIY5xUMDMnyhdnkiJsqzCC7R+gdxFtT
DYwjz2pLJk2TQH/djfykQ6zc1C9BBTbceBaS0sgXju2qMZqPJErhUlcWyYO5IkKH
Cw1BkpEPS0nWgCt+c+PiLI7YhvBWVqygrHu166dQueSx3NCPvpSBLGCYq+7B4/9W
80UEangAaKPZBApYWBuNel95NAdrwxwNhR9t6B9TTAxMB0inQ9rHU7HITbt1Re0E
NA3eqlglnUqcyCsOdJHJci23fGaCPiaaCih/GjrI5/6ORVcz2FtsIi7j7uYjhrbB
Pu53FWEBB/az8IoDHRpUhoR5QadGoVcVC3g1uNtv5DcLtzv8ZIB85gH3LQ8gKy2u
YUIZO+Abw6fXZ0aCsrTKZNOe7lCtczfCQYnBnY1dEt3tjumgkZDTuuBQ/Rjg2/g8
VHZOHLMnz6VqsZ+2MHA0NgRiaqYoUHkVxcHNic6synIDpBWK/ksklheSjf61fKPl
+DKT273/CV4BEnf0EPnnAdL04Hdcnt1/HoaZO5jhI5rbHYuPQTzXHotUT+b5x6Xg
zvuKrxR3Ca/NNvDICH81oNiUpdxuVuSV5+9Qcp9SkdAV0ruz7WlHYTM3oNVxvvb0
Sm3pikG684qZiaWEuKb8plyDcVQkVsPSi0U9tRtvtaZrMuXl2CEH7SV/7DVchuk3
wI13EZbiKSLpkCRGJe6LXIvVjOez4Sr+d97G543Wc4LTnjxLN8X9XniZcLLalSzp
XNQNgtIHA2bUv+l02JFiuUv877Ysm7+DR4j2ZtNQ+BUfSU4z4bKHdwcbhlEvZQdV
eghH4CTCEbjZwROQDUGFqVREsk1dcRHdzKoqbGOsPm8uxEGYP33a8ibN8sUGtTTD
2kwBJpfO7eefOZyHEE1pPnjj1h3E8vAcojBTVhdnv4r5IPghsBHBZmuf36sCHPUw
CVnLmEe1ZdcSRtJPN2MVd/2Q50lvw0ZIW+SEx1KrtozJc/tE+X/4tjGkrE9GNitN
ogFbMoDBKR9v80eRslGPIlGRwfAND6+skz0uphvR2KTTLhz+FQUFTf2KjEDcSP0R
07X2R5QrTTjX5EDgz3uVvR43u4pDKbb1y1tGPqKJDh5OvbfQmuphBWCLmaY5n8M5
/iBPFuZRD/f1w2CsxWJu6bnL+0y3O/NM6A3T5xD31CabckgI/RxeUaKKath1DCw3
RyBNT7HL74/z9cvnWUi02/mvJzyxTzPOpifxnolRqWIIuchM70KWeZhkPf91SgoH
gl1Iuh2pZrDxHLyGqs7y7Nw0jrj07yE99iX8e/pyRYKCAVetUQLh0jgBHrtMJpIu
w9a4x5YxssPqyLM8rUniyYPObZnqYctSxj1qtYSXOzC+61K2wTNr5iX+a1M3cCz1
6KYksBc3KY53/NgiInHrpI1D/AXBA9EwVh4AfU8ScJZhaleJ945fYZvh8yzPctNe
yQcFwLoCoxt9rNv+8g+vE3faEM4Sw/y5nGgjCJ51nR97fu/vh5dqiKlKoN6SQwvZ
zdJZUx8K7fM2KbRvRKP3JSgs6wS0SCLWWT6wEsaBMS24lyYH7LH+2MJPV8IBQVzj
Hp+MUHXa81o89yWS6HApkrFi0ija1+9Wjl939sf6XGcjjrx1Yu04dpfuo0NWAQG1
nEWgfzdrLCca9GpNFyO3K8yXkvjsPHzLneBv8DGPagpUQUQmX9QdIY2LUvq980Bl
O1B54S3eze/GUGlGRjLwKIc08TwP4aDb9Yb2AUERSUH6GMHIhHSXzeyLQIMPkehl
CcFII2Wi9yurgCMEJcMzwG3Tbrlvszl7Zqy4zZlUxO1x0rntaszESnK6dd5yN8qo
i9YgqcuTH1M71SCaRqFk8Bfdr0vIS1JvAI+uGGchtd6sR3pA25r3hsw0deNgA6Om
HTAVkxFYVuJCZYn3aVy7tRANsC7n2Cq0y/q/sAoZeuRLkCb/d0ciELYXu01zyDWP
f+6SAmzDANtetEx8/0ZbxxvJk/fQWWmUZOkAE+Hw431SeFKVMqp5JxCOIdd9pedn
FdDUb2yFH8SfPhNvz3A4YYvBQuGzUrIYTYIsl8FagKy31agjSL4e3Mc+LEgXpHeT
XxcTHm8O19j584x1rclKQrNHkyzeKIvkjJwpnEr1TFldMdGJAXOZ6aLc+IKLUFmc
CEDuS56473tUKuL4OFhFooRRRLu4zK1apVQbmwmcf/XHirSR1vZegkfvDXjaNFiM
UrdU18MXg6uO2Ru+meDSyTn971ipzLR/GFOwzRPqVZ1Vtvti3/BpH3dYU3EIcqtV
IewjKHL4L5IgOYt9mxI3S89csfOkKJiiERolsaHf89QV8PGIYd4cFoXuN3I9HG2A
qqVFuSQtYu+DZHaipi9wZX0xergeMrgA8a1HOQrmfOZ6KOwbHv9gH6Oe28qQOr9O
n7p58XX7CxrTGVaLNwASvngMewFEEncLE0359QK3ocQivfgmh6N3SGnwxlLUX5v3
FWY9EilBEiAHvac80VwAp20+x97GU7MBWsv0zILQgRZRfewQnPwBUNLsvA+VVf5p
Dn/7v1vaRM1At9fBHEda2BjHCsx84Vme1mDGnxSTiUCUSD4EISOqaQjyTba3rx/q
pAI8i29cuOfcFVBFnIJgPPSj0Sykbz7VqJ/3+fK9jSJdPr+CIvIPnSdXINUGTQn+
ZAlhkz5gI2On9JkQO8XSFfkbu+QbALD49Lg+eWSEIP6Qhl+pqh4fjSTRtfqW7j73
D064tOXWg429jL5MPjGTSQiz8zF4nGvLx52DbGXnA22l7iDoFj48ntnxpSlUCd95
whwcGhYHeE96MLWYfA0kA4QsfAt9w8mybtHvBk20e6kpAC+8XRXdpFg61+W5rjDr
XWlqOqh8rv5KrNmLxRepdXluEMwY6+lhyjTneExJao3or07tkxU/tqhEObSXzZYY
1AvzkndLsoo3Xm3Q90KKlANO1xOEMIRveArGxoG3FItEODhKY4Clt2lM6eVsIni5
/J5FIB+aOD8Rk6qIYHPHAdmPOJK4ycX0tpPjY4Ggh9/uox+1eqtFqnwBCygvB4qS
4AvYI6OWH9ZPsxmwwxTOcqOILS2bPS3HWTr6GsECwnQUFWPkvQveLm0h6Jb0PQic
g6np6+k62BCHemrfwJMdqNknEFQge7orts2+CR4pbVSsFMkXkN9aJKOzZLzIoWIc
ivllk0v1ydtxTTVx6WrIRYG/zvRU2o6PtmsKmgAoe7634co9I/x6ZCHcE/DeUR0J
RIahIwdC6KWZOiZiRm/WLJkQgF02qHoCdAiEKsblONIAx9XsHenZQXLj7DQBsQvS
u0CvtRk+WYilbgfEB8q5WHBest0pRfBX/9B3aPa7jqZYbvHLjUXr8Iq1tpGCI91/
lknZwbTQktgDpQ0eN6a31Fod26O2KUuXorBda95hDzCAY9Pz8XS7tAnPPIzYsxMu
kaWdO6vp8Ctay0VhEw+rlx5q7sQOYWYjjdurOu9JmZdM6eezQiBMWqfTgppwYAjL
hlc0MZdd17tAaxvAtA5Ur6T9LbOJTRed1PpGBIQ4S2096QyMlmyx1Bq1d2eTBECz
ZFa9rDeIph15yaI+YmUmXaSf5wmGYDg4j3GDatJaYzT8EZMHac6WsmxEdmSTH4Qs
ntp5leipUz1NveD+qAp0ScvnDD8acfYSAoyftiXxEzb05tGzKG8GzhCdXagNP5JL
1HJ2RunOdLdymuYW6/vW0pHNHLQGcMvpm7x7wvF0xVStDf+6dmtfyk/m4F1PxAJ3
hZ7M+czttTarZcAA0nK0mcpRxX3B4OvbQpcflRaw0hOR4iy6VrMkaU/dzMcZyVCm
/xeoqynyfqCB2Ra0dgP9ROt769pDMUMQGen/c49LOTqX5V3UYPuc5vtks2hYxZnX
yP89R8G80hSG8+MiBjRIfEo3EJCqXLJ44eLPglK8i9OJJ22hEWWScgTGLugCgixg
V0RiY/quqhmj96s66v2o4ABOypU/D9sPqFmVLd1QcvJKbojO/oiT5X0LPrYP6VDD
cn9T0slOZSWCEkXtjPRX1RkcMnu/v1FLQxzxeF4dcRJAIH8iU1zz+hQfXMozslBX
J74bteFXmPQHYBTlbI7WhpzhBNHwuDEMKQoGMr3u3B6au8lhcelp5L97szyftSDC
gqcgN4KcLClOdf6Iz4HHf572Kj4iQo5S5bj/gDxjNB98J7R8IotuB9Wgl8oUA2Cn
f8qSm7u9ntlyWnG47EseDqw4U+CMafFaLcmnVMYlWLez4Iattnwa0+CkrrD5ZGjb
f144qFz9Ks0oBlYuoX6Iwu+xLefnXXtCM7GqhLIFSrvwZeasOi5w/ZZDcwJAIPbb
kqdvQibt0FJPiyYNEYOe52Ogck654MYRPSfWPds1GMnG3Z3H0qlbHVn8dg385kSf
xsXQoE9pSZtULOupdqPXdoLYOKGpO2f09AE1z/xF2zaoDnuidA8kUyx+v2ndfKSK
Mi7rRE3WI+jWoNiYnafyQs+gE8qk5wP2gX1o9b9LbMvPDCNG4n9zL8Mvhc08evzR
quzxbrPcVUOh8O6CYlk35ooDGJ673SEdcq9BZhCad9oG6ieXyv0wrvqCeo1D/rWc
AgxYSy0lSIpBrb9iGnBnK3DxlxAISwQV2mbcmmp/O4zQDKRo3LOnFdcrpaKbEfoC
LfmD2GIgWtgS7TpDnZVGyKh2ztvV9RoDGAZu2SeBRLLSzFmhHWTzXO8OOLf6sJ+B
xpxzBJdBXpLL4n5Pd46ZQjt88I5HI+PDYnNY4khdMw3Iq1uUtMHkNdCeSEQP0G0K
QeMmYfXlUFQr+H1PYworHAD/Ks9U57232VyNhwGFjGneWOSXGjAFxFKMC3MnA2YE
fz+4DRJC8X3pryYHMm0kUFSjKSUGSFGcOEfSsqJzX5me7jMxtnZnXmPsNkQn5APe
7jUMaHQ2W+a012ehqhAmX+5ko9fF2RT7X+AgSasOz3MMpMRcfhcgt4OXLOk6cuW6
9RGw80zODg+7vHkTns3GU15ki08YWV8IsA8Eyu2YfAawXnWhPxm43EJuOe6KXBze
vWsjqG5zK0HIddMyrDa+K3rvBl1DUIRx++r20FMOinWNOqHuxAtS2SSw2AmfDLgt
BndKGwhEy16XNvFm/e9WzZ6/m2pkqrjGEnJYjeT6lOBCObs6mBwI9vhySPxmhDFE
yqSCtxegzz7slDyK7CNFY8tJuErduhU6/RVZfPNjzvcUicG2/a6u3ECSzhFYg3fV
8z4xzV2pgJmmYIqfbUO+AMzPd5mXt+KmrQcL2HJLCcMfGOMAyDM/S/PfX7AAIPG7
GtiyDTc7QbOXljy6IYoMKwV3jYcRBBUH2uoM3/itpFEm1/QOh4lPNN9VUYRFDOe2
x3Xe+M+UKpTTtBi0mDaTevs9cwN7jRZG7cvASh5jxEZ/Z9KZe6DaLif15oalpAe0
SaXtgG4JSnEvKRrnQuUeKpOiIUS2YhGZxWyWQYLw4N8iBiGhaQWteMiVVdASZobq
WNK3T5Fv2BtrknQjk+qYPJ8jE+4jpqykhr65anKoKYwMBWrBoaY9RM2TDgJ+9I9n
FNMGgdJMCIBjpzihD0LwZeiyKDfuDVZn1d0BMwyuX9R1/xPq++K/Ga9t/HJqF44i
rXKAyU7oUXEVCwhk8aiO+n2L2++1H1jBNVPV2ATZUwg54lYuEPq2xR4ofEOtL70N
4r1Ygur/Zg6wjdCHRaqGG9LL7T8eSGqE5FRNkoM53hmtJKJYWDaiSgKQ8OruHQZ7
nNd6mq03XbHsZmQDnFohwEBUi6I9ncBaR+BgMcZ8VRIbD+wfpF/CzVEk+tS4yPFk
krI3fMLz8z8dvoeoMvYZooyn05tuD4G0IQXqfUbLoNGjQ1hd2dnlyUvz07N+1j73
fuLMyt8IwNhe1hWyyBiOl0ZW3fdIGXyJpR7XRCu4jP8HeApJLRMpgBoyReRNtaNU
bS7+HbG17BI0OBUWey5ayfsbwfxArx1foXIpNQD8Zgob8QmMpPxkD/WQVDtG+3it
eep6YBIU8pJieI411YP6l5ytUDcuzXm1W776uz/plfKZdsF+EgbgLK7SGQfB+tz1
mzR/jOFymxVWSUSr4LPWA1GmutGwgEbzjrdNpsSUnVUu+4hJ5C1286H742mh+QQ5
UaqPbLL0AS6aJFotDKKx0gfFVBpFfqoF5F+NVecpu52/5CRQFgwrAidiqqPxegWc
fgO35RjLKMaeE6LNL2QzN6J79wAYsLj2Ypq67nxodpVoZ9ilxyQVYGwp5oZ+8gbm
bHNBR2b/Aqiqn82/ZgSFM8IjhgRYRPitNyKJsuGrHCD+snwOk+zDGluGdmvPJUE6
nzAkUd1WyVL9WMNxhr5UX6je6JX1FPU6g2esDgHHPTMNPGpjINKKPcvKWDNRk3bL
3eWf/8sq+zpMcEoK4ECyv2YJybEoAU1+nH6TbaPBG0srDVAeMty6JyTHI9Z25YHY
GEj6cxeEtwZz4pnP5qlPRHmMXoG4zfq+KasJRCKoIEp+k5Ydnlm4wrUJ3cZzPboS
ljkRZFwmPgLS3RaIGfeLytb3RHV7KSyPhh4/Itq4Q1d6LrKHosbqK49x1LgRmjia
RoiuyfEebWe49yZdX0GdkN0b6PsDlol/SLfGYP9tmRNqKeVZGSzoPPuvY3hqcuxa
WwEYRLphvcSgh61nomlK/7Wcjim5hGZwNdq1cz9u51wAJZOci+t9dEZ1EFDo9zxD
bERUqjvkn/bSPn50PHCIibq5t+sazItZGUj1SwvPRF3DnjMUvfcq4ftnVSX5IWD6
pxKaGWZvaQstD1I9DbYk9qPeqkMTF6t4MKycl0ELOSx+MjXfXLmGfOitMs/an1gp
wxeCyCNe19XViCU4BrDsxpg959jzFde/b0EurleTcZQE1KqTddX3zZz87iWxPggc
a676MO6fNwLm40gOlZyK44jfLxeClQDgOhVNceH0w1kXiDg34TZNy88VnE8JHj1C
hhrRNLLI7PL6+p0qk50seCnv+A6HrFGd8Afh5zlEa0vRWgfq7RQaS3dpHdXvaSUh
8XrXzl5abVtQI9uA+oT1mN+7ims+mQauxBosj+WqQA028PmuUeKISm2gpKe9t8fT
vD7uesttBdSiGegTMVPlUj1KU4ct8QoNK1rGGC1Fpj6tbqrr78APe4xnYVHlxe68
2BpnBYCrsOZ85yzxTgYWWQAUjUoXgAs3WbfTxTkgIhEzMoUmkE1IdSX/xiPes/4z
hRBgDSn2lq9YH9hUyClWypNgLGt2fv56FAu1IEDs9IbhmiKidVcBCHGHIw54F3t4
KbIgpAz+lw+Cp60urIGA2MMjoMj2rnre2RDvT/T/1DEMdHwA7RqrArxrcxsB8n4O
6QDwTMvhOrxdDTkiz9jy+UK1x4azfKBzHvnDO1vSllrEK9Om22Ihoi0v+cp8ooiV
wc4oCiUgY3jAE3dCilve9P3Q4ziUDpNtltGCyLJTpgwSXz/pgO1CyekPdMZ+A/M2
xz+BDoSxzEgFvvGsHBQu24WBxTJ3YoEde/JpN74wNSseuVWtLGbJtk5E+DiPN1HA
90uRA+9TVYr1EIZXxD5Mq01FBrLsrmLnPJThYPWu1zof3dBSNCQ/S22paUUuCnnu
JLs4XxZCllfIn0y3siyc5N9B71SsKeUDFe6MzoeMnZiF8H2CJBpH5hyydvraqCAi
ZBEReHPsnIQVXJ90rCCtS9HGPYrQ6j7rF892sY3xNdHjwf8euXVEnZPfF5pPCizb
hb+E4Wb3V+y/oFocBlN+UaiFvgtayNoX9JKQt3ah+ofk5NUn9bDX41wCVDhYlBAN
dpVNVDx6n5oGZPUiUvf2T/yZuXENCBY/WQtHSGOTVBWsICWYxU0I212CoEAMVEtg
AVIouttJfdMOJDNl1WzVwZiKtSQgfVTlAHiPEul87fPRJ7BKMJ6MTfHLjCYvK4Ft
YfSDVWd0USiZ0ClZsDrESw7BuSMkz4Iv3wkXVIzg7deLUG70FXEhUJafaAM5yIPd
sZE8wrzjUvXrD+vhfdk+34JzzUqx6MAPEwBkLDELr3y4wr/kKArcVS4xW+XWrt8c
x6ycUdtQVs8vgRiqpb1C7xV7FEEkzQaoBkN1VpOyM2P0qllbtuY1U/m4v42T6Uhc
UBvxbzyvawaq1qoDNnRaDxsaBP5/P1llAL8+g9PC6q4uAtgyVw37TQZj2Xa4xnZS
of9bGDTh4gEjlWrl3URTTl/x7AMuhl9glSWx+pYUR/syDP80IIvoqhHPgOv+ze+0
aw0sbsZE8fB3oJNubM4Fj1l3EBLcgv7cxdrjQNBBegTpeWPGqE6ieCLmYwkXKHO2
7UNmQT8JNCRA/qlgkRvZqpquQEsZtyf79R6N2M48ahgV5Yw2UG6xCXggw9QF9ad5
KVIos3h7/RpXCyz556Q4F9IFk/soaK3AMJyVXOPEGIsYhw+hcBhhk+7R4+zQmHAK
5zkNxX0/Ggj5riUQNyTNh+3JdcwOBdC5Tf6sOhvua6JiRAW4wRM9U/ZhW6LLKB7O
XefIyhHK99kK6zWbHHk+UuCr8PtO3C8lIqYSWBUedhhWkgW45WvUQPQP96rN6/ea
PVD4fZuj3+YjGmTDoewiwtwoPIFEjWmC8CaTClpcZwNQq/+R7oEJba3ewX3irkGm
S7wB33/pARaI1R1UE8E32SCe0oH5PTH5N54fhmB5Pq7JIur2Lyp2PUH4Y0qw2fuR
sUgJI5uwfkaskV0EHVrJeiBJVcoVA7fWm4tfTVNvja9p8mBnqFfsjOlqp+B7R/I/
M6FfG6pCICupxm/271RchaxxadAoFfQ+rApPy/SGpCLMx5cgUcUgIKx+LNe/jpYj
bwF5PYnvgz4dIhkIc8riUP5wrgTMMUJMNq+2jem9qnqCu//YprLnwWzn2AxEf0WW
hgHnwxrWWbw2cxmrw6B3Rt05WDuI0ITmMokhxLcfvv0zv1YbdsPFrYTqdWasY7wL
pB2SW0jlMAvdtT5f8I+WoDndM3Ljq2Or/5wmMx+KFf2p+YqUZl5l5NtnX1/ZrUTW
K8ChR6z8sDvXHit5sd8i9kvpe+i2J+QSYJEKD+mkHNkmxuRGMPIPwv6jIjOPeISt
K/iJ3leqqjuOHsylTv8qGqXRA7wG+VLCkXaPBSNvRXpgvGyvP8TBkzh2qS1vL+Zh
QAqWJYef5yLS1qbtpuZv7XhgAIFaIEQIFZAzsLjQly2pwDi9OCeyKAxsh2W0dFZI
YhljfN+PH0oCs2F+8ud934HR/YdYb8mnuKEpQwXFPZLgwim/oRXiOUyXmIwhw5mC
aVyWmuR5vaUBxuPQoHYmrs2aMs1CctZZZH8AVF7PyP1NuHbS/Wt7QxFJO9bqclmb
RAImUIlv6fykhphdv9mngFl+VhNtU8X9RCvbq/zLSpLiIr5IZ89KL9X5MgZYZzjO
s+z8pCiRY3fHBE3/WPS3cdNgvIvoSdzrosYb/701Da1/PUYzizQlsn6oSzKVtrpr
OfESqZWawcbzVvAuXJXbBtfwNLxJeS/oa6DzUGyc/YfsyO2Qp0D93HRkqq2V75B3
YF54q92AXVt3Vq0WBhybDgbLSvskcPAm2t+IWoVOgL0k5IeKy44ahf5AAr1YnbSI
RfACqUj9cXJezb8gutLjsMLzzwBHk0D/ktwhgYOSxvLIP1NLq3oHt/tkXlTQUP0Z
6JOYCJm9mSO6iU238DUcqrRqT976gSSozjVsvohJ5j6RNfCFUj3KhkzUHHQrQaIW
V6aZ7fPusyNGvYaW9e3yQ9qQP5WWeCUZq1xT7mtx6TbBgQyR+9+l1XaIHfHvjwaT
YZYKnU12SJ+Hg7yRiI8AjzObTlmheD8t63u4I7zNjf3DnemO3GeAuryKXl+p7Z1k
Zewr75jINXjriQb+oP7XWdvRqFYjTjidwaU7Lcm4MSQm5jKeX6obbivAmM+7icm3
Yf2v+KuIjwlrFu6+T72jHsUMPst4MvEwdYkpfP5xGq/wzYA+VbVCreDi/OHG00Yt
xzPgWhtGu81rrE1DZCCMKolOjyvrhvQgaQLxfvIpKZnzT9EzAdV7bWAuH2MxDxzN
Ymdlnogd9sZWpYqeraWYQQFzQ/pcQ5gkfy/E5lk6CPF0DW2Tx0ciPFXqJanKtohd
VqMeoe6jDaxnnkF26u1aloV44IMzDogPUgOHyRdfA0Qv/hvF6apag/nrOyD/XRAz
omfKAxz1bqNrT/ukhCLDFZTsSycR+uUOgax4R+yNhSLLEuXBiJ9dt12RWPVJFVh6
rkR1Q0dFQ1qKdq7n/UeYRH7IFb9VzwgdCP0ui6ESGJSnkP1ZdtumEoC2Q6RLew7Y
IYiwYExwCRuFz7GQnMpGe/VYjRZBluA49/grVZ2USUOrkivRJ4+yhg18he7Gejrg
cXT99kWWUsvx9bbJ+Y8FzeE0UsZA2e21STY7wJH6qxtLofNMDw16ViTEmS78PoHG
7wmM2rTuf8C04rkZ/gy+Lj0N1yECBFI1jtwjD6rVo12Lt9KjhUMvpokCf9trsbIn
SQwhnfXa5TnIDwiuoHLv4O9foN43K+IXIW0JRvTdTI0Hm54YdM+hRzy05TffxUIb
D1woul3FGYiLBUg1dV4I27hT2LKdZrLBZO/U+GwWF/to6R/t8ajDHtGnht7yGE3/
OJRrjaV6JIterDhDIXRHSRur1+8T/9nLETBnEhHargZgltAleZHYzRlbKShmZwAj
w4GGrWL4ApecKHwsm60ntrOrrP1n/FkGjZljvJPxBaH0YiBu4tR3GcPMD2uztaBa
5cu1VqWY9Yh12W9bHkAvsebDRV8B2DmMlWUEegPB8HfB2ak4E3orYlQcKRkKGj7g
pwtmx5fMOBDzQRWIQmM4B869PPr5uyC8UxDDhk68494R2Mmct4fvq/wVrV92S49n
Jjerv2eIFaQ6eDOhdKGh2dp6o5jibAOOm30/Kmj+mMybHpAcyIuB/l11Gr8vqjXC
/bz1JdBJVeEXa2uLwSk6CSSePAchWWyuN2bKxbyk3GFokIt7P23vorPgMT5/RdxR
U2kyJOAgrYTS2oFW8Db0dSQNdsgJfm9+0rYrIqCuHzfHcQvz+ur8sw+lwru/IqEC
Iqv65Ngr3J/i0YmZpYgB28agErcLnyNZ4IHdI6B5yEjxzFz7Pgou9HwDe2NL4nYm
9FNYlLUJ9njAXn7cnX56Wua2qlSo9WYXc9VOwQh4Bfixxs3kQlA+jfKrSeSWMpEG
oUQqKrNHK8rMHonre1jhxlUA53VJ6v+cnsaT8W2I4PZYpImQugDBwy6ncypC6D+v
3lpHqhZAsRaJcS16qevelpUdMxBmr04TaiVNeo7Ve7iT6PVgaadJ/OeczLG94KU9
LTPSggW2rDV78M7MsdWYSG3RND4tYen8wCGn0qL5073JGlUFWHeFxRVW96Q5ZzxN
4LIqve7ij1toVx7p3qjbG/Orr8ysmEdaLGzTMwzimQVNRxKIrcNoxWifbNm39scU
iRpHNZ2Vb3jA31SpmX10LQSL05wuSL6IMsaNGJ/4B/0vAAErT6+Ft/cuh/T6ZGWA
cP1UWNbStQtUiZb2OCF9c9Mw+XuhtrjCtL3avRDXgl70ZDzOdeNmmuYzxW+WybPB
aS54Cnz6tPQJNV2AETRBF47P2Z+4AEI/bqdvXSfv5vD1njk9WXHPOVIFubABKcjX
y+MmdvjuODTVWTVDeYPFqykcYTUg+8DLU4bXCsewVNcOJZZZ6vfw1ggP1ww4S+iB
PJLSFM7Sah/f90GpS2QMvDNwNcDU4hBW9K5v8lYn4jAMsCpI+TzSeiBiY1VGfLhp
l0wIPlVdqiiUUTKviVFQXBRRooLJdBPY5rMjec7I7zlo0tsPZtVly0G30tZhYsER
vLEoE0RgPZA9fcsy1Q9RuWbhjTfS48Fb6rQgieCpZ+ywvFDUZsSnFIkhAbBE7vju
SNp5r36xPudWwVLH8vFT46dKT77SGsWUHsJsWiRgYSdpEA3tpSQO9NW5Ti0PpttC
0hzsdB3akaIcyp25n1/k9WLQlfbqt5K2oKeCZmqzOOn5gEheTLvxnHHby9IpJXCt
hFDXCMEieorBaGrY+iV/l+Y9qGS12CD31WYIa9m7PluYg3tjaBKR6eIpi+76giAe
uxj33Fy4WurAAaW7h+bfvaTNB6T9MIptx4FGHu1N/5ClnBmiXMv3+A7lIjAKVrZB
HZHiuaDZMsXiXC94WHJ7Em5UzMpHp+Hxbew3XC6QUk5DnHaJfz/VMsfQSv1z1Pht
fkXkt6Vo5eciBufF1MKCqkEL4HbwGeFKU1X1dVDFx52ovyDeA+YUZT6fOtG4WCxG
YXps1YQfCpUhGfLTv5B6Ph3aDvivAQwCzq2tw+aizwgq+dvxcHB5uKIz6g1k3EZ0
R0ybDc1xorP3e27D50vDfMYh1OB+cAerKCIc0XS7frp5pUO9yJOIYYg5iQ0Te8yT
rp/XWpyQ50HvSWPP3FETRH8MPZJEt3xqWF7HJFO79qFc8+NyO5Wy80PvkcRqY/Fm
EZCniuSRf04QNSE+gmtVlTK1/xiXn3FOkSmQHjgcPjF2EOAACvzNuXAWqrHkLkUx
veKOE9Lz6NY+np4pjU6O4uaywp6aCdRJH9rLzzN1og213g9y1Y1imkQ4YF1Tw3/H
qTvplBXOpw3P0Omr3TROhl/Vqt2vw0HMUBUkP/rGJoefwFaWLULlprohW1t2jNuX
vgsf/hAphrM/OwZdKu9fL9/+39wcBWMG7bti8GJAvxIgnHarcRXZYqA8oor/Xr7K
10XKfJ2anC5lrX2I6zjaS6NLfSshh/+ahEth5PcJ0PXc3fX7nxNLLksWY2C0TwYD
M5t7CKnJurFPOdBrXe5yIiQaYc2d16UHQg1WM1hqZ51+8WsbWOjMo/fUl5p50jWJ
r2QWPi/dSn/XDCvxdj7ivYfirlrVupkR36h7NgWhuV+aaGHNM8wskYfsfhDiBoC0
SrXlKjcL+uj5BMg9HovAdslRbbisE+W48/Ufq3X1CRArpKpcbtoI4QFeFzhlH1D1
GVk38LIEmlBHLG659xq2khUrZk9uobPoK28TZHl16wsxgRaNckvNiF4QyxCTGxM7
UMBR5gDS94lCE94jVnzK/bcP57ncphZdcXgfMs+Di5l0nZ9rxU6RDUUZhYv0HkdU
FIFH96IOioX1lTjtAEakZsW5YMB0BW41mwbrEzh46AaVF2Le7iyZeKhPcprTnnbs
wzFQU0PUdIByQuYKNaN51n5P8gs78clTIFAMiwzdAsYVO0rI6do/HB9+6GzyAnaK
M4KfdouhUHfk/g0ca6Cwrps9Zea9iZcOot3buBLliXBBP6hnmivqKEPBIlfAwFEy
jH/tDdCe1rFynggwMsE7l012G1DKIss/0e1FCJ++9C0ehLhjScpCRJ19NDhRVzhM
4AcfFv4vByP2hijBzF8fLkYWokzKO1Rq3y7QqQnhKw30Rp0PQ6HTOl8bSG218Xzs
60pRcIrIQLm7I9OGBHG0v2m86UeJPGBfRV9x79szRDoWHC5+U5vLlhbMkGasWHXd
DGM7L2iILYyWjcJV46pnHrJLNV7zeKZv78gzJKkm9isbgQtaZKB8L1DANCdHhk3N
PCe7Ue6zMDiH7I4cfVpkuRXB1rwhU1MT5/gPzius5HcM50zP92LWj3ih4VFTZ4in
m0+GYo1TquwNx87wfu3frKzbLcriJLGiUbum/2itWVxHNEzxGYD0CqK13KLY+GDL
vLCAvA58lAnR6nnOEN0XRdSg6lxZotZ2qB3To9qo1DA+g9PmsQuR6kKk4N8x5Z6U
vLxDawNZjVDjEWaCq8k0tKOWvgzCIVAufq/ohRsK7mgRiOZ3xS1iB92gpcU8yoy+
4B5mgiIDwOyk4Mm3KJsh7OvqBs3cEa+6j5FsXX5k2Gl6Tz5piQux8WM15FaajSFL
cpHKhDk9jaJ76szhsv/64ny+73DLBwU/E1q8PLqVBZuFN8e+EAxe2YBj0grsBJqd
FqftVl4cKBnMQCX5YC1AlWZf+Ek8OfUY85zd77v6pMH5eFZsl0A2EIDWK2vqYFDA
hWjiSl9FF0/x47ZFLOa1WAEvYQMpqDGV88WnVZzMo+KR0/qv4F3lXU20TG4pYbkg
EUe/6dmckZVzrsCI7yYWvEQPPDLz8xf/O69sOUbVyM3TuRO11giwZl7go2Go0zae
aD3Es5/ZL8/wU0mvtpU4Ohi2VuGp9RdNBNKDfk8oQBdtq3BcwUXWDqgkWfHQgs79
qTuitBNYRPEDSJSAoiSdPDYMSw0CFnJ5QdnI3YOGkXwcdJtwMq46uNanbgcqMuaz
MUVOxZf7JOnRuBbfKeZJbMkN61VQuCgIKCsZv1TJf7xpmhhzUL4EvOpa3ImjHSvM
q1d35ippc7WndlQVmACb/0gd7rynFSj5xoHfnbOwSoemdpbhQ1sDGCD4nlmMUWUT
4scVmhrqdT/8c4hRvZj4qyqrsehspTkrGvjv/RLhOWzz59VTAqnzgZBmVoZLlitD
9GjdlF3DjO7NPKpLAy5TfOioHg/zopZZHs1JxTEA8g+3852zOoyrfWPEhkURZIbq
HDexkJNLjfW2U5X6ScQX/5A7pdZKW1NhVVwJOLHfLVMAJ8o9muFMfIXRE/FpMXWt
V6sRpva+J3FYKQIksKhKvyG77ddjI13fwl7TlKpSgL50yWHARxBEmHKMVSEW+V78
icANXHKSeW/1mTuB/bMzZ2USutAGbmp2OSpelyzHpAw5RXueAd+RSVm6q164OQtz
uD+EBPp3m3Sijez6mBdD8EZTr1op40Xjww2O8f3gzJo9GjppNbl5Q42taXb5Ugwf
P92uwNXLOmYfy21wRoFSoKDYGCxZWH81i5PsJP+pVWSHB02nEd0lpMm5G8DAg/GO
J5kfRDcpliRqn2H30WV24vI3fNwuZCguvS91BkwcThlo5pJKR38cNKrCvnTfGsmv
mwnCiBXCURd3JVIUQuSswjMKNlSM991GLr1aJNeGaSEGDbzzy8q2r+lRnSVsXdcD
A75YN9yRoekmq/eVdkjv2jWpxuBWsa0ebMgNg2xmcnL3V+0u4aQm3MFVeXY4QHqc
CEaUeXQvNAE7vYVJIUQ4n3yHvJpiw7Nilx/VohbzL5i6RZ9n5kf0kqm4cRLTZs7e
bRuXZMiG8FWqqpMhUevfry3NGMC390eqTUxcFhpwS09m3zjfttFbZPr/AtoIG2Qx
KPovu3Rzrpu2vAahlUFfJES2YAM23AnlBPRV9PZvhp2LX068cO6z92dhFuyPXbei
QtsWQ+d2ScLBf+gO4clG0TB0wrUWsdgLxpc1CPHK867tErHeVTruB6CLre9LW+JG
NjS9uLY0x2cWsx+yvTGIyY8c/VRq6jG43bhe12pBEEH3Jx8his5syI+WjzxnLZqi
fW6irz0P57YZZkLU9RvfTCTBZWVU9uSACDQKzYrvKgwO3fX2jBmnJmLTDUMXwFsI
8uet8mszuUn//yPk3+m1FcKlj3vfyn7p5cerMOS/xgRbZLfkuyuEwqJEPkLKa8s8
RmB+1WUDa2DNJtEHRAR6LiZLxQlyAoW8b66/REA9Aqi0vf1eV7oAnKp1ljVOw+io
lfBX++NxQhHyiXI164fWG1Nn1ryAEe7B+e/oiM9YRgbm2gDZfwKWCufvWGTjJhw6
LzKNFfEaq/X8SLAF2hG/egiIHI1SkxT08TmvQ5qor8hQ4wJkK1OzU2EhoSTUUZKH
oHkTxi9NlTASOgfjxcBe3+9yTHx1/Rd0Q6qVCZtUsZoJbQR/Dyk/M8t9NUm9p04d
Hb1yVNDHFuQHZgoQzv2z+34/54OsyesX9N+GcqGWnJk6YRjjpYDwBlmxr4iGePX7
/3J6P4Kl2BGpm/EvrIScaBx6RcNDUZXcX7M1S0S1tHjTfPjB4+FyV5QC9cls9PGz
bHoGUiLpRqpbvzvEaB63s8LqYnGonZOu3D/seo7w4SvKZrCIvTp8gztuRmreOQJt
YEl/G+zlXHM5RYcF8fRKTGFmcE23LgYwK0kc609zymcooAab5p3C6hVpXRBNj26r
R0TxM8QtrWujb1cj6yrTS5hVInMjThqd6QhvH07axcs/WsFDy2ynooxiJUtgfDXv
vuBQCBQ5Uw9jEouWJYBa8M9RxZHIIeEwC64WE+GnVN2bGAFAEdyXwV6PsRGrxXvr
V8q04mE38s69dTCzrnZnZ3A1ST2PDejUg2bJF+Fu02/3AiqK8TomTcZ1e8q4xl1o
5mJKFoBf3KzZFirhAJ4zDqSRdKabZWofveT1WcYStS9AZpCSQtkJAYf3RyQxoSQU
qXe+BT5vVNihqz4m5j8YNXiG6jGLFiOMy/IuMqal25SDBtXTMGM598bX+dlce3o5
lzrwYL1mMWBRGBRDZC/j/OGRZEEIezOLluUWXF8WAs7omFmBO0iykYhAnQhT3qCT
DTDDO7Vwi54uKUuMZc4BWfqbGWgGeZYc5EyHyyNB5HDDeMFa4jDg7ykWNmpzsVez
nDYxzKcZPq2qvGq6cqnl9K9rpwEtu5ETlxb+3U7nNEdUZe9QtKcuFMKi65jp9us4
qG4uqvRymnh6iiFH+IIjCTNDGPQqLkUgtlCutUi7W/BzBW0oy+WXPP146WoE239I
VLWB5Nfmq2SdBUN00ciZ//sTlYEaaoK64MJmngujrJp0yh9cQHQl4aT+z3lAaY+0
gnDoNNlz01en9yJoZ4h5yC9DXuvNOD31SIxbQhBq52oD4UZmch8TuNxUgTaccBHI
XC40PxOweogaBf2Oos01Jiy0BysQQ1jQR7U5TA+YtgeJITIkcqysjOV8TzmNW8o5
CHhIHLhPl0QKLMysBcuK0Lm4eu/FxZFYLFkpSfDNTmZOOQ91BuUdPe2QRyAJcxrP
XFWq5IftW6rt9OuM58Gx1AZVKERhBEQP3XA0iOcoluDuGHK2D6gtcTpFg+Uryj2Z
XMA9ge9PSm39euHlE2woELb89CbOe7lIriXpWldMWe+39Z4zAIhbFeZz5YjB1FoZ
RNAvLLSo3WPsQSa0rZtXZlrR/5OygV9+tLyVD41QLVnQxSudH9sq7Sl1zb76mc0E
TnmoeKDf81HizEHCR7Tlsply3g56tIgVcX1ZxMN1C9bDBiFMNf5Wv5iCVZrnuAqF
cwHzBhR6dBWhtIkfwNrFKMgoQvPEGHIOcCOxKyRqRO+zcz/Vifv7HaCuGe1tJfVk
ITvS3LpJ+X7HyZkzy+auuz1Lxzz/rrwqZNhVtLYfKNwZZwTHKb8uNY/wO4zdlkJ8
JO+lnZOIaaHypZ4FBH5wQiwLOF4KVuvzAZ7LrHwrDHef9SgxVTOhuW+6YSpte+BN
YdJW3vqVuWMMSg6/6fI46TVrPjqvAq9oJ+jTe/FphMXWJHiFhsqzUITkTz49xBDM
5Jtert8EhRprTv8UAPeiX/Ddn8gYeVB4K4jEgRVOlpabcuoek1vGlH+yBUN2uM2F
A3xsKpsOYYqqjerunJM9QeaTR1XPeBStNQoHjVW/ipDVnwivR7LlHR4kqab1TGDa
kE63kmIT6C4P5ONfv2vdjvzhrS68sS2MFeMHMJ508nAY49wvEZ6tPgZEj0tl0q/T
YoXODCNLqMYyGB4xk5CwqytJY5H8mqIKpkzD/xZkvOPOxXE+5qF4RUviWAMLZd10
MJUxfh24nircOl1r4RFrAw==
`protect end_protected