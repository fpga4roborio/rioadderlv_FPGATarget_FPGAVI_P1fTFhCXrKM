`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
ddtXksX2+yylW5zu6QL2Lhnb2d1sD00763mmSITNX595NcHTEkwn0zB1Dry37fOW
FufOhVzEJp80NC5qZ/+F0Vk7Ik02dIR0elf3clrjeJRK85K4e3Hoo4xn7YbFUIms
l/8VZSb14+JVGURjfswrIyCUotIzlzVYZ6gzoZwDXIi5gQIBf/gI+KxNXPaKV+PQ
Ufys/12rjO6aI/pPlqSm0hCvftmBcnezN2hk1UeXgOIuKZnogjOsf0iJVX2aOOWE
6pD/psybjbnsNB6kH5uFTA5frkzIzkzl5d9+YDm9OyC+k84E83I/7/j+rk4L2dah
QJOvksSIzN867/4Qt8qYTQ==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="MvBXkzurAa5VTw+1JJ70nePUfoQXBvZOku/SMmg4TwQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
oRtzZL4VJ4iwysPsC8SXYCzXS8Fw2gtZTOskLcDV+1B9Nzn1zTyNtlo6lNICRmmK
ZRVu2BmCc2G+fmzynYlNTnSa7C0Cuel6FYpxCBlOuk3OF2tzAmLAuDyOH3Z1Yjzk
a0aHuoCdIRKv7BrZCdALt03JeUmXKPdOmIlkVGFl8yw=
`protect rights_digest_method = "sha256"
`protect end_toolblock="Jn9CQpRhJt4rnzZPRk+dOpzAubz7omckX1MrFd4p81o="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 17296 )
`protect data_block
gD6l00tciPUa6pDNTk/+t0OO0nC/UTtBwLB41d4inuAUA3i/ALrNyoJVcBnAmEQW
ptbcNp5fxEUJjnOxnedyZEuEBxWRieZFQnkRdF269oNbX3CN2hPF/Lrg0PkLNAWQ
cKfPpHaAZREmKVXa5cUCWhqcrHpK68uvbbPr1lK+fr3atQ8E5A3VM3O8ud7DC7dY
9z8fxMb39a/HmRTAjINEQHW4Ywu7+A9zLs8iMBGb3mYKbuYhH/XabiWwxvvcl7LB
qjU8JqFfNCOtBJx1CNsIHWIZOfcdWHRUuRqBZNbsUVnUs/Ko0xnt43FbA+7LmLIR
c92/bT3Us5W4ImZPlms7DnojD9A/cs8WVN0bvrKLCs+FQ5d/7BjyBcDETeCbCmFs
7CFV4VAGS92v0VdisYpEAqc+5YX/MNyxBOGaWJmoCInncYOViBMlLEkqPxh9AxTV
kCiCSGj2D1jW5zmLPM9/2jWvBe/4NZMM1xjA4vbhi7k1CDF2VSb1jyxJzWcrYCRq
pH0CsOBqRuanzFyWB5bD/p+3lCBf8hlltDJDu7ZoMPUPqENHAPIWYqxwalxKEbQA
mVmoZD3MBEj4vaDmiT6utTSKtnLyASz+NHcAf8EIk8CiVmiUYTjrIJPlBxl5Gk4J
MhbGkDPD1seYx0BdQalN8zXUjS2zd1EP6jFay2fyvsD/Y8hdlIYM35kCrMeetBi3
5i09exdpUPMqxaPVQFxh3JDBU2lDl+tQYf8a7cz6roGnE0JUtmHR3kEBV8/SKKy5
kLbdYMJuK6SRfMZLtms7DqeSOfjM2ZiQj0Cw7LligOdd/e4s8hjVAnmhmHo0rze8
zA67brRpTViXA/+93ptwjwpudgudeIVyWxO3d/eh1Z76o+Q7fyNa+KqQ6BZWmxMy
MvEeTrBMLkdMLWM3SxtTc2/EAbbe5GmcQybsVxUhdgcCS+ajKRpyqzDlqIgvHvty
Vk9+f3n8Lkvyc1Y8TZr4+5Gqumz8/M1XDxYcwlvKod5CVRghcgOINgE9EhjwHR3r
Q45PF3E6hk8aJZc0KkhwWC4XHP1lTizMHo6jhsyLOn7+rj3Wdv2NbW7+E5OjL2RS
rM7AU1FpD7/bPv+H1cZKfeg+3VDx2khZy09xdjGr0iLH3biGzq3PUToY2IeLaRpJ
3SkjTJQ8nqpnM1lyDAKFjXQjpawOXcZOBdnDqN/WBbhqWIArZb+75DUCBBIDvwkG
ViAwcsbXXunpsiAmuqtrKRnmYpDFpetXndwqoDhHVe0pFVg8JdAatAMEScKYMleQ
+T2Xf/tPwnS8ckYNZSP0DQrYQH++gyOigrspCpG8KnBRQCUkHoEAxbUTqiPNuRpA
bA2lhHIFgnYRjjyb4ML6JfUFavmDXKLyZY0kyNCxYvRWvuhA7vCSBnmknpauFKyh
r3ORQYZpUCDqYmGZ1tIAc1sUXJFcUosxf2VyHQAOr2LVpIbkIDaxck6Gc2qVE/xO
2nA/zpJqNyg+sS7XMJ3ADGKXBY2mhKM+sRQBVHLWmRijHZqbhX6tRZNSwHVWibwA
+RCjuw9ohx/P2fDMR0UIKboVxmtmvi5K71djAWA/zGv8xfEj0N+iJSzGCyuOcntX
LtrOZPkyisvf4joHH+mxFb/zxgJiF4aH6b35VuUW4XN+wOxC4o0EnbmxoNkbn9JO
KTyMoaNTBPed3GFpQVBeEfrOYzkznaQEnKeEHa6Bhx0D2wb5w2m8AdbiskMZn9Dz
BKfXJ1hky58Qok6QkOX9/tN3IOn4GZcNOn0k/jIV56zgGoYZD08dyXNZaAy4Jz4D
BSg8SRsUhKgW5ye5IL2c8HIAQZVYR68WCi5is9Z2kl6DdT3Liq9DYAcIXpuGsKd/
kGQO0AjHmTnO4eQ0YK7Dg+jSZ36n1DdXDZv+FaMDgo9eTRIXWtlyCxF/8lWEte/g
H27WRlFpes9GrXBMYsJVW6qcC15M40V1vsCLGB6VH9ScsYyBXhttMAw/KECq/r2T
eDcZf9KWR6X0RFZbZHLFcWiMhvCUVRvAWlyD9bghh32sSp+u5DILnxkP2VlHJjen
PdnammkUOLq4Umvq9DkKYShnM2IlFtZKZEd5Bkhv8Dwyhv+WaNCvBjnLhfRTx/2m
WZkjwzOuXR/uDAI+l4cgrFEwdx60X5X5MCqC+PhoI2b33zMzg8vqd1mOQ7HwVM80
Jo1fYUY2aHWCPB8IlKy/COVWA+RRJXeCo19+NB/0Hwjo3NWr/X516I+PJEktaJbJ
l/z1C+WpooaZFhe0C78Hf/mI6nOBVZf4/4b+lo7ix8o4ZdtOMCRswMvxseaxzRpb
QAgNZc7GXvNU2b9rKoaeN+8c5qEJ+n59EC4DORE4c1DWB1+SUQ9tj2+dO9OxkycM
W+1WCDb+QQk6PHw5mhHMMyWbXvP4iJXBn4AJ/Ka8GBJvlmqbybtPOGldH7PILjpQ
2I1r4XNIfnfcEV1qMChAJf++H3ohxthVgaAtzbu9yB6lLlVQnwXdu63LYFwMNgnI
xj3GBSa1XDdIVYLwgKoPKQvNwG4qq0sbemsiViuAHhDpzXRIzF6+xA7i9nsdFVmx
qe+Ez4NRAliPx1BAEu5fnRv7MhjQXNEiOr3X7l0qCYJfHAD4EO8F7cLKqA2NeZu5
6/Mmxhs896K/o+ejJHTCcDHPCOLlt3cAT/0GdSzBj6TLdBq8C+G3kTzs9GYTLL8I
pLi3h6lGPEb6Ew1UAMp+J4SYuQh5w0fntpysU3iGC3gg+ykjCCjcFwI2Fw9x0v2o
0cbWb7vlKFKeWi6ufFFZuSrjg9wI4dGdM15wGC3WWMgRch/t7JtS1wjlyGG9SNdk
sj3tFh5ZLc/foBDHAWHljGMhXCW3Y2DsuApPJhSusBPKZwnGWJ7YwWqVFpO8SCDY
B7E1BlUlqbnYaAWxi7ZAog+mzE70NNGsOD0hugflCb57fSMBBjLDCQQvUpMnYMRF
1/9JXLAg24FPWfJpxeEJT2ifKZIVyCCsd323TiiSTPZp3WoHuh11/QVSsOjQwiB2
niO2yxMJkNK77MVCPqWww/U4PSvJBl7QVoXfGZujJcT7xIZ2pXSDlLmLNGxEFWW8
us5y3ciOI3h7mAAkuD9maMnRFcCAAs2STjSSFgNXdi5+SulA9aJ2+PmJDFQb3aoO
SsFJkg36wh0Uh6j8IcU/1qrSG+j3pPb3jmDlrLHJ6MDcX8JfyQGFSjyMqs18H52h
3aDvXo1emwJjVIqBButvQaI9QUI64aaMie1KvEZ3XcN/O7uUPGIpxDhoIc9ePqk3
ohX7IOZXaloUIPuV0Z4DZGK35/rhTuk/t8gDWfVGDt6ZTBr3Ieblrrd3rrDWsLlk
ZBeWxz8djhllbukmeCzEx09fqWVvmOzGoqJOYtbWydFoHPP9ai8Y/FuKzlQsPSWN
YTjLRaRPbr26eKVqxmg/DxNWUDLqrWE4uNyW76Y++Blf5soTwRS7LmV1YideVRRx
m4bYpXmJrmwmU6gKKyKrNYD07k9G38NiRYLXOCf5Zw6YEWtfL7PvgLHvbzL9cBgE
XsiHChQlDWqP+t6Lb6l5nJcmvAW/NPO8FMJNbLKY1kLV4JcCaU9fOGbH0nWxLptF
9RfnC4sEA2mOJWVdYdaZe8tzT/h/uxr0lJ6oNPJvyDuGqRCZhyxj/B6XOHwpsY2i
GZ0es9jnJcus0rVLc5RnJVueUaXj9pQBBWdXXyCTwHu2Yy/tBdk31/YJ0AAJ34RU
HaDM4su8u7NL89QuOitH3HXMfQAm2bP/ooDQ/25I6MEo5BroDpq5MwJbGCgTpiti
/+8oHy+fPDAIf8GxPIlXITMpGQT4qWDRhJGvKc9LvVrhjY4Z6PjQe9dbok9xAX1o
8Crkev9ufPL2ILQzLFrA0ImFCKlzpPj1t26cQj19rD3xFsiOH7Mx5RlmuJaUmwuL
erYlA5N1aNve1kuFi7gByzudxhW/SsYND4XNbI65TzF9To959SusAp+AYEXZWi7j
Fwe4ZU1h84P7N3+AThVOn28Cjki8kZ96Q0STWLMBHCaBvVZpG1wYUxvLYrZXZAnJ
cBzYzeOeT0LK+U8yE0ZBWiVjTCwrMDGoJpgthTBw0HUc5/P0hCaKELpBLTrJEBuk
kqN7Q6Houmwfq3aGo5u9u1+yRkv5cPZ8TlJzVtPPbinwjfNukPLE2ttfv/H0TqVJ
UP0hMr/DvWp1YvSyz6SZIvIaTUjv4xokRylFX/AVt9UKuPmhMZr3gFaQD8K+x2IK
bgw82HB6MdAMd1IR6aV0UFBQoLi/hGEbgLUC/f/lOd9+V2bgNq5fXnNh8Fa730vI
7sk5nky1HpnW7mbJ2bp6Z/RZamxoCqQjDu/Pqg9fU8DCzvlIPvj7/QZy2tJhi2pD
7I5KUwXP3wAgz9R5K6piM+o6JmujHODF2vRnQHpEu3w8hAdWrKKnMfQosHVoreCT
x7FDpruK9z7gABPPK17SnEFLQSGQwG4ZJ3cP3fGRqQq6Up/Bxb/weXTtnT/xn6lz
qNWqjz0FzMrVkHQ1VsQaf/rfC4U3ZEPR7eo/NSbGBHCwtUWEvm8OBnwXjH5TrtZM
XbQrc9FqPblkSuEcQPFHhCGECCkunqblYoBCINc/PWuTZpCTvG25iJ/Rd2bAK6d+
nGXHOAjwbpWCwFv88//ab7wtw3i/VxNTum3K+bf6cL70gQJakcu99ReADe70Pkp+
LMffMDDnDqQ2ZERVuYYZ2V6V6mmLtnZxq5BnyWPFpOmb6GaD05ion9F9yRqk5u32
RHGafwsSz9J6Ld5UPOHHTpioYAsRO+nfqe7lpfWZibSFWPzBrucRYnAU99odirOW
rfNM/9pItZOMOabIZVtH/BW0aPjG7TXIi1QluJb3UafKDgrXkkH7JEFVP8MSCgqr
mxTsDKEh2lNPyiemL20YUymdOAzUmxWETHIhe3Yn8B5UX9SyDfguXc7PWtGBUUWa
7Ct+Y30YGc1cV5qCvzwhfDESpI9ZgCd3Iy181vcSK4AoJPWlVRmE2XnMC3cgjwFC
pkWPBCqBBGenfxU2b7lGqJsr6YTZ07r5mjJE22RvOSQKL2gfimXtJHiCKP/Rzd6X
ze0HsWSj5nCsIyrNh8GAoFyp4Fv2PBe9RkY1NGMKSyB/vlrEMXEKvOvAlziAGUWE
3/FSktluzdBcKiMUQIxkzC/gcn2i7qFMVriBSebeq9kLOzUtZTqrE6JUn3fwLqTb
RHAOYtaGKxbBRK0ox3hdIJnNfEnjA84tMmY4JiOG8mG0PmtqH6P7GL3Mu0mky/lL
DpzB45ebZ0aC77D1DP9lVFyOB07BRb6P2Rih53a2DjUmxlFSSFDvP1xoqgWIiSMR
lbBJ+yU77+NqevlPXe17Mp+uiNETdL1ApZtBn1aaOw6KJjP7nf347TbKzRcQRxPb
1tdx3xtzCX0mpeFW1fLeXR4e2d+70M5SaivH2LAh+z/zz0qsiNJLkF2PPzOuXvxA
bOLk8i5d+MQRIiF8UUd13RHbakg7ibHiqhikZVZ081fnYxqRwkia5YWWFYzabXA5
mX1IwTYrfw2yiKp9iyyOES6QqOPmZuyYxglH9VBUKSKf5+sr4LamcnAI9hj6HH9/
gCnGvAM2WGUpl0NGgZ20dNzPALYWh/6oxgpCTAY09lyevvSQ7ic2hDtSFFoIzptM
R8ObIzj3nmSDq6tvIlK+aTVdjNmZzHHGuQwMf/sSrlR3ThYdVAiLrXvrR4X0EzoF
DBhNP8wXzX8F2Q1u9qgahNSNg6a0YigJpvQahPBrlhUwGBTIgYLChRo+C/8g+a1I
YFpt4kZkeHBrklzIOxKrJLMKrDaOPT0gSlowZlJ0oQP1QvKN2Rhcrnst7e0Cn7NV
3W00F8r0JdJzeZR+OaPsL1sSYzKs2NKqrgyjn2UfXH55Z/e6bExNMyRIUJPM6HI3
3vdElG9us9a9chve2Mun/TgANULPZXlJW2F0UWt+Dl0IAWClk9WCMPFhllxXGlGC
evARcSi7aRIIRPLq1FqSAuVmNnZobf+Gvp3B8EjH9p3xfr7jpmcDay8tTvxyoFKf
M2gAMxRVQZzRYgB7NaH44pO54XkhWP7FRWjb6DcVdHnrJcb1OGvu/lXfnYlAtc6W
FnhxtEu5+6y/Hu6rmfNAYbMZVsIEbyB2SDkDrdEkXhWor7sXXi0BK1M1ojoizza6
Ea/DL580g3gfoFZxrSbNU6eH9rmIwn6V3ikRD1T9pvynkA95Px5d3TC0nZhsbSsi
83vX5ce60FfXx63jwEIdZFTAWH+VD+vBOcZk7RNK6thxOjEjWjJI1zly51EwP491
LA5nX8/WCQgmwjYRLaycBq0KqeYXU7C3ZOKKPlAsZ4ItIhk8vWu1ZG7dIKfKS9QI
z/ZhcIDsppW4RWocE0oxDsP2m0QC+X7Ryc/8UcbUwjwsY6AAR7IYfr6zEKqtCAzK
p6JHdCuOMvrk+3vazBtVBhGpRVj4IZQC3GIcdVv+PZyItTOJF+A7PfTNb5uhpnFP
EwpO+CtqY+xgQkX+b2Mf9nfH2yTITs/irh/qyUy+WjL74kOEj4MX1U8oVC84OJO3
94BwKStVsZWySfKUg3dV5m7fmUuuR93PocKVNoGv4Iv33Md+DjvJsp8iH8tiO1DQ
LyZBGfu1gPXx7Rk5/trRVdft68nhn7zB76TUY/gVU4Ea7B6W1KU0ePi1jLECpncj
VlQJLo5WOj1JxI9dv3lOtFgKYEqXgoNO2Ev1Vnx1QNfZaV39OJfqIiMLNRAQ/O9M
httbUsvwCy6pdaTnoApm5Hwl++h3jr77wi2vgjisNYECgfM7o//DzpTYDMJaiDPa
JiBZh/h/evFhcki5sd4vqkdvyt86E56fz9N87IBF4mwhr/iaeoboP4Wclo0exioK
gAi23X1pd3UodDwb7pg3vdEEf9J6g+YOg6flfhieoJDKaetsiMt1UKyG1kYiTmvu
wVD95QUQRQwTlWxNJvjDyD6JQHekDjpsJVGd91F8t4dNlsKNn+QvIGosrp30Dg+e
3ePOHdIT7PXUPvr89tO9yye4EDRtTbZ/Jyu5C6yJaZ4FuZX0Jv3R9GUS4md+DhXv
HJULo+jnpn/S3zA2GfX1U5WVP3DOLTGAripX7VUgsHa7IXEZuIWM/R/jZukKrLEJ
63u51KidjYyy9wqVkYtGF3+mlVJNqKddC6br0tPjlnN7VRfX1NXQGvp7sth4y3l4
kplFPn9Ccvwo4gN62Ds5DqrK2/vYxznfYh405LrzUCxjyOE++lHEn8cLImwVR8uW
ddwgdjQlpIj4S92pbJNMRv4rTNyisAj2QcbDPixBF2z83V9GLdjxL/J8hzDaL9Ld
PGNjyZpw2M/CLLWDx6o+yxMKoRB7fpfUaq1CqoT+4aUcIkhjF89E6E4+c4pm0B4V
+rtuRilQ2v/1JXK9lD4jR21KjErIVYAvmBgLF2IIsG1QctGsOt2Ck0dz1pEVO9Bl
2W0xReTe7FQ1W0w19QuP+sSrQOoIXHAKzAbFYnaaiAoLtYjToEsrYBNEEsWlrZBI
1kttC6onyKRqBex/JOUx+q7fIy3qjpf4NcbpGOUHrTzQM1GWDIlAsHLB0wzXjl46
arU0mV5DA82K7cyh6Up3sHnXsJX6csvV4esOR1b6Ilgvld8KYCaVFrbuBilGjsBZ
DTcG5b9/BJLy9G19OUWr52lkeVfhtq9a4XtcPBhs6HOg6eHvdyTC67EyO67RhbyS
EmoAhOGwq/x8OMsugswj+GTI7Nm3o2Wrxs2ut+mM0ujrUt7upMW/gbu66gHRDVel
Kci1GxtlRLEu7IGv2ec6i7htL73H7JYWgOJDbHCVvH5npprI4SeZLwWVoj7aADG+
q1RsD+0NhJecZ3VTskxphjwh5JqHPCl4VnFm6CRM93EwDlPbMUR3EbcOBHwu4VHC
jAIrI7xpL5gQFvgQqw604JEShwHrUxr/VAPkn39sIitK0UZ2rnFGtTlsO7ZxjkXE
ki4S4LnNUSt6K9cWhbxc4WWdV4qQAjASUujaFU1Yrc0eGKkjmd9EdIewE87pprpK
xgIEQYfSv6k2sNmyth5HSSdHxI2vLqtRgBS5TCcwtFC6FAlC9hkhcfjJczy+Re8J
5JDZX6Uvv9cVi95Gq1vY9haZiNOuKnqWrIsZ+WRjNzuiMzRfDPHXHtreeEzfd3iq
OJOVLAlFmwJH5LWBgWdXucQYwZamzVDd0gqduhl++96cwMtBNSsv3ANuaDqVWv8u
uw70Lb2453czEII3C5Wr2aJPmx7+2j3l+f3gWNV6wto9IsonWhFUsOR5+R/W+iLq
7n9PT89KKFWX1c9D5kEUQo8nNae9ct5yUsYLoNtC/TqE4Fnxho2VpF8V9ZSNDTBQ
G+2LqKKTkz+EJhAviLTs49iP48houpsskFEXV4GdxCvvB8jZ7ZPk4BlJnhFCust0
IgpD1UZHW2TBQ868l4vtrDtv1ClXx9xju0Kky+zO1EnPYdu5//LvZ8oiaVWGDPY8
3wYsuulnTBZorblyzo6HhhKq60aoJskroLIdK0z5xqDYJCaRT0fTWXdLbvSLHYDB
d+3LMsT0QubKrFvN2/zYdunlcbhQp9u3ibGE4e13HpvvzkZASdlMtfdKQf/vY5JJ
7y/7YQzEOqH48De9h/Dr+NtjJyMMsZxVgUJyb1Z0JqkLEgmABp/DkOQUfNwnT+Es
DQsAgwExLUGqsgPhJNv+E4NN1M4J5auUlDoDzDVExgkzWt0ekjsYIvpFL5RPQtGL
p5OxFbiWuTlAYXju1A/kqjLUl2TBNdPXjN4/dLvG6yAHqtVdtqN3Fm+NyBRr7MNb
D6VhKoBlv598rFwOq3CKYWLjjcwKf9Dov5m+JjUB6gjnu/J5Njc+Wjk3P+rLdqTX
Is1rW6mojVl64ZJFRglZ97ivoJzrx8e4EaO8RXv1dqOg5nWj7Mjv6IvJiaLZwWgu
rwiYJwsveTEJakQZG7anVoEjMmfqYZJoUPh59oPPCo7m5DbrIpbBFjBqx+Ka8CRs
WPeTQQW0FBRRbZLpTk+U1mPZhwNnMvwBBAfh2XFHJr6SeGrV0SScWIY3PcbW8lxy
nmJ0t/Af1CxpGPp/rx1ptXOpEz4u90XE0QCcGLRWnT5aMhfmGs5SKzoJ8c0/Dhyz
AA7wIjLa4FsPQusHrewo0xSMuR7qfCZdb8o0rDG+c5oWU2JQYbexGFKvIOPjicoi
mmkf74iMl8/QOnt2tGd41hNS4zDjQaWlzZFQoglub42jJ9XAShIb/CHX9C1SKQp7
04UWXs/FLrg7ONy8Afcxq3InGM9LEILmVzEVziumdJ+wM0WGqMh7vQYSxPcgzWyO
L+97jPFM2Du0aIcIsO0kEKlVRG/7PIEkytfhL3BW0xyXVaeuAj4VDHN6wWyYWQfb
ETmDORVprOcao7pVgqG0NR7E2c4hHvculZOQPB/85y5gQOk4H+08RSF1Aj30zwIu
9Oxtm221hl6pfPssPzxIjMdRf1dKEdEAS+XDHH1GtezXUD3TbomTtiMSbQF4b5Up
zdUdEXXE7hZCa4Yu0PaxNd5fwlEphOCHVpuUQHcDKkD7ulOHf716iLJacEiGa7cY
tjPsM4YN3BC6d5aOkZsrpK1ORQPTetWEvvsE67WHpDBWhab2Jei8nu4/Hx9enrAe
75kuqznXXBPZo7rtmqqvi28i7/BAGgdXW1u0YNVVG3+Hd2hvS8om+8BxKUYR+Ca9
XIvJ+zivWjT9JVdfgrfIlZftVjVp/pweqM8rzsZTnoBKPUyDlGBEiYDjdjxMfnFZ
S36PPKKHosKVzQMcB5bsRszryFThbyPwiny+3NQVM5ecDOMOp+Fmt9g1joQNjIsE
2+HKhCewUD92UhL/wlB+j+ICzBq4c59JvmOvu7jf9CTeTMKGVQrdLfNEyOxtRzLP
LVHYbLG9v0L8poQMFzuIwSBZybFx8JObycAjkziVo6MN7mCvPOFGvwn+OrLArG8W
pLCFJITP3zuVt0hy3i4cmxPirAyYLw7Rgrcj/AhHAss4lQIeq7r+5r0MOzD2BcDl
vcyVd4sc5+bjoFdTASZFf5Wg3D64bLxWKP0Rg7fyknKi3r3eN3aMVovW8y1cmRom
MY9Q44wAh3krFFI2K5+M6VZ6UfXfL5f+4IgvE2lWMoMOawyRcs0luqBvBBWMtu8D
uWYuRh44/uIewQgEw9UVTOeb/JHZJZlN9byVFAz/Y3sNxevwHsWKW2VxwohS7UW3
rEzZPXn1zLesMTup5zQtESL6I0hydrWBZTPqu/33beefV8gqf81inkIFY8Qed7/b
ecltOO/9KqulRa5fFWu9+3r4kWCIJA8oIlFVKXKiP6Hy3H82Tc6XSAOknsc5mCzN
grAaOww+EN8V7+y6s7Rm9NDyzDUc+XiG3fqIgESKPZ9fRW+NV8OGFUtB0E3DLEQl
w4uD4ACVgVlCCgL3kjMp0FE2qdZq6QxiMktvUQRYt/6C7XUZXS9A89gOJOgvrySI
zw8xQ8KesaIHDgpJW0xiWAUXfdwLezVblIAeZ/FUi909wkPhpSL6UNfahvpgm+LM
C1hSuH3L7fjlw/LQZLtvGPmIcYK4yoJo1t8CWooQGrvMDaeSi8cJlxZ7F01/whEO
QBr0HMbxU3CaEyQvHgUUmXRbV244zgEpX7GHI7bNySJOMBXHkj2JCS+zzpikxzlU
hYJ0JziertziFcIhC5oa26nshDdhCCCS2u85z791soO69909SducyefcYmIRQ5cH
7xNhH51ZIEIuW51rILU8Lur9RahAuhcUQiuaIJuC+1oViDb4dvkFJpfVwH8MO6Jz
3ySNOMmWoz34rhcsBM6xnQj0BNznGcGoTv04GNPRKyTOonIw0dw9UQzjZYQn2OTJ
6/Y5SHOuq+KfIhlPm1+ZvxQsEvBygCpXdxAQSIVeevWlCp/oNavwubG6nBh6r7y5
2hrkiQV1wIKcSZyLOIyB2oHnwTBO6ezNFjuT6/UXHg2D9MnDNrQaWhWo20fImu0v
x2z93XNUpCUnPiwPtVcq00jyL2Fw3Py6nFVcv6Zk4hk4L55xr6QN/RsdL5JGY02I
GjdoODTwwIEG+NYVO+KMFQn05mb14duysYL/mWt43gxEytRvFNgvkHKCIOvjqKL5
ocNMt6CV/NLr9P+lPSxD35ejX0TDmzehkKPJH/M9KsEPLAP6BwMEHbctCE7Rxt0Q
LI40uFC+8lh/1eX+rYOyJ3k6nIv+laEOfB6dhMO6KDoGHGEXNL3Wb+ae5x3eZzm3
dpBPrOwmo5SmMnwqHD2FkLebat2BaZNj6hz3hzoSszIUxfusA4h9W5+GAtgkQ1lK
ErKxJdlLKwOwjrqHIOjw8EFKbNQNayHfacRf1dBDl7uGp5oe2KE0cu9tsEvxfsIC
Dwyujab5yGX8UFy6+09uz4gy8uhcyTD9kYskMwbomnJnFfVi7YPCjzRuC2kydDAc
MKbaZab81ONsji90vgYVWX/LYj2/DShZZLuy+DsTBxP6w0FTVkDXGsno929uB7Zw
wasEEwo2/kMzkJkRXws/bB34l6wIaZI/AZAZXMbTe7D8XUmJ0z1zKf7NkoHIo0gK
zwU9FV0FNW6eIFPpjViV4jqismv1k/T2NbfDQLx+cTzbf//aSI4zBcYWs17PMQgU
Q4GQ68bOQB84xYSEcxbcAz6K2ci7ki31kDJABQZIOJNzY4RzUp0RaO+6ka9tck6N
MyeMf3MTwUGsYA0KsvkBlUVWGE3yEsoztq2EnBrUH4wn9dYES2ENypDZUQ1n55bX
pE3xqr3zkmJ6Pd/nqxzCVjUxjJqaenOxuOmL1gqllUm5F1xfumAKVphrYapeAvPS
LYGOw2NE8t7O4UiX86Y6XqMVYyDnXiSUeaGjmirb+JxzqJq2AwsTy1P8cdVT5S6Y
d7wGK/HJqmMDvgII9R1Q3H3Na28mfT64Bn32y0Cmz7iNbejoQ5yWGm8kP+60NmjL
nx4Y7czD2awFfgVWUYVRpINcW4MFpyCbHxyBt7Osy33eYlRbt/u44CifQlGbFlZO
3RB8hylgdZ6TQZvo+XsgiiGge+CEYb2HVOJeCHCIPZ0aqvvcJd9kPAAzbop0IZAD
1YIgyu49GnAtGvuYJJtnbxJDuLMxns0t+VGPkDp2skmpWalSGjlTrIHcbXvGG8/d
6nLWJVQXVtBb3QK+y1O/Kh0oMhxT7GBlo2lN0FEiGnyqCJnZpKjmIcIRFgw9vIyC
5yONysjtLWOAzZyyRTIrE0hHpzUTA6jxBF22ztVa4ZV7ooIK2xWE5aGuIX7TF8Kx
Z0qmvP5lAEDwIGPt26THkjjQ+i0phx6hW+JNaEJOvxZaVRpgCvczHnks8lf9G4y8
v8UQyBcSzzGtDFBiKhRS29aDOfL27ofnynz8VGtwmCjyyXftSk+PaMU4ynYJi/mp
O7CNnp0L3LL8wQkdnCVBO6tQRonQioBeEH0SEwU9c2VmUtI/HOYue85k4Xh5POaH
WVSFS8t6fYyTBdZ938m3xnBmtdYZ24ruHtA5oz3v5R3wxpEKsQLKQsul2EXOr2/X
LeYdV2VTIEXoRVvtL4vucfIjio/aC7duTakVpIweRFRHapVEShjfmEHlpIXeM/Go
Gk+GriOIMhOTKs9UF9Ri6VCTSj1a+LVrZ0DN3tUWujOiiQbT5CSjoqVCk3JjBLz+
EyWORuEgGKEGfBzISLQ1/sqUgEGyzvvNkYpCeM2BFssYMo2r8c/JPSas6W+HUlgY
Ok1Ctc/+PGpFavdOBTBOl6ULdt4zVHwACnY2CTcU5S+Ab9dCptQNAbC6SIzdn7aG
kK7IkqyFqRn6CYwcWnDjMFhCnIx5HWY/s86RyPgRyJb4ytnNtrsPoIC0ZxjsC8Ea
6Q4WthjWbCzS61TLEG0NwPrFCGiHSRTEVhqnup6X8xPJM2oNCmbX66z1aVcas7Zo
jYx/xLuYw4mgkXeJFasLtDuLvOC8ZmHjft8qkQRtT3HWp4R1T7iHMYLWHLFAR5QI
QPMh9Kilcv0xScvKRnC0YmtX3a5+pF5S2DiWYizBklVhVKPSnc4RSx+8E6isOt2I
cyVSF4n/gnj1kT6qDrxOq1Za62rh1UrMe9wjvBfg6Dx4SXx5fi1oG7peW+t/AzVa
mNz91RlBCvi4w/xXdTDH2GOWrEBwHy33rdHTa27jZ+yKHDW4AezPocIfLRhTiHDE
6CTGjahgIZp5XmvvNHkw64Uf8L2HibZc2s6lsxzlZeOEuniri5od6kEXXTDNla0I
EjkeI3WeTDEH/VN2rcZ0OJc7S2llxfYtvBMpthWZww1kxKtKtQsnxeUf8xSXT8N6
xsJKihYkUs8OZyp7+eSTKNGTdtNl+Js6odbefQMqFPO7tZZg7isHRCSyZH5aWwSK
2/4l5sL+b8P8e5gTxNSyrX2yBKzUjdpluzH5I7dccVn8P5DaUteCntquxPo5ax3q
RETm1uXyXvvYojRjbMQ6KRc+cao7JkTN7YV2sJxpJD0/KM5xi8LpBCz2ozkQSqAp
FNUlejCwrxxVLZodgHHa5fbz0EhKtBMIiIH44ivBGVntbu+AY49lGyrNmXlsenVn
WaMKX8EqYHBErWX/SwWudUSq77qSCRsuV5w6nI0bCnV+guE405F7Z8dJZoyHLjnj
Xz1VegH1lRN53MXW1vQCa7lwJ/DJjQIt3W67ZBm2RxqAusFloQs6m24gHS9s24p0
lHNRkMxCLDZ+EU0lb2HUY0dHH0SbGU9rC9/fbK2KJQJXGXrJW+nkfp/2U7+1kUnP
LQZwmzBhfKaOz2H3dkb7Ya/3khpXoa9BO+WHgeHNiyJCXy09h9bgQM2KF1Izm0M0
jm85zqrtzSFj+eraKMbxIm9d15VPDoxPeJakWHzSKwFYC/FCxfm1zJNJ+dH3H63D
tSs9ACUMjVFVHR+i3czeOzhxYLnMSpGexwH+bna7zHIBjX31GF+c4nMoqJLfDEe9
fL16l8WVurFyjVYgyIz23LXj0wyspIlkMeRylzAd0X6BFRTwWc4SAMkoX7npsXbc
NCYzZo1Rme/xWDlijQU174HwdPDpvY4caGuhyENNF9PliH5iXLjuGZCExtyAOiY7
x/BdcA1nv4/0OHvCyDHkWjyDtPyMkYD3lQTrZSkS4H2q/NTjzS/pij6S8nLdnxTy
VjZ9grcNKnFGEcojJcL/MPo8nLop3w/0dNqcCLyHqI0MKd2XMSv5tiGmsiAJKawy
Xeh80EYWSuA+gsVlhvMK6gqFJ46dcujg/EfqDRfzEsdS2mOJSurlCs4lKUTi061b
jRrzrZjbOVDW0Gk68TBKLNNCJZ8y0VZmeTbliIy8JJ1aGAXZD/DENL6S0fNBKWE3
g8FfM+NlD+6a1UzWo9oIiK+m10sHabje/EUNdPnN9F+GQ4evgju1ImwQztAjiJsk
eQ6RAfLm0P/gU00aRqVTBb3r8N2db8MBlnr4OaiowYWNa9fABhg/8PVW9dKBUPdK
rSU35GUDCfZUSybeU1LEssAJGqKcD5PYAUJ/r6+egf9juT+//ZXm02QlzOCZiPkc
/loCgi8WYc/Q5skH4rXrEMKyZDUP+vO8SUJpjbYwQj5MaYOBUQHMC6d64o3gs2zg
nVCLtQxGQ4ODxbnOYCckrvjNRdjRBUwHvuq9t9jrhbD1AzQP23FzYDeV0z/O7RKm
2KhIuJDvYzIm+n6UXAxa4MI/QSx0ml5PFVcsvC5ZkPnM7LCzHoSN/zyfu2kV1VN9
/Wi14IrXwKDIi7qykWxVhkMp8JKNxAUwAHu4jSB8uMQylyRUd9anuTU3YWYxsGpI
uqCh/Zsm6CSB5yFFvUVXCupbThznA3XFdlUfHDl/dh6OUJtwTrf4yzz1s6QXZBd0
ad7i5uKCPKE67ajjiXeQS/9x7TdbI8DKNh+9k82inarPRJCPuLBWrcedO6wT010i
TyKs/jMA7CjLKoEznQaSXGib97rbQheoEEAPCvYSesK73gE/n8J5797cnO9uhFO7
nMj1vs8DOopJsEFs9GMzjm72uBBldE9tV7tyUvvsl5N9UexnHJqU6rJNbuqMmzDc
F3DZFFHcptpc7MDPSNIDksfHXMfm6oEdFrrKCxbmqkFUQL1GRhNJ7HvmyD+UPiyh
Czs5rgf/s5XidLo/9Pfs+/TKfFL1mkuLY+0AWXdk9eHLHL3i7SwEVrH0vxhaKUG3
s9tsIQ3TZyPT+BMdJ/LfqyeqSi/CKst3wT48QxUYOr+KNBMLzaw1hDjSopgBS1nz
a4waym7MOAE+VVj2jPBAKzriaoB/AGblbpzOKm0E0Rjc9Cir40I2sA+yiz5yTVSt
oGUjTUJlh6dXrorJv+y6ytICJhA9d+8bAnma0rgQli26x1txK8AD7neYSebkqpkU
f4viAq8kidM1dsArdf2pA1dndqTAG7mIyBxuZmUrZxrXbI1Xom9DElPtspHYynfS
jMCaCsK6NSWyAYIqUlQ9cTt5XVZzyvWk+2BQCHfWHkUean/fjEd6CdHH4A7GX7EJ
soCjVNoCTsKRBoJoMxpmhwT0we5zaAMsAQ0zOseS6FAFSSyCOD876TeP7pwjA4k/
Ib1454YtGyVDDbqZVBXsmm9Ud406IoHetQtwRTF7GIfg0R+HiTQN2RW5y21iCo/a
vwnvL1f3tGLAvfAHOIBtpbH/ox4yQGTVJ6SI06CAhAk5zA50cMiVXkXAMvU4il1N
el6Kc/diYWxXHsnj8FbkpTJbosK7pCPvsG94Uf9PAtU8niJrLkmwtQVoSfuz1Brs
LlkZ4WnimtnnbaGNVoDZip4e4/R3rlSc+KmmKZxUA1S7pTIZnUmx2GM9Y3sYknpw
Tanw5QsNZaSXOmaNcqpwrn/SmZH7uG5SpjPGizV1RwviSe5ZK34TCWwTld7kgr41
G3GwxotQyT5o8LINIeqfo+RoTXvc9VAnXSQ2+QsS8KAt94aA3uDl3y/Rdps8Rn9b
V9gC2rodsO+FJzwvDh+PLcfUzFMQ7z9+NkWUJs8LZP7YUoQRYVrn2e3h0FPyyXQ0
wdzwRNVkSw+/dfcrqqCGFZz/XlXyo0HVz0jJXuWRZDnBEsYoRu68uXM8jbk3maWz
OtHXhC6FlMBYnY7PWL9VPhxsHvWXMmxRQQpSyF6KHxcC+O427hMpi25CMHr0UwUc
tNMn3RRoZqAg9JVh9pFDgc7cWfDNr5Jxz8EDeKKlmvpEi9DpIbOBxARhuTxQT0Py
FgNnw3L+2ViVmdetdbbXNiWfhm9Q4Top21p0q8XsLdo2HOEHMEFsV9RJutwxqJc5
zGJB1sDtpx4HBLXm6j8oQ6a7LCV4f2ZG8n4LHFY23lraz+QHAIVaWjqxv6m8yxTd
bnTySnFMdCMWKkQWtv1A/TdVZ26WByf4dOAWKokzNOED6x4LYvvJN/HGIEM/mTm5
tLXmMKdk1ok3+QKYyiQ+w+wUxmny4BTIiy7/pSdTinBnlSaCkI2ttlGSNP88IfmD
lRIK5H+IXhxMZONV27aYkjetf6X91SLNP67HZ/vzPQGbGcEX7I5DGqyEIGnVwjV8
QI94mCq1Pyx8BC3gMcvYcYjCLdL6howBDkUeYLnX3LY8ZfSoFeGLOKcGEkjnIZoH
XEjSQU51jqusNPbgKzOCTCAR9yImMH4qHarQioC/u/Kk9duY1vXsz+RCXPd10XCX
59dQvcxtam5oNGwFbgYJn/meOFgIFuom0jeiUZDM3+05feJquol9fmj9B2cfReMV
B2yg0392MQoeDXaS035VCAF45lx8gfyjn79cmYwbhu/OFc7FUz4+Mmkm+JkP07VZ
pEPLTVPPTW2lmYrP5NxM5fF2l3Tzg8ZPBLVNqErswMegTa0f72d/vbcwnp3wODCC
zTAJXz0rOHdNTOmQsg3872XHQQUctTfHeBUEO6C6D+Yre8eL/W4ZSU/fQnNCQAgR
+LnGL2yIUN0NeJz/Pbl4TJaYax0svJGJHturBpIbTOrFn3US5gO4dE/ZMDdKMFao
PgsKgvmDEr3rc8Kyl+uq3OpaL8kygH7E7G81ct762M4UhvMndadS8m0B6j1tTJTf
wERiLSLlU6DPUENWzieuT64AHVQqH6+mFOvShpvWQ6I3H4tokrGIyn9WFj+2rcTv
UXcFdvdFcuDOmGxys4dWdf5LkcAuvupCArjNVbkhD7NcFKU8ng0cfDMlvQLe0VgC
JrSFuFVuHlqpl0DJtsGpqCHktShcgcXbZV+CtfCSjbCbBYZ0e4EX7xgrM/8HUcmR
ursvuHSekQ3qp3+sZFVpuXMPo1gL+/3cBfCVax4eeHCD+IVlJrmheuwPeCFXOS4X
7nXUntJOmnaAJh+C9Q9uS+MNxv4xr68DRTym+IL/VsTwD15qqNFrPkE1nkyLdSfz
R0UCKmjUr7+JBz24GpgV0e+tEDlR0q4qWH6M8G/U49b29Tp461bMrUyF1CECwF5H
tThGhnMco3SxxZ9Hx/26NzwlrKnEyzGLlzVFQMR2iXimZN0renXYcKFYmHpVKI3+
Ly1B+fHsQIsdBj89YYCpwsOjAtkFNkM+V3YiPcrpToGzj78eQu9+eopz1HBjVq/5
FQ4L48ekNU6+k0qR7glvOffy+7wW4VB8HM8Z86PRkc1AzU6Hr99LUrofppERCCbk
Mmo7bztNWFaNTAuVR6qvFTJACgDLIf/Zc9QiN2Ui9FM7auhfspryRViJ5Vah5JWC
FwYeqhNmsAjWH8ImuWktlHb1FbsY5P6KGijNy+z/cx+70nSY2S8Kkne4fOV7IWnF
u3accBJvka21ubdKlpzOuCDkwl6bwETPPsIIfIHFx8M6oXjWeuUJfe3VkJqu4NTs
/lprwGhPFpK5ezy4nQBwDq5uhymHqRNbfyzb+13AAfWjqokIe6GRgVY1BH52Jo/4
HZR/9sjK4JHZ9ffHtghN0VPOtfsMMs60hFEkp9XSgJ0V/fAJxeEz6C759MGn/eV3
k2Co7fCmAdQhCnhjkKRd0unMLWNFafNs4joA0oeMzDVIxi9qnFMkZHWEropTAB+l
v3+pFD3/cVhClL62cxpu/UUqeSX1ilEoWgsN9oIpqbvDTzkuGVqE9Nt6nqfDYPd9
mN1IWHd8KHx1RoLlxK8yIKSl4VdOwT1nCVh5TPeto92pK07nniI28nNAoKIKZb5O
HCexYzYmOg0r3W0fD63kYvesZXy0qRxW++0GnHMj9w9odIarIaJzStr5daPyQ04u
lynv4B/AqyDqEFx9WA4pB21ASMAvlGJJEp2dyj5B8JiE1VW+q0NwG5M2O5mZF18M
9EVg8PkwP6drJRrCplWjX55e39hlI2Wyern9nbQjpLJ+oI1ATCgXfJHDSMgAd7JH
70U505Ua189Ld8FjboRbqkhV9rpwx73rJLf1eKlMvozKR2LiAoId0TmGbh1U+610
FLWjqkK9ugXBNDvnuN9/oR1+b6gOpxZdG6TQ4ghX11bP8u4cfcqX0xlVcbTRrOzp
GBOXpvtOrbEKVyJbymxhOzk2w+fbUkb1xvt0AlPzjMxFbNQe3FPrT6m3GDXcy1XK
cqosOQBB+e93+eSo4ftx1Ku9LbghZ2AQSfluKSrhy/4KbQ3/SrxSNutEChdsC950
PMwh5vOcPMBbvZgIZu6lJde18U16Tymb68hktN37XCMClSIuSl1mrSLsS89bcwKX
PiX5Jc8LVjnLFtO/LSgjQYIFlK79CDL6gCaC7z1zb0dRoC4zJCAOH6OlMqU0RvMH
cVW9y8t3jbN/o1XLhKh6FRm5J+fxIFSew/SPNLT5CwH4BPO999rN1C9kLiaLDDgM
hiQZSfkWYrbwaHPNWnXjectHjdG0AmcZFP4X3xysz9FUhbOeLmJwW5VjaGOjhF87
tJnkvvrnW1bissltrUEZmFkIzBBdSSVN5m6xxSzYmFVBqK/ZI2eVB6Pq5myIVK7A
qAWn5XAxudy/p7aUbCoiS5GdoCUP/wDMw3RG1ONrg3myVgyaPu5XQobwXJVpfNL1
iZwsldhiud0Ot5meWhc5LPK7yfMCsbopRMZ4OongiWzaA8NCHENJ57pEMjJeVqb5
2yBLGmedMv/tPmGBJJX1eajVpaGkcRp6jonqmdrzttcgxIXNboeWq0y7jgu5PSYy
pUrLhno/Fzz9CTlcjIzPYJlOr9JOLxBicyZi2EYjklCVcagcyBQkNeRDNijLkED2
KZ4Ccue/X1GtXzlAwNdUnEfPqYKIjK5SAXk1YzNECkD9wkQVgoKXTjqOq+tpPUUG
FpB8iUaUQPGJgtc7s9ajEVtwwrjmztkIs0fKVnLNw2iPxa/Am+dP0UuMftOxHYtS
llDfBk1nlLqAIjE69xl9jHO8nUrp/AmyagaA40KELLUhrRDTpB37d5bws9IGrzhB
SzLgnfiOsC+KopnoMImDeOxn32gFTSpPbpeqetw2a40WRPogmqqhDaIL15Q0MD1m
bRV6LdfTpP6zZPet1inNcINnE4GnFJ6ZAOLaHXplEYXzNUAg9tJHIrp/K99JgIqq
CaJdXAMKWSBH0OdQLM3fjEZVYreP4AcH0+Q6SmLWV7TtWWVD6L5BjMQNdtW2c69A
onSJF9+lImWNJkU78ld4TYUTsG4qNUJs2hXNl9czQpPtDdfKijSmZreFBDzZLQ9J
d3nB/dDaJOL1sPRK45FMve6kVdUK6iECZetxe4UqxC/IcVFVNALKg3MgKyCA5ae8
Pa2JQQ1Vhtpb9GVtnTvjzA0aKQQSHw1RdYO3tdxvyG3wmrOzky//+b1QYvcci2l5
n520d5vH1NjLZeGor20iVfTUTSJ8y3IBjs2kIX+CF7nzafYXq7P59ZtpcwMK8awb
iO0br7aHf+fi6P7SLOWAVfmxYrj/5tlG4Fw+4actfda7od9E5eWIA6vIfPvj9IP0
Dody8NPDrBrMPO1z0uldBy0VR62maV5PTnGUCrz9+1tNzPuMRW1x+ImTqIwNJCc9
RKyD5VqCIF0ER/Fgdm8C5qx2KoTmS36JsOq1RsHnsgk6y3fYLikb+zRYtA3I2Vrq
cCDA8qJUw+fL1Jr6ARIAX31bJqRd1+rZL1uzk+SpQYKJYHLlXFYRrbE/tiGJI/x6
hZh/O6S7bXWNRHXVp7dUzI15xFnsRdqMdrDV/vykfF0BkwVJUMjGx1nUHfyt5SB6
qefGKg0S6nMHWl/pBkOclWMVl4iEYK3m5SfpY14MTGIbVN2zGlLIghV80fHMg6Ks
A8Dl0AhoqgqPBG3p7CRhHcDuyR9owiqceRwMLABVHucyRUDgv+8mTNmVdxBOeLOG
bQ0hCs7DhZwrKFpXtl7zfedV8JWfZPm4nPL6AdhJ+dJnsbh/KDoHLaXWYprbdeLW
JsuHzXg8RsZ9hBFDvIZIW4heNHGVLtv+FeOhqTcbX+bZbKUkhHTItlEo6J7wwREt
n0o/Mzkw8AmecKhTXGfPeV5unB0amLKwlas5bkhRsCJtCa1ohKQ8XLjmWi62nAUE
tsF5lknei1d+UKSm+PEqt0mfYldWtWmnda47reO2z1+LZKHb4lyY+W4ZRdI+72kv
o3mGawIqooUoe76pw2CJOv6MwP+u8nDZUAVEEVnApgYA4IRTTJNPJzVX1iAWRn9c
k3WyxdfWPSrKxRPiNpn7X/LryG/lzKd6mPlH5bOw+ze982WSjHeduaLWsfK12XoS
GzehQpVmp5hFzBa7WHBmlvfPSknciiQ12d9O4mVVAGz3WIQPTMUZHzpqBfcGg5CU
moGQpEWF+Hp1/u3Kyy6VWEYhLQRrOorwKMkh0pNzocmDLb/0Ft1hJcqpl2GUQ+yf
Jfq5GpdvHXSIcsbJx8B16SwCZMmTAlS+3cv8vbK+UOSfERzuxDbld7/C7np8xEHD
Vuc7CvDJ8NGFcEhb8IQoHJc2XfWZicDvTvbhwWapS7RSZBgSHK2fsrwe9pkzDtHd
Bt80H5xg2F5RpZCnX1trpxtfFzBOZ+eR7Ytvhgz1T8NRofDct0dQivXxENM5zIlQ
wNI4jc0nEY6PTLnFuzqp6c5AZd9fasb2dzpJAZyyxBd7Lb3qsADcAvmgZW9XsutQ
9UmG6uDgoZZL4HF/A173eDkBBWJFbiNlh7MlMiHpjPI3Vg8hq5IyqXD20psj6pv7
5SZZOjRX4EQH5+XXRE27fCkAdugP0Xb76TQdYbRaayDgrtOQkwrYwHU/bTkiPvk/
2ieGZI6mNDoFRjnYPvileOy3AOdVHCU1KHuCrq0vF142LePZjwjso4AGkYj1V1dW
yNCmT/wEC8EvpjGqxBaSQDduadPZDHPyEMWtXADR7jEC1Z392JwlGnlHfQpRc55C
9HYGY8TAqRInAzzOq0KFEuu9DzFj1dzAmqbY1a3T6q98GgKQHGNyaIBo2DpA9qtj
rSWWdX9ojWCqhn5WX87JZk30rfXI9VryCoUPC647fip3PJtuDNLv0O0tBioIb7np
+N3dUHjB5RCvyqn6sNfUQz7U9MZckUO+GdRMMSZn8vrbFaU6y83YN1JlDFtHWtoX
Ki+aJZ827PMHBzI/njRnmd1xhtjyA5Romv9mvkr6+qcNmSW5DKdhYaG860il9UZt
L0bZF5BsDg7R+3KS+4r0Zk7dxo0V6kgN5va9rxuSGbLCj0ruZuUGlxtGwqbktRwr
pMROwzPWU99ck7jUEFIlprKCtEdZcdO4pDYEqvLZwnEhcPHDD16IhVOaC2i7/yfH
UUgah7l3arq4YOu/ehu0Xuz7KlPzzbw9KT68Uw7gTDxF5n7v+YxmBz4bhOHT5bET
Z2e8i0BcmHMa/cfgyVJ1iiIaBGHcvrooMJdcPXxylXjclPjSAK2cJPlG8q1TfCUl
gAFWBhDDES3vXd6POwJ64bhHLUDg+KmPmkVwUiShE7h+K6EVjEMf4q5KpCQZSfid
G1goc/OpE78kSTDx4eQm9X9HiJzWAgGRk6yzvPJGmKmgF5a3OQo7ACIpqeSQ0Fs3
6ARPxjorqn2dUSwMgcsm42/6Fd5VS6rKlvWnojs5LUBrjLMN8KCTzzSaaE5c0tXa
6cF6W8G2yqwhwI7v7q5r0blFbuJRqqVPWgbIV45dieu7WwkaTfxQjmRqJmb38uFh
WIzQDYU8wF4NVo7x8xJYcfKXtCRO+HBuO9EhZyvWtOPgAOVS7c9yUH/BCDDz66XP
ryulz6pMkeZ1vTt0dyRj10zoGFMMiovBgFuGkv0aysaLNAk5kJfGRLe+mVmrGMQL
D1KCy22BuKtBmRBqlUwvX34vJAHDsoTSsLnkL1FBOwK+vY8lc3tES4/wWwlMmAPV
VI1NQ4iRnym0XTzrZHMMPvJK2wi2mPdIWu4qPhJ9VRZPIQS4Gm/LcUQTgMfflScB
/lP+3ncDx6CwgyrjBV+RdS2oSlbbmMCdv9pbFHL3PMGuRAORYrba0ruRFvMA/zLP
v9shVIu1XIkQYbfp+6JwJ4EoexUBgS2bWB1DLrKJOaYbGnqjqZNkhZlAto3Pt7Z1
REUZN9j9M+BdlMAXrs+KZSML2qGLnVJbJcvvP9eZxMGsHib2YWoek8lI/t5IW3nr
LAlYznTXjVgtgZ+XqoV36r9EjiaXEoydcfpBtz5SYta2UCwLxK/LCsKizfK4bHmr
Bq2U1QvsZEtek/jet994WPVDKF+NuNeRUmOv6KlkYieyd1LFIKsKbq656kBnqmTA
D7DlmT3Xi1fCrK2TQlg4oDA8oT23cKfDU50GICYDGbDIKBe2YNeyde/EPrTli1JR
npc1meLAOodJ4u6Yd4Lbcm0ftbO+FZ/TwXoBm60RfHWDbQ8/GZbLJnaWJd1mNkqV
fmVMUTdsuhU39crlbrl5YWd4o/6BVsXYRYQvBqxZu3fcsbO+3p7GjYcjcWcMpPlF
mz28lC14HHTvmkf99n0R0ZH1bIPJ2/v0tKVXJFgIgOf8yP67wPmLTnV3+QzaT54+
LKnZI9xZ6rSNdqOx7piIABagpou/ALPFjPu/+iJ5acBzQOkHv0bn59S11nHoWLZL
dlIjtb4WKHR7kis5qreEagXvzmV1QSFyo5D0rI1MjJ2+ZPUsII2TLOa3TX8XoMkq
/ZSuGis4SdakPtS9IgnabThYTTq18yhRISNa3SzkmX2SpukhswEi1BKJrrjmgQBd
ht5f5If7FKHJQXlRz8Ginrb6Y8SwNqWDfiJtMQM3jFagr1qQTMUmQgUWFtlXbZep
5VnbSM8BzUii6FRVFHoJpw==
`protect end_protected