`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
ddtXksX2+yylW5zu6QL2Lhnb2d1sD00763mmSITNX595NcHTEkwn0zB1Dry37fOW
FufOhVzEJp80NC5qZ/+F0Vk7Ik02dIR0elf3clrjeJRK85K4e3Hoo4xn7YbFUIms
l/8VZSb14+JVGURjfswrIyCUotIzlzVYZ6gzoZwDXIi5gQIBf/gI+KxNXPaKV+PQ
Ufys/12rjO6aI/pPlqSm0hCvftmBcnezN2hk1UeXgOIuKZnogjOsf0iJVX2aOOWE
6pD/psybjbnsNB6kH5uFTA5frkzIzkzl5d9+YDm9OyC+k84E83I/7/j+rk4L2dah
QJOvksSIzN867/4Qt8qYTQ==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="MvBXkzurAa5VTw+1JJ70nePUfoQXBvZOku/SMmg4TwQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
oRtzZL4VJ4iwysPsC8SXYCzXS8Fw2gtZTOskLcDV+1B9Nzn1zTyNtlo6lNICRmmK
ZRVu2BmCc2G+fmzynYlNTnSa7C0Cuel6FYpxCBlOuk3OF2tzAmLAuDyOH3Z1Yjzk
a0aHuoCdIRKv7BrZCdALt03JeUmXKPdOmIlkVGFl8yw=
`protect rights_digest_method = "sha256"
`protect end_toolblock="Jn9CQpRhJt4rnzZPRk+dOpzAubz7omckX1MrFd4p81o="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 3504 )
`protect data_block
gD6l00tciPUa6pDNTk/+t0OO0nC/UTtBwLB41d4inuAUA3i/ALrNyoJVcBnAmEQW
ptbcNp5fxEUJjnOxnedyZEuEBxWRieZFQnkRdF269oMixu/P52yZUmVnpAzflxBK
Vqw7DmdG+RlJk1dZuLsYmJhACmTPJ43aZ2kecylBA1wC2wlTkhT968n1LFtrpMpl
jt/p4C3ZWLAn2t2zGT6pplthnl1tvufe9fNRQK/xPYKbBb1Jd4F5gUxsBEBJ8Mmh
MrfsxUxgdWy2In8cc00aPZXXV7vqjTODu9+QYJLkNF31jJKwRLhZbphl4Ja3WjQg
1gUgupNKBz4azGluZ+S4SznRQ9MEo52Qg8RDz1/3Hn+PJo1AxKeW3vAs1bUhnxa4
kLoA8QftBvhhsYVZ5/CrwoNt/ouGWkrrw1vfV3HnnOtUszptND6Xg3D4Y5v2zJMB
qnM4smxcrY2ke79rVMUwOf0cr3EqP+4CJobAH2WZZgcNwOwlyUvbeKRvW3g9iXXN
PaKQbTniObX/5N9fcej28BWcaWsItuBb8l/+WP8arI9fWWwQXG1xMxgaFLXSLFmP
EhpBnwBR3/9p8diQJfAgSma4EWIl+SAk6Jk6MeE7PMIItAcOUbHjyWAvr78rCJIb
hnR+Jk0xtB8q1RJsHnKL7iaC8bLVBXPUy6z9kuw1pMd8YIwEgBgYa4SD0c5Z4Q0Q
mfK+Ml8Z/4+VxWYIWZ4LQG3VkmpBbevGjbOeq6gENaPXzTDe1Qflm4KyQIU3Le4l
d/9DbC29lDEvEihoSRwhCSyFRe1Wv9eLt0ez2q+mmsQynlb+JWEbFqsTcfqc/NGJ
Q5VW/+Sz//hh80g2IgaUTfxAkET/xn6t8XfEyDYXvlecCVzf6Owt/wkLLu6Q4JHK
wxK8JJgmt8MCRbmV0bGbuf3speCgTc49ddaiBDpDWAljA34t+O7iIoCrdEROISo0
vYEbRp+9SAjx6IHoi05LhkQq+eCM4mRdYh3+UqDAjm7kRS49bK/2CuUAxLib+ujK
488HSKkFOpK5KztLTIdJyIWwKKwb3qjx5ysi0ninYOlHhFyOMDG5ZVcHhnger5DZ
lWZSlfR4rryLTcsDQquAImiEMZCl6Oh/e2WzqHdFL8At8hnQDnoHsJIVUt7Cl8sb
ARZkIl4t0KLdgzgc94xpD+pSMwzuJQFukw+1G5+rLWtgV8N7njjVX0poZVcpaXUD
3HaV0XfUVeTRzFuiM9nra/Xj8PaBRtE6m6/jB4NREHBcsfg0/KGzcv9TXhAGH2Os
RTXqyUc6wN1hJybhrunMjph9HwdBsCLiRXBo4kHRFsi4Ju3sHtgFnux3hekZIPn3
o8DpMN7LeNtRqJfe00OnEbkU19MjSYmD4h7J7R/NkWH2l4RGE8U81LEQ9GE5s4ba
dlSXlk4obA/4vCxTLSm3GsxRjYUytxVn6LkGOnVCvaxV1GdKA6tNaMfwRvb5vRhl
+hqNyoo1o15x+9Fx51OJxs3CfnljsUal1U/hICc4SBR3LLHVKUoar5KkeHD19lKv
Ol0f8Cqv6iJQz7qqIqu0MblbP0bUBX+gSQ0OFNAQAMtYnXFWAXl0m9hK8XNy6Lb+
rIQvX2H1FGMhyLCAZu9y2rjyrRNkFuPILqbHXshisawhD0No77Mt9vhLlEJA8t48
BunggYUXQiAQv0H45iqI2SwHAP3e2q2cDhmM3o81EwMvZ0Mn0oZ1X1ncsxRluWfM
CXToIPwkGJeoFb9vhRCPG+YMrdN6O00Y3h1E2oIKYx5Jqdna30vf7hUD8jM1Erlg
xbiLJjjFcQBOCM6GN64JKY0+MJihF0Owo739kqnL9HCD8SN0FqGhgNXMb5vmiLOB
nRmptJ7Q1vfMvze+lz7hnaSQdMrEl0G7tL5yToasZA/hNnyGdly5tEVLH5wR9GTW
kr2DxwQ3BVzUtjVXOfdgSy30kHPNBWt1W599RAzNoFiddPV6kX8IdiThd+Tp4coa
FzJYz3/HaQliUmwETKQRhZiNuw9GbOgmi0LwrXUIXBvmnfKYOWMBUtVn4jEtyK6Y
4Mmmzo420cpIfgAjPjh1/o+ZGk0FyOMoDlII4gTcmzt43uQ1bVNmRpSEfxWhSd7l
2OaTS68wHqB4scQNYYr2NH1wtJZJAEj/hhSwGJPZvXBfkovlUv68Yg10usQN/Dmp
BxVhaw4x/Lm6PX21gOY9pa7R99yjXNxkG20d3VDrHHUfW1S7VnGPuL36ubfCLN3l
TpPO0iqsIrKkeBpAE1Dki7jHViS6xxqCQJ/mPXnM7BuSv/zCDzy5++akrWtLi+rm
EK10BZEZll3CiwOZwdcjNdGU7i5vzFFTG91SRj4vwFg0klsPddqOoKswJGwXrNyB
jGd/WiAqIWLBJbto9joMtf34pd44BWLLrxMNK7J6cM0cLDojxLS0WqeJlEhys0gd
SoWET40a+AP5zr1/a9OuWPd09j+h0r/mmAIFyopDCfemhEn1sOr58vVc2LmYlScM
p3hovit0MzHJrGfd/+Mrb41iRbHlt3MUDs5JbVgPbempZQJgw+tFjrM1I0gZL+TF
EtFlgeee9kOrfmVVvXAtvaTpxef0oUO2Uf0PIi81vls/Xy+6cTbScE8DnJNpM3jF
knMB71tShFcgd1w+y6ndzl6BZ1O+98jvPXvXxBJbOrbVd55T+FioaF4wZfbSgh3Q
yN2IUoYKTTmqlGbsA0jQ75dg7vBTWiez7gNSVMbHHy3y/fKBQlcyq+8wB1dRGtYh
mSVZybZGahmJ85GG4NYUS8lwqdI/r7Ro4Px5/1ho8DNOUT0IKR/bqQ2zCqe3p2mK
cwmRGTupSvnkQbXWgC5c4LhU40j4BuDRpHBBzBJfTr6kkG5PoplVv0Ub6bdgJ2OB
EDjZebqHYImJf0ckU7GNOqMlaNd83PEmQzfTBJ96Rf4tcku4/VCPz1CpzzsdTufy
H8h5qpVhhIJ7dTUCbIK0ryZkIwkcnXH7vY6tuenD5lzd9gVk1nkJNTVaip4ky4Dk
ZBpZo9Ujo9VlUUMOqYGFsgE4WWr7tq6Zr1NMhAb+heILjjPDpYB1jAyOPx+vcKvR
JEArIj+R10kUpmlBb59K44n4evktvksIunBF/0LKimJWDw6m4SNMpNSmGWaesl/P
90tf87bGX+y1nTPxcuPBZ2vsmbzFR+eM8TgbGtdwMyvB5iv43NJPVFEeJW+nzjrB
Wrshv4SJ1pG743O0vXK5OszN9QsYmR2rt5hfzjZICXB6msqmnH4CY4erysbOuYpu
gfvh/g3eIpT/fhXRnSkcjGfj1Jxm8vJd4tf+VrJGGkDwDg+oZHr9ukUgShYQs3rB
DPORTMKgkyBDBffeWP14WAz67f6kB+3UU+gRcUO7abzrVKsoGQqswc3dUUtzeK6u
3uQmPx/IZtGUMlK1jQiPxtkAq8q/ZJoJ7JCKEusAkJ3qyZ0xPhrWKEaocA4heQ39
mQzeP2siMrgke0K2BOQ3opDUhz2DwB1RTusPVyjNN5b1DhBVbT9yW0uVqDgvUsmD
F5b05FkRQaFHT4muxrzIHmDwDke8Vr+HSreBo20ZX/HXOo8c/MJeuUopdepP7JtV
HeHh5tGxcEHGT8Cm026cleZUriTOe19kD3VL+y13v/8wKurQVztJYvI/xyertbb7
Hb0MNSDttCvqvUyMhSwjSEbhsrLnoMJVHkI0We7/a1S9QG01Iz5NpCG4eRWw1fTj
6OV+UNPT/u7QiegYGONjGMhi6GPpx9CqLRd5Un3hJrGIn+vQ0F9ck8jtSXPRjoDH
Rz4tHPuWiJYXadNWaxrZx8qUm95JU4MinJhM5V1KmIxrecJC8yb6ZCo6+Bk6PvKM
1XMMNvZqlAkC+GWlyCaAoBHH6tvxKJqVSQuYcv7JM3qu1dLPRUln0I3rZov16Byq
uns4GK0rYCNNWeqrC9rJ/ts8Km4TcKND5qs3fcWh+InMvrCNRIpMT7SKyGEdnyPQ
tItjO/GV1gYmi1EaCumjHWrsr8/ZHT14zLH/Da4r68gt3WLs8fxTZLyOAwOLpKoj
EkfnV/RSbzA1jxsSteSEf28i5O5WrEOkMp6Wmhy1z+zBEwWlxKEhkRueMs7dYbJg
Y0roeZqYxysJ6sCxzA6ZQQEU7h+eMoutQfuP5KZ4FpNvdOGewxAKaDlyKhHXa9pS
XzVTAwSOHg3GxGr7PFH8iWuM0JATnsyyQat+MHSWAHIFVNbKDFDJV+QKSg6svFP3
7z70rEfTWVIFAN0AAKskDFX/IlSgdbIwkFkz4jRVhEuvLnwsAZVXvFYuqF+RW7ab
Uyuces2KnCyW9nGLTHNwAMFh5KCyHzF/bPoRkNWM8ljjfHGKSBn42zT1bzw/NyT+
kX7POvs5nZZpss/Ey+7RLCBbbHDHZd3SIr5MQhMgNqlh6vQY0/z+3aDVh04OaJfr
zbT7//EWcsMH4i5FtJNzWxb3QBK6F5+th+eXlCeSkhlOkdqb/e22JpkL+MgM5sUk
XXQS7f70xMPEe0pXyOBzuAQ5kTvpkpxefC9REA87Klzp7Qy8QZzAuxq3yQehcBvc
KofL87ErRcEhZ1wA8K0ZsRRCeWHapLggcaxwzK9k2bhelHmt1IHeKwUDCNM2R7pv
9Rfx4kA4TXZ26Vig8Lcu3howUou6GjzAbevI/wgRy3laerhuuUis8ZYdtlvrem5Y
`protect end_protected