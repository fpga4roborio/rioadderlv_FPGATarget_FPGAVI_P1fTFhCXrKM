`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
ddtXksX2+yylW5zu6QL2Lhnb2d1sD00763mmSITNX595NcHTEkwn0zB1Dry37fOW
FufOhVzEJp80NC5qZ/+F0Vk7Ik02dIR0elf3clrjeJRK85K4e3Hoo4xn7YbFUIms
l/8VZSb14+JVGURjfswrIyCUotIzlzVYZ6gzoZwDXIi5gQIBf/gI+KxNXPaKV+PQ
Ufys/12rjO6aI/pPlqSm0hCvftmBcnezN2hk1UeXgOIuKZnogjOsf0iJVX2aOOWE
6pD/psybjbnsNB6kH5uFTA5frkzIzkzl5d9+YDm9OyC+k84E83I/7/j+rk4L2dah
QJOvksSIzN867/4Qt8qYTQ==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="MvBXkzurAa5VTw+1JJ70nePUfoQXBvZOku/SMmg4TwQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
oRtzZL4VJ4iwysPsC8SXYCzXS8Fw2gtZTOskLcDV+1B9Nzn1zTyNtlo6lNICRmmK
ZRVu2BmCc2G+fmzynYlNTnSa7C0Cuel6FYpxCBlOuk3OF2tzAmLAuDyOH3Z1Yjzk
a0aHuoCdIRKv7BrZCdALt03JeUmXKPdOmIlkVGFl8yw=
`protect rights_digest_method = "sha256"
`protect end_toolblock="Jn9CQpRhJt4rnzZPRk+dOpzAubz7omckX1MrFd4p81o="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 6400 )
`protect data_block
gD6l00tciPUa6pDNTk/+tzLxvdHE2s3DQL3/JqqujQBC/Ei+vcAB8wM3doqg5vTg
mdfn9XB1bLOis2CVSfu295W2DNwHfMSTc/8BhCDRnTlLIX0UCJs9Za0+LoM0rMrV
T7EjVWppbP+Em6PkVKCwlmIQ7JKaifJ+Y+kjw9HCGboYo5074hY+K/CBbfsBQY86
90kqG2i6SiqExdCqs6kOyyyAZyadRJXQa0IEjvum/e/m3/ycJl+JUddbEB8nt7q1
GEDpU0ZgF+E4i27gAaHN3bVktY9Ey7qxDN7RWnc03ia2+SyGdbwosBo530DXw/fw
/iEg+c03KsOPY668YGX92VdlpxalTw/jReeDzPyaOqZ53LGgau/83KGeWl5w5u2y
TvPjaYAbl2D96do/yZdiLjsPzXwCWkjISVrRQb9+7URzd/0SsSFCYQs64z3pAlo0
iEOleV4RZezhJk1RmYkUj/7TkD6PqFWZIk2KvtKCn8vwenAo80AntVpq3wAtdMi4
S0OQMFrJi0wTukwNH73TSvch0sy6AztsUMzPLsXUirg0jm0GzC0gBHHYwXNHHwa6
oiPJAVr9JkPqos7IZTyg0JLY5N7w2Ot92RLQjhw0r/Po2dRy50xC1NlPl4wRtToX
nl1bl1HhkjaAdVq3Rl5ozgsSCGTdcDBi9fLqbjw1UKOuap47VrTd1p6PImyAZEGp
lYuoU9a2U79jgTQm09nwwGJTo40CS5dohlBlo9CHz6mCp2rDsXc36gff/AMujhbW
QdM/OI08PpH0/Gy/EpFuuxOXgYzBhFuIQC5zDILFtA4TudoDV3NuIR6XIRAYxIRm
f6SmThbay/BPC8CHp1LlXPWP9gAJPPMA+y8vdrTW+Z0H5bAvud+r+/Lazv2gfYHG
tRKM0kAdsmrG3WwP+oi8Hc2atYEgudgL4C9mHcyIKjB2wCv7sidIIu4+78qsN4F+
STXgatpYM586zIQFcpbNO2aoeKwww6MolE6qgYZE1kVv0WC/WU1Qo3CbXMAOORT9
J6HWmW4vrsKQB9dJBVwPPvGtESk6WzS8DyoGFqSrIyo05LUzeYwc/8CBx1vTGAzC
GAMvuJyUnrIc6n+nQS8z4lqrkqnNpYlyXN2K7UY7inoKwd+05pN7pwkN8eI+zbXc
jGD4AJlZDz5kJhnzYbu4zDwOw4MX006eZ+48G2StxUs8IHzXYx5+DAtpb7h1ML7t
DGm8H+sAqEFDmPgwpOp0YioVC4PXgQZPy5SYzKG/St6PpbgVZXdk19FdQySHyIEe
JV+ppcI3B4mg/VDeM59oYJXapSifnO5lbS6dJDPM7GnEKm5+2t3Ni+EozaCGkqXF
kegCmO70dzJTdPj0Vxrf+PZNMOdq5qnu0pu+HMOAJYWQejk7svdQikWWrroiVfT1
KRJ60ZXJ9DKoiy1KWKVLvYPUJAn57Qa276jKbpL6Z0zCsAsK4HCWsC/GO4XclD8G
BJW378nUmLEdeIoGKPqL8EmNdySnuhdeh9ixMytZfEbbzHlcS0aCnHi4lOAZRKZA
bF/rzndDrWaLIZ0vhW03xZfnVZ1FmpgHbyh5q65EIunZlz+MhhYW618loNbo29xR
aZ3QcZHP5gZrH4y/RVsCmCG0/w9UA4/5xbkaQniuSVfk8Ig5A3mNsbjOg2MgAOSj
PYmiqKigpnEKI11aWEpHIY8FcUq07wywQ6HXEjsE1SaWmhckyUx4NdkGdi0ZJynB
KXPOdZkrQsUMXbZQsoQW2GOMRnrYvnORvH2INuncLWB1wXZJ8c1S6jpbnv+pNzSN
D12PO0ESjPM0a1dUpiDGQMfM26BfvKhzuWetT/vG3X2tTg0SdxzrygGHsZGwSw2B
Ibx9dAPtLSo4gql9lgBauucqXWJKWM79CW8L8LyaulhUbBFcrR2m1s0IT704QcCH
Akm6lHX9CFfOM//Hs0+4vVzRzcjAtAqEKfXctRsk+raec/FF9h0IM7GpGhNV5Dp0
eB4AAYjQZoA8KNAHlLM/ZVH63UY+SSvHXn+VlcAQsBic/UJE+W8FxeNVi6Jy0LPR
6BniHn3EJIhB8CdXg5zqF+wd/XYaw4bGFv5EHV23mRDB35ATRzVBH5JtYAH9vvoQ
wGZF+90tprzDB80TRNC3Op9aABiV/wFqZh5jd/XRWsPqLVMOxEEyf9jaLdF9wYwk
frAsA3C/USqUUIF9+KdRfYE6HSeTVq4bHyLO7HhILHzo/iFf7rBXoxSUltscOWMw
F4kk3VHPS7CyKtM78NkW+NouP1GQjfCxxAX0qyo6m/0+J1/EpZIoXsxfQK4b2ZKH
rQ5eeKSKv7rAC7iIXOoC++Kj51CFtAx5THvfWFHsIhyLKKjSmMqRwVKkVc2djz3z
dZb1etrfUczpikWnSzdYDoQKgsY9w+5DhkI32Q1Win9A+xzhZPWhSoB0y5aGRenC
LPclQK/5QCRsWlDjxrR0JXG0D1fPh01XwtUtVoh4DOKy23Co038LYdVYTn1PYtEu
qvzx517LCpmQgy6QC93Ui9sBM8pVZpa/1otXp4PPzqUHFELCVbnFiIBn9vbZ8ZoD
YoUIUmn2Uur2+GmDwjiTLPa34JIXecLdhwuoSl2DIZQ/Kwaf0ZjNk/3Y7yl2jkWm
6VhT6RkTxHw5ckHuTg04nAGc3LDXW8zx+K4VJZWSX7pyBr7WsA3AeyDxd+wvL0hz
s+94u9ioGnY/aV7dDvScEkYUO1pcf9Lx2N9+hhtSlfKwaxWaJHa3YsWfzYuU4xKS
ZIp6eGb31iUt0xiHyLth+WHBXR7eCdCsQI9SpfOc/LGQcVGix848Xt1CUKtfYDmS
UPA6jimXRkpMFKtU3yRxbRvU4rbQF7Ur37Cyx0vBqzsTWqT8eV8xKEsU7VrLJmwF
4gcNKRciLImWk5gL32/urXof7CABkRWm6vYinadIM7l2HV8AL4+WY2Nfj73ldkp0
luwK50sOGChxTKRWO62QObJfAnfCwHO9tehUCruYkAz/WVCsk3UY4euOgQUk8XRj
NeLkmvz4oBsbJ5+gB4n5XMcfJPyRWKgxTE54whG84HnQjeC2KFLUhxo6/+W+rCuH
/OKKP5S65/eJbrWTYw4OO9+uz3I66rqlsXM4w0LOUmXe7xhdmxGUIXz7FSBEMEHI
qZfsYOMOz3CnrWWDD/e0L3UMrj4xw/H2CMqz0ULm/HihgQDjgSiIbn/nYPz14yqS
vFihUl8ezQ2E8xzwySKBJtn07DIvlb7r0IBqkSdBhzrbqt6H6+f6JeLpzE/7Xjji
PliCfUp6+sAI9znTaEWowgYiskRKnbE/ozTKfIQVjvACyz4jAeA70TzhuccRxKyD
HItBTv4wewmfzM0VfyUKkdZcRwe99TohH7neTw3z3dld5e902bBH1OEyHK2bb+mw
nonXyMDtUsJoMEsZC9P31Mslk7cCT01lUr9n05cB/ypnm/0OfoVEzIPKrpr3IAW7
RQHthlSpvA7N1Bn4PTrplw+Fcf0ALA9Cfpy5odGliPauY3S+4xPw/LrttHEXiLBL
OJhe1aVt1k9uQEhukU0hyP5KOgbIxEAGm+uzeAgkTO1sIe7TQAtsHc5W5irF0Paw
3hmdH4yyiFFZ0mIBBCFC8w2CAwX1LQdkeOKI2QIt4Fh3blgx1AHjZOQ7T/7aCEOS
s1yPoBgeoh6HWlg4ydk+WARE8ofu+c2Rz9nfTHiOFo9IbdKOY8UJa0PzmHUBhS9d
AFPyaK9E07NzUH4UwpUCIzoNCZD8HxLVB+fOU0Dcn8D5JFQZArp0ItEgcZkTP/En
fQDcfnmEUbzOWe73z5YpqfRYvKdAzLx44QHkUaRMdIeO/1BWYk76kHnU30A8OH9v
6zE5h3eTNQ6sWSI5HsbN4YAVygpy2LaGudgs6iRTSJFOwxWr502ZhQRSRmvVEXYo
ryaFf9doAmMGkbWoCMTJSqTHwcPwcZYjii/PtNJI9RYUyIkvxWi1/dVFZIdK5Ei9
jEOWhbf0l3mn61pKr1/R6CCrtvp7srGVFCKLmTDWo/CTbDBgySEV6hifB70uvr2E
cBiQcvrkIhIkQsIUA/Sqd02BX849sIqUOA2fYqgtSbGGOUXooF7BGBYp8xMSG8s5
xxKQyUyCI2oEZtK+lDeawwG33wRZrFwR/mXwrd4NQZs79anANPMX64F2aef8trBn
0x3ZgrDjigjtgX/Lz2WrbqtM9NbXnvije7Mub0XVHrpjhOqpjNq6MKNbmbb+17+Y
ZDE5sX7Fp47hrnqn/tpvgwyKDTNLZDsmw4kPkBJnqUokSxQx5vXFjcdeQEURUpY7
vPoN79GXoKfecDNbAKgBiuT6xZu/TerEM7QpkHrNoosiao5Ihk0GEEhiupzFSerN
b5x+mG4rR+yRajMi90V30/JdeItooADserPy3Ychcr+0QzST+PSooaVNPwZ1wAOg
rzVfeNubl7iZYaXAL/IC2oiLDEn2nRHVen9HpZPm0gREl6ZFoIUJGg5eXbnVuHLl
UgqqWFiPqF33gZ2Bnfa7LkYg+Ihp4r+affgpg6l0ZHxwScF+GO/DY02J4zTmpnGg
aedIsO7XhC4ZPIzuAwUNeG4SxoXNC8mo/d3AY1WFFK8e9H5xdMcaij27Wmh47kJO
97Rbvitbqm0NIO/cYPzq6n32sHZ7w7NPndf4Utno2Z4/ewOIn9h4/nMiCjU9SZL6
UAJwIbUdKLEdLJ0nDY80Dbs5ugGRsk4im6VntK/Eqv7vcwdddYg1jDcSBihOw7BM
sPuwcMoCeFlT8mzdpL+2Plo6poL5zyCQkSyGJ2kgjYc0vRtwDaqB80XupLdQEBHB
mzs6hNK1hSAmHIVDDMopME62tKw4arXfrdke5/mUeAyNc5iuN3ZIwR7zLPICBg+I
Mm4q7eghNIRfDm0Uh9Ie5ZXVw5Vqch0vW7lCGx8Etj8X67Ay1LEEOruaaw2qZ983
C113uK1552qJrVpvDnsuoqzzeyFGRT5mb5bPVEHMhPjVqg+G3ROVSTXFOm1ItgyJ
0xsjgmcAPp961Xg/gXAzeZHw1FzxgJZYTTk9Ale6oeGqlnZxmZYOauQVI4gfin2M
evLIAehN0duyJD+QrkAv1PwJcsx7e0U7B6IhSxRD1b92xtB0l42IoR91OE65vmUh
eQCWuZP041yWDgoo3PYAX5eCDtm3fWwLGvyzpC+yCVJ3OAZB9Bd8IzKYo5yc8Q8T
cAIqfNkhh2tkqJ8gOfGDFp3AvmqJxDLi7JCg9L96v0PVSrpxAr0bgK5hJ++ZHnLb
e9Bku7JK+rXXpDw7AR/1/e2IOlQV21jZTwvk9JCNvHRuQ6gNNU/7nR4kLMoWQRDS
9KSoiCF8bkUxr/W3wja4wKmPRSjWG+4JhM+T/WfYek9HzyqLwTDlvk8l8KoIZMo8
+mdf1hsvvWUJ47DNPK9A4HyfjKlrXmekexvlZZgLVtEWVYp7UWULXCTj3k9t6kHl
rqj77aIC/X3AEyQbu5OQYgWrgQ31X0BKu+imRfLmGXkxeNGf0cWB3c2UgGTFgA6/
2GkjXbThMg0cj0jQ7xxVq7866vdUsguTDlBJq73hyOGEyMCrmDAkKOK9bSoOyntA
1WXdIk3Yk535v1DH/DY5o3x8WL9lIy2R+h/ZOGO8giKZKWowHaNx+y3QxNodSQSq
wWe6wbZMdODsTQCuVPT8eo2ehvvidgCV4zRZ+NMMzN/RoKkU1xhXWLumE4aXYKnU
uz1hrIesh04DdM+Kk6v6DgBg/HwQXtQV0oLs3btGJlj1Ao8VHobTv5oKR2Yw1qOi
RA2a6lE0SJ6vSW7+TwBxVhWF77hvD/8WN2jl/scLMLQPRN6DqaJPkt2W6MoRWzgs
A0uIpenYRvhalD5nrTU4qCD3oCkP5XScXkK3Fo27ijuJHDiEN7viS26FdPpf/2lJ
BZvKn9wyAIuN/Wi00W9PXzXXLVk3mPCz3VtNQBm4Jq6gsygvi8BTS8JnahJV8SOG
RDtpKzzXuYBlGxtucg6ujFWF1XFS55kWxEii/L6ZO6JFECRoHkoOoYnNwi0uTPgF
pFzrMmTheJ7JB1KAee9jWtLzTQhR2Az+SMGT1xc5nPqumyEnRwtdgRL07fFS0r+x
P9ZfWc8cgd+xOWL3U+LgabpHEmzeEmWUEXnMj3nDM0iHyFlV70AXkll7r0sl24Ds
nPrenc/Kb6+z/+ZZJ8LgtMGyZEhKuvo4oC59NG2CtXvhse51D8Zm9XP8bHiW+XtP
lV8Qk/X/q000zMMhkZijM4QuW2UwhZCUR0BBjU3UL3LzEn6aCqWGbroeECFnEdQL
JGgYvLNmb5MNoLuh97JocfBfTKrfwlOmVQ45+EhqatE7eubiSo3CZ+BaWc3S8nLx
vfOYZMkfbuOj80rlEsPpyqOYDRx5W25nmLcVG+9H6/t18SYQrkXuTeneSbWcsw/u
v6Exe59zEOAZKnZAtnAFF6vX5k3hxD6UNrWbhGI1aJewS6V4MUOm/iATs1gIemVw
zgSj5wqHsOhm3sUmVT0pNooRlLwqgmf5ZsQVZJ/J8cMHVzu0klnvzKBenNnxJqJ9
Oa7ZfsVUI5HeQ8fiu8gyA2czIzTyXjCSCYnw1wfbxOx9RZ35wvUnh0NP2YzS9Qek
4fz/VvOpshyl30zRGNrbCQVwZKxCoKLHbZdIimSown08OPbb4e82hiK9STP+EKpa
mXntxia0+dUpOLhsPw7Rzw+HafEGr579Uc/Kf/do6Y4Ha3KUL6J4s7nrguwxGcbD
arNNrBooRJLnhOvnppUAegDOxzE3RPKoEhChl/1hqWsvulbKMc6hPQ5qBqz9kcpO
OALZIItAjb2syWerSyuNs2QJhU0FGTRpmnPzRdTYfSnAm5n42mZ/RcZ49VAC3u3P
LLiPipmVlPKb5UI2tXS/dqiG3cEl0vcUJ2OSKBzupJYMfF317P7k6fyzPBuPjdfk
eYYWGrtpYgx0mxQARt6yB1kauxnZ3QQvr1ln64Y6n+B2+rWassHkBmJnXUebfV4B
2dY84YeLx31JoEr76bnos6+l/HV+1eISJJ9SBLHmX6rI3hKxdrxjkAEccK5b0tsC
en/I4T/m2PwMAyW7j4HIG5BG62cTLD6f9BGFE1X8uThoE71FV0VnRk5xj0WdJwAT
ao27FHvUO06Ug8VAXJo+SpPUxDCX+f2nCylCcVGzvArVuVvGiq4xQe8UfUI8z4ZD
1hSaQ4htZT9NphdpEkQ+WjSVQnrx05ikOJpOyLrUBMZdDNbkpfyZf7bZeEyW8m2P
SY7qRyRvzYNrVFFJLabr+XX8G+Tn4cvJRVPDqrtdzgnXq6EehwUcby6owGdl4UEH
ONnvCSt00kO7GUqKIgnoFDcU6xTaEbJaYPjaD6vz8V2tiYIr6NXMwdFTE5wbXQHa
pp0tfvrkA6sE9aEOlsqTtKU0mf2PYNIGz5GTTq5QbZwwa9FUI5jPh3/Cy4pK1uGC
otV2LJgzV32X8fBN8elJHN11StG7wrPtAbDP6tqfKVMoy0MddcPFqITnDRHsph8o
+U2h4OHJ1656tJ9G00H/IfJ4r13v7jpyV4xkrIHr1vohC3OR4ebc2+2dHciGdFap
gNsJAy4VXIBwxVl/luI+i5tAw19mz/zGEVJp+WZTQHFvArBpc4UZTSFECEmcEl2+
CsI8Fh2DaWMVes5moFV3+AqYtR0DPGTabk7qaobgqZXJK9g4UNPmtyELvB3uClmo
ko879tTqXXUQ+tmN4Thw11S2a+rOt4jYh7eFOEh/EP8vtYQtlMOU/ix+e4I3+UkE
Nming+r77Umw/30DrPy9OzQM1JYzfTHS/MPK8bK3txtJETVsXHLY5cneeZKGGjBL
SQWRf2T7tqyJE5P5VahNZONO2KLMpw2NA75ndadrYw7kQP2857swb8VAnO/Qext9
K0ikGu0DEINeY44p31ZIRw0AJT4XxThQHtMP2CFigjcAfCFr84bYryc1Xm9kJbw1
5zHVjys6qXj03/m29UaK1UjhCmkbXYXwQI8Osjfl5pHO0zOx7LEnxNzgyTj20Ce/
kjtgkxjApXtJ9Wo39pzSyn6hxVPFzYvZU/FX0YslknWDbJNsru7Gk03p8DgRr0sU
pyrUm5brw3H+k7AE492a9NXlQyEULn5yXlnMdP7Xdor527UDPkZlNhu8fVEpKuJD
5hgj4RSBHZ4q/Gumao5Rdaj29PtsHUFqjYO+7abwxMRFBFeMa4tOv5UDmY0rqAoD
CFXK7qvvwxqjEGqS45uydDjpnayW3urvH1hk3bisETzEGiOpnS5cI8dQXsV+zoMO
zrE6kIYwOD0u6lc68bU29n0imilrPD8bna/grsZsP/vdT+rIyrGJssqr+XXlfzDN
n12sNGGlKaGCZUAKia+9uTtpROtXu8UXgvSVos8J+w92P+DusG/r8VloQYcNq1Tl
mEqHzvyBehuW5UJu+lLiDRIJz+UDw5JxW6fzzyJ7dSs+G2m2haMwiOhlcTBJSMu7
m2HJkZ7Wwt352oiIJHNSXYiSzGwSsk4yZQN2Xc4Q+utmLY77tG03zSsT3jXURzvh
h+Ameq5MgUaeOOq0jSNMOQ==
`protect end_protected