`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
ddtXksX2+yylW5zu6QL2Lhnb2d1sD00763mmSITNX595NcHTEkwn0zB1Dry37fOW
FufOhVzEJp80NC5qZ/+F0Vk7Ik02dIR0elf3clrjeJRK85K4e3Hoo4xn7YbFUIms
l/8VZSb14+JVGURjfswrIyCUotIzlzVYZ6gzoZwDXIi5gQIBf/gI+KxNXPaKV+PQ
Ufys/12rjO6aI/pPlqSm0hCvftmBcnezN2hk1UeXgOIuKZnogjOsf0iJVX2aOOWE
6pD/psybjbnsNB6kH5uFTA5frkzIzkzl5d9+YDm9OyC+k84E83I/7/j+rk4L2dah
QJOvksSIzN867/4Qt8qYTQ==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="MvBXkzurAa5VTw+1JJ70nePUfoQXBvZOku/SMmg4TwQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
oRtzZL4VJ4iwysPsC8SXYCzXS8Fw2gtZTOskLcDV+1B9Nzn1zTyNtlo6lNICRmmK
ZRVu2BmCc2G+fmzynYlNTnSa7C0Cuel6FYpxCBlOuk3OF2tzAmLAuDyOH3Z1Yjzk
a0aHuoCdIRKv7BrZCdALt03JeUmXKPdOmIlkVGFl8yw=
`protect rights_digest_method = "sha256"
`protect end_toolblock="Jn9CQpRhJt4rnzZPRk+dOpzAubz7omckX1MrFd4p81o="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 37376 )
`protect data_block
gD6l00tciPUa6pDNTk/+t1gcgy1iCdpjTkA/bOvU9JA+cpFEv5u/7dp25hHk7lLT
6tYtR8HgwcLXTcx68BnPlzdPHkVIv0lwXo6yhFVkYlDWBcqD9ubowgKij0UjlXmV
p4anbpVt/gKvAYRDYe8Q5F2CQ8AIsxOuOcJ2vhCPchS4QF3n7+oG0MKU5ZyzxTu6
UFh2tOZ1UkjsCcDisYgJ0hj+N+AkaRyAd2uuv1L3cIXfBLvhAch4KcT9WdUgoxxW
Aqd2+wbPsg0kc1wT736ZJ0BjMQOgjXVpEuBr/hQ10JZzzsPEQ1iJul8x1b9BGtEp
x0FHtxnpf/zJmq9gjKOX62Pqrf3ZKOh/aeBxXvzsc0Qj6aOYgCRv3P0/K5hbLzul
cDic/f7QJevMNt9aNqTT6+6QzvUn5GwvnUXegxRXU06a9q0Srn4UIqzGOfzIGi1y
nr8bp6/tgy/Y61PV36njFylaq3o5qRWunEep5wX5D2W/enMMXBNHozXnkDjn0iY4
s4inHYt483Hy/Brgb0we12k4RYa1EScQD3jTB0zA3YkcKyHXpOBvsztdfdC4eRLv
TF0/c2TOKQU5RCaMPG+DMe8WNq8z9556nZdU1+llHbe4z0sJ16NoEI63LVv+9Q87
KUWkQ3dT+pJ43+hxH3XXvA6RlAUaYlX11FNICqMlyApHwVKL/jeW684kF4ffJxeY
BIpPcBsTzdvCpG3H8hOZlEbTFPWcsh21AWqnIBu2TQuqFAzKAnD8x1B6kgbZbnhx
iEIWr0R0LXtABRqEmUNjYS1esKfcOkJ4tANH8OvyuYY7zAfh98+yHcPe+kd/wk2M
wDLMvJkGlK3bvIPpv9xCsM3J1uE+rspuzzE3x4JultyoX5whGXUpD4wpAGnKl4vf
yDKHTOPHZsvHoSxRMPerjNUahI8tc+q6271YAOsl9UsAL+JZ8fsqQbVIVMwiRQqP
6HgQhjP589fwqP61MtF0WAUyJGyrJinrGc0qh5YJSkmj4qspXVrmQh+csoBiZ568
iOQKckydmK9KvI47+GtN1cX0s4L9s1uA4IyIzEB1Nd4nYpDo4Ps1px+02zeTL8Bl
ldw9OMuJRn2w2o6Oy7SYqSXUmTnwScsygVEHbi2z0vdJ0H8Zdhc0ED4UuOf9iHmg
YlYe8JVLOYok259GagXyVnptsyPP2nshpOeHpih7Cdjau/z/AKncUuLGaTRQqJBc
rDvStxf1tE0ZIWVKqQyaUuti79Lasl9TBXZ+bNH7LhEEp42cbGlQLNgiJbmzTjGm
Rw2JWRLNdscE/YmmDv4FFCnFtXUSA4h4eIbruOA8CqCpgGh/Uuc76g1uaHAAK0Db
TDx/uIEKnv3rV0UPNTposR7W/8yYuCl7a3ILtneJxgdlI4heSoOsHhkymBiQfd1R
R8Y1jdzLV+AU41d4qy58ITJKsNbJEG7/N200ZfvMZm9bCPj7NndpWqUfildutut+
/L9coWXWiPBFdWn0fiURowMpGLS7j/WhXuTbi7Z52GeOptDzgc3IiRxKOnOdq+p4
VZ7FrnZq1+k9oTzOx1loQqrKGRcO8xSiDfG3xCSs6Uc4a23nEWtYjxZKCdcwsd4d
cELHxFaOr4PTsiY8zFz23GaLk/AavtxkcxWL83iFKSV6PvDYR4xj47mxGQzzuVAJ
i2x6ClnPreNJNbBSgQwm0wBm7rh3eGx0VMFpWR7cL2DDxu5qYxjwN/DmZ1vkuPXp
RwtJ4mYWrV6nz33PjvHXTxuA5Yw5XCxtkaSDta7+NoyrisdGgPjccc/S60vsC45J
Y/E7nOIgGspmXvDBgztCaFZCnvqkkI0rdW3ofdQEYPWCtn2acukze+BTR+LafuBP
GWmpZE7mABn3OkQU8pkooGuQxBjKk5/mQJ682B3cosYyV782v1GOdsX7XFR4Fo5B
39IgiFWv52iY5R8WPoH866C3F5crfK+JFSZPNzlNZFZAwD31vxWGvPnrjMQ8ZdyY
oBS43UDDH4WE3CMF0ZKHMWKJp/+xOxky1CPC8y5plTu4RqHmLKMQVO6JGrgRwflV
AzkAviEIap9jD3tuzHkuxMZZU9ARmscPMx48aBld6chQW7jBsrcUUlpcpBTyCrry
A3oL3kxYnkNHSdgSF5EHh48SGU5XIfDMqqJApA/HgMnGoKQYhyhEx+Zdy20/BM7k
lR2AocZ2xqtaEkywv22tDmPR6iL9FW1Pq2dPYnzlGm5ckrhY58sBYEXVStDfhezF
76K9ayTki8qX/aWR/6ofBooI6kaxCMOWIAi9+JvdThDbZrmhYvyEYowMBRrIAGRL
jVL9DXuF4DpMJy36+GNt5ESkLUQQ2D0ymABI1Zc+iE2wQ/FnzKAofgSiFtGjMjd1
xiox8cB4IM41NLEK7yc/D5+wpcdOdudxf7mjOEgCbWefur2HHHedroIYQ/jLcifm
aoFiib5ew5jvmBC5wgMKJUak/0YtalozxU27j8AvVJEgB9MBR5+EF1cxkDCg6dsi
qr0OE+3+jeIoGjtXPze49d3rZgN80X3O2pEgyUhiS1sclOb5HlZoRnfdL2Znk2J2
uW8k4lB4fO/Fn8nXtOD8OXMWPU8C+vo4ELUUqclPiSN0kNymAXFr7infd8DtNtgt
dg4w/UHYxIGfb+VJ/9f+YHJASWsJaHyBw/Qt4e5v1XSZlpGLmEGWnlTjO7r2gzAz
OYhJ9GdNHXvOuflQ4oG4CxFikzaiIN1IfebQcxD4le9YLL24D8bvto2XiOfvM3PB
iEUgbrgIjKfBtQWz7DfMsVwjtlauNK7hPw4OmfQzRe0tNlBxrlEZ1lz4Z+OU06fw
GPr9HSTu5Ufei6OH5xohJkOnrxFS7tAE0Bd8oEk8dONq0ppVGsldD5ucL7RV2lzq
QMzTY+pnAFOugb9Oxs4i1Koj6UGFSsA572mE22NKS6FhbLfheu8cK6i2lATMmstP
j9b9C91k1mpNqGLt10bYAVpga0ygrgg+BhXjQLVUBhRuJzISPOZ2JwyCWksvjks/
RPRoi12oRaGlZ2u/CG8XIUHXFDkI24kaoqWttM7+72xcDvhqmRUWNfaVTsflRXoE
lLcdmnhBgzOlZlsOvY4ZU+xXoK/gd4Xvxsd4DkxeBIHRwkgExM4WwoAIm0U1jIQ4
ce4VJMFts74XtjZFcXdRN64J5v7f2/bST4+i7IsuOA9xxK5IN7u8lL5MIYTaGdTL
2dE4gtcU+YRnzfH3T6mnhq2AHrwzP9SGPW7RXTFTdcWhudpvj/ARqJOgdMq7B8QY
WO7Kuhu+XJxl7XEf9C/d4xkSc/hYwfknwXxUFf5eeftWpZ26DiE8aolpt5YxKIZ9
SJgVxnxAofJ+Nh6WPd0WsNjyyEtAkXi/Ob3vIN1VqmiP4Wrfc8F3OeV2jXiwd47P
EB097QnH0064BN/D+JEL9DZmsLImwjq3Vqigr1ggGN+WLXA6oOX9r81Khpu3bbql
041tqB3GcSvewmXQ1LBzfYhkz9A/ESzVsbrz9wvJOwx9jhTPSzIOtnOCBx7ndbzN
mSJXHlFZ2ORikmvJdM92aYIWIL4ui/hKCcrz+E5YP46z1siEzePHjl8/XJpFppWr
U9NJZrNBBgjdVvTEmvbY43uU5Ai6dM2EnE/PtnRnH33w8M6KkDx0eItykUxCa5hL
jvR+h/qMcdOWAK8hgmqHEnOWb1HWktD8rmUsqYgRWleTzPLN079g0tkklF3fBh16
O+PKYfV3BPTn7urRj+0q7yTpgkvZhHw7AwRabIj8bTdU1xoaJBkhbDW0XJkVpa+S
HYRre4QPaQRKoN7ryrtewxc7p/SAHh9W4goseGphxCbvpV3+EC34wzEA/zsfaYzK
kUdKJSF71M0bW3uR3uqRoEVoQCbApKr6cp3s/hrCrmhm7Zz+xDsSfDc6WS2H0zID
kVEsjKxENsOYbB0NtY9hSmfQ6/tsM26PHt2mbCBN1rwhKYdKNMQ81ezQH8XAIkQy
FDLd2Jb3Je+O01wDY0g/Vay/xmebPBI1pMHD0zZwu6GZug7ry7SlIYaJHkJcDABP
6eGB3HRI4DAJmY4gQoLEi+75Vt/fimHQZHvoXC9nwa0b43z/3M5Va7DrldhuDfJM
/qn9CauBFXE91xjV5cCemO+TOiyyiSQjoX2qAxWPqWz/QFOsTJwi2BesyYJgJswr
uXeVPUj13PbdL7Sy6SSJE3Op1wtxUjZjpxFOJoEiMQFGAlMvEigdBPVjc88E+l3Y
DgAbY+5GlCsasPXgXewVi523f1unNQ66RDV8GJnTwzPON9G0wamkHrxERvqGn5OX
du04GFenlrLSGunx27Qb0M00WM7PXEI2kEbAqugEyr8iKFcfEk8aseVPK/83dnfI
A5Lx9f5f6v/KGY8HXp4dCEHvgJyuhhhYvvJQTCSmMD2I3Y50iT9SoZoxnZUtr1ol
7pN4t2VZ4rPQ+UV80ONsamh2EpqTbUJYaOYYf0CBhH91sPXB/YMs/cJ1JR83UhJM
rCOB4HtiQfQW9J1prvBIhaHpXkmBktSEOiL9t+7tm+1NLYYahDBGSun16USsAzhM
5/B8KRSMXxu4SfO+6sQ7lYOLq0dzUXD2Y4IbQo4mIMDW8Ay9ekziXK+TXaQjtl+7
vyt2HWHFwkUORA0drrYSBjxEnH2vBK4cS52wfm61TNrayNTSB2/rPKlLyCgNMY6/
rTciO/cDTMmLWBrODx9zuWSIvvI7JAhYR1U6BJI7/jrCNQie6GFuQjdB1no6oHVp
+elUj2BhR7pTqG/NjYoyLSDnI3u04jHgmGQR5wlDx9m4qMK7YkpDnljWsnWmxmwr
iZ6sCmRVdoaeXBtsRyp5k6NLrbHyD1Gy5tgeInry4Y+UGiGJxkDAIqS4jPs0GWZn
UWLFzON+3gXryVIDjva1rcUQ/+bZyAkThlFAyl3ABzqPMYSF88AO0uOcLKrGer/x
RqlXRleg7O8/q4Xc4BqKB4I13LszuGNvogk77MVV+I/7csYg6cOziizoTPEeou+y
D1wn7HjPWzdvENzXzR2RXbZL6V6T3nHj7tpyVNRh9fuWqE7eEqzg0/Ry2aIL6jOq
wVXvtFdL16dM/1YYtRg3IRAYRKg93nvSNkc/jGbs/txpjqLPA6Ehxm4eaZFFYH9i
cmjAjzBoUFYxicIbViEJQpN0yBpgjDSpargEtMAWK7y3jqHGcboXpSwBUiRG9LCi
OUieXBLUp4weBw/YUgT4m9YSYDDi6DOrUgeCm1TtQ5t6hl/33UgBKMxG90hZyM+z
3KMk3bK1Pze4DL2eZBYMVXewkZJeT0ok7I/mUKziLVMJPbsZ+JVPzARDOs880uEM
bANQieiCXj6WDSiCcGb83aS5i9hUvnA5JyVJyX785AAMo6NDEG8eZp1hXd4cWH0X
A5oEs6BfPyHB2q4XKEQaE7EI6KJLhdJsRmSliwT5HOYakdi41CBrEL/Anqwn4vdH
IV+xoBrhB+i248KMzHcGVAXTbNdWoTBCLm4/6gPljrNUwOWwUNhhzpJYa4yFw865
eXA7rYQWRYOaBmCQ6khvY1FMnfG4/wycQQIE+lXg8rEgZCIXPf4jzp8skg32ua6z
RCd1Nv9af0e1ZqN1CdP9BSM62z5hD2CbrwJR/nLm1FZy39Jz52REBMe4boxYjsp/
hhITGwVCogQoWuDEEoPxaT3FONJsQmX+xNr9lXAYw8121xHJo7d++H/nwl5bsArb
/mN28a58dqSBRkTn8MV6bvYGvAS9nkkGVT5xTrZH2mBI5SDmCE1e1QyZ+kj91/wP
L/GkNjErB5N3wvrbd6a2+RZAi1CWqbo02YvUnarFnH7UVL4TTB24A9YLwPDjls//
+dUxbmGaJjgVyzmgOBXJiO0Lo6Uy3PHLIH58HFGzYHkpjoExIS3fMLZ4e2WmsGAB
xQrgwj3twMYA6u0atbjlZW5R0I2y89l9SAxafgQBbN6n1ZjfC7qdLyzpZUzJljnv
lJTzerN5QhiZ+IvlPsibJiGx70WubDgHsBU5OXbuN5d56J7pmSGaSeSeKn3W0X8P
EBwtSl1vkpzCWdTubs8vpk48z/i2tfvMn/Sc1YEm9rb0lARzIg04mkS5lYJLwKJR
NJ8a6Lp3aUuAUQtjRlQawn1KtqZliX+r5R8aRR7KkrCl6KS+odFo0Bp02+mrTRBI
hbUB64CkkBIAaRXKPaV4vFku7fejWFRyXEwA/YCAFHRGuRMPAjhYl7ij+CZcUM/h
NGhavylHV+GrXVRY1gHMLkLqymI/oWCkRmHG21deOdWLvFrSUwhJIoOemef81s/W
9kH3iyF6Jg4kSoWENUnPeaQcgwMPeob2C2e0vl03rfaVJUzjAZewMqnfttN9Q0hF
J6bwyVET13QlAVSX+vCBwH+lvkwLS/JAhnDnfCggk8ecTtkyQfw9xpa4B5hpoiFh
pLELK8W29B/LIwtp2xmFSropbvhJeVkzbR4YNUARLmGxVIhL144vlUDNAWkv0Uuw
IufUcS24wda1GngbbGHrgZLHs2sxriVpVFEj/t0oU9V2HdFRg3FlXT8ohxEMxqJK
lujqD9NApdcwnqkM4X81locrksoNOkXrDXLtusEN0MLiF7k2l8TACGy3t6aN6H2w
4wGpTxVsmyRZW6o/LHV3bJjuDSFoU9jU5Seqr/u6kmbta6C/Vsjf9+h2YOerCyCN
rzSPN5OyUxcbNpDw155pekl3H28eoX8bOSGHnb3hPhE8pr35MEYo6p0y2HZq+sgX
/rTkKEAkMQRm1qzBSitACaptRXf6SiQiKlFAnO31/3Be+yjVHa3krzuGrzSlO6sz
+8+Gpqw6WLcklYVNBfZvmS+3E3Zo+MQbYlmg0v1Y5NmesRfq64uksyWqLwcmBlIC
efxeSNAlKOyeDHEy4NGzuvpKypWliHzl45meG0glm9w83GFTFwv/nvxow0hNl/V6
ghQxFEZNMSbjQD+T69qLc2Zp7BnA5DdvsF/vyhP2WDIkXIBMgrZ6Di7A3n7TdWsP
jynEex7QbTiwGa3kSzMvZnNMeiiFkvg9H/9K+B/j5P45M61tA1RCIna5gGXmzzB4
W7FJLKE/rhV+kPwa9mVo34hc4ULNzv2YcE/EEZDVbDfV23DZXdrRG3ymLCXxWM0t
wKR0xRmQYUAk7f/j1hjsE1gneGE3T5+KNYw/rNTE+VhFgVIWoBEsmtP8ORbZ/54/
C9rhA6bS2WdWNcvu3nuvM24wwkuTZH0lZ/zmxs7gZs3r8BCESCGmrqF8YSgYgZn+
90U41B8EZe+jnhPK3V1r0qYrEvYHItmbLFCc84BQc+oj7SCiq3f6q0gYkLqa7EPR
cVolMaozcBlI9tkzlm57JFqtCoznIAKt0vtgbrejqv2WJsNGf+ek7QQdkfc7Mahb
sSFUaAV93yh9rsg6VeKgPJ/tMFi4qGozEccbYbm6/8DDnDP4fifFO85VzcwpG73o
9zVCl2uHBMSXHicGVlyRqsTK9MdR/B4+cTS4HPcwDILqtMflh3v3dp22mrFtif9t
mCyqsATk7j5h1R6FciFChxtdOwx7uN/c5onBF+r6Sk6XHc823/uEZh9LBSvHaJXM
8LYOuHyWQcIfedlKHeDLgiq2EemHH0kA38vMmrFiM3U5nXqTkb8rwMLBwz1x/YH5
8dnGepD+Z960p+g02+Q1+/MHQJvRmvZwUGSKkjLwtMxjuOFOrWG7cMzZuCSvk9iq
GLnJ7RaSBgVxiAy3D8FsQcTWCxLbXoxXbJMPhIzyl0ZmtgUX2fqWWgM/nHMhAWY1
35RYF396pnL2XZ3oQqoIVCjKhQk/QT3s11+9/HDCeKO1OJPPTB249h9arMJDX6jY
ERNV5qv5BCISepcm5qS4sRCGuyUnxhXohF3PR2wDkGlTlBACfdULvXPTwXrDSkL1
GnZf1Qzru/r/T/oAPwSN1fH4yN7mo8/WP/Mwi2mbRpIhVRjKVVjtpqpHwd8aLmUj
GvEr6lDaD/MltAj3cCMvuiooo52sARXiJIj57rWR91GCfP3Yk8NH4Os/XxPX/hWx
kRi8yhZSgx7TSZPhyy1Wn1mZo/q+ls1k9y9aAac1tUnPj1ZxcC3RJw6gYptYfHQP
C+Ajqrf7D4f20boqLwgaa6iDkTY1HlTM6xnqTrbq5bzp5kIfja4ZHLQtcaKCkeMV
1KLB5fFrb1bx0YK5PFZekXgKGYras0QjJ0dcuVAx5dJ8WYw9AamTRraU1cnTew7z
HOHURhDNMBqIiTZJ1u95i6UbHw7hx4x8CbSYFTNC3/dmm5bjtVBrJmbhCxBChOTW
Otldzjd5Tj1iTKThTMYSxiUUlLZkydWBh7nGyBzzXDu+mzoCRY5V0qILSDQLB9l3
clD5TwTk+wJU5ohPpWVO9zBKSoPqqF2instBsP4jjr+Wu4qnJs2XiVmg+H6um/Mf
dgCP7LDmYYn3XuJ8+xNvppAZACOAlh2CS5Q3BRdKThYq1guRs1C40mBd2qHt2vOe
3IAMA2H3VuiSgf0IuFwbMRMVN04y3KSYqvLaoPorUULIcJltO8wgL66OZfiLE5U/
OMzAHLPk7Ib6nbfp/s348bRDD8Zrnysy30xT/D1vwDicQDCbsyCyDaqnMGpBvglq
g1H6iz237VJgO28m6qHkYfBmQ/XzF1d1ZXi7r31R5SZ5ABWyIz7BZjlPkpwCQRDg
hta1Qoohyi7SDuQE2Ndr/UayQ99ecEshvU0q4z17/+pC537afvWA4kHdReE9OPDq
cDYy3kz8AicmnKCFBRpamdbxb87Q1eFLx/aOYiW5VQ0zwBWUMpM3qBIaRZ3IEePd
cQKHflJqrw0up+rxDRqwOo+C4yh3PR6FeQ/GnjWdQoOKBgRcbdZtlv/UdBoCKba6
HbNP7vkZUG5zSshWqhChlerF7WQi/CCOECArxnNaH+Uls0Rl4gW+GdQjIfl/Ir+j
Bs8+CRkMLLj40yqRY+5r9X0EfA/s5h2yzM2Cde76oVzaqGAUCu2+7LvMlpsxIXWh
XqLBhS4Troqv1k/xa6NovfDb6G2A9calNOK6LdeTRrTCv5aVhHRlgVE6tgyx9xtx
/5lA8mzpob86ZgKRs1BNZSr+9+txLgF8MSCD5sP9a2mn8bRUfWxKWmfPHRZZw4ez
7cB+AzJGecMD9qPh+oveP00B6DUjkfbuKNVmjqLF+iGipiOhXVt4aZPVeZuB7dSY
oe/cfCd7lPJlGfdrgg274yDTi58naDI4pwwY99HyE30+wzCJl0jvJVOfOBKqg0ZY
AwJqRX9oTqh0DyMaIWNvooDI5BG3ZN9d57PvRRH3qUTzbY4jKIlNukGIh68qhiNy
MYCXOk+MgbyWcJM/9nqBUqSEfzekN5eJ0CU2sDHnx+SmppvuZuforqjnmtVT9Krh
UyYfnwqzfwp8dB0Z1YPCBozM3Pjq8kq+lb60VjRCG2TuUygK3hejr1qPjZ3VcuVL
8t3mrSBcPih+j+DxvXNcqhFSCR7XPVptOhXsxKuaTMzjGjpFgeIMKVec7Wiw5NXy
wj0rZHOCujpyhuUKL4ydPf3tqEOmTK7ay9QnH39OZOLyvy3HbsKMOAIM2iHkB651
1gJXhV95GrgU4JO+rAR94n+BTgEKBBFQLm05NYaXmwtVF0E8CH98aQ02DpnsiwFG
r5baww6daB7uH8pN17xuViMqtoeb4NgR8nj8c2segnXIsrFyuxrUQL22hiR9exqL
NSrkAdWCaPAEGz6Xs4SrfAIhv8zcZ4n0Ootbt9RDgmyfItFeXxbRcuukHh9Z1ca0
C8tY2OPcNSuSHEwSq1eaz8ERF3j/BlH98t1HcxddluBog3moI2NOLh+OgZ5BffdV
sl+BHzQV3owp9/ykXUApm1OxaqtkBJXPLJ2jzleVK/4I537eznKAVkNjS8KTKoRB
gCPp+qGG3PcEbkv+E+wWnpi2rYdV8LGGr4tyGyp+WR/zCNovZbKnooYxTn10Anmg
3Cs54Ls1OIriF6i8m43Jprw7Ksm3fJ6H9BPCHZnBJH2K7nH5Iiy+D+c2W5eAWPBT
k0EhIGxojkMweY4WgI3tBaJT+xUsanH4aaZlFCvhGm3x9K636cg3p3VZAoGJtdZi
/5SA+mIwYMtQK4m6Ds3k7bKPA9dror9OUU6OIZ7IWMcuDg2pq4Rd/8nYZB1Ba19F
8oWqY8j1bCIlGEteRl1dy5jzZxeThiLsQjDrm7qPzJKkFBbqtESM+vBTZMzuR7mE
MzixVem5KhOpr8wLJsZUFrMD6bU7I3aFaxAwLyQIxuV44tXkHAbSXaTAc5fZAu9n
g5U5ouqzc6EBkFmtD7FJZYDPIVS+q3dqN91HOcAwf3RaNva4wPzgE7lOaWe0+j/8
+nufdLWbjGZ0onqAmwdgQ5olsL/4aliHDDLUbA6wN07wLIWwe5haaDuvFnfLuQXv
jP9ZWckyDnoOedk0Pbw/DOsInu8TrReQHQ2lzR4SKo3lZXvO/cXu0nObS/o1UwOo
Xos1tHCV8JvTcMNaVLnFzj3lNdVcWeF1c0h5+qm4fw5GXQRB0bn1zkZJEB0mrd6J
Y4ke0tqfbEs3VGHJ0chfahMJylBQkreSA/ZO03WG2cc0C7bklBURjeYyw/DPJIPM
e5P2XE9gQEWmUO6vn63ba579zDeMbv8VSzNRbH0vPCKftkHRAOS3Urmv/2Y2HttL
ixYEOTTg8CVL+dcVp4Cb6TJk9tsXCL0C2wUvo/1xmUmb9h4khdTn4V0hkvqNgMG7
x8ScEZKmLPSFVdPRIXYRujis/sEfoz6290T9aW8p6SllfHRU83J4v7DLqfYyXoCM
r6TUbSmabw2rhbRr9b+Bi9NJ7WkvuREYHVGENdS3b0rLOQN8MGPPR31+pPPUnpf7
es4DOTTYuoo6pW4hoylE5E0SP86cAug0gKdJnkUat9Q7t4IYIpv63/T45YPI3nSz
47EaRO91i6EOxaenpOF671/7idsBE5hMlMNY4W3NDS3mylYDnvokEfjSkTMqYQFu
jj1fZYHZpGqe8RgDCl2+dltQThclCdUi/A+tGgUPeYplvLksv/ymCtJ/txBuYVo3
lP7t27P1MGyPuw7vhwks/ZkhV1y43pq0IUFwt0+recHEe5z2vMfap3InumC6cdMu
2tkXU9T80hkhoP4FEEDWzYnBnHlyMM45vFWOZMgU/6uaWPOgq3qPxmfa6JjDMj3A
TL93IJkMUetRo/stNWVXPOw+ZiK9Tw8CxWmDFGD7b6+zhkiG5Kx9fIiuwQA57LAa
vRXi/6lCbMmoLT1dbt5YlyBD0paOWjfQNSGXXB/gTPu3z9TQth3pHFj5EQOqOeNA
OJ9An5bh6na3uNZaESOMKkHrqglr2coFBr43rdD2QKJqnEzjkww8Kx6uHYvXNUG+
qGOhtsCtltx0EAbeXO/vyIQLtJp8ohRj+j6koNtQyCuLreqLT1y1lWIBYdvK+B17
+hnkjPzfGZOLS+9ATPRiuLUErDnF2ukGxN6CbSPXrNTsgK5XO5Ph4CdjiG6l06wo
NUU0xB30nMQ+RYqfDWvY91xa35t11duzjHwt1Fusntw6kOqkIVD3leoQUVvD/XUn
KzZvhBx8+JqNBfB3sP0OVG/xk+8FyNOVEE2p7hNsPtp27pbCNwJK0K8cp4k5aKEs
9JGyB20tQsfK1yxSemWX1Eyt7WFh7WvcWoGd2oZ1kPuLDa7t6aDNgvQ7Ws9wBN7c
kvQOeXrMCwN+0+/eV7lxgsHEFfTLas/AkPs+J3QaO/7dw2qcMOSa9rOxfGmmgwdG
Vu1fhRi7oxQ1sS+UWh8hasnf6xDH/w55VNUQr2/c4aT1Q0sk43F9kUV+2Ge7PZzI
y5ZDM4e87wIpsMeB0Sz4tFhkl+IYkqyjXkBunu2mNIpghEOgKWsOuKO/5afJQonh
zbrOMfCyzg3NcBU0CbohS2Kt3bdOKwN/NPJzhRZQHU7niDxguLp4Iv84VMSt46Fd
NajNYJfDoydqtylG8HVMv/IDyztBBpXZ9ZilvYa48dnrrnuUNcMkfGSHCZaD4oZA
xEtxLrVvyn85FsOLOrK6GJ0y6QAze9+UVVSH1LTL5DvFGcg8j5pcIlQUe/yLOTV1
DJSYIlZB9YRxuihOcGXbKy7Wtgaf1ResK8LC1ub9zeq1dniPrXhuWGqTI47CCw+d
9GPWBaylgaYBtozs8kXbF7x7KuIYn3eK82pkvihIFLfoOTjZMCcmI6lsamgRJP3A
rH96bYD343sLbHe1JZ6IZwDHNsmSLdPBZv/P+d1NBe6VvF4YQ9fEZWFDKPnCBfsP
nIy1/mhbF+N1CBI7u25BXFK0MJYJkrvFm6KJhnag0R7VhbNmfVfABMvFlLEIghaM
1LiXaN3QkrwrKRCc3UUjYr2Q/5AwTwpVeOPgS4oP76TXamQPrXrUM9Jo+0Uxeepk
kIyvO9FKFVhRHqCQAwYIOhSMTzxOK2Qrv8TnO81x8395t4r5+EpkyeCgVAqRSi0b
cdCXk1jnAKIHh524FdqI6N0A0x1HmiSlt6EoeuYhvbbdENfHL3UZ+zu7ovpVGWUU
9vaQgzA0IxYIfS2InHnZYuB/C8Dm+D3O+IdCyI/GnEhqatgN1gqT5z/f2u234OVa
E5pJKsHa0YW+AlzShnGq/YjyEdQ4HOns1DHYPW37MkMEX8itZJ73NFQ9jmIQSQb2
pJcrhMsHnDOdvp0ElKT1qL+hHzvNHmNusPHB3/QJxopz4yNXXeNhzqFBoTVyUwLD
1rLyHVyumnqd95mMXiTj+MJBb9lfvMTQeZuZz0RCFJBgLBQ+bE7aEK5eJs5/GGjN
gLpP/pv13X4V/ktcxfJPSGS0xlUdnmKnyct9YRh0+lSDJcmDXUIuRMvvhHAmW1ha
rplXekALxgPrnIF3nFeX+czqmC1SBXVqUR0hWEHHHxAcs7rCAhp61VONDt8Om8QN
gLEd1B2wodwqFCIohGjeqayVA15VIHh2JayX1fUqPGTkE2zISdq40UBz7/m72yBw
/0pO1uduOmDaGiylQE24kI+zn3G0XV1wIS0e4X75XxY27yaqbcUPHs4HerRyjLhW
XUsSEZL5Rfwxh+ylpA0VwVJPJOwrtrRv+VwC5bEoooxO2UZVrbfvfLdTdMyl7fU+
yyZK5CyYFIgDDihg2TtFJB5F3bBZqOIvkZdkijCct0T4Z1xtrLq4uerYkLMH6S5A
PFb/p/AjRH+f87zHL9t+uiRMg8noHcizy4nL6HnU4jjm0vM4E3drfGWOzg9VEHrY
XyOEwrW/8vugoglKfz0c1UlRf/ypulkrbsJOeiscXAPmZr0F9vLPhQeX8cddMcL+
AP1kLsttcqhLv8czlgeBEPRS/Yc5DBQr4D+2njxAvtXcgHJf4GqkSKfKxZd4dydc
VdEF9hbz2sKZUdByT+qW3VgDhXUEs+b91bFwLUjiL5NzXKKmIvkTe1kuiGx75VFE
CdbongJSEe0C5TNgQlIUW+cvpda0dRbBekV8bQmb/d709mIQ6mHqvCQgDbrrv0dh
4+a7iV0cT1v0q2iYMaTjnpLEO2Mjf1bcsbKXafA7zR3ktdbvUjP+ESW2ljFg01Nm
te4Cvt1iz4+baqTzYpcx8MjVOIst+rezB9MEAV3cXfOd28/WiJrutNN5WyYyzka7
WJDbQnTIWOoD9cgWnId6eSdGjhLBFcZkH9JuQtdLlR17V7AHycwb85H1lm74kKqv
gQrTTL3ICoSGwineyJ6BpejxCWtTsDW+ALkblOugH0aMQ28j3oFW4z1FZILMAOgY
vLcuxZkPvs4BPFj72MKmHA5R668YdcmEtfI3v2gOPrVyKuV2RZVH8auIEBLi3Ltb
ZG2+gTVCeLgvoN+t16h97jP3eqskEyqWkkxSrW7GddZdswUl+9t3bZ6KLVptmWs2
tnEL7JWvx2gvTVPSTcYMr8aMgQTa6SjMvA3NEQo6dlK719LIv2zlQMNK1NSoClRt
zA3jZtwMI7ZhRXJ+4UzSrOvmIcfMIIcfbuiJYqxei61bbL1rEEfYzQySzIMAimEc
yi6npOdm+AaV+YZXpqr/ZVWrK9o8nmN87H1B68YjNPcZHKuswPg195zm9enqSe4K
0rI1Gg3v7MWf6jcAxB/yfTvfrQWm1DF9rqO195s1W2s5h5i0NAd8mStVhHqahDD8
fMcxZAcAg80nvN1zV57lBkxpVEb0pdW5Q6l5A0n1R287WT8Z4PLBTsr4YtMJz3Gj
ec65sg2EToE8oGNf3lU/K8nWRAUNrGn/boaENmz/kq+Y6uG1eQe2JCKo9Plm+Bxp
VAfHxg0aZzkeSpzEtE7gFPZs11JzCFD9UOKVVCDiMKUPnfzDeHPxRj+yuD05Tmq4
uWxpS/HjAKNPECEu+ZXvYSpWYyI7xHpgs3bFZXKG3ymPJasImkrbiw9L+KlM8Gb9
qxvl4KPqt4QLHUQ5nRE8UNNrab4HJNiRH06q67ExKFx3jW8Qxej7osmoyna94IBg
77aFqdnwkexxZmYwPAKjJTee33oDS62xXlspj9GlLD+SbUaiKvQGgL2BzwpfxbFA
5YFY6+fat0mjNdvTMZB5aGi9DtFvjXjC8vYpOxSJW7Bcg4P1ckm/c3Cx0hbsV43H
pqBFXEGhGfN/jzzgvw7fGnJS+48qwaVM8Ai23bQBlKRWndveNmefKPFmrqgIQERm
yODx5GmTJtQuAk/vCmS9t8Bv7jyj4DjXe/blL0Pp8bAU1Z71WdhI+T/+W+hpaiBD
6nbeWTmktULXxSD2P8tPNBWkIqID5cUIA3iV1R0zvL6iAHg0LZ04997IWm1XUSA7
BwDXMeZrFTc0OC0o+RZ1441XXKP//fkMGi61HaqtB/AHcthuszF9pUnnwoU86HH+
pe3IFUeZPiieCV5bW3HhiPk7S0VEKGGEp4IjaDOjnGhXFF46tlV87j4zRSy4qVNb
Bb9ySGSmaPOYOk5CMpn0+q5uUCap0b6U7CQP43VWDwQzmYew50PfEGtJE0ZtuAbX
qJh6ULe5Fc/VqeTBEf/BjbcpnTiYfBpGqpMhRhwDfA7vVzhi9HM3zdV4GGdlf34Y
W0CvruV7zhgDG7J7+VHacaLAxd5zF3ML7E3oC/LxBBW5+aV9ghFlH7SLGiKMOlYN
WRM6ZrgSluliLfxMCmRsWaCeJudidQuPGjI64wY87ESqH5FKFSzsQUHj4EwRqc+K
4n7r1S9WPL3+UjK8v9Sb2VdyvfXX+GBKZgJyqXhkXyKvIpkEnkEhrx+1vdijNaOK
Z4cQ9Jh8XWd2nGcTfBV1nTlG+0gTzsATX4dAkwKrY994Yl4ew2mzL/bvFAFLz3HR
FQlubltYNXHvBDfYWKq85k0e7Zz29y/L1G+A3f/QpEMDbiIQeDECLqdnyzWDUdql
4B2HicwbT6FM7v2F/xQNpvKNEk5AxnOhO258uvbT7Uq+cO/ANde1oDxiOk2LgpQG
RFHGuKttKt6YODiK2Vkkr98ctC3Cxwq1KYfShSnTmBOYSZ6Ju5UINtHg9iUTiHca
DvKPmYV93UQxsu3YHRCRYkS6DgOhDwY7EoUwD90AkZxe+e3/5UYdFk4qU1OAraxq
0bO9e0PyZIgZcVlWqcQeoGKM/6m9TOkH5cZx+ar0ZRfeqvG/MZdW++57vy+t0UAX
v8YwB7rd7dJYu61V1jCTHuGbtk/PHgtPC+zFRlKlVL4nnBpNulcnQBnn+M+ciI6p
ERt0NXQFMZfM3/aYz6M0MNHwGRW+8C6MxD1haG0A3Y2b1XMOrgZrVgj0/YT5U/1u
qHWI4XdGiUWY9U0cmy9hDYDim4I/8HEys4R7ndb2ySG9VygwXFDaeuDLFCkdA1nH
VFUL6gis5oK8a7f7Z2B6Fy9kZ6vcEML1HxH2xQ4FV/lcoG80cnUBtNU8l5MTF3jT
4Dyo74ZnxUIAPXIyRrw7RFEBc5/FxM2TGEp2GEFLcebOkHp7CLv6rN64yBmAhcQs
9BTjj3imOUycnDx1BL7EeEqijVObvCazAqMm00OXLsaD7D80SFguuNxPV+GjXidl
Fzkklu4WOKObuo6fYS6k5wYzrb35UVb40R38b22Q7rJlxCcr2UPEQjqJF02i4/yL
KcvdK4m0Wkd45JQ8BIKT4q1itRZJFJ3lmZJ0hfLoICJjBkzBbKfXX8MmAgg7BPuF
AcI56/In/0CTy9DC12lNJdHYpjEW37KPVziME9OvaJrle52lLKXqb6guN8ugL43T
sBPm2NgXGxttzx1VRckjUi8KjGgJ+oGGzC/iP+eiI1Yeb8TLufKjSxD0ojx7/EWL
SmGKpyQyQcfarrdUXFbeGihSjjmpX91Q1omRI/yWbClKLExsyuQKe+ZhJm6h9bIf
ymP09QuxCop1A41bcbq7EEkQzyegYOtMkItRSvHX/Q0GNRc7xQosdKyDFqV0tJtc
LqXc6DdfKQ16mFJjGVHOQGHF9xnspceM7ae5r73evon3KmZaWpEQ5YozAAfNkYdW
zACM+f55EXKagiJDK4It29tQu3MoHqTsCD35MUDMehSFKCclEp/c7uHGsS7liE/f
uijyIL5pWmkgxdxrWGe29F0qqqI3vHEMUiIRuy55vUjfGcub40jK9JM2/ebqRgEG
5nPLd4TWRNT/2UqEQZ46JyFVHAaozjz9Vp1rU3VlbhuB0Ng/atCfo3/am2NUXII0
SGi+jLUCoUEvFaf1NsCFC66yeJF+zfB1qxmWcxIiREJq5Ibl08hbxcry/4j0D2iW
rG4h9K8qPAhn+XSgG5X5uvnabYNZyIc5mCrpTyfBGbOMh++Z8ID0/AexgGGQkq0Q
Vn0EFPUJ5pzv1lcG3fgmrjgIQZLAUvs5yv8V0GaWBnn93MloCv9s3Ay5hiJjYdvd
oVgiD5tYTIwPmtzDvA3Sim6UtFDJjP2E4LdS0ItRyH/QUvzHX7LydXGBsp3wB6By
K4WiNpxsQiVXQ2BzaGhMeLT7eJ31pZm2WVvKGVD8nvPXMHKZo8UjECz8KsUEbZtn
8oBZxJ1RJKKegIQbdjPSLLYKfNXCbrwcvz2V9ifHRwLxDGNkxkczrgHC5ITtFkwy
hqNzIhQzGSf+++qry53xdd11AO3f+ekjYU8qzoQsAd3UNYvHyDStd2k8cExID24f
XV6uj25frwoqReba6G8EPifghAmibx7/KtjuXjGkpTkwgj82IK4mVok9SFAGlqkp
fpdyB1n1gsurosZ2US9cyABHFxV6c42OLOOZu/Jcktdofwb3RCy2qy8/4yuQHwxK
wcmx67XnlhbRzOFIOcJNlKAcLckxymXUW0llbugqZctgEaPYP80ybcucSYuopw0T
5hnQAr87W6PA+giBzJPm1xysov5p4zec3EAfaLjxWzuiQZruQmLk91UJSVm+S/jO
4+4ECQhVv+GEQ8ZQ0sFH3KolpDDOA2isdgX35eDtUm2qkXKGNAQ+45jcP7w/pgd6
6848aB52wzNsxrBdK+8RiM3mkrG2d4QtDAPWk0JFH3KtOLPKWPrZb02GdXImT9E9
zY+LRKPdG861nJTcR9xOPUOwdHqI6xA9Ort1Y1HdaXUVZRAz3uld7NRomPBxm3Mr
AIj03NPZEBb616sF8q2IVk34NbyKRwGOZwLd5b9z/qja8QGe9IoHGQrxnlSMkto6
t8vfAAjeuMQ6vdA0MLCoHWGJQJDLOj4iaj97vdrv1wEnsNswy4bGBvbWOAp/XTWb
+jnD0Vsx+R2qnQZ3cXofTVK35SvVk1VWNgBq10SoWqKsZBVHgl+CW4O3HF9QH+IY
8Grf9SdzkBRl34Nl1ErWfLWeEFabDoacF1LddTZeYsSBhSj0TWkXSAlrL7HCnL2k
Nqw1inBvEZX3dQnVCXE2gRBl+8xM6W7KxsCAidJdkslTmD+8bH2eN170cjLegeon
4acFJlPiHLxLLMET0z3YK8D6AETSSFGCXmEr1nWmnPnUkJfb8F+bl//eZm+l9NLq
m2bman39IOxAn26mmucqLqDgEy2NkL72U02jw6syd2LpEqhgAjUSm5bOkaX7Yzxp
z2a22RSHR5SJLyF96X8bCNIjbVX6XG9Jt5Fqxk5kMDApu0pZ9KsBg2BU8VRuNaZy
Z/YFbueljZ0qNCrNUeYJFkqBz/6RwCpp4haSnUIG53iLWkHCYVOivy72yiIbepmv
bfEmpSatNF/cvyTilrj3o37eDKZdWZGgXVPtD85CogIUkxW+dRIUrBhoBCET4Lxs
t+oY5tR2dP82CYvej9+Pdu9FrWCuxh/GRs1hcGV66KwuvQg0e2prVbHvdf4wQlB6
jDhUpg1YWZ2dLVheIfVTD5F/iwKRM5n67Q+R3zWRKA7MDdnkInhxp+CsiQrvuoS1
7aKVV7wH3yYcyniKhQzf/h0i1axp+np1pnGSS8zg9rYnJBIyyBleARJgP/8wYZbw
e6lIWs9xdAilr0gDBkQrS7JRY2ZK8DlEn0hUBdimMnJKvP2833LnJT5j8HjRktJw
vqMbUc+U7yV/j46KtAreiCj1NntIkjAcyZNYeyBvBFd40sKioUGrIjvIonTDahVW
sD+NonfnPb7qIP7LQZEyJBADJz8ZYoJf5VUDK2xVpF/hEXxCvp41kS5Z7aOIELSD
VdOfVz0SwrQJGsORRbIIX7c03D6FGFxiKORAxq8oMcdOS2cOQtVRbcux3VhI3tAt
CIFgw5N3OLJg4TCxyWHCKIeIyjYeWrummSrTtE8j9OUvD3n+/ptIvzsAgTKVfOjc
IEpMhsrNI2FLOD7imcr1nnHy2RerMjTqD92PGPIeGd5A7doRpTOTm/jUbH9vdQsi
WYUjNGg4FraiINURsL6iSNn/fXR4gXMn4jZlC57zqpzkvGg5uPeNeAyVMQdNUOYW
CTT6pnmk89dV3smKG43TQVOLJuyqxeE3zofqNvQzafPUXLJ2h4b/z6c/CkgXQrBy
roqhezgDGVjE8wgljyf1Vop2+NcFaYjeKRp6x5gulfUKMLlrmke/sImFm/l1cIzR
YOODmAgozQ9nyZJaDSP++ctwbvZmwiV5SVqC4Xl0tNkMF8Bmip+5TObU9e9Dg562
u+lVguFnoNpyIobWEzvWyWS+VFxn7hSErJ1tMuvbagbSl7YL1dzre8pe9vcrsfH2
MPjshe9Eax5CxaSRygvctGJtkPPMWPFiHk9cqcaGwRNkBLZQx+eHAy6IzKtmsQqj
lrEr0Koc3iLllPb/ZtFAIMW7EwxYgye7MVNmTd2qCKIWhQKDbTgu4dEnlxBqYa47
yuown6lkHl8ms9fiNdqMfQuRoe0EooI2t6zVq28n4UHRy+lB2x+LjytXcdEd9LlF
/hMt7k6OF8ZHPiKBlVCyS083ocgObatnut8bpSEWXS32ShZzDeYcYvqaP2MxR9s0
XO75eLguFXVljO4CTHwP9a7maHfSwmHzYJ0DZJlJ1M8meog0WthmAr5jOz27+U6J
C97cRgoGU8RVkzi+g7gqZwLsCLJSlv1WagnKifeknXmdVJY49Lpv07qqVBLD8X7s
GGUHfXvNkcX4HKdPRpfUrQ5jVsvs4vb4UR+IU/2juVUFE6zGxLxs7k1vnO64Cb+K
ovTJDxBcfQ7z00TSO7cNwxo1VtVMl/ENqtL5szDEIJj4lF/7xouCkDQrMshI/Iez
m9A4vP3inyB41I0ze9NSXcfOgEA5w4Og4ESkzsOvqYd8EpcEiOccqK7UaIAn8/Cd
PuIfvpgx52xb64UoQJYc4tGVvdWqj08xCa76ZQHwcOmSl/EFvzHs3LKpoiTSRxxd
xa253GaitfoR7ywKixIbiYgEMNPqX9Z44NJ1DrfGLYYE+zlFRtl6mxxV7fq1tKV3
itPTcy3ULTH2NOVKI1z/15dwch9D/k/gMmZmEsJZJSm9hTicZa8BwBkxmSWD0PhS
TmuywcBFv8bMxQXixjTX0wmvG6pVnAfiKcDMk+EMe94oOtbtD60qu01LNmYMd+5m
7rnjtL2MNiG86IECbmeG3VpKJZ76fwkBe+ZGjPPBkZdIjRE/PpmsyNS9fMxJ4kZu
q3ycL9PI2MNSzk0QPn4jN15C6G0ycyCA55YBNU3BjV7L8QAaHqcoE1yU8vBEWltD
Og386TLIqRPmoInzKK8YPpD5uVricxOUYl/P0kyZeVCPSeddVqGgrma+Q8Duq1W4
omH7nkR4C/rIMRxSzbbBgPLCBsHaUAQMDgAqSYOlxflMvhB63KhVs6frQNXrg/+N
m3AYBDOCSpVjOkjP7p5NUqtPzppz3FU2xcoB9NRIbnwRkHhLoastQFpFRO0msIK7
T08Qh1HzyMkxafb+P2afaWDfAPMVGgoD66bxKgxM/EfUFgl2udXOhIljiZR9GaQB
AmESVqC7kP0KJVSb+rUGoiK02qPycuNuWwM907OARXWSQTvoiZXLwzUXff6SedpW
n0KOzPLcfY05nIWvBQvrzaz87Om1WZa7GTFL47uDZtMYBmGgiBzCyLHsCPUlUO4u
NZt7IQdKFmTvkYf2snsfJr4G213+bN3h7ZYbD4vtEq/VS5nzHpJgkN0sJWlngBZc
WpTS7N//Ls2pJ0c43ozuOaYqQdVpWsYDGUyGWVT1eUcjY1XgY8nTm3Kgij0/svqW
0BrgijBeJqKvZIJ9XcixePwfobCQqngJY24e89QDhA9oF+I/9uB/TJOtdAlrXYXg
FqSZdAArcXclXUULf96fTNPP5UXO5xSvHer7cfxD7nWfED+RBEX+Yv6UWms8/KPq
/KJSOO/4pTwMYnG839ZoyMZv72m5EHanLQZPNOerB1i+ZnaRnMkk9zIE8xAthZRt
1vKazk8sH3YeRmOh/Alj9Hx5EauK3WFM9v+JrXha2VwgDfh9uJl6U8UnWjAu/DcS
dMSHDJ3kqtVk0FYB0bJGwqQF4otnN1QpE8SIG99v9kWPZkllJmJsa2ZNMPZAdLad
BEWfkwoUz+pg1tn0EfRn+4mKnXxC/uxC6y3BkWK3DPRGfhFHkhmBOAWCcCd4th6+
PMNDtdELmgp/BYTyROgwQhJDcayDi6zRq1hxVTrkQJf5Uhcvh6x3hSqK8RwkZPg+
gK8nDSmO2eHXlm0lBGAAyRXSDXXYydoXjOQ6IvY02e1AMeVwoEudPK5hQ9ttSRkJ
PG72/l08aWM7ZdvnfxrrG5pW3VQmScibk4tm/0wOalmJX3W+2TUALEwKb+5oehch
6aMl4OayEgA/Jk6dV9BOe50dWCWz4G4SLmuCNrFBYhHfE/EZkjTg2ZEebpJ4Jc48
wchZMMQObUM/KTDExqDwbPQBPWGPtQLsp7pHrC9PiBG9MqWjJwp2WUZIp2cSsuA5
vDPDXr8TXy09uGY1/fvne1QWlJVhIqbs2nyNUGVuzuELNTxZ8hDiBuEu8hbl/6ZQ
RL8mvdulG4hrta2fMvrsRAxmN2uHBMvSByviCLpM0fxQfm7p156eVVzTPIzj22iY
Q0wx2rGBg02Rekj20cRYOmFbzQS0jRalo/aIkOIiLxko6wOJX45fRcwit2AJ4A/Y
lWTpmtYiDAWHvejIh6InXMistqA6TyD772m+vW9x7YLCaxv9a2x/cl5o85Nw1D+G
uvCbs6vyNlnQtte2Ds4p+UEXK5mp5VwMrlxU2jEBbt8fi8mcKR+sNrPH2SPBj96L
RM0wH8joSgTr/KOKjPqY4iHNQFBJxoeJj3ALnhX39pUe7fMCuqCDZnnoKfwTpOd/
ytUPztfU+TSXvt1FN850sq/bIOJCIRmdRnm6sJix5UZe8WuxNloyZlMU0wSo1ISs
VyN18uZtjY2XhbNWjZMDQAgCK+ArtwNTb8+9cdPGB+P9XFwiLJwEbb/q/kyQpmH9
26qufH6snv/xWZcwWsLaJ1ksR4ZoJpuMG5itgMSWx2oGih8cfFSvjoHwCR7eTm9r
ts1kJPFBEHWANc2I6tixJBwettBhssQjQoAvOdz4mtQRw4VEGbOYTk6Bx5Mm8ofn
NUu6WdOC8+h6vn+/P58owNPaztFqLevFt0BbOaiWYb5ByNCDyyDTd8mStdkLkIcS
uUujo27WsFGxXKSdDXmbu0nmLQV4PVjDM7S+V5syUrXcUGznYrb/MfpT1uRLLaJf
cdriWg1cYgzyHPKjyrhydhO/vgGcq2qITVlndkf5Sk9VLZVRlBsy5diJMm/xNHYv
ogcfAZyrZAyy6fZ5D1ZMoOarM57hdjkX2rRgrrjPrcvlFFvPOFPC56C1QSxXnk7X
vEJbGj83oNV5Tc9Ma+ku0auGXDsLo4ShGwfNfDY+5xyVCh6Ru/4YQaMI+2WCDC85
wHrJWwFTjhuXeoHQMevpkIXE6d6g9iN98bHNctZwGrjTaMqdqGAjNQOnzinY7sPZ
/mBOXt/rYxFSI2/CgIfvx71u0PrOo5pTj3HApE5Oq/vFQV7Mn3LOk2Bu3MVr55VI
JEUeWn74R8kCG5nk7ly4rOQZFFIhbbbjTehLNGpHPAH0Jl8kZEfA6AqaeCMH3o+j
19f0hBDS4rjP2S5vBHQ0yiosufs8UZRTwNlUPkgRCbxRGx8AICN4HfXVx2hJZ4Uz
KQ09YLCUNGA0iXBkQZjlwj18bHwamjQuqjNR5SobYsgEInPLyGAgjEsX1au/gg+m
7tUDStVXdI6gM1QfnfEVnfhrmosCh2Hv72JqWX6pozzoQ3s/eumI/rk0FRI0WiAc
HdbKwL/kifyztaKnOdspCJiajNMpzT7fCzGmtNI0/D2dDmf5JRdIVRT379LTEvmw
7UzIZ/xsp2JH+46pqqo5+okz2YBYwLOdp4ItjyFujGyN9FdNNRl8bq8zSQQqEBM7
z6IPL6Ny+Vz2k2Bg4qtlP6PXlZHk6zEP9L7l2wVkG5wwx0Dfrot4iwePFxGVUdCk
y18zzQNQLEPF60b2JN7mZ8fitoZKMl6j83JtZyBpfX88I8LXyS+XxbUrM6aDIOfs
Rf2/421BgZUasq7qTISTfJKGt4PWKHvNTKXa6p8GzzbaI55t1hcPGEv6iJYpLzOE
n6Xd58NWKJH/KMVkTErXJol1rWiTs8FfK7JGBQ3kA+8Ql7Pn+Rpzj6hD1iS5zIxP
+/p4GNA3jRg9X5DPqveiRNipX0vUTJ/SpglStXc4PFldt5m1ivA5dDOTr9wLWN6A
18OVVaCGdJZXFp7gzQLFVbVBBM+lVptQYV6zZxTEbvlrJra8coYHOrlXND4NmjBo
pCB9SDdjsrviVXGev2lzIx6tTaSHCXbXMF1RYei4TUQ5hYMHP3EO0CXEFlKjlpMM
vr227C2BMbqxdatttWEymePNeiEbWOhozvLjGvN3j9fW9VowSljWUD1TcDwE8Fa5
9bGzTObXWBbHHoTb75zW9Yib04bcOq6r7BVtgrwNhN0NyeYNe9j9/nJHKGMK3cl8
HuzqfrHgV7WXAsgzYYZBfGpC7VplWPUL3bNdRYXgIVTd0OcPQ2xdLCuN5MkfcHRJ
DRtYPhL9ifLkktJqDaIfD6KFHjx0o3oXpJhAOCXxL1FX4mCoDHdUorQFuXhYcSBa
lhug3M/0f/42fRV0pprDPf4we9KNv7wLO2YUCO7+vHcY5xLsIM+oYe6arGlUG4ZR
PsiSnJswYf26g1ZPQpQsa5tvRQNO+Hs91cv4wfL+4UzKAk/uu5BLlspG21cSxpZH
d2Fb7/VTz81OW6j5u1E0Kqoi2IObbx0hMgVi+TtS8HYqC++piiaJYZFr+aNYnS88
C5pilMlf/etzIiBCu2CkIiA0XuWywo18AEWOBgLUR10CQnbiRVy9hECEOVWjmKQ/
gMD10TQ7rimSBEAsdS7Rnog/NMTzN8HY+UAjwrHIstWgtNeMazzOSV6ct8/UodKn
RYRmRgd3yF7vD0NhHQFlqtdEihjUG4ctX0FYMA7dJH6DRNNAq7hnIVtEM+EeiUtN
/jpq5aIKFS1ELpYFPfqxyra18BUEYCMomRLQIhd+gm8ecM+weDNEuarQeKcp/M7S
+yuVcDacYyzAKZxMdOc2WSvX+VZ1uWUv+jITBkL81QBEWdvm3S/XKKLU5cWWJyzG
ZiGA48iHDX4s20pwj4fhvdJNB7ia2WUsXmJaCgeSro7ULdLBk4MA+mvsIHrSNy5i
jNYlxIP46vb1cGujbzTPPOzeMi6VStURFLmxnN07EtaUL61DZ8IAbKN9JaFNzb/r
mesV6qfn34AJWM9xcYNTmwYQ74ghJ3A39fvJJy0p6wmppT+DFSl5beNuKhNMtGNr
VGh3Gc33OWZB+wjjmFMtmXbdqgMCQirDGs/+7Coy+tU7k+gAerMk3f66ksjYCXHV
e9+oUhyEIrJUho8JqpDl5BHc/mlzUc+UGMJJV8edxs8Jd1FUx/evKU7f9VW8N3/5
IRZr0P0ZMlvuo0nSADYrtp/qSaXq8Tq47sqJSahrc+0gBBdo3h25HyR1tLmnY2KP
0Tq9bZPEq4P15+tDkTDO6Erb1FqdHsFpxJHlruQD6B25/RsJnnk/hshxVYxgyDRS
RI6GCJEaQBTBF1JLfWZoZTNeQONFiYtKWPILQlwMkNjNEPM0X0Ic6hi0qWZ8aM9Y
tMPUaSe2fC20v4jCl0Vq03lraeIWmCeQ1R/VZ6qbA/KfIrmm9Wm0i4gaQS6zUb+q
L5V9Xe4jsmtKNluGR4ulgHy6bLX9+fC9HsAE/jPvYBkvzM+wkTZhROi5XnTUBPPE
zOjGv0aouyZs0NVnAwrFkuN8u/x3rL/p2HAEG6vWZayey67QK1GM++GQyFRVmUCT
o0EdNmNrHEbi0GDUUw3u5WpViAXPr76mOVNKgmdwcved6ZNBPhSzBMnlFt5kzPH5
4TYtXkxZgtMAyUBdAFZUiIy3M6qdmOAXRicrfbM05J9d4ghhvSdaxKOQlFZ9vV1O
MadaGWwEqOwZvxrnhr3dQPQn69SrnVszI/UBzRf1GD52kQ4v4G4TjH1349cMXQN/
OBwIdEABVZkTOe32NUYa+oJpRp5UgmVwwaJf2exQ2EFr8gmINItIGxfS2nMk1Fr8
jM058r0XDXHtyEQv8HSzgek12nKdEaAqagDzFzloXiPYFY3pQWxdCvp+ieALSarx
QGfZKfzioQ1SJLaPzuQDLwO40jWfCbycW2rHjP5/K1rC6wCeR6f349DI2T6cwTSm
kkwMf7vOmn6HucD+FJuQN3Mf/XyYLw2m9ahDTyNidg/YojM7/azTn0oo1Ohi7GS0
fu73DpfLTjQJyYI08tN8qjoDPUmj5lgEl/tO7lYWu4vZv+//X6l6FLhd+PHKXAbM
wCputNUR9TJn36Qa8/g28slXuN3zw4dTID/1bnkK0nbpxJunyHFHLd5M3e5mtpWP
3mc0hGZgKDTa5i04BjPl/TWN7u4nFXv5bbd6LaMhV2KNTLdceV8AMwzWUHdtryBy
xOXa9vFwA3VB8SGwgLBDT2aJUl9wtJlR050s/BHHG1MkHyrsyrsMxXlj6BQP577L
lnWu2XRCXsFc1SjlllhWgGmFAHljhy2/cnJaKhmoaoOy72/PWW4QMsct5BjnlhHP
Dm/hkpURNNPbGSTWX+T9RRIlNlxbER6P1/OQqCXT9jh7m5rlLmH+Xr7QeXsdBooV
eYzeyte2GZOcg0FgPSLC6lwl9dF1JYXJfhFu46H4hKuXQ7Eqe0KX9hAkbKwNOkOY
6Qt/o5+lKs0jZz6+4P7bOx2E/Q4mOSbIN8QS++XrrrfKNXuhgpZjDPBzHnrSLpbc
pWnT2SligUMbe6pHlJqX+hBCXk760ginUqLdahDwRZyJvyzZ+c2tiEW6GEf+ZTW0
Yrrc7Y5uIY22U7/JtZInreX6AYb9soRia4bbL45m7rujjxe8hgJr5rE1gQIb6/Jl
vGvqen174vDhGNvnfZ6CWLTN+rzidCSCNbXPdenF5cn2wx/gAc1l1Xw4xuEoJrBo
xoFIaePg7/inPjMTHsPaTLj99TM5GpKevNzTpg9MHn4ex5OD8SeS8mkYvUjNC3i9
iSmrnQxT11gZLlDvbC4dWr4hQUeL3zd4/WdksgjrLkpe5BwXZ+HuwQiooevuW3JF
N5OwdA5ihc3W6qEcUv/94JztYbl/nM/A+Oo4EK2qsKfotvIWKiYArclvDtWbCaBZ
8Iou/rM/IEshSlJj9JwwyjB6fkEDkGhYOUgWXqDJV8nrLNFpHS0i5hh2pYjUt8Ru
DWR+wystGRH7UxO3MOwa7ESQRlTiB+LaxqezD7xVfyE4nART7RmPObi2/e6x8px5
+qkBochrd/rMx/A83TMNxKnUqClbGuHuOD9pif9wtaWJIt89LLLGpcsEU0MWwDiU
yUrixMuA9SKpkkZOWw2tYP/YhMiVo0Hb7pjXf3+6/mYoVYx3Q3Dfx25z5k6UnuOD
CqoII1asScND5OfL/NjOBxPJ27OMSIh6J0/13Dr0tf6f2yaK16937JMswEoE4qd5
fB1a/rSwbGCF5o0doPtpmMgdxNjN9ijC0AbioAFYgp8ffLiqDG72mVruR7Ewkk7h
gbbZ35zclc0QWbnCXqFHVrxFVTcG4Y0N9JGw46RnNpwcGdQkU1lGHCaVcitO1oxL
2c64yA4r7Fio3aH3UO/6IdIjn2h2cYaoWKKr9OlwYE91k4W16zC6Ws2oe3b2yBvD
XekOGQKw2jwTkLehZ9mgubSApqFHdVAYLmzTttqysiK0H7p286S0J9JNClQZuveA
0bgybpu+vS2rYgE1xqG40de8LKjBdi5r+ND0z9SyFjqjCKYn4whDh9Ty1x2f17Ol
/uReIBVof/B11iK5x8qyzzM546Swcr8NKs5uZvAuVB92RngmwfWgw3UxTKjyif1/
P2XMCIgS1Yc2Ds1F96dHpRyS/H87eip6CS8kWUETaj95kP1GAOCs4Puwm3QD26Dl
THd46+B8BSssG5B9nxPspJQngV+ISAzI21xsHPCBVcaPQdavI6wMaUVGEQ4l1AC4
wwxVSkilSjx1OH86BtoSfWuZPhL91ENqPVUpzKrg2n9pxhJa1r1XWvNzLOdGQ5bD
X7cf+or3L4SUNTK1w6Yjf7Dth+e48OTAnrjHxp0YMbwUM660zhijkDYCPRGJjAeJ
vqnmbO00McNspmEM/DC1GfdKMygndpIu41ZG4ppBoJ16GY9l3Twi6jBfOGyvU9Lh
dqy8I2lkpNj/eshA1KVpmCk0KV3VA24//G3NpAvir+K+0Uszh3D3R2Z4MUkAWGIc
VyHsrccBneNSPxCg3EHw5iD0WBHI2OxbwC5USoLOTanRM1BgRonvMAHmqp+kO2gm
ane5NvVNTyGD17YVb1vERKkPgTlfWg9gQTlsVIkeAWQpYFBK5HUzyg4Qd7QLqzQi
EO1xd/M3gDrbCcMctFZVpQhumxOUpYiNTCEYx0/pvvRWOlSU6ilmESrV5Zb2USMF
gz8y8Mqj/PsqpqEOgk3xZNK/mFVjrwG2HkrtUPUbCfbHgnrJVxUTXcuqjrQrzcpR
51yVubv94eMtlmun1Uldt4wvWNWzbvCr3JRFrxk1xLGOywi9yMmU6Cs0emp0pvIb
RsojwyRdx/oFc5XFliUPVTcSljJmTb9XpwkYiP1C541p5xC201GQEEab5WARMNrg
9dmDpoV+GHp+gcpZpoHt/8nRzV5EJZ69X8MXk1hJRChEygX3TpLvdH9xnLnQwidp
e327qygINrH45oQ9Rlgv/wrIHwq0cdQBvwItS2YBsbA8mOZJI7o8udogwfjV8XI9
/4vFeGWVNsTu9G1WAdnG8Lg6NhoIm7SowMboHL4qqIvRTZ35V2TQrR8mxvyAn10V
BAZKYSd1PKUEMwdM54Vwu0/VXRj/L9xJO1lpZKucR1pwmW3zPug4gDvBmxbEnwIw
RB1IeeJW8/JQ/y4THbwh7fzfTKce42WWGhnx5uwV2nnPdZtFDx28o1omjATuiAED
SfAQaAgaa5VsssKGVlHCweKl/99hZ9KJxoSS7gqmrLK83Zrk6e3mxQkpn2vTr4aZ
ZlWGNOA8Y/737rfOAqrnIlKhAeBEQi3LuiyHD2xDYimf9hUd1z5xzA/G+uK3SDK7
pUEddBlVD7juNVlEow+w4Prc6IWQ7gwAeCfndogEk0BKXtS9HpJowkVfh3T/cDjv
E6np4SnqKQi7ciy+RjH5ypinFX7s/6sIm2UUDdIg+OApjMHM64NLYEQ3jM0R+B3V
sXvAKZm0ct9Ei/f3rTy8vWjzcw4HrbPODQWZ7erQi8Fu0EciSAN+25O5XvzPsGRS
G57aZUk/n0vmTtMI809xowrw85L4/Ui/e9CebaktdCAnyuV5Q8lEY8SC4lfdBatj
2fshNmo2MWkBq1kK3E00UsyLPI7roAUlITgvfeGQ/RTuNVZqTsMnz5tCE1CRgiIY
hQv66rKq8ibyzt4C9v2uL/79+Ygrk39GsH41YSHGFbNq2RfmXQe2ujn8j0A61PMY
3fJAmCfSxhMnxuoJhO751kuFnqp+OXUbjlWBUVtlnoJ9MkyeBU05mmS3X95jSDeL
3F30MZ5nBI5W3fDyGZjjYIM/fWG4xWiVojTLvAuCzdGF89bxO4nOB0H8WXbFo7xb
IOVCP3qYvVmnP6z+/7juA7iSVxL+zPQXbk0lmWRMe7G7n3F0DdbFaSv2hLg8Cy0T
yYFqu7xtdV3y7JvFgc0lxJgup1/TrF77CDw+E1SMX2BN8A/z/Ow4zAFa8niOhOg1
SSS91ZLB3om7fp1FEOJMoTgwKc2s4SCYSzqokoIPje/r7e9fmj9nE/ExKAoogkCv
ZKihM8gfSJ8zOIPwflUzh8+gs2hbAIhL05KlN05LgwSiyF4UPv8HIguzKroS9YUE
AGSBlofUhFBZa9psgjmekR/bJRL3BgjfA8YeIaA34Ob6/HLobaFFK/VT3NTrgUEl
iWFyK+QFlVvlv6O3Aphp91Ao0ZLO+df8JSOgSrgR0KlT7VeeMNhEvd/lFrDZpfHC
+1ba9IC+4mQmejhVaL70onlaJ65MR5S3G2j6DIrRlgInfdGqyL9iNojWtg8V85y8
CJcNFTbpm3RYqKu5wnfukBNMZXuMCwwJI8Tm1wC767cljp0QbI1CH/QHedftYn/y
JCYtKILqGiTzkyGoLbzvssaBjnvB2b7Vc29oIIpjdLbF4tLPjdY9UO0QQFQb3JEx
IIcBesbzHyx5wQcspBEUxRTfbu1WiBlLIVUhlLK7XJsAXF5wSYFr/rX+qmCQnMpm
KotSbXIXJHCxWCnNMoV1FXhF4Jw6XwCexhhDc2o1glITf3/pVi16+wJPH6fT+eoL
rIFZ2cveIkeG1mtkEfqB0jtwTlNRehMsIzLe43yfF2TdaL3+3UZb99UDMaXXZW2y
sEiJTJ8IVzMPo/yfRD6pvOh7FLCsU7WpjWFPSQ0OLjCE1ZsV/rVOBOs1LPEmorwZ
vQNl7vSeF5euDkOcoYBXN+uiL7MuV/wDco/GtWA32YVGoliZlHQ2kFeYvRq34nIq
IYnxi2Ndk6rqHSrNq39Nr7a/F+WMteCKPnm0pLHYMbXLCF2CSF5akSCAaJ2Tc1+y
aVI9LAdQ9Wzaoj6otv49EWGAgk/PBGLNbYWqgVJYpRNf2bVhlH5o5uT3EFCAt+xP
S5KDkzFFwEDkB486dc6HHuOlpu0UUF7AzZgPC/xflz1L+T7gA5u+ShFPJqNNNJtL
Sn/kNbnw0+WxH0oqmgAlXdq6EEEDSsTLw48eEGOVP2BmFsme8VDEcIqroFJGECLx
MBSKRnmarOma1nh5rk1F0zHsvpnB2kPACjOsF41NBWequSl4KK/hz63KtwwCLyZ9
IXrXN9rDWgT7RaufF4C2xQGoard1sqNpvOjBDg7viqUKeRIl5n5Il1HehQLg4l1S
oDNMdw3Q4BCghD+VWsxHXyFWMjsid1LblCRpCpmMcKSsHgJ3WFkS+BevBpswJKad
jE+Jt5LPGxxuDYBpQDlT6wWFbj2Avl516X2qiCAyReZg/9lJJfb3ZvuIYaFXmZ/9
ZpnUAjXpkeyEUkjSvhcUk9F38gAUXjrVg2EzazGMh86WE6VpbDgwWAJqwsQLNSLk
98MliAUU1rwh81AygtjxnJ+j5rL5IrjOB2+RuvHCsYgjmPQFHm6VkAioq0JP8QTU
Tn64l/KDTccQGruj9u4ywmyIXOasltV3uhjo2yz4YzVM0ZKeRd+oH0j+nvhaoeND
0oHtFixwjUrd8uItqEQsVPRxlIL8pjpWSeOgdZ7Dtf2wOKV4odqL01/LHtZEcGu8
6qWnKrwSr3IaRpdPBlNN7Mv7HcSRPyNU2G4EB7amhbes0sljJVdzXrx3accgXedV
EruPbKT5lIMRi0AId34aamWXU9VM8xgh8BDqH+7PB1oRZR0UYsRdc/QUskcaTZOu
Pwd0e50g2HxTVLFqbFV0mujzdUSAwrZVL9SH7cItsTvsxnkg/a5A2J8//HGZoFrP
PjbbO5UHkdRYri2VlzBwJHQdGJHu/S92i73FKArzLJmRFKFM/8ErHcBfWyBJBLi0
ypDygzfO8t60Gv6B8mzG3X8nKOLR5hhWWIip8UPm7DDU+x5ViKCRvD+7HmOGqGid
PMl/LI0hFNs/6mhm1TmCbJygXQK/QzKT/u6ZL/62CuMVlot3XzBENus0RXhbtONp
QJopVGYU3kA7Bmk6W/AkDjKep6rrfx9XladqYDposH/rFcYokY8pV2IAMvZZOL7R
zBbL7AbK/iCM0ixjPrpk8H6l7SIaAFiSgGZw0qjJPiQCRgG9JhJvlKOjabKICGTt
TEmmveQvXcOMAsoYdnEw9SaXw0/TLp0mNGkddoB/62V7/k9jgtMZ17R70+u5KJHQ
F+OuZtfwlEk84CgrLmJUkRYw2iZWyYZpKN8mp17DPO9uLW48lrXqTHh9naAiacIT
s9Qg6qKJMIWywustPlkhLQSvF/l1YFFj0oMp+5fwlhgKI9Tfwz2oqldV/m/488Jv
NupPxmv2OhgswtFV+n+Vw6/9e8gf3gqL7V5dlnvB5gdkr0Y2/T1knFFC51lE9dOl
3WtPh2HS/tkt+AxFAh0zNbKL+/iG9FHDX7cevkdUUpTAe0/DMXQ9DLamtkwzoXsz
yolhZvwNU0t+xmibjpFCRzRMgHkcq/JdFMYrooyYJMN9urHW3c8IN8pukd1Nvw4y
/fDaY9dtpnSAeOFDwJElJ6L1I6lxZJzPlxrV8BTuI+aaum9mPR/fH/7/Bc1QcdKy
ohKncf7Rd+LlhsUGnHxqOzdxRD99ydyLBbUngtEF249MM5uXzXku1Rc8Vnfs4qnE
hAy7dlwp/ayfo3TCE2LkWhsKOzeCw7MwOIC3JffK4SeR1a8/6HnDL6tCP3KVx1Ng
D/7xJDNiLbuTlbWXSHVIWo7ihclNARLtIBelhuEp0ISqhnDWRMivJQvJVsj8F6cL
tiyBO/RZkpOdlHcgHJ3oV8OHmmnGuJnYssT8FOeOdJSInlCI5zw/YXfq8X/VOjUP
KPbYD0m/Knhgm3YNhNPfZGkJbIUxScDFh+DzFpxVMgbpwYkJItT+Xoia9bUtPliy
iLrPiXNwAQVuaNWQf1r+m5Tz8IauWa+0tQS6Wfor2ueIAVK+6EHdpg+INizFQ1b/
XNSMA1RrFJGZ1S5Y5AI9BOlbVdbWhWp7pa5A+fMBl/Y8QAvCW5GbLMUWfS3BLquG
DxBcdJHK/sW+u3ph7jtZ5oOMbI1YwMESOcxizw7OVKaJP4scT0PhS/Qzx/aduLXZ
SpTI7C4K5kdirmAExEQOn4jrWbNwbVFPcjWrKNcvhEcFq47E5oL79dFovvUl1ZGk
7VfJ/nLrj+iVKzIiXfCHkjMurZWtq55MhQvWXy/fH3QWQcmFyL4IX1uTkYZD2P1f
H9f9e74kXpQjE7njxcqOnNBAwG0Fp4HyqG0jdqdwL2JMeaFvu2+ILvQdZe/tB5hW
Fi5guO++qNUFocWL2p8T9tvmXGQtzd3JXoTI4ItfQsCe0N/W+k5H/C4jrWFrcQfN
tmZncgJziH1e7UkDRF2WK7hGM3Uk3c3uRBc9tbvVb3XaN9z6KATIDJ62f6ORBkZc
RT0U/5bXZUrpKCSC5/o6+cRK4L5wH+6DPL7wIV/+l0m4qhZCwJaJ2OX+hhu/46iM
WtqWT4hf+aq8WDhwAjmmdKusQG7vBEdNxHmkueck1GfN64jqf6Mfr/EWNU5eOxgi
EpCA2oEqeOqYttwaxq36JG9iI0XPBHIBNKOkTtPB+ybJCAClXH8edSAPhRjXtuKT
GR5GvrMyCNCWcCqPNJbWj3dzcgDn4eqioqWCEhvumzOb/x1dQYozhwAkAt0olbce
VLEhmDi0rZv6KUu3+HQ92SgnaWWKLlFwVR9HCII8fGGnwpIhdGBAb8pNrSTofQry
Eq3Y+uloxNdXOrSQU9H72v0RCqyPStD0kq6AW5kzh43+uZa/YHzi4zaoY3tuloTH
GGCokZfoOHMiVj3Saf2SU3KmbAjFhf2zFVBeg8hmzkF+T6ke794Qs9HWD758zghe
uRdjMTIFNrM2oUy6E2peKt9nA94fju1RE2j+tkl+cRpTFtL89vuhkPiR2qUvDRLY
KUsgpPtoGqK87ooYFvAlPnktF18iohi8xR2l67mZINgsNiuKEBpwqAvvrO3mk9sR
kTYr8PiDY5tdxOJcelm7IkHVPlomHzG2l1NAFJ/cubXfuQPRMjQgA9qIWqHWghZE
YRnUDFFT/jeUZTFZ2WNPHHRxWSvs/xQXQYiyWWNWvEGmREhfLmc1jpyyUKwEy5gj
L3aqO3qNH3eP49olwzKOtMAwcC24AqlufONNSpsSoS3gIFejvmoec0+TEvwfSK/p
+CD+7GOrzW4nZ69X64cioRDsh57FcYyGFn5MXC969hT7jImxcr0/yicOYWoi4V0Q
lSOYzErwUw0SQsD/zeDTaO1PrPyRxoW57gco9VDXv5cEfY5iu78cgZVyJdJ+/Y7m
gZGngVi+CD9Z8HeNHeY1ULnATOtHsxa5Vr9jgJRMo7FGTcDsmK4JSc4kGou6LYsw
GGB+spzizQJZAcTzbvcoJH4/VuutCZdlLWYy6rz4CWsVXeNsS+au4StK6/NPoa9q
QQpMc6C69yRWzVNt3tlHAdQNpq0tasZB7IbYR1/QNYXSurvLCif1gJyFUTCOXIum
t1t5MrMdvAW0FKdDLZ+w0DwGBgsUf5G656EN3W7Y14Ntu1Gg801Ua5Ifsvlb+vY1
X8f5QWfi1M9c25iRxrF8RqlXPrrxqOwHR3GyXNcW3uLvbvXlnCUfjwLj8i47GZQc
QLsokuFMP2lIoiSrJg3w3Nw6dkBdB4a8ngXvwUY2hEoaXxwcSjEyNDbzIPiizw7u
kQYDINSaFayBH/ckWXc731cbx/TunmjPOZvXhkGgK9/oFJ64oKkJ5q/cf0dOPnFG
w9Qa7maSbovWKwR2IY/1O241K/MMyDVUCA9FWM40tZwbnehWSPwhoWRKusmB5/Fg
/4pyV+eTesPW1h15zUC4FW9SciGw9LM4LF+p9e6s5PKptgOMGg6fU/HVzgIU7Pd2
gZ0WIkTNzCi3HaO4/ZnUT/iBVJpADPVGn/X3kxWzMokGVJKquwmPtEPMKbk/STMl
L+oNyGXmq4DoWYblaFsFOig+Pgs1cn9rCFNJsEip8sp9VM5e2MecW6fFHOgeiTXy
qbbBzbsb+NRI3GxtKRRass36Z2HHOOECZJtJMYc+EmiSdjanFNNeQq0mcKuPEcQ6
on6bbwfWN0VUbulI36KkcgtVqiKwD24wXH2d/pP883NmZvtWy89SShTjnOFK455e
LkfevV9k73fbfUOsSwl/L0zydJfotFzOJivscpzfG+zoYXvYwGR1FDCT+v8TBUDk
UT3D9sT0LxcD0RnB+35gMjRc4K1Nq08oaJWneis0jT8T6Aaqhu8vc5cLr+zr3fnA
HD+5ULe+wfAI/B7YddEC5jniW0Ky0LOo4M64jNO4C0EPCbwqwpY25/I8QLwCY330
P1pXWzt4s2x/RR0req1MChiZKTFEUkab40y5K49Ej+us5EtkYxcpPrY2PZG7AGQG
MlIOQSiJBTiVTxuwo3Ys5n08WQIPBI5urCAJlYNCrf0jtIZ5iHZjwr712bNXhK6R
EXJcB0P7PJfSqw00/1kEqX2jFbuqAoiPD9MKRK+Z532CafriVqSv6mj3L+d2hOV3
izjbO8t7qgvwXRjaKC+fEeXYUe+V58T0dzBfyuZUHKL5qnJSwL+NjRB9I40y4pSu
G6/fR/GbXUf4ImafHjpr0wLLLfaE2x0X47FHwPB+Ri9kMbxvRK6SVJ+8ZbVYtqxj
5XRs7z4sAXLwlbW8sdRZIRI2mdCEq+si3MqI60K6l0sJiHfpm2wvDDcTTD3eVKPP
MWZMzjA/wofiKX3fjMtKlQdLPZevsa0uFTYp57NyVHhUw3XnbrtfdOq/ChJ1nld3
0izX33GOkSCcdChpVpXo/BmOJIusA5LGS04p87byOja6jtM78j/pr1fLOvKJMsZw
e4BCYVsmBNvvoOVfFay+EHAfLYeMmjRkvTEBzXgPJ5WRM91s3Oq7WH3scAmYGa4K
03cqBJX+TlL83r9z/eksY1JBA3811OtzqPTksuBz2cpVaCvSWNJgYWuTOWOqk6ay
XLf56iLsjIrLyy9bRKikjNt5usEnVjOrEEYi+0Ot0CpTnBFy2kY7hMu9s+iW5uEU
cdFhuAdnppq1ipXb6A1H+ahYK7gzcxntEAihqokPcXhtUf5j73wtd2cLinNTbz2q
tFWy5VRR9awzkJZ353bJ1R+tJhdUUxRgeN95nGKs66kVBXlJqYChCu5BkJOoaWYE
1W/OGikUeoZ7ytBnUr2SnRAUwnKbD622aryhiMtf/vsekN+yOCMm5TNP4N/HkgEQ
UpiWZx/Z/uh5Vd5gv9++ZeK4QPp15wrDR4a+IUCBAKVUg2HRz5JtERLe49QyB2G3
ztDtcwkzakHFcOe2SCEPH0eYrZS0uN7ksjxsYkruLhAAbpo0b+sWCuQNNc77hx17
e0mX67RxQIgbDStdGnkrx6bGkFhma+mGqxvqPscNZ3LI19TBHfzzpeMxQbvhqXRB
EE2Uu8kcnm3XbMv3X0GHvVC1HpPJpTCXMArT21cRL9RUYitsCcg7c13t6MqYY4bt
PhI9zJdzWRpvD3znrlk+GPETROg0q1T7BOzC8PNCJxnh20B+3B33F7cuBfG35g5o
R0nyAAEUZnIMSf3GOzqtq4Fk7QlKCxyeynNGUpoTR6b5BjzO1TOegvAWej6AA1y+
rTmBE2pRDyFZNyjxxzg2DYuRwwq83p/rlvNzH3ezVji8KqOsgCdSmbwfT73adfEy
C24b+3j7a8MVVSg0gBEXOkaeZNWNZWZqA29uVctCPuWhGnmOinK9wzHvEAgyF/NC
2zDmZ3FTdwn60aCQVHX/3h9NEMTJJeJ8Skg70P72CayuYKfnVMFV0Ao+0K0SvfZK
qvrdj180AMpKoiM2w+rVBh8ZVw0j+2JIl4AXnM/YvjKh4dbZxW//+FVkXLEDZ0zZ
F/fqM1oXfvJMtbUVKBJnjIL++OqtfVzCDrixcvYvqzRGOllJhcz16GuLJPxCQbY1
rUBTXhNvQe3EnFQ6SUDE7VRLVaeiq/6o7AjsqsAUGNBv+OScQE68M2hClu9/nDfC
ckhrsDq/5Aie+nvt8AHSo09XneFG/uXmR5L885ddx3ZlsP/1vGpaiy3gZ55h/RlT
j2opjupOG7vSTxbwnoJ8debZjhKUiTQuThni4DfaEVjrc3177FvKiXhiicsq2VNP
1h/wvUN7jA/60sPqEAemtch5thaAZb7BZ52POCFgBWWg2QbJb5rhufp0ryivdA7t
29uZ9b1ACElVzhxSoImVTgL9poSnYIhBur5x6cRgGsM4KXzYJC25KucY2cCC7IHy
7eW7/JFwThFCRJgKGnGTJPMQichLgDtMqJ4+0Dj/lgO5lX2nRVH4IYufdHuGJevV
GAsXaw74llXnipSn2xv0wwejJevdwdchXexitnynJCp50iOj2tvLC80xSpI/RxDz
UXaR5lGy+xGT4XhihYoOzmpsVzzbd/uN/JFBfkOuHdKx+Z4UQ/mMbRzf6apa/Wkb
TbTBczpOI8znxxJohwcOobZrHMQIDzb3aiGzZpY2toLp1UzAhh3juM0TP1HNb992
9ZfPbZXfUKO+aSkL1yt7ZsiCe/fil/efu/hWSXG3nlj+LwHdQQ2+dWqCYrnTQO7B
f+2GELrcaKF13GFTjeYlyMBb7zYPoyemd7tHv0chD8ez0BjfpmgW7ehGHymtCI2K
izFOIPVlnW9GThe0LUldbH/PVMKPvEa0DH7Si83QXXRyZ+XDFxfRt43wZgTmzZ4Y
heWYS9SzwISuMXf06+mZo9M5vmsulVyAG6SDrpwst3GC51lKAkT3mJ2WXOB9ARHa
+VHzkGHoakrYWEt7LKCi9LAgvSi1v//n3Fcp93MYZ7ofPC8xZ7dl2GFyCFfwVu6Z
sGdoqIP3MKaIbnQ2vvhwnOptKbwCkr9rcj8IRzIF8A1+xgftcXCYga+aPXSV7bRs
+vF7lWGaC8uPvwTV8HP+OePF1HMcV2UDCpFDTxL7Akq27Z/U7uvwOo1I4QncgxC8
hDQajeGDgMwU4xsebqDT34+kJiwrFLlHq4ZM80sDW6Ewj74N28cyw0706yj8bIHP
r6pSgy5loTVXkHKqyzLHrXmzVb63cm0pg4W+d0dWvuiH2vH5R95jFz5tVPkkfaEZ
SDH1QmkjrEuXpuW1tt/XXMZ88RM8zoM6qxWUO81aGfa3kbEb+1TqZXasBzkuVOfW
NFhHUw1+0Tdng1rYcbCPT61aCIiPort0CVy/VYUvyz40WlAAkwFHAfG4rls3MyC/
Y2QnodTWl07rRa040qFthgggA6HrOXMLfvzhW9l1dHDb0/IGxdde0MdsD0bqVi5L
w8MsCwgfBfikHe2jlcrHpcgqmQfJSBlE4FREvdozxI5sLWZeAIYIcPNY+y+SGxzs
1xZ1A/+HInIV7Q7Y1THdD+m5ZpoSKmUn+iZdKLrZIUyOrKdmBuzE7ehI3f53ERBH
zH/hkKbWebH3a3RigI+mzUUsp6E9yVCpJygdZZg+kyImc4I6oQLvyryfLWTqeXEl
ne2ayPNqFKYJwVWGBAp66X/gEOMcXaCrg/yknXPk5pxGcIro+y/tQ8ifBMVniedT
E8Sqm1xZplND0LDfATSeQkXgGm1+CX2E+d4+wfFlBaBCSRnh1X4140BVq2S+dmgg
f7ejPV3k2OCzYRVywffYhpaoqe8EIQMqi/sH1cVujHJTWLltJnsaKJrvGnRXziSk
+L8HxO1GVPOC+S2T0Eunqkux1o/9tiqozUDQwHrweuoriFhq9wAS5E/4G4hkfh3R
l6zUYi3xHkf3/j8RGe/mU/KXkLBEoTob+3XsKO2Sg9hmWoE0+UZ9h275M/hSY3Mq
iU1uzOfd6vzcXuVhZJ+2LnW15vdiWYDTvHxexrNNZaFHPRpxzaEhrZoTDAN6JhBU
EcEX2qqqdDA4ghs8LqZivTlUwlB94b7DOxPZmI395UYY3PXQe5TXfqn7M6cwCehE
wdQA1U1ZWOjJOTtQ7tjoXUHlfvh0G1pgUzQMmj2Qc+iik0E6vWYRa/4BFqcn/Jl8
MgDAoHvURdgd35Ar5PqzQL98xhzzasObosg2FjiQsSXxuq6rSEUfsgmoYM8mKi/x
vaNxm2VuQlHMvY1BmFCyMws4jDOroakvLoGXV1gdRSS0qxdV2Azt/0Br8qyIjFgH
waNmBOxZwTZVJ+5rAiz88F3aUUcw+ajc52wSO8mbn0bp75Q1nkj16816E5WzB0gB
H/W03oF0eQ8Nx1fGdDHBGCfL5R04d+A8zxNjcPKccFZvwywSOdUM5hUE8zI3mc+E
hYKn2aDO0RSVopvxJHx961eYtEGnvp72CsgvvLtQzG1HoOnwkk5/M89XP9la5S9C
+FTHooa/rx4uBfv3Pp4042qbYsHfd5Sgi+uMA8GH3f3g8MerNqqtphxMjt+IlODD
b5jLKvYzu38L1JoSIdxxt/M9NyyMamoVKoCiv9VXRS/rhBuY8kbwWR0ZPs/9RDS9
WaAQPP4xDHNAIzzG7EUHYZokiW76eM0r3NR3rL1bB3CuWEVGCloNHkrUClzw/Cou
3rlhT2XR1rk8V2DDkrA+vF6IksOGwZnQ6AF8xve3D5+mDcnKCUzW7RCtuC/UX3bL
14SOaXcedIZxEibHZTAh8QiQRN38H1bPhTDml8Xuj8PH9/4a0XvcJjWz4GrcjSVS
rGyuLv6eFYZZtFwksIVZP7EIXwjxi6UIifHeAOzMUWuBfoMyHPgM+CUo5Fyu0ya+
Wcqwb1m99qVf21sPTMxee29fBphppGzH6E54IdR2a+RUFV6IxX3XBT0kBw4dBq9L
KNueut4M1Ayj0uvM85UfC0apE6ipqggexVX6o1tXFdbIjuuxHvz/1ax34Hr+WADr
gMjEiw67/H1eh/1i8spN4uEV3gw47EpWGPGMKBg5CfBuxHekwUvrVCXgSg0X/kt+
pHVQ77UTzofH/lTyEWqoOOCgziPHySNsvGLz5eEmiMsJxBaDgiMS/IfaMOpIK4UA
TvnidhsyVAtxrYWip1LjitbfVDWKtxjol3W5AAdY61cb7TAq2/ubc63AbfTtdClM
jK598/JXw3UXD4jYwbAku++xRoUx/rLPp4ay/aeWz6IqgClduL+IjK4NHl2PTEj8
RchNas/7T/Hf/257MW/ytgrUWYESvpzUT5pcU4sacf8uKtqwwDVV31Iwq9mEJcuQ
RpoAfQYjf6qAJS01gT/tmuL5EJV6GUSr/5vO2Y2BnxOuLluowVTm+uYbfK796v4E
ROEYq7Plt5eA7n91fjlBFT7ASjNMCW56Y3ujUwGMxdntSUOx9BKBH6lweeSoz7Ao
N5dlhOKeAnVVrKpzGt+doZQXhW8gHmMDXT/B+7K57Oici8/66EDp6SZmdXBvEwgX
PTcQaros5blz/1sYCeun+m443ZXk8eXp+9li50KRCYLigitU6CZHpq2tge1ZwMDD
Qe+i6P+It7xa24h8adGFfbxQVAA2Yy/LABBu1zqR/0YoQkGyxviRPgHrmFDHLhIT
zs4c5WKDRaYEbrYS96GVwwYIaGyEwIWwhubmTAdNmv1BzHrKmJLKpTNXpa4EKV/h
2NWds1wxJ0GyUAiuAgREv1veLkMJssW4wY9HE8TiYrwE42Gi/uCrmhXoj9gFOaaf
USLo4pMX62vF/vbpFbNGjRwDgSxinyhCPq61B8a/ojwDWLVdznXQElVgIeXrOcKM
zzXqzqrbrxQMJ1oHtW5STf3qxAMT6oLtAX5hZ+T2XMgR0rjCmc74+ndwpNPGIABU
gAuVZ5IDYcwsmYsqFq67sr6rFrwQ2HKTzX46+R2ZxuJy6Y11QqZHX63sIJ0Z3zzE
8b2q+65Gj5koHOZgmLBjOtNavgn5j3jS67sz0mEF3ae455ExOwJea8C0Uvgznlhn
gFLnu56gATesmHn4XeuMMWJxESHJDyLGvU15QNMULszwYrs/BOFxDg5ihKL1E53T
9NtOHTMSTfIYPJRbYS+xu77wkwQqOFqItWhkWK1Te4RHB9QtzWHihGs9fXWeZZGE
ixVWNr2+Ngb3yeOu5x9sv5mp52P0TO5rzx66iE70Jq4DvuraJ7S3ZO9guM2irmzO
KmbtUgBMARoQFoG/gVXB9jZRYH7IY5J2wtCj53DOut6x7vMjenGvuZDHhPXWrMXc
30joZuM+YMw68ztnQccWmZtUz67781rmvEr16/OaaAbpVUT/dMRlixqWyNWRsQjl
Rp50Uxfo8fUtGS/g7X1QJQr/RGyYrZFvoc1a7BlMUXNWAzqB2gAl98LsQ1SnimSq
L4CxXUADsNXOfU39RUPW6TJ4TiRM2OHm8Is0iQxDbj2wtMB7/EQQlG6lJ3xufy8f
mrHTuLLYq03dO7XdpVEBTIkB9vhpqSqDoxp00OKub9ElpSfYu672BekWTW7Bgkc5
4TK8MtoqArbxLpr+TEz8859420JMP4d5wIu7EqB7I2/Ltv/tysgf2L01ZQ5tFm6w
hVVhxbzfecgn4QDRq1iXJz+GRos/bm984+AFT6a3OmNFMQOB+WYXO6SMM42lXxtK
N6T3CVPzzJc/xI+pYLjUHAiIKVkGq2PFRn2ZDa7Mj4WGvb07horYhmHyAiZZqUHk
aEv9BYwdve0OQWbXw9qQe53MHb83B4b/F6OBj1gve+VFrMlVUJz+aUkITGm3Uh31
akDqCIvjd23CNhAQEMitoyag9iEiA+k4OXA+oWgxm+NuIpaNVqo4XJ5Fxtq5TaFS
j3k4faPdtDiWZw+ErviLzTUo/SSmiv5iYiIlBnSP14tadpKX6tvgNL113fH1lKXK
NlsPpgttVLfIHmi9btQeP+JdUMMRnIVmEBnPVIUc00fW+7MAM5lebGwxhCEXHjkj
0QwfgCTK+cd+0PgQT39pQrGX6h5Lb0VGzDYMj2qENQpBaT+iaZ1lWqJabQOZD2TM
hz7WpQ0a0hZbzsh1v7QxwfrZn0VdHcU4M3Ni4kCgO2Vd4n3RfYuFLtKriQavjrIi
j7omLUzDLsg5Q7PGRodBmy8Q0ZMGcpIDy61j7pYy5tcTWENfhq56vZ9kPp4Li5Vr
sQMrJleaViry2GGgC81ijxdiWd+GnbI5pUE6LZtSsr/TIfxdgcBlxEeOKLpy9H9y
1u/Mal8b+skCB7keokvB0yg7h4rzl+0RBK0HnfxoSrj//6CzDCmVKn1EHQvccl8L
2IweazFV0DYqBuqNTkR99lzbsa2qDyIm69iBjRo/xwqv3APTEcTAnyhFMwPNC5/Y
wRiLOObaPiVI2cpd/oCu9LFHdff00yfbJyzR9Bchk2h3DqEsNSFa2hhFR/zMcG2T
7f0v9bjIj6D8HbXTeCdG+ZLvBEm6cl4TJmMM4R52chJfkdXXQ59Pr9qMLpgrY8j2
+2jYUbXxzq/KvsMfGssiTFTPwx+7bgu6aK4N2F9zFN4LPseWEtX7cC0oUaKL5K6t
heqc+sa3if8lI3ycSM2hyzoCRz2KuqmbZNllKtmVPcJnDT5rEhr0dY6glE2/Ea1z
08wIi67w975SV/9l67RIP5m/Cmn3ix2Q80TLmhrXtCfgarcXAF0vyXqpL74e0Ubf
uQiUOqcCr2SRaYOVxubWurreWiJ/ydch6FagjG96w3u1RFYInCjBavrHdaDIGOKZ
F9yXjnvfBR3HIR5NnNrGiWqgbVklS/FXqI8Fw4P0xzQrtGxl2bAwvweJlgCEfNX7
w8ygLWqiLyV0lQynCJApzMIB4QRhgpaVi6udFkhp9+jxMyasKGq7xbIJWiYhpCtU
hZeVU7rXm6tW/AWP7t89udGsBA/lOdvmj6mMczE7P2M935OEy6x8Eh0tSjI4PJvd
R/jeBysPD0DlnPt/X8ARwEe7K/iy3V05Q/TZWguk1ST14C65ifF9Us4cQt5eA3ZP
CYF/SSGoCWL0YX03J+vcxYGuBK5l4+IsVcpoRlKR9HeXZHeMAgAU2c7o87QqxNEb
01usYR55VdHn8hHZl0aMZhGYvbaTDL/I31xip1kmmG46mxZIS8J0twea+BJenqa9
vE4TnioQyd/E8nRr8m7FDlMiSVUWJq1qHkqaOv1k+e5VUvUF/EMrGmh4ms702mDv
Y0eJVx/TleNBOyM9/b3b9SxGNG9A8Mmm7gcysG95ev52tZGTFzqileamid3akenP
9KGC63R+qMX7gqeKpMk16UxaBSxJut86SQXIZCRalDQEKu7EPxHkIZO/TuDzAECG
vEsMh/FQGlt1uoZ1Sr9PpHKGJvVMG9PpF8xAsSR+QU5xRdG8kQTom37qQRhtm387
rjGQ1JlLeF48AIREST3pmFmpyApqxwNSBRtiK+va3bKyc2DsfHS5zsed1QGZwVsy
0/Ho41aE+KkBluu7rh8CX+MdRZ1ORKZgUG3SDEmRnR7njLliqWMJdZ1tClp6V784
16pVRTVvF8TIcilqFcMpAKqMj7SBA2V9UsmPlvYLiqyKzmjwt+QRFocfdwBnanyL
CQmAid+/T8D0d6qVEeimNhjZLvU5cQ7ArqNam6R3ABW8iOBWHmahKWjhXnEspyAc
++PBadIKAMzPCHdYLfsQmDqzfhcXyhdUWf/sfQsOqFleFCHIprK41we6s2FZGymm
tgseLt0J+Xqqk0BUwMjt8VzTaSFnZjkEnt1hHXXQDVVa8WTSebZYRrU3QpTFYC7f
q/75Z5WbvUURZwJxyugY6CGQtMMWyLFM8OXpLZADRAPeccBdz+hX+t/ixd7FuAig
TLeDVz/I7eK/gjoyP09YMjh6S8vX5+W7o5agDPquzCqU53GiX97xCs9Ze1U2rpLu
2xu3DOmxkQKZ4Xgai2Z+94D5ADEDKMtZ+4hT1vf3lFxU+Gam+BGepUm1GUYBa8Lz
VsNwuRyU2f8gUY58KV39FljDm19duKYlmZ/QzGMGExTYhALK86n+W+hJJYIhKVny
iRihrdiSCiJAyIUqnSd9+agylprMqieswsJg0wDjE8NQ05vlvOY7qPaKMaNe/DP6
n9C+NHqtHCz0LtVJhIJEnfjnIM3Wq0HvTJ+IOCvbi+U4VIndfmOBpgQBRTROc1vG
lram7lOGJuWYh0reXOHpiJ7liw9oYspyvy3UHO3GCTEMngd5YwiFO8oD8N/e5Jz0
Dq/C0v3Emfn/dEUbGtm3pf0bgNonI2A4zlSnY0ZiuL43CXJgZ2bohJBMRCXIDVRs
vBQR+pLk5L+kmVG/uv6HTHk4SjPkmdRycuPnVDuDTgdzf96+9i/IlvWEjLEiRZzu
Z08J48b3+hHaX0uKtsHTvh3G2wiDjnMLSRZb1Zrrz4Vx+jBY69kL7k0Z/JyvfIjl
9EJMtH8CGxxrwgGYBBu+qYPfgueZupIUWxwrHNWb2krRMgenLO0gDy5I5atecYaE
VJDUWASyFyP93xJ2d0iZcfUigp48Ssg5/J/p/4qE6ZN8M98wQ31tgsn1NNPeH6Ud
iWXHTR4UYDVCopn2RzXWYwJGs0Uti2bM1bNcHBjmShgSaLEBTgDjvgskrlwg0C7y
sy4iCZ2f7P9R7YeQKibNq/hlLlhsdDq8hhQY436PtdRZ0CmBT48VxtxzEt2bXm9b
Nj73pCEVyFFD+nOcCwpUCvckb6TQMb3ta8Y9GnXQTi/trtsyLDxvG9WlUmnuGdG0
y0naPalkVAWB2aXz9XG2la5ukeJHgBL/KO7sUuc1kYFUrkh+imrKRtwhzn/U9ua5
qsV/D84mZ9TMNajZmorNeX5nbj7vCIPeYOxMEe+ZFZ2q6cuVG+DjbluL1knGbgTh
aDg7ZAjl6PEa0gmi/F3MMY18EfAeNwDCaz/r6b/Rjpmf6GNgAz2C3p3gxL59Hm0T
mff3vTr3y2S/3K9V6296lFF1NSn3yrnsUWsg2UVgEF+oXMTqqwXWdeZHh1q0zGar
9aml72HEpdzv6X0vIgbOrOkMtrJdDZz+tq5/z2qEGCGwnCGRT0TBmwHI9ob1eNwL
9tMmFtwBLeZnSfHHn25khdyv7tgAxIM9UCmfd5J472TYxq4DGj/+a1WiYSG5EDoH
9CgDjsMa589NqRpCFIvBaJESY5uR3sO3IkKB5g/DnIrwx29m73gbxgQzmiqDnYy4
fR/lDT5h03zwrXF116SPIuY8heqPZreweDbXfRsy2l2pAjy4bI32xvK7Ptj0paeW
80rNk2T5u8bU/XzPqpf9o+Z6SDZzK7AMsZ/MekRrMlZvl/ZWQQQJgnIm1T4d7UNF
OgHDE+/9TVxCewlkBjQ5jFr10RbgLLblWLtVC0dIlEaTCGpas+wjCiS0o+/ALfhP
iQC/WfsibT5Ni35idKhHxfwX3w8u4/was5yjwf4AFYRYp0JUMUnm9xDkKx4pZmCd
fd8FY+YE1pkV8cTjzjMIFvQfsWG+0UhacHqC0BiIhVBqb/1PBm5U52YhNoRJ93f9
f6OQXkMlCtN3knpQ+xcu+9b9cMeKiGRWJVrUpo+j67Kfngg9gGgRMyteTW+vF2q8
9LNrdlI53GaAHQ94U/bXJJH9yiduIBw62McqQm0nU24bHdAlfssnUDX7N8ebSwEV
d7GxptZG3cO7Yorc8RF3YPTVaHbjKzmukG8j88W6Q9zKNlf6sVCbiqs3Wpt7acaI
U6tRto20o7H6BmTiH0FRQ0T+tgUtH4M/aWxT4GNrCoFgyNUCbuaFSN9UtElt6KOb
lXhFKzYu4tZQ8np4ZPh058vLFPY4x/27c0SvIInPCWZER2ZD05m+GKykS1WGjtk8
LbHOCJZswKEerrltJkLC/4khVwB69bL9JGzXKVHi5oqVtkKrBERf/G7OgJ5oflNi
0Eu1uqlixEbFqvIKUm5bvq3nzeOSyl15rAESz/uiZKJLyBHUdwRH6PWqKraw+yFl
unQeIJH6G83Q8SVqdgo5p8jps5BC74o7mDOaCmPNnDZZ1+J0cGzR/pMsgI1KZ+b3
8xnDss3eEJanyTJtaY2KvrKEAPYnGgqFaRKwTYTENznTw9TjbXCy0LKA36UUR3oL
kIryjHoPltBB9I8jGbTilGQKJ/G4PacMmKWr8mwHbTRVKBpZY3ARf/7qxbdWF4DP
xxirnAF22B+ck8aaJqMrrWzTKsw95nB770Ol0f0TnRfNpRDBHFlbXU/f0bEnRcfy
hI1jIk1Z8rzzgCSUSaPMN+VBN8HLSIZDOhhofCDT9HOKqaudGgAG8+/WBiA4fRUJ
aXEm9eVLCjithpz+qbcjtv2y1EV4UUnUK+a70c8YCUwJGgNJv3RoSYqErn2hbGtq
abp/v0CBSCJCk9aubZywL4SDmVXb3zgAfjmrpFxLeetuiKMcIpR1zTiQlCgRatEt
9idSMLPo3e2ETxKALPpvbInBfqmUIgh+pcfPldwZIow8RGsXi3jGCsWa5RRtJTR9
tze9dX8et17V3JWBVFzpHQDQy5+cD3WXPA+/5luEMM2VqhUm6vr4EPYeg7MNQGWW
gKdYISAlxnKnUN/JaK+ZEQ41H0aOrfwr2g0+Yj4KUBRAApZvRqtsxQC0yzmhMBs4
pf3KqQduo7pJj8C5O57X0ZdLMGcrF6S4Ui/ajH3ZhEv9AVdtn7WcF3tGYtEZXuD3
FxK90B9rjPV1fgRki6Vj2C839VZ3nUL7wEV7N2DMJcMGkpe2bjrzEoyVrGhyEjbX
qMSEyN5eI6YG7OM6QrWIXoO1jv2zWbS+7nutDIdp95BNyFMxA3+4FUJW4JLT6o/l
LlbM/tjxNntycVXVIy+nYPR7FaR3c8u+PT3YPphKDpRFRCG8gtTBh6vfJyEEzvkn
Hz7mPSsk6ABbPX24ichbJ76lnNc5SRn4VlntNOXPnHQqrbv026I+wpkuQyXpH+K/
Vl8XqRnOBS6Yx5HttPVTbtVgVME0H5vtulsFDWZ99yRCxb+PwYrpTmEGgJY/KRob
13K32GG3FkwKHLC6aqcolsr8D7+c4nVMPuEDvIfAavJARcm+77Tj0sSLMXS1CT4Q
sNcTmj1j8yhBljjCxLLB8wI9gbip6dPNAbJp7ZIW3XK6xyr8j0Rk+T9CWrPZKxiO
VN5oSCsx1mqL6RYU1BvmGxNZXa0LHqmck0kyT8ioI0iZQ93eYIGOIACUMSr6AcgS
VfSU98ko8qpoH1svcUG6mpVBPlCaoiiPVa/fduQWCCDA4iQfFMK6ueIqL6P4EXZb
zOcLERfL90yUPoquMkWtquVHK0ckD9n/yMOJFEBWlFW1tRM9sdFlVCPWL0ch5dJn
V3m9nNZEmXTpJ0GU8pIK2mzUzQob0P12yQ6+vxwkAPzHcn7NXYU1EEdeUIJO0PMS
2zLIS+HOoLaDi5vRGfeVmiftrr/Vnka8L4wbo+Z+GZJCVzIUmOltMYtq7mH9/zeq
m0tltVy+g6Uy9zy9meh0Rx9zl68Haq6tp9AJKCq5rS46tJe+uTvSmKao7pu1bmRZ
xav9oQyeEY8G4OmWKhQjtOnyfmttrud/SJJggUAQDGEL3lzOhuLWalQ9QxPAWiXO
2z/vA9kI/Cp9enkXWEW/PyfbdPhsXSQOtCMLlLF/ZPU6aoZvh8P3CCbiPwlxJA4V
BRC1gtdg99EG2a8Yl9UDfyT76FEQ3Gw8RTQAP0jHHLp7zSLG3YzoyHP4WCx3UuXI
5mSFo7TZW95EWUuR5n57w1sGlDuPiXMhb5vandsh2nArTbhCDkgGh690zq8E7WOi
vyDx2bRyjxRYiVVvWHDaD45u6uKgOHOHHl43Gk7P3myCHGlCQjKrwvuVN/WcEXKz
EDhxrcC2aslkYFgzHv+dg6Z6nN1M3aOXT66HqyxOFvv0Y0KLcfAeexEP+ePcH97A
9W3ulS/QVSaD8m+fFpMEbTmxGelh0Ab1ErIllKxH3k1Jz9JRSfTYwHy2TTWfNBDD
AvbyT/uKZK7oLeQIGe+Nz+Hbl276PvQ6VEFQtsSMIGhFiQ00uYk+E80r5Cjh9VMj
dQEytkZMBZ2xJ8eE7FedjF4JR9q5ODdvG+R21CMPzN8zWI7G/Q2YpVfaHyQ6RIa/
dKx41VB+FNNn+NPDFl0oCf4qL3SqHGWFHxecgZKTncT8UVk6A4l5QW/zN9LNmrpB
gLCVPFg/DIOZ/TVoV4K/xjibpDY+3IS1nsFmW+wjXYjv5ADOvlWbz6F5PcQ4OVqt
9ZgRZCmB35MB+JeIhHydWR0qRwI6dIKqhRBZBsxfI0e/UlrwP1auYRCqwyJrME3q
/Su4t42xXENVss8eGpjDr/uQRmBen6CnTh99rs7brOk3PmvL/FAPkuG7Fey2kbZA
+AZX2uaF6gadfLqRlni3Z9AW0lNvj6qg0blTGBcDI8xn1VVSNMF8Jb7Bx7hslIdV
rIhyAff868wNAlLU4CPsIWsvqWLgq0LUXNWPzk4jOCeqFDz3N57gMTV8Qc5pZQel
apz7zlhE4SuqL+GLwcQWJ69xWNtw/MMXl9UM99ffJ6/oBqhSPqyvIrVGBsKMnDnB
ZXfs6DIjNO0CSN4LpzIh+qIYr7oo38cSXS/PW/u/8tk1fhea5eENhbgvOT+OTrBx
X+1F31lxznvrvFBySCpKSbkm88ORurm3/3nDSH2ZH8KqX7J4iHvir6kOlnh+h+hU
rBWcB7Il8e6nNfxM2Ofk2evvR5vXQiiBEJWY/YSU/woy3rcV8/MBAcciUp1kMBcq
vJkKThi5dPygOl1eC2Cuu2S4b8B2eLWlMlo3b6AthYsogE3jYpq1tnv6iAbt/v57
zzRWm/udq0g89q4UhnfIuGl9TCTs7LgBX16C2GqOOysRTWGAb+HvPYsi7/YVRQIE
ciXKzhAWPZ39jGbYe8eFZiPM93t9l1y6sIBnpw2TAWI+tTBlzUK0HbdQ+PSKxe+U
nKLy3f2hEQkAith96xZvhXyPzYBYDZ+5luUr38DG8orlAgFB9jNiIyWTfTKdWCuo
DzTTrDLbg4usrV9ynkMU5O7y7+ZHI7UMQog86grmskN1GsZ4Vxvsb97aN0ZvOsHb
Uprnd08EvkZj+/0lgS5NF+3j8K5JH0TWpiY3BYAi4P34fnpQ0kU+CFkSeLQ5xIZ6
7kys8XYnTapOWoKCQOznLV9mD5dfmy3mUWty3Q5wW037eafYpnvrNxvyqKSDOwcV
LOWAJiB5STTgPsujPKG+upHUgRPETgqCOE53dMUOjPXN5mbnb9s+I9+NcF9tYNzI
2cOcq0UEXU4sfDx3/f0zHv18gdu2QHKoH8t7JVtZc9PVvt4cmFQxtqixXYB1KVe7
5Y35n6rEQb5+8zHueA3mf83pKbY0DRJAy5+O2cto/pSQ/SyaUKYu+k9B1EVGJj+h
s/FtE9naf6wPkzp8CKKzPJYWFt1GGUWq6aT0wsZbL3xXuvaCcYJiMjwzerv1STdI
BK5ibOgA9KPKKjOih1yC3uYIyIChEajk/PqornJfd4CsfMI1LT/wjdwxHfa6FiUB
jYj4AhYrgLCYgqQSMKLDWIdVFXKD1JA2sEWasw40z2co9b0ocTBvVk6DhK80L5+F
edza8MZHVMKfnwgjj1hhX8I1guLB4bDP4XxO6X7ZyJjEk4ni8PXSJBFsrWjsZVhQ
Td6JCMTZojymKW6FvjkpZN1DExP85Fo53VNMwf5Jff2T5fWMBjvxjFoYxaimNoKx
jVSvt0rfbHgwMyRgbTSAiw+Pek5vwBrSmQGD7cRsKiUuSVy4q/UZBUhaRvstSbmf
7/IbwYuw9J3r0tlq2igEm/l58jZfK4I8GLtFufGBW05Bm9CzfnD+B5tJQm5zOUdv
QFwNYCpr8vXtB2gx5q88Zad5GW4/0jfGYvz/kIMSiVakpijS5yNr5DvpZCWpP0eg
MJ9ckw0MpSc6ilusqSWXCUM3zV0e9Px3aaqw+5siEJhNDfWq266tczTfGf+AY7/V
4Qoh9kjWkQArsKgRVqUfo8RK6bdWpgURnc9jCfdtR2Z201UqDZcMlSrdlTx+LxaG
LyUcR7MpvOSDXRp7/FRY0B15M3HyZRpkRC4kFi23r2wRyDo6TeHgvosJ8FHfaQsW
T5CJ67fe9pDhGZj7dRXmn9iN/HbA+R7q8RCFSdMWRViElbU6rLkvyrXM5WsxvjMX
OXSnDJAclH8CJ65oWo00wlbX2QxB5rKA2fSb9Iz0xqSKy1m7jL1D7ZXuXayi+ot7
2ROEGVIXbWogExwbrjvZ1CMHoUrPj5bD8+ntndCNY0ZMwTxe7Vv1dtXSige8NTeS
IKn457whEDkrloRxYSZAoy0pVwfOmtjwQZPbSgatrZFtkTd/iZwq8/2fv+xsdPpz
6aYoMlHFJWt9fjvPsHkFihci5y+xx1VjfqFNtRvdgg6oRu7cYhblY+0WTw8H79Iq
I5h0wt74nz7NaKuDlwJBecGEbdOGQyAknartBpC9UMweOoBGbAdDw3UeKKpFmm+b
WbWj/KSypUr1kyGeTw6xi2OJHSfedp29MOFhi4XthJLA1yM96vyhv6kao1Tl6ETt
JJTq/ChNNs/Gjut3COUvYs2w3v4L/OJ17jpzi9qyX7n+LlOpOzVW5unIdztE2xiI
uPzYN+yT6jByhmaFmpELVlQHZcsyZ/0hfyHKvrcAwQ0Jp7wqoAA0iTICUKTKRYuu
AzA3JPAqa7UapaEmI1g0RBccztKVCfqcd8WYfKh684U9gltS2oTugNyVBxBn9vh9
0ErEfcq5rGxWuoB16bghvlElQnwvTeGMXhWXyFs1GCNO9neDi05xDEtbyMPGcUDB
5nWta3SknnVsVqXmhXPBS3IgmEbGHPks3arFBi7RVM4m+EnB6tO124+ptE/zwaH7
IfcILigFuOENBlRQWWNlzQSmpg8DN17i/fY1w3q8Noroqcq07Re2Vvninoot/wCs
K/6BgbotX2IjqCPWZgH3uz1t0ejWoLb8mQ7noPknz6eRsTcxiMohw0wu+GpAcSR3
L6rgDmXfqTsB+Gp1jaFEb7AVEm7AsC6y1YvLrqMNLHT9SQLxnyX8iiBWNwdwo4Lp
8uLXsDkFMGfdtYx6R/8jIft7vITAdVNgo637bnDZCW3jhN3n/hKx1zIfZQ2vAq2n
8ekNMIDAf1ugX1X81os4wtoOMJ82ClE94hPoNuErQC1sOVJB/W+PQnOglM8iOZA7
z7FY0FRsjl4qq2Hf9F77Rux9tGMEdX113yZwrrnZLqNzto5StYT8vemURcLMH9rH
SWsIh7VpdtG8K6H5LjbL5ZWY2R2cUtWcRjIOePVuL3/EVkIl3SNwVs8c2vO5Aeur
kJgmj42VmK+hMGMK3+qhoEuJwbZ/WRvjHDPDQToiwt6Djc5PJk2/iUofqXza5Qv5
MP2KMkNrU3/km4tFAvyIwCe+GjKoyIQEF/342DOC1TsP5gNH1CtJYDQibmtUggaz
87ZcQJACt7YTPEozsrp+OVzr7skyR+AeHUp1zxjzfroXnkce5V3GR+AyDEza4MhJ
UgURE5Ws8UhabvfEQqyWlcn1zJ6k+SuODH1IUsV0PgByJ+jHu0HiwoLtS4G9w1y1
rYmWy4/4uUbS7LwQpnBoZMR5bzxFHLK4RhF6/8LDUeWaENkWFf+2cMEjoJ70+2s4
ni6HHS/eUkiaIwzH+p4In8KrCR/3CsLkWX0axcd4cOM=
`protect end_protected