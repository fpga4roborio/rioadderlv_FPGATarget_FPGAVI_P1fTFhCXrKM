`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
ddtXksX2+yylW5zu6QL2Lhnb2d1sD00763mmSITNX595NcHTEkwn0zB1Dry37fOW
FufOhVzEJp80NC5qZ/+F0Vk7Ik02dIR0elf3clrjeJRK85K4e3Hoo4xn7YbFUIms
l/8VZSb14+JVGURjfswrIyCUotIzlzVYZ6gzoZwDXIi5gQIBf/gI+KxNXPaKV+PQ
Ufys/12rjO6aI/pPlqSm0hCvftmBcnezN2hk1UeXgOIuKZnogjOsf0iJVX2aOOWE
6pD/psybjbnsNB6kH5uFTA5frkzIzkzl5d9+YDm9OyC+k84E83I/7/j+rk4L2dah
QJOvksSIzN867/4Qt8qYTQ==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="MvBXkzurAa5VTw+1JJ70nePUfoQXBvZOku/SMmg4TwQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
oRtzZL4VJ4iwysPsC8SXYCzXS8Fw2gtZTOskLcDV+1B9Nzn1zTyNtlo6lNICRmmK
ZRVu2BmCc2G+fmzynYlNTnSa7C0Cuel6FYpxCBlOuk3OF2tzAmLAuDyOH3Z1Yjzk
a0aHuoCdIRKv7BrZCdALt03JeUmXKPdOmIlkVGFl8yw=
`protect rights_digest_method = "sha256"
`protect end_toolblock="Jn9CQpRhJt4rnzZPRk+dOpzAubz7omckX1MrFd4p81o="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 11024 )
`protect data_block
gD6l00tciPUa6pDNTk/+t0OO0nC/UTtBwLB41d4inuAUA3i/ALrNyoJVcBnAmEQW
ptbcNp5fxEUJjnOxnedyZEuEBxWRieZFQnkRdF269oNTEz69Jmt+uvQRdP9qAmxm
C2beqHDsKYF6/baZhUd6o1Vc4J52iFanfopAjKpR5INVlv7dNFiVh6fJKBWfFI49
C6uwxRHFRWpoKdaRIvrLEBvX5B4WpIshp9/inn6eFWvyvjPmU26Xlsoi9rx0ztuy
07r84SYoPf9EoUYBH8e8utkpLpvOEY2y0hSsg2US2ZPAB3CdaiClKOrZfo/LQiZ3
O/r4Zjpa1myiHwumL+I5xSSwXB7ok7TbYZstTXmF0uNiEYGECkzborARcJCd5EuX
LPE6HkOW/SaYb7GVU39SXjHwPhiHtoZPtv2t3euwDSqOYKwUWP4Ijo96ISgRffUC
FUEachHu27gkpsEdTXlXL5KBFSZ56heKWZyq30pOZhJYbOT7ZoG/4GpcdZdDmWYo
/LHzpXY2HZj3dnVLHMSyqYyd7afHaihssSkvaOQMh1GYMA5VI0pC/LI0UYD+iyo0
LskIG3Bmiy2mzwHgMXm6l5KnPKxXTlQcShybA3L+y0r9Plj+TdlMwFT8s5ZuGhC5
vZRukHbwq1jdQuChOjDr0NBIXLvJH06qiCqPkMw+XbgwypKhDPT7vdKTXPGA8Rqk
NEL3mNxDHsKnkXKs3RULa1khLOERT9W5yb8nfe9SQdcZ1gSEbHJnX4mmJpbWu7tG
oWnDT1lxCe67uYE7QWwxjj0B2HE28CxHHahdEHAIEm/Hix+Ura4YVIbJ9dP3g8hG
chnxZFlJlMzwV3nqPL1FaYxTKXCLFXZi97S63a/APtqR0lA+PLkbugoHIqc/qAtS
Il26Fku060POWKNT48lxQoKtvASvaIE2QjrOtli4YGPBxHvCGtaHxzKTMEAiUIpf
gnxaDc5Bj4k9KGT53KJ2xa71fWm9mK3RUdAC/15JGleVwAnxZX6RD8MZ6/SV+qCC
Gf34lcA9L4nP5r8ttVgcQr1pPoERwcGMpnaNztufW1pC4pOtdkbnQ2HLQLaze8rr
uu/eCI4toJiPhUeq+Hwx03+akL4jLo7D0rPrTp3xhpickxWJvqNs6GSDuDBVKFmI
CnlHOhXvu65/So2+1D32fcxZPzKlINqxdsdYts819bV7/IwncUB2IyBIVm1LxBqk
lty2G3dlerhMu7x9IaiMQk1WsQwz3lGUxCCQkWmIETA1Ybe7yqPxhU8ka7FyQIds
hi4OFQN19ckDqRssZLYs4/RLNYtTWJFQHB4HswgNtIuJGM2eZUGtYt+mmAqVbEiw
ogWNBBvz/tseV3Aom5CvgXN2eQC2oMQYudUhcyQrDOZaUXYwJDpmDtAusGjaTEej
J1ThGGPEAfsA0yOnEV4nKY+YW9akK27X6saxxgVdyjBa0xwJ72EbSlQPec8SkPWZ
5jDqrbkC+Um0ZRiGMnnaK+lUf0MbDXvuI0Nu/yl6/lwQa9f+5yyXX8NCfGzWjwvW
buAOcC5d0C1R4HiYpuuxsn3QTumdjFj8yT032Jw9efkR26zyWMgr5V8uTGMtpPS9
paN5to3aIsUnF/GT5muoX0+San35Uj9O3FY8SP422SRc9KtYI11jakpZOYCgW2Ah
9K7KeYvnfkXHyLaP1y61CNixWQuGGzcVUV0cdx845Kt6A6kB+bAGsMxS/TI8x/Tb
fMemh6c5mnFeujDEEIkmAGrEXRZr0ykvgrPE77ScuyO24pXC1l1B57J9Tynsm+W/
RGpPREUsNGxZHD/DV5USr9BvfDccgm8qvRuBhJpEWwlsjT6YMKL3LzJfMUxT8d2u
JKWGjym6GFJNhQgZ3GGiMM0qrjUTAcYZRB+t9tWwPmTQmCJy4xzlLzkcv1xf3fqM
KDy+UQRhz9kKAdlm9NU3zosAGDb9QCVwTqrONOlN55wnHedKoKArRxWpmSYSxzRe
XIl1qdpw1zI8gOyRSuCxKITw4q1lkwWwU3PXPw32ucOGIiZjQ21VhDwNurtX3fBt
wESjeknva04fzuS9mDL081h+vqi+Ur2oTziS2gJ8yPvlmgeMAmSzAsoJhzNC+YZt
APIYjPQnmDfjCs6TCVOgmlWqPspxCak73ZmEeFUvx2QLoWJOxpn5fZduE8a3wceX
tR+EsEy98/i4Y7TWehpEyOMUwWWPS+sPyCrzXOfVvli/ErD85sl0obPhqy1ak0Vq
0nNYAS0lpw4rcTlbM7HUE+z4+nwIlSH2Y5JOb0xDk4xmFNchhAXDCX75zj4tGFoX
yUm4dn8NBO43JAWxFU8+gA1WtjBMdZ3DWuFhCTndUvSkhDNEjYqBJT7pOa4FLmcR
/nCkjJUya0RvxRT7P8Mt5Y8wjK8EFJrUzM8Vn1xCPr5jMHQ3NE2TlrDIMoti6YOF
3tEa+AuJz6tGuHkQbMY74okOs4qp+fNttHGGcJLYS8IbTgcNuetMYCGdqUs1NsTe
UNGtonahlJLAfKC8AvTAydETyb16UHHPs85cjiRdQBc+B/r9ADKPcieW5RJhHc/C
EEM7aJgc9LjZebomZmEAIB4R6o2YK6NEDnMSx9sKPs2ZJURRz9D9/fvOUHVj4Qtt
4QtV9dN7Kt33xX6qrXpvgUd9zKtz/EyMAoXd+dMZDbGe4C6aS3L8CtlD+ipCzYwh
ZHIPrEmb/gZArQoxKjINoxVCsCWYsd+nuiF7VHEdbYV68rHmDlpMmsb8ODjviXhI
cl9zha5HCgAbYIoDCCpzbo5FGRk4Zi+bSohRtTPWrM6nRUiQlu9wCbMgOS70FQDx
e+BeMgnKE8Bl+M6RxwqyGaopoFtxb49CmYN6h6hbeKkl6VY86uhkNx91qigzmFPy
rQxsmh3AWRP64IWapA3Rx/+VjXRSaiyIpINwhyzNM5i+iZEMVJyIw6pUTpLDgogq
K9HLDIPQNcA+mMw0AEycjESjjLm9hBbNIbaaJth7YLGXx8b9b145c04RgVnxcA0i
g3+j5OKlz3kf/n70dE/CDYOmjtPscXjI9UOTv7bCs7MYRH35NEI1u2al/b2ch0f2
6ev7dR7CVKGFVtqQYimN0Xi2OAh2GjhK/ZoOAR3iCA/5BK+cwMFx5YQZhDNjBBk9
IqHP1YlL48VvU5hVuCyDbgZQ/65Qs1dLvxq+op8mvhzqn7t67s5Mpw3J9mZd82A8
UOGNcId6nT0HFJ8GBsSSv5+wQrzYIzCFR4/4fx50e0NgK+PwRTqEbhzaH2jmiC9Z
NMMXTlDY+9a2ZZymELiL5wlamM959zBHS9Kl0gPjz2OV1PtMUFpSEkELn5yGLLUX
jTS3gAPawzL0lUlbsITqsv7DaZYYzJvkLMn74QSazEV79BgBgnj5s1MntgwiCI+Q
jNUI3ubCT1sdl3b/N/uTRa2qUmuoR09QfUYueTI11IQL92wu1t3ZJ8GhZCmYLBFt
ZVpTYDpHZr8+ogOqLuuJep8oPcEGJ4rFk5oN3KjQFtdAF6WAIeJ3zq0NhjdIQ8wb
M8vP7jZ+l0Rg6dRAMceXKEBiIw7uFpVobHnZhmwuihYBICphxQyGFimFjNpMOZQX
bNJQrYteELiF8onrrTs3z6Gihr9SZIFkYe3HE5dIaK0uYt2HOFg9MJYHnFUqEnim
pFpi1KrjLo4AdH2YMSUtdNXOPlAANAAakyPJv88tnJm3lHFkQnxwCXgPjLnrpqB4
6JYGV789/rpyTBj3o/1ey8R9PEertArVb+2L0f8DLNVPmvur8lXvjvwWG8k9ZCzt
Y144JJGOPLBxAzgaJ2JCcSFwsbbr1H1K3jSD+uH12CXPCbzN+Ik2MwCuW6ubyotU
0TEBVxEFmVrfYDCh69otbrMmjgW0sd10VnAP+6e1ZbTwGTZYe8xhR6g8WUNpwGwP
mfy8DxoG/EbOSibrqBsFMvHc31EB4lN9urWSQWDIBhD1T4F43FzBpFKQIr+gze6G
U43wWzzKR2Hlrh89gD+8k4AlxwEEhcdWdJFylVyy69hOtxFDgWEdp69IOiWht/4Q
YK5FZuYhtjsKv0ZYhcnFC2G6FmbDw0SuQDZGPYiNfO7Yjw+cj+Ef5WUhlbzMX03o
Bf7eMKWAuHS4ZD/Bvo6I9vbbeRLGRayC8S+6NKF7u/U9uIJaR8yAhKx1wxWh535S
OIJO6s+9bm71cg2cx/2+YGbvhjXVRcA/fgSG5MmcF+e6g++VqhtfU31i0Jp3xTu0
S+brbhgxFGcuN/YoIaqATt9w6NMOIt+w8t9VHEaTT4wqv8U36hKfKmaAs9RQtYxZ
gVU4ccZZGnmPXL5MCMu7kxQV8rwN6taqMKvYssf7tjszEL4zRmt0eibVFd1oNWjR
wWcaPxGJr/5ndOBa6Fb4XuFkHb00Gjpw7991DE1GPA+iKvci2/e5TmGsofQLLBSS
Cmy1/zo75qDHqmW9k7Y3CvskwiGOjtam53PLufhfAHPnfJmrsen2VWfdi1UilEWh
/FRrivOY1UK5ALdBL0Ktbyo/bZF+CTx462nc76WfU2mTbakv8jL5mmX8U5hkxSym
KZUEcauDlp8gbK8r5QkKrH1wn5G94eW7S4EcsjXo7WB8pMFTr+Wa5gRqxeTu33ud
CpgGYpCVr9TrHIQf8Q9OE6YQ3W+vVDxMfBMH6HKEr5zySVUeI1PgufK94kAieOWy
06ttMsjpCHaN2pZLMta+F4UuH6Lz7CQzGI2UecX9uAVLLZG4EbC6Wy4ybX500LOi
VaMlAEsame9Yg9wh+QyUXabi/hAxOJJyXIC8n8pbg7So3ssnI75YQbc1bzjQL3Mo
bHkMduJEe6FMmDkYHnMxDDm6+jJ9JYpxwmvVVyUGgzko4OnuU58RpXqUomUkqvUG
p3aB3vr1X4cl8M2OtiMNPqgPTK0zLCHKZthldZkbHiCUKuX5wdTOnIIXGIckmDKg
/rEbRDA9JWRRAdOnhtMNtGjCD0LDa7WyA6pDnxYuGx0M0kIlRfMOJZa6syyko5WD
CXF/RLmxPlu7nZd70zMO1tTZbg39p2dL7zxD371W53FSfoOhybwUDoNkrZ6okYGJ
H3hqlhu6Ix/qdKeCNAS2xmvzN8tQnVGvD4pQdav4FqRhuLFPrqrJrb9+s/YsQq03
i0G2NZr0lARhK0St/aOAdI/qwcRX8WSSAhRZ7KNNVYhQoRJJJBqlNKrnIj/Zvxjq
PmpQ6QBkpDGa0gGWksl+LftXDiFh1rUdlamcjmVdKZZRgWlHZdjFbSNyH7ggJS13
1o+b6UjXOp2U7u4FkkTG+gw+SUy//gqPeTxpDcDqRKx1llcLHIfAPkJPAyJN1CWn
M5w8JyovNTj53t0YW5iZHwYf/pARpicjU6gm1CZJD1jq8UiO4lQoC4S3xZnpP+k3
W5sbw3KA2vkdkAe0JUVheSb46BkRqymeVCbPLxuCyQxv0l2wRUctbUchZRC51riH
7Rgk1tBRCwzrewrmnFOzXj9CfRDIGHskinJlfYbKNrzY43rJR/IszszdEjXETRPM
MZjP1q7G8Y6tS7v7cjQZZUuXMSLhVxflSjDTBERUHMTa49ov8L/a4YBCXNUN8sHH
SN8I8NvWUPCeQ5AEzLiXCsnkVb/XsSrqow0NbNcyHWm8X4qrkqO7VWXW73J6GsE8
gm2XttEwbyvy4Sb24KWLCm3kwn4cvuDxoFtSQJhjT11l+erPNirvY6C/YJsTWb+u
RUwITuNTCxsR4vGtx7Xo6+Q/i+IEvVl8b/gYBguSvOOc5+oszH75oiSZMAooKMJl
BfI900UgJrltQIvVeAj4DrSbg5qsf+WsBh8zjQVFJqR11YO0GcPzLSE5HwxiEBfj
d/MSaxVs9jzEWFJriDzrDqJNCRzR5FQgeHAmZ9gCaWX7XADw9dDDEhhnQq5baNWj
/MdbWepsXu4dYbU4PA2PSnTUvN3c7M0F6g/0KbYJPG5t7qOBFHNhzAdSnf9nHrV8
psBdfhEGAxPbupwnTmWMTC910C9Zr1kLeTOTxRFX3+Oa6s2IKa4Mxno92hKRAwpk
FO59pZZX0Ri23STo+AYDj6KaTNwmbA8FUwTDMqjeYcwDp3x/q/sAvUzlnpH4Dx6d
LzBJ9Mk/KWFG6c01uJqD2g6PkSMjbUt44Sfh94zujWWZRFpGtK5VHMkiUJSR6vDK
BAV/L11bgDa5sxuhUEJEdMmev5oYPACiXH0tbP25lusZsD3AGUooQfbuZkFv0SCS
SbmtDsh2LlOzOl4pbl2m6L0bam8ADSjnrYnjoHDQXUALf/UMXSDgPWzY2/vbR53T
Y30ekMHim0p3BofZXSoMc0fR68GW6000xjJdcz4NE7z/tfPfhZLFNyOKz1mIW6rS
LISLu3WceRr+Zta063+pmyPIZoo3Gn7YPVbzzcjcYNrh3cG/NWwApbJBqI+f6211
D1rKrngnRjaP4YHoVTI8ijD4gg02gi4W7vjnvUOvBVJTep8B/XN0dD4oQMO4Q9Tu
TS7vES840gkAjGoxrDzsjpF2JJ/LjlOZB0Fi0usIOvSyKvYH5Rc46dGRKWxc6c9k
Qi5bFZDTQKM9/qkkP+tv438HH2dKxSFg/6QD3FhjdepS8nC/0L6UTUo2MTT9zlBX
U0i8mKrAWb6LGwOrI+UFx98KL0ipxGBA5qe/mreV36hTn2FCzJ7TeJifOfXJoHUh
nn8ZeCV/fmSpkeSRXKP9xHsT32mSQ/UvFmvHZgmB2feNHn7Sqmx7OyrnM3TEi3RA
tkZhQtkPbwXpb2TzInmT4kX1kcYZUBkPD57S6PNZu3YQWpITWBU/9PYRgup3CkA0
jL+dveiY3kJxsaHwc4CdLKhwd9LhNIScC8qBovJcE1a+Zq8cH5Q/NqHeG3xVKgrr
Q3E6HAPa4Iup0WysA+07Aj6mraJwJIXw4FGVjau0J+en6KyoZAep8nqr7peXiGzm
yGkUQEMe+crvefwNI18lEi7w5ZNnwIvl0dpbsJX8p2GN6JS5ytlwM8kKPnXOytFw
c3SunCU2xs095sa1+/N61K9OsKXpl6rhN+tbTzxRK9+tgRqIZaZ1WR/RuH/NukSP
JzjAwwBDL0OsQsOtXofD9m5v2crykDUvKIRFvsA9U+MujPXdUJIQkSdpiNdmVUY7
Ed3HEmAyMBTbm7mlgKVaqq6PnVgVC6iYN2NI4OvsETo94HcxVxL+qnPtU9IZY/Ur
8XqhUUx/GeTTZft9WM6Jo1cbE7b6ZqV61kwZc0Mj2OPhU1sIimuTS9mbb4iLnJCZ
SoH7DFoXD7261X4Bl8Gnr2PxyvmFFl00CFXJ8VliPwzKwAMMCjkvYoLtaxx62q2p
7Df7ddhnV8Ji2+6wB6b7nfaosboMo0Afv0/QK3eoNp1MteKn1YOhNzKVXNlKtAfg
MJ5x/+7yl0za8F3VWikp5p83YJv+yjf1EXYFLvqXYriFASTHfOgFyblWzVM5A6vO
0zlxT0RrUBSXgj4FJ3jg67HHwmJLWVhzZZ29aiW2DapjOjHnWigf50+prAvo9LSN
+BSE9qZRn8ECmva+p+ysDVmO2q5VeDXI9lhVjA/WmkN5C+HhIxcdZpu/ygx7w6Hv
bd2O1weJkRiGK42Om/rXwFGgzp8biv75Y4ESPMkpisY3o/J2dCdCgvdpMFu69uYN
cO5Kmgc0PTZ98NctKuptj7CZaOoTh03pwqo28yr6LoCPtxbw2r8WRXL7mTtw1wYM
OoU6mNdHnwlIGN3Du6MwL7JsCr1lvPyA7z9h0dieIuDbHl/iIUxTV9YSavA+P/Yi
dR3ymeutN7DjEmqLEOS0pKsMt9q+a7DkjreWZ2BdBctg9e/jfG1FUA7+pkVTIflf
usHqLnyOYJTXTqchg5vjzT8QoXnHEsC1XRdPf6GcT8q+LmeixBBiYPJN4SfMXujl
28DpGkRHua/6/vsmdkdx/OOnJaG55JEidOB4A8N59VQinzT/i9a5beeES2v1ko72
tqzBVGokQyu8sSXPafY1rQoit0bN0qcvEfVqRvFkphOmDtS33PI7bYBw3wD6TA8d
3ZRLB5mJdhf/ABeUFULLycqPm5NnwB+suloKnCQ0HvVkpZdO/PfVQ+7X0JQQd2M+
wSAnlN3K1Mv2BPHj/vCm7WZJEB1lKfL/+iqBv+Q5ZGI777GmBkSRiAlVak1+H7u0
fstOTPTmJMNGqZq3wgl8IRny0rlwrrzupFxPM8xJ2Ir2PVncBFFxmvx1xyQxVU4z
cddkXZP2dXiufFYytAJRjFqZ+FzyNZoLDVfd7sC5rfA+wqFms6vDh5nUWsmhuB2n
V7OvtVuvZRqT0lhlGqrzZYmOfxfC0w+9cxYO5Iw9LAui98ik7ZMtW41Z6sLgUDFh
0aOzjRXM3zEYDPkNmiHQQ6QSQ2WdMUntbXEbx2r/QP1BqTTV/aLWE0T4DJoV+EPj
rR1dXCt43IjymfULCGmRCrFFd1YTkjEsuiwSFxyF4MJtVN857La5LOjBN7Tw7JF8
vgeiu49H5cMH1xiy5jpdeyQFVO9CCcCGArkX2lOb2+zjF2mJSYXeAFLLp5w4RibW
3yaSEatZvUipX2NahRDViLQy0v+rEV1oNIdN40Wy4aiXhFelTB2XF7u/XhvYlIGZ
5t7IEDQnTeKpKGq4jMb9NVU3LAmAFjkRf0UA0w3Np8vTL4Qx0lKOZQoQeTGaXHNo
dgQ5UoRaMnT6uqxjWkuceZjCF9IpxhyjabETgiIy7h22AWozubbiKJzbLdeHS3T8
rOGz4qQfESehSiI9OmrGUsT09JrpaPnFMKMmZIItnNdNGWcuChCRj/DxnLEQZ0EB
1KrhXwAoY9hz6f0S3Uxvwrzh32UamGj7PbWt0y8J0uYSF5po7KRZq5+CLqVQqvNG
1+II3rNC/fw1enGMMlbW4GQP7zxMLt9Ehj1YTHBkRAGzYj68n/Nt0VsBaFa42NEo
YheApxL+XMRLaiW0DFToscZRtckCHTTtMVFDTSf4bY7jV5d+DmvPg8UlotXQbdLe
zpulwt0CCIXK9zFft1XybV6G5TfcoTzn/C1r6moOQDZnwwWudx5U2rgjdZsLuQaN
oH8mpz/R8xmOwSBm7o45RVTBRo7r0aa+CMyuEDH6EHQsL65WG07Ofsb7hun6ewC0
AE7gmP41ccDR4uRfA7dskqnmlbvZoRIVc93BTNfrmtAbV3xsSEHiprUd0oykDrBv
JgYr6EgALh31/ATtrnqci+FvukH+vAcsoPatAnryLA/fdVOZYoh4/qey00rqybcl
LVmftJZl9F5t/y7ekt42zH4jN6aJ8Jau/KUycTljmHUEh6GhpHGY6I/rD4xl8dJp
gF3M870FI91HCN5IJEhlWydeOdADQt25txrRwfHF/LMy3/d9EyRUlqckUc+sU9vp
x/5nKudlyBYDUhA6TgvOnpDharxucl02F6MqQQYwE9h7Ef0lYWhR6bca7/nt7HLw
1f2FWF9EL6zakoYoH8U+LHrtguoPsAfR3HcSqDMdrs+TBWW5jIDyWsKfktCv8opz
DgnuhU5+/rBhcyPKk/bOYlNMuONETVlgbtcXZKubLRFKoXPNExV91ec+uhMeA2B1
7koL+1xhQ2ABt2eNSVBQg9hMhs1NS8VZk/dX6JakKMMoF+2DBV/APM0MxPzw5Lsb
9Qq5dSxz4vNWiXjv3iC0wV+260ybhSgrrZOghjbnk2kU/xgaqLQ/DbQoX69TIieT
2QHp99v2KQRpDEIDp7+9ZRyTli/wZNQRgbvb+6ORBXOyJ9J/lX3KRYEge+PoKu/K
kiRcf5ZD2YuRPii1/iOO1P+D3jJvaXIL7lf3WI80vL5F3FMV4VnBxaF8bMCEflLo
7UmIIytjAO9P0qKLRjtJEk3nT8VCiERhEz5Bi07NYcb2xI3uvVMOrvYV+kAjqszM
hxGPgfm6XE0iBpd9eqh3fgvi2D4qlP7ztuWIfih8Nzq+WHFI381yWAgXoIXApXMx
56SDJYNW0dm7t9iZH9iGEXj2Uy5dNmgCDoJF02KpmUKszz6kqJptgeVCza9gCD+r
tOq7RPuz+/ybw7HdmamlCv1CV59S3r8/5BEdXEN2RWhVXPTiNoubBTCrVRUfXWJX
tSiEWL9NnFwlfx8P6t7Yb2qCePvgg+eAi3zL5W3+yii/eqvHlk85Czw0vKHe2IXA
tttKYTqlwPrY6/l0czWIH3VOL/V3jrtHvBybkdQ1vdN2KvZ87MiXXhZPQDVdg5Pp
NQGqxoDDvs98nb74kKrMUb3+J6HT0xRDdLFzmWbbjHAcP3cMV5iJx55T+dZ9o0AU
/CTzGiWUPnDMPOYK42SsmKaMBZKFwVzFOrlUMHPMPCTqjyhCoSy4WmfkISYD8c2o
iua7xAgG9gc61NJ+PAOmxWj8t2k/w57NNSkKjmPdmET7Nvvlj9jJv1t+fO8SWIZh
rVqkz7p5l8mAX6D1/lWOeZF0xbJCEVduxo54LcgirTGmnSTjbnffeuZbgMWwTzLU
EFaLLDrcnxhDqXQ9gIzwCm0ArAleZ98EG5/rtIJxL6k4gQ1QTAu6uYztFMzcrm2C
/7IyZjPEJci14yA10AEo3/EbPpwhLzi3sVY/L5XytxbIpPIA0u2CeN0faLiIduwR
5Z3kWaS0wn5RC+b/BDxLuMaffqYFpPYjM6SkdkjXSg59PoMEUqwBSiJvC7PnJxlD
urBE35B7tGmTd9CNUhbz6DTPHHmVYDeC0gjy6WGYbQAeU0BDoy/kzA346k6SW81e
0Ww0UAqR/itBEcBF44SDpa2VUVQ0Lm7GCXUam3l6ltNxse8w1mHpqgjtBcw4xBg/
x+DzbGRxmNN8FoeY7bm9osKSV8XnGsCR5ItPXKg4WpPtGf5mXYq6nqsmWG+6edTi
0Q41+ApA3at8mIVCh5dZ+o6SrEYvzG+Qh0vJQdYwmwlEyWL9oOlJzvtFH0reNR5U
xZw8hXVCVpJWtT3NyFIrBrH2TqR6t/UJZh+sPs+B8V/qXxu+b7RLkt8bOIy1FfeH
JMpYV3wJsolHY8cxdm1V12cPPtcNr9WFCTfqe1HCmQPZIM/Zx6nmdBA17sDrUFln
hc0u59UQi2DUIDTHauYwwZGZAeK4G/hvuOj5Co1ewdQZAd6CNdO5NK7BfYFJG5tJ
T/Mb67NLho4O45L79tJgq6VJn7OGBOY3fV9TIenF638CsDAU9Djt6Xfs8oHuuVCE
OV+jkJNJzNrlSMhmjjA0+z2x/drI4A+EWEuE124CqG3/yUrAszKPVqGUKohk34LY
5IVaXWSLjiVjpUBFqq5LjWfzZ0oWOk7F/Rz+N19njXMd1a5obHNz+jdKJz6HJHmY
CRjNs9D9TnsVBmZe0Zq2EasPN3nQ+NJVQ+T36QFUAcOzmfm2mVqMa2acPOD6Q3yr
julPxjhYZ2xbOrz31P3T5JHoDnrfUbCqVwB8f6aiSChpxejdHUch0YDE1CVtWMak
dNiMzTPtBh6kheqnmfL5sowHYR+26oHrb1sqkKi1yXetOBkjzWwoBtsRhSJN9HTU
hYhMF6jskfyVWLre33lG0tj5U6Wk7bmc+2QyOzWRMSw3OUXFWCswXniUfPc9/mIM
jaLeqG5AvE5+n7k/yj4CaE3Jl12Ud9TPEY8JDzX+VID/BMf+f2FHrnXgkYmYCGDf
XSA0Umv7xuwVsZmLn3DaDq9ScSG/UaU8oW4F+binKRKI4k1kY2Lzaohdfs99HXKL
8r9Z7727vq3i8xls/1sgpWIe6iIOSVhvZDtl2fyosT6fdOoQPMnSiwdvuuxrVe5f
9vJhqzGqKD5rLmymQnb13m9MLb7LSDtHYeSFm7WdaSbWOI96UH7c9w/SyT6P/UvI
4O1HzYyn+JkVRdH+OEWD8w3tAZoBQqnzJ+B+UvvIs3OXWA6T3yFRHRkx0d9PR9Ug
jA6okHxGkqJY2/qA29F/BmLE/W9sZceGhWyBbxf4Mqhp8x7r3Cpv6kx0FzFCNN+Z
FKHejt0N6sOIsFJ4mjCoV0cTBmmI4iL5gnf9TO190IjGG4UpZVzIb9seZBEhSup+
QjtMxINReafm6DN/NVJYEeQWCz2YrY5cG818oBzeMh6DbFOGGnF+CnSDsmjlK/YR
qbbc37fpK+Y71tHqGxM3ubo8gn50kAzD7/xypyALv2GvMRz8WVvJLMJ/ugDJP+Vs
t9TD+VcuQRYhaboje5MfTpGkIffZWkTub/MEYTe7GU/7QxVvHtf61CYoQdZ++Fbu
q5OWPjQnWbaJ7Kr2EmLoHsgPTSkA2MARwvN7qep6uqIPK2/Q8ugDuuerBLssn+wU
bEU0BXAGSaFjFo4XWVx/pTHjQpaeF/fkk+lq0msHYCBqec/dr8n3Tld7LWls+3g7
cIlnK4L+08O5G4bOwbIjZG840R/t+Mzoc/L/k+QU7ffFmS2zDp8p3KK5+INtTXf2
8WHKoZ4izfEJf4lh+qGvzO6n7zWAlN6/rgz7IMWz7BAUsREIZDpwh4QxL5Ol5NDV
tvIYH1+I3a+q1mKursiPtXtTknC0dmdQmKAH7ME2NIwN8xFaN9wlTEDdQyaWBFzA
gtZYJOR/L1HzK5BtdUSDc8BBK3YpAkydL4qefsAYxcslHxeLX6GuAz575qb3i3EH
pm7rLc2W0vhSeiCcClwcVpEphqayHH/UpS32ppf1RdQMn1HKAbpjFMkQxf798/3w
J4uDXv8J083B2ZzPwZWPTVOx+AZhSY6/0Is0z0TAhe7TPN3RTqN4Cx1cF5D7dHtI
m9XmRWrTX+6P/HM8ZW/qg9umqskEZtf+F5lCUSQcyd2PM2T57ZBGzArETrlH4dQA
Vj79W3v8wyHa8lsF8c1YjOrx0QwLszhxCooJjpXWqJJQq6slcQxyazKLVDOktAuX
XKmoWSiamcZiWmAre/wEQX5iXGGxotDObK/UA2I3DKnOhCIb7JPsOLYWf+jbBm3C
0ZTPxA5MuAAl+h+t7e9xeNkrCFDxN5BJ0RM3FIpjqnsN/oduJ1sYuVcgAgmrp9bQ
QwksPwnMs5E5xH9gl5aCzpeF2T0Ok/Qmzgmc1RUA7V+qSn6TzJjkfO9/pzd/VQtO
snY+u06ixc+dX4C/BghpJWzvp+T2O/qkDwiuI4sC1g1pLiNabz4kB5nwM49yBLcl
8Q1Ind6auHXTG3g2jvkbAPJg7S+SxWdNk170hs/K7Wv0CyA7ElP5v/x2jNuRjX7Z
FQoJ/P1BDFS19AxdxR2vcBiJoqStx2TwDg8A8CkIxbgS96UmIrKctNKwiJqTBVIc
fqEMAYhO4b+IGMum6OUGUvMV8b3iPzSpiNRh6VA8+afRu9LeA+nKVCSb8c52vSCQ
KajfsK0phbHADI5gi5+/Gue994nE6ZGw9bg0diXpom9h3NGE4DiHbRCCMkczEodh
raCp2N7bpq1Y1QFiNmzz+37yRLBIXmOLK8gpVy5swDMFhm1WpVWQysEyv/jRgkBY
HRq2lcwNifKUYDU4kw8JlULnevFtLy2A7vcNZtKD00k+ET8ekiErKBIjykjMZxrR
fH5gEyt98rQXMbRGNyWA3UIKpiOM/D6lechJgOA/il1gsDgVFYy2ueR5JA6q9ay1
wA60G3NWBaoSPLnIe4n7/BjDG2Fnk8tB8I2jsY5BIbShNTW0ZeU4YYToqUsA6PbM
9AMwvHbED0FVycV+L8rzKvCeGHE9OUfim1d5JmCWeAx1DxKxg/u6qQUk5VYD/Lmc
v9MRtMda8otUPYvywIMroIewseYLo9tkUkKfKGE+BF9mMXMMnCt00st3VJuOxPfr
JY36OO6xUpmC/pXmPXqTsMIoE1wPLwZLN0tNeaT/aNWw/nnQU+G2tYLePGvKIhYs
rZGwaK4F15+isKg6vdBJTkMk8K9IKq9NeS6AEH0lRGibd5Gqsf5sjo3PISoXR7rZ
lzOeQ6HhFKFou4g/c4AKhQNCJFlSxjb3ENgA4sEV/NA20HbDSbZSgaQOvwqevC9L
89VNsywvu+SgpgsGikZXnVzO9Q4/JJtMIINDLeQZx73358bofJ3iwD6nSy8ETuDj
O73UlyeeAXHoSfSdOrejwwgu6lualYcPgH62t1WtIfSOiZctag/CgVG94N/1/GaY
10H4U4ZjAwPFpQ+rzeRsEx5RgmmfuCRbERZ/bIjpeqI3wnneU4UEW6iQeHSRAREB
gby09/4TH66Vd5hLphcajQUa6Zhv/ZDzOiVdabZtiwO5bFRnn1GnDUnqPqcFt2FL
KeJrdIuNcHeJzTpy+iDqw8MeIndkGHejhWkx1NiYT9fpYZzW6OIwVaX/ZXxW1jay
DEKv1PxbSqxWQhQ56vMOrYkTqiOaqMJbmK49F4XYHGf3MvplBAt1Vxq0PQA8dTlD
vA1tehdSVz4pKieShM9DAK5RiHcE8pCkbV68QhSPGzExbE1ASgyitNT13CHzQKYN
S4ZCmc75s9bzS8wj17Hu1VzrJP7bPyhmWDDQZBF+9PQpf6xbq/9F9zs1aaG8vqQu
IYHt0N4qhwqXT6Wu4ghGWnI4QOi0+A5D43Mu3Jr1uu+lZRazqJild+/Ri4GcZeTp
IBvk+O6QjbO3xdhap2QEL3VDNe3CGjSyRcCxteypZsqGKgP6TCY6aRas3XYIBSw+
B4XPm7jhsOwkA2J6J8Rc4qcto68xPQVQeAzaTAL33QJ967NWcMO9NF59w84O86H6
WgL6QeZ5GNPUxWGUudxgebwzlA01MHUn4wgPZy3CIDm1FXwL5ztyP9pxi0XcTp15
FBrPeD28LL2K1aZxq4NwEbPTSN7I1aC5QbDbSFU03co=
`protect end_protected