`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
ddtXksX2+yylW5zu6QL2Lhnb2d1sD00763mmSITNX595NcHTEkwn0zB1Dry37fOW
FufOhVzEJp80NC5qZ/+F0Vk7Ik02dIR0elf3clrjeJRK85K4e3Hoo4xn7YbFUIms
l/8VZSb14+JVGURjfswrIyCUotIzlzVYZ6gzoZwDXIi5gQIBf/gI+KxNXPaKV+PQ
Ufys/12rjO6aI/pPlqSm0hCvftmBcnezN2hk1UeXgOIuKZnogjOsf0iJVX2aOOWE
6pD/psybjbnsNB6kH5uFTA5frkzIzkzl5d9+YDm9OyC+k84E83I/7/j+rk4L2dah
QJOvksSIzN867/4Qt8qYTQ==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="MvBXkzurAa5VTw+1JJ70nePUfoQXBvZOku/SMmg4TwQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
oRtzZL4VJ4iwysPsC8SXYCzXS8Fw2gtZTOskLcDV+1B9Nzn1zTyNtlo6lNICRmmK
ZRVu2BmCc2G+fmzynYlNTnSa7C0Cuel6FYpxCBlOuk3OF2tzAmLAuDyOH3Z1Yjzk
a0aHuoCdIRKv7BrZCdALt03JeUmXKPdOmIlkVGFl8yw=
`protect rights_digest_method = "sha256"
`protect end_toolblock="Jn9CQpRhJt4rnzZPRk+dOpzAubz7omckX1MrFd4p81o="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 15504 )
`protect data_block
gD6l00tciPUa6pDNTk/+t0OO0nC/UTtBwLB41d4inuAUA3i/ALrNyoJVcBnAmEQW
ptbcNp5fxEUJjnOxnedyZEuEBxWRieZFQnkRdF269oPlciayv3n0PZT/+0sTOd1K
SoRogn5AwfD70cFZsjz2QF3chqEI2bN/2NwruARVS0lye0KMLhDCqXNNe7Hn64YN
HXJV0OOSJouNQqQWfun2S33W9AbLU4JZRwVSF3faodGZ2KGM0LUiBGvmvKdx3XFj
sRr2pK0qTtqHeKxNjRmdH1NU7Q3tpJTbYyZOtOoJlqB8I12YbC1p9nC3Ik47+Erf
ezbP/yMDZJfFYc425+IsWZ5Xmpu+p8JEmG1ozBBs7+e7m9aVzcHq6IIpFC0q+G/x
tpmA5fHXfLdnDrtVgYGY+8hL8CH6iKAbj71QbTMLARH1yc2jSs9ykzt9aHbzysgT
9hfdWM/KCkaSWIPRTgXEuP/ztQOdARYWyh7MP5F3CmH0tR+vpaGuNa19CFCUY0Tn
Hw8kEZxAmI8Eh5oV0+ds3Fy6fjRGgZPzD0yNu71C5n7Sy0SOeGhJMKztgehyulba
wLW/yxjf4dAo+n9mXRvUug34mZeShlagb17xeQZXCUdbGtm5JSl0+aArMHS4YbYx
BPp5bpM3AvzbG2KMMLhhXj38VAwBf3LZLPerhpMlcQizTj404z2BNbzhgXm3Sy3c
iMPHSW3iuwte90Xtr3tBuhgyQdYsjizNwli6wUfe+IJRmFSm/c60zSDOCheg/EXH
841kr1fjcJkVPYrwhZ0XFKpStVNNBUgd3Cp1XZuqE4Hnngxy9WKsAVZjmifD5+Ah
sI3e514ayGz0pYQTyk4St9vwqQDGLwVuE1Q5PsOfM5ps/3i4y9Af13AV08gzLqk8
4c68iyDgyeb+tjSaKFeVvEjMfLl4D+97DJlXgYaTveUMclHB0L0bKQbDIrUh5+pg
1yH69/etzIuvmy25YzhQUJXk1demFAAQc0+TOdItNu/yCMWXjhlsT8QsL7hrLcNd
ifcpSnuoR/DdpZtwYZ+iU7GlXM1vmNfzQftsKVfmpU4xev6yGL8aIQYouINe1gtO
BIR0bi0wFBp4QdoD707kp9qV2w9eX3xV4VCfHdtK6EGrDau8nXWAjQSQSsUWRXVw
ZoCS2GRX44fpB51uGVaPg3xHamMN+AJr/MErIAFX0kMF3Wz4PjRYlA5ZCSkkz2Uq
asxNa80i3aMZWSq/yV3620XftJ7ym8CBng5IWqdabNIAbk7mthoPoblNuiom2Qpa
Kz4f61OG4675rnEEuBf/7HC2yEg/vgV2Zk2tLNc0tg4gDeXVV/rkrUhOW0Ex6xCb
YEU09ES10dv47Usxo05HRaoBGd5IUP6IgoZ2nlMFxICtgRD4BdRb3mnIIG1AhDoe
xXuE1Qz+zvaOHIRQ7j3P8U3Y4PwN6PWHpN7t1WC4HTIQ7FsEo6WnwjO0F32SVMrv
SJ6K1ntmAGSaBSWxhNw2AkLseTX3zpWVauxbhj1IUXNcbbx6uth4QhsIoOApSPMc
a7sy9l7tIacQ5kXUIPYGZDPFxCFpIj/bfXSlcpZYypjGRGCg4riy3zkHjHxEOJY9
+jZfnkLRMpjIQu40+pR0KAXX8ru1u1nAvtGtUIUFLVySiFSycnaRhL6+R1DM7G0i
3c+9QYhMdnqqmTUnVf6zZ46W8oNfoxyUQLL960cMZNz03BudJ6c1oh71ky8pULep
3vIHLNlcR12Qaw3qTsZtbev2iE+3Ec54yHwPGdPz6kzQxKLkNysEdwIZ1De1zPF3
nCprLQrggw9nA/DzMg5LZt3c5JNVhaN+A4sSPjjJaiEcN+Il4MhyPJx4qKJDjDvh
r5rK/ru/O3SohbOXZB3VOVsbbLOuY3HB6tAp3ldbw/FK/d1AfKj60AOayntDH9f9
FTYN6yV/SmfbGl3JdaHQIm2Xx7pGbIMFK9U59B68TvrRQbjhln/fJhsa5Z3foc/t
4oiA1YXHBBO1eqACtxvDAFKD0e2/NSUFPM7TdWIPYON8TaYIo//1UnjHf6u4whG8
doffNT9Jd6aWjekUc3oHNC9bI6Okk/4a7r6SO8oRO0Id5GMSLyWgH7xwlBCOreI6
wb/GCmCRewxtcMDnHJHwSdNLxZtM5SPiTvnRoNmBBjWXViGzqOkXqqFcxuexcwz3
QIjfenV8tjFeJ30h1WHV9b7K9O7kDamlTA/CSJWI09fyzn/mooHxLYVXEzbQqDjj
JDTq1iD9NSUHhibd2u09NYa02b5eegH5s/a4BjVwOFs/C8fPCqLAEhycMreqGE8g
URa+rkX+2v/+8Soo6KCN970CC3iVeM+rJbFsLG/lYHbKD3MJANA8Gli8T1XgQraY
FHI+fWlFrFLtcwu0ANYih6VJ4UhytaiCsUk1H5K9e6r65bNJlvMpiTEeH2FhmtRw
V/sBSvwRhlQrpX1heeX8crZvkNpS4ru6V5yTE2ubEF1nHuhA37/HhbUDy1tILkZW
5RwfODBx2WzofjIoXdPvwn+oR2D9dEH/kaWdm5cXZXrP1Uc2ryyP4o2CFovnRgsn
BK/vjLrBtFNm4fLujFlEntn8H2HxsYQC7z5w2uEekuVbFXJXmnqahcIHaW58Ys7o
T7RQaQkYph3Xyh2DGdx9DoGbGsJPkRbHa2LXunCwHDyJ3OHi8iv7mR6HemlD8Cym
zOwYC25/06+ybcvS76mg/09Tq/3FF6EWfkFQeXrkkTnnZHnLDPLTiaKStpWqmPUO
O8eZR8WipuNH5JldMANUVwRsythYZgLiMLSF65yKCY3p3bamAyMIKHqWFMLkV+w4
hksbfRuA4YuF+IhwaNDHN5kLP4efBIlcnNnw65YYc235wenh3oy4EqNsSaddakUn
vESY+7Rn9kjnXYPOhrSG8cxxOLFm8Dv5y33+nWJB+edU3dxwLKLuNpImqstGzEiV
0qmiyQZ3M6LX70Dn4WGtAjaSVxqlDgWD/8kO4ktmkQyeyYQv2inU1r1F5nK7JwxY
9GgLzPhRVV1dITx7QFy9q8U12LWrHIrk/BE6LsQhTodz+QeI/kW8Xd7OG0kIJ71A
657LfETBT9qblCliVDI104IAs+fGgN3WpweXf9njSyf6mZKkLChoWj8SM4dcRbOU
2JMUFzKQYPsbnjkA2dP47QWSRwKCNYg2aoMdIKc+PWn3YT9dq5G4AviiXLttIwF8
EqOIqaulHv76132049Por1MLcM661TpYbqW7D8ds2KLyGAlHk9ySgf7C46VwtbOg
UrlEkDv8Li2W2AWhM6ASHqAMRKxUZzn0Ck0ad26fyIjWHUBYfbQZmg1jPqPFpxaE
c1CZ4Jr3eV4oXL7wL3Hj/ydLNcBhX3ueqZHAFjXMIrKHw5CiTigLUGJW0y5hoQN0
iUQjGhy2g/EUZxDvqsdOMPWv9BmSetKhAIKAV6gH81MbOLcQrGxnSM262fXGgdDV
vMSO4eivZQRsk4LVUFI7OYjmlqq/pWoLbyKEhQWw5gLNiErI0TkTTccUuUI6MIGb
lm5vTPqPHVPKB1ytDE+LslJS+5I+7TIxQ5UGrL8gFa1mFxW+UTW+Pw9EiwBmBisZ
N9mxInZn7qP7sCGx0PC9d6l8KQGgLcoImzVzYyi6HbBjo21ASStbOq+sMOveHOKW
kHkEx5vaubDdyl7UsVeBh5PAnO5f5S/dL/lsmf7iD0ujRzvXdy07RXU+4ll2UEcB
l+yIIjtJU50geKvvuhPGhhFojW3YY3p3fIDxsJNb0u41bvSH2R5NmeH5ZOZPrZrY
Lfihk2NAk4/zHd+COdhWyS+wrUCfVfnoxYFBl9bng+kqdB/jevgJRcr7qo1eDwDS
y52vgvBslvLYGLWXHisIMH21QCej1uiMmLg35Za11meuPVuUPSYX0/H/bwCWDQb7
1Sx83OG4SWVG7i6qzBwrjNDhDvAexapTVdESCHjK6mrRfRPXPochqrgY+WE268mA
rnyf8J3Ws8zV5F0JxgBgr7RPdcDi/EmkyS1L8zGLk1/DvFJLyvW6SkgdKfuidU5d
H59K1VxMpjs8F81i3w+0cD5JDyH/tYbg7NYmTqMMgd5braYDVpH6ZgFnX52AoJ6d
SfaPg8LhCQodJJlazRhPTBBVoTx7SknPqCGApmMyUIZMITBUtL/pkeIEDKN3Sz2T
8Bm/7MY937GhMJLIkM14CrQ9j/hwS+Q7KeNrfp+Bca5XVzM7pwN0oER9M6UAhF3T
GdRQ1pf4bZyhRmPIyPCJ1VUFJNNTac9s/SlouCondE/FMmm7UIEsdDBpjyfw1QyX
6WOTk71GZ2PhLwwbYWwUGe+2GCjrGDJMbKEp5GfgyItMaOtAKrKPZxNAvcaF++et
VMzmv7V12kakN80dfQ1TjVk55Vzmqd1dto9Wv7tS0HTAn29/lN29r+kiLIy2aQna
ep/1j2pC1jWFhkbaNtvgPJRtuq/OkzSW/R/rEMOnluNz5NEU/Dzcxt/AuqqNewsy
jf96y8PxBPWzBZXxg3NociWZsouMi+zkxLcVla960Gx/W73zhne/t5jTDAlCK6kZ
ULmJkuwsr0FNDTDXHVGUiItPEr4t/Hf4u5YxPwvBuKnp6lqUMg+sN44U3ZWtnefT
OqvXcN+nnocCu3boCF9rOKvy6uztnp7VYReV86ZwEztauJlXQxwLVaR2m9Up4988
6SFlFDbOYmlB5w4UDiD0UnYdRO+2IKo4/wzxOFOu19aWFJ/5mfxXv0tnufBI9Nc9
qu6vCOwHXA9FUqdXQylW7hqIl1OqxNySVsZcW+bLlD4yHHmEmOPPsJT2YDrq5dny
U7cuhFAI+267YVthDEoKyH8feQH8kNF9LVsClm6WwVYh0cHeVTqJ4pTHHPloNaYJ
54A6HrfU5v7O0l7gJs5UAl1O7I0TWj28cb4MyB59rnES2/XB+yzJVFDTkR5X26Sp
7l76joNFSE+Z2b1vjTnwr+gqyQaHvveWLDZfrePloZNjWZX5y5N8ryUJOwHPDs3y
Jflp2BcutYxr4BR9fjo79u0gcZCwJyLFrr4UurcV57rF4g7CAKYeGUZMykeUy2K9
YKSN+j8gl40mvyxsRO1WUXNLodxhgUCnm9jpPXklAe7fzOG1+ZuE2jJ2sa9oc9R6
Zc33N3k/XGqSqqJyg9+zrk44Z5NavI9dy7u0oFckA/GJbtVqP/Qrz7nDQc0uWNKb
ZOci8j1KFKBP+AnpGUauJWP508NnkjDQJaKQfbM/FSfpY3+bNR0agSDmtOL52LUi
9wfsPj15WBaNFda0lfUjD2QjiV4EdFgFjKvo2Brtw3zO5/vLHaF//chtV5PGSvO8
ASi0GzRa7hW8H23eoJnFxWEeHvkiMW3/s2cT+m3tUY1ln1pzmvRenyNVU3Z8508M
lE9gXNqmFZna8/OcCSYZUrtS2kF/UxU3j5GMizannFOGJGAHxy6a1g/+KKW0XWBS
i4/zgCm+1xovhanFxvi+HZkMj3v4vZiuva+xd7NY5Bcmc8CwCyrCZoxlL6jtrdVs
DMlwytxdmP7CthDOBuqxpbyUjO0wn68ELMpjm1vUbV96a3nRyTVvafCIKDXgX4GZ
xomfuDos8ZwgJjC3fLsZsWmFBeJoSOAUYAiSXclSFCnb3j+yXb1Ev/+MiKeUVVIN
Z6B9hOPdQmtZmXdYyD2DVx1nk4Wq0fHS+JBRBSaJvSlbhgm1gQJ5++5dAFtBrHEV
mxnXkBw3ciRnDJ3kFg4az6mAkv2xucR7v5E24cXZKiQX739s762Sv2t/6fSDFCfl
wCj+KHRkIuoWh4W7FgHSnRbl9P1oIMcgsqVsigi64LbbINW5ebBu+g+Xz1KA+b1C
Y05Q26hjISDMSFi1Zmsd439MAohVwMV7/nFRtvuX/jbBS+Mu0BmL0apyg5ggQKn0
u7W5d0xnHu499vh16YAlSzHR+ZiHi8LfB++ZZPa5Nvdqd25eiFAjDokGMFktNFy6
8ojpQ/Gyx0sivAeJ2KUZ0/A9uxoVt8pbuH1GoM9fA/BMt2+0HFXEItJgb0fOxXW8
cLDBM6E4UmtscOuUdZteOWIGNVrcy3654iy7pTGUX53ytS8oD5Z8NSItJ+/ot9Jw
9i7E329asAWXog/p7dMsc6Bb/QrdqBjECVAdhLSWKXRtbmzstIbKGkvB4NWobtjy
oH+ghC+lrFkvmj5/VsmvSTUUnntJkcI6r5cdfjoPKbzcRvt9NFBe+bmjKtDA8Yvr
d/QQfx7KZz1Lww0KqnlrWM3Q2kiaIIFAd2jJukUEOPuU6civQtyedlnS138ie5LM
1nI1U89FdfrhsI3V7mqqVtTZuZLUZ7/jW9PZ92QbtXDYMFujZBNQzbU8Gc8BMV8a
feaQ/NHeOW/GV0eUb/Saufcio8OhDvMzH1F1N8vKT2mJLPL1a/ST26KYi1DGYI0D
KGwqM43aNXPr2L+8yZzCSy0OP0v0uEHpzB7aJUvrFOqlNbLTnXXJxPLMnxAUzKYQ
yByJX49QwlJSa4OyhEhg5bk3lFilTlPHYskzsCUDOVYom2B4Y+ij5PdbDIWwRdsZ
9I8An/c7JJf1KvVzcMpZGRDyNwziYH5QEUjyk7eXOl6bu2HXVoQvoVWxtZ/fvTOQ
pFONdYRFl9skmHbys4GRPhezg7JerfkyUBQ3aU+1XWwhh8+SaMDYhj4ZD+p/Alg6
vTGjU8rZV+fzMQ/+mevwU3MPLDDg3gmbA5FTRq1OwHJvBsUMDn5tKvMjx0/vX3ro
LN3fNXIi2+6NrybBXRAJt3m72AX/23bE8Rcs7OKjS7AND7cZo0qfBK/0KYVzunIj
d9BhLzWUiqoenm6f7tEuwriNb4rD8Sm0h7X2Y3iXFJ5Mc8HDvr9Wxq9hyar4WaPX
jIMplAJSIwdqW+X8ozzej39Tw+0XWCf78g76MI6K4+61tuOwr7cEL01a7liEQpop
zzFDbEXrVbNLlYw5+UI1/iv3S0lLsUqo1c9HZgDV7bBVslXvzGfYFPjdA/q5rJ5j
MZ8offXZxPXTihcZIlUBQF1hw0ip2Tm89/QWUdBfwkFJftQvzruIiFS6zZeZA4hV
FpBoPmQmqVpLlEIuMgA6v419AP019pp1GI4UC+iFITHtqPxdAupJ4paWXCbXug9D
ae/HKOev0Otu/nIYklw2ddX1uFGGIh0zo7rmG6VIImhj7o5gIr4SM138E8L2dCTw
t9cXIYNIdJGI4+BFCOjo0gy8NNUMUo658b9gsfb6KyZDRWCS5V8VMLO1GX7x42xy
AXtxgbTNuIjWRVh1E7tNavjTMTjMZUZwWApAUtLPvlwrmeZuC92HssNBl5+Tocul
F2a1I2rlsS8ovxjLMqDlot6996+fvDphkicR4bQ3ig1oDSl3/1FsDXEZInvfIb3B
jmZTxHToNl+tCMIgMfZJeXwH3q5XEtlK9Rd4UgZKXhM7YW5O2f8uNBRsNBBm554C
LOQnkAJr/89frDQFXXvJwt4X72Ok3GrVYRMPGREcARDvfMjBOBTjImWlsDu94OUW
bA/bu3NW5w7cPI/NkkJc+L8NGDfXl9a9xPEjCxA1ClaiZejNBsUordJQicNBifOn
/DearAzOIX/PvzpS0Ii1iD/Z4HM1XbeiNrpH3Z6dacdBSTWxvNxzzaBHanm28+XM
9qUbFMheZ0ZR6aVR2J4AootEyaHcc+X+GxbxLEX6HtEjhZ2+9bSBG220P4FHvPoo
+KFJ14/1eqcXNTMJjaIt+yUKCMi0XAKPr6sYzTzaOqnQL+dxOufUqYdGe4KQVO0e
BPQFHtnIYFX8PVjdOXkOZeOPbz5cU8qLOLa+zvOTFmoGR4anekJt81U+tfQuqPZJ
7EIBY3Iglgs8N5jTfZEU4nQLCw2S/p09lRqikptUSTcRcVvDEfPl0FMp4y2zfQA8
sDjUHN43oJ2tP//yBVi4oHSP//3HrP3vH6uYhhYw9tQhfOdfCVL0IJ7eyvpIi1uf
2PcvoXIalYG+IruPaXyl0mMc/Fvczkhg5XMMz0NzVZAX3wIm6hQ4YRLJzPtQ7viB
MhR9www2JLC715kycANdlUHTcIZ9fept58Eyyfipkx3/MW3q6SyB0dAujk3LeTmW
gSH3RT5+T//1g1vYgKvdtANbk8DMLX4h+Iw7mQpGiUvCz3b9MAzsRa165B4afm42
YxV2qFjiqSUSrkJQi+Ewb6vFN7WTqaCLZO64W0eL5bXQor9V+5RM1pjrJX7yRXKV
LNjWYKdLJtr65svj7mgJHRcDSyYY+Bjkzt0DhDarYdxNbp4pWZXZirPw0oi20d72
Sobf6P85q81/pYhdN2cbEkDFjLj6n4YY3nM0LzQgmnB/bOYN1pl24OmyGmaRLsYK
BkfnMe0BVhCVRcwFKN/S73I/+xJjxW1x5yEM7+Y5umIGvM6ZeiJCarTa+7HCIRrs
Pd7HG4EIxKwwihq8tXprZW9RO4hikPePRQroYFfcVX2tTVyQMFHNgltItDe9r7RV
E9jXXJ+6PSTi1HXmv088orQwGgXgDB6nRXjGcZb0BWOfkZTFpxvtcCDhejuFcMfs
JGXWSURCBvg0w0ho1HyJTjhvCuqUby2OcmCO/EjBiPqXts45d5M5SkvK1+ZLC/DE
4bRqNqxnbzNDwzZaWxo7BPCs1NNEeUtuSEYO6l6rI2OO6Wbvjy6iM2I2tv0qcq5o
s3CyVNWVp9EOcsZIzAXmZw5CJAVuaoNvBKvJ639fIBfsXZRt1Wyzh02aIqh/drk7
1NXVeSDbbljMbBLUoyIsQj66CwqHUjvnfsaY8izg/KLgaykhvtfaQPpV2+bKgy0R
MFtzxdjWMe8sJqhB/JzrKdVY/Xjo9mzn6R2QkscCPBobuoKrloWiCKv/m2zI3Loe
dTkjf2Ks9LOmui/wkiRYpepFA9B070OywB2LjxljdnZ1FFNx91y/QaO7ySkP9nHS
Z2R0ZNMm88FJrqpi0eq5bEuqk9B0FbstFWpOeQL7uViMMme0Bi3bObQweeFlQBJB
v6id2+gxS83GWCQWZUk+tUF/GybOkeEJtEQbJog24J1Zvz2RAfYXCMWbyLy6GjuU
JcLSTVhUe6o5OqhYogrjMDi/2fQgFVqVA4eVy+qjfiMMgGG/yQe7u7WaOs2JQl7p
a0ByJVm/x9oD+6W3RxTUG1HJToDNbIy0zi3o6/c1OcABD0VehwicpESOkt72r273
rahKcPgnOqFyFNt4+n4R3gBpoc3++eIBC6h0vaKm+HNjfLjAVF0MUt+J+aXk/f9z
6rBHGYha6G1B7hyvucK7SiiEmPIPD0fTUC913YFQ+QmpX3UGEodHn0+m2+E3JWiT
nRub6r78LLZBCuZDFflXVUhxmAC3rZ6hgiHCuGSf0p9hU3DOQZc0YhASB/4ZMBGe
AKdKdQ6Ls1N+OFn2tooedCclIwwNcQNqBmxPyZ6yGx8tW0bThvPfwzULsgLVdUJZ
etC0N3A+fP9MwmTe4f+PmxN2Qh402I5S4a6zt9ddBfES+GdOFdu2PDtM46Y7hpXQ
CU75UjRAajfpr7GsOBHHjdfI4ieIcU5PnwDATCNlnrGSsEQSQdGISkpCP5BSDxVb
2n6FjIN5wLlcf4TlAdy/0Arjpcw7Z0mfSlomWlmzFIaj3vUb1QgQWgYIw4ab+wya
/YlRwNOW3sA2zTxYg6ibPw/c2zrskp7ddeVfK43l9Qg5+fQtWwDgnFDK9HP3e8nT
LgEZz0vCozpEZuvQnvKAu28odoH+W2BL3cr1CbKfBIMT52bWRdMB7zygHr3KGi5u
Ay7vsMSbpOIKyNLwVQ9cD7IFHuLUTdyh9/xihnBi9o3iJ41oG1+FPO5pnVmBgMGB
EZl33+oRmufkQu6qTnL8ibs1Nmik+gDNolwvMXYkMKOSyHQjD26PM7PdDu8GtuHD
15JN04e69qjC/pwiSF6B51/SSYQhhal9ZB2w1XIwZgkwqvgE2VopUNvLHYjXa8hM
ZtlbWKQpHhJs8WZfR6nofTaez1+ROH6HjgXXYUy8mtTXyNd186w1olzhK2wftaRn
rmt4APZbig4ZXIMHqQPDl+L8LQ/j8x0dP/g+eJhILHRXacicBAP7OuqkpnQm5v8z
8OYsIAHyBuO2vjHYDhBpQRKrHMNbUWHfvLTTz6MJvmpK1312ZqLwc29ECRSfJFTG
HbELSH2GrA9u7ueE7W5pz36pktnAT2r2zELcg2jCGs6teL8JivjJ7Yp4jgjAZwqZ
hqYlbh362Xe+X8t2svxi95GKFfnP/lZc+LA+HlRXF0lzLGgXK5GVVVVbry+Up/zr
w5/HL6w5Dl/Mnh2c9+PIHXOD2pclFP3F+2G74EmhUx7KfVmpjCKEFRXXsDQoA15V
gvbhQwXPEmvsKEbstInZDHtSPHOfPTJqPRsnIkjOq+QHLstN7lRCEwQGNzkIpumf
b/EVPvBEjZ1UXWt8lb15VhGC9IA424q2I1QIPpWDBvDZSbGZ6m/REkTMRj3SaNTv
g6dMj/KFHx4ncBpkv+kDmOzJjZsm2kmOf02VTg2JArYLkopW9vVvbZwtXjqPr/1g
Fs4rqAIE7wFn5d7R9EQFwISrtr27Z3zgk9FKHw07PDUMT/U+HZgyrSjUNq3bFX4R
urvbHzxXY/vFFn1G5kuX2daNY5kUeKfOFwzLKnkwFTxOfgQui6ZbE6Q5C8paht6v
6cJ7nO5y9aO1RlShEr7nD5Rz9xUG05vO1W++JrjNCeQoc9B4FLIyDXKJTV5XE4ft
KCTk5YF1yY0tBEiVXzG9CjhI+uUl41tNY8esSwSEOvRNMvWbhSczGECwftTd9Sof
xrmEE51fXd1Sbwzz3yn0E1S4tM/yHIDdqHRhJdCejjqvo2v5JCINpeDAiHOcYEC9
MtC6If9uKCGNDIAn4nbuTouKHOouJsi7Ld45AGDOAhxkZcg/16JHSrwANHBr9/pF
v3DHq1Fs4/3DA2WdN4uROoBVsX3aiz9mFH2kQaOc9oQ2r7vq01usPNLNYrfI1fJc
Y5VF4KSNE9B06cO2KvaSPsUhc33qzgZObzPwO/gOo4xGMeOEs9t3GCFvMtubxqzL
MeI74+N1s5sRTtPQJY7Dca0i68phtDPKX8JkFZohXAj4TSFkrrfrqb36y+EDYqHQ
eZgKXH8XZtJbp1qKhKxa260UKANI1yHLZAkg2AR42ZqJWsfu2tj8ZVQudEgo9HTX
1ZgZZ6xoQ813M3ebP2gW6DJ+/u2v+Mn/yLLEUqVktkMOFc7l/5SUCIbsKSQoM6Oj
PBB8P2AiUCM2+abo52rvopjbVUcrgvnN5xp9NdM5zaFgxtlxyJkSmonN1NdrRUbd
XfZ72dh3qUj/f3RPIRpM9lWwZSK9wMjEVvgCe9KU4VVBrO8SR+Y+47EZl3exKvMD
qTUYuIgdpZK+yLVLHEHE9iPInPkwROqeUU+3DDfANdsxXeoxwg288aVA+uwwdiru
haxA0ZCI+Pag+4G0TIr+l2+Sn6aVAKDT0oqPaouVJlvV18S6pa12XjunV4OVgDVM
x9k3rdX6fp6e+VHD5ikLxo3B/Cb1sT/IVw3JNbIvamNO+gXmpiRH3vlo+tMmVMvw
AjCUpfU8/KsYh0s4X10UsmyRJ5tB0p/xnY844mmR5t3CeLpX03xVbteX27WVimd5
GK5mLDdPWBKBoVWavdwDOht1Lwul3RveWBqmb2TiAfn/jsfgZRsC9OppJQpGdIT2
g6gd8qjOkOckqAhjVoxGDVWWtOcxkRz6qyscZi/Kw3vX4Ejs7sI1mjNR1tmCz5Ix
VDDsYE2lZAwYBM3CiIURmFGDbwFzTrLhrxDJ/Ot8u2HfPoJq1C5s7lEKGW+aE6ee
hstQXiunWZ09s+gYW79NaZ36eiRGGTlf1D+Gssxi2zZ3C8pS6kDFsr2gaOe06tVt
K+t4szQMLrmJYaiwk4ZtwGWeXo59LfE0xYOsBGVCH3Qu2RFC679X7pBNGeRErsuS
Cmk7lisz0qBzvOrg+gCfjycCuMNJeQg6R9moGhg/1OT1gKSc71c1H3laEJ8RMVou
hG1xOVRbVPdORRnSaAH/dWbk4+eqUkuos5cY4vMkrpQqPh2zhIaEMuZjPqfOYxLa
skKgXW4MDQNpuuY+UcaOQGpSIAOV6Iuuj7HPUmgSNg0TvJtjoepmb4x+IKWT13tt
+oa0K3PM/1aO799MFE/NTlYsyw8Udi8oqrFWKUbSEQ9JF7dqVOwNdzqVJOdS5zxT
ufO3uWPeSdep/lOgQsfT/TuOcuAXPRWje2yVweCLxGGB6iOuRVQLaHYj2pPSKOW5
cGCfSEVuq5ckXaOH28kNXV0Qm67oNre6Spu5ADueOW8sSmICf2s4QRdETCTm8wE0
nJECcyRNEtr3DFSJwmT+wsaKrysr+eibB9fvlxybz5MeEWSUrk5IVtQIOXOGlLtl
H/Hf/D7Z8AJoXTR30TiB6gQ6yNKI6R2y7q10xKE3vKnvClWWI6Czl5EbZPrVf9kQ
pSvL93Txq0kVkne1IFMuW6v2a9I5uB08vNdeAEOEfeifXekhhd4rZZJsEKLxooMX
1wL18vKpJ0cXgKlYgilu76ZI3hP6LEClJfVeNCtm8wVILnpcLSWOa482dlMoZwjH
z+z+Ue7eVjqEYv9SGuA2J4AkEgj8ysMyyxzfpraAny9Ju5D9IDlb2+rc5R9EJ9Nf
E1yvXG9ni5qGARn7aVpkeZ5JzD5MtKIjLCOp409RXuOAA1KpwQilTEtRTP05lY28
7qDzguudNfnIRP6MeyCtbw6hLKbqKENnzuUEcZx5PKTgrEeUX2L3EMpUD2A+lV7d
I6w2P76SbOo72tfhOgCu7h84b/BRovPFhoQ19GbZUVbSDEn5h1w+hOqEHUnglNOO
pr+fvMo4kwmD6ONSFPSN4vqqL0+Ih+a3KbLK+UVa/buXIMnOO9eyVCB6zpiUu9Wo
oeDs3VwqW42fT4Q/1E2Ggr3afrn6gc2peCIuPlEkPx1IpgwM9bc/+8H3Dcp99RbN
ByAmv37piJhNtbSNV/xoURp0qzfIQMKSlzMp8OHHnvVbcYUXKc3wcCFrY/rjYcCH
5GxlWtqOUL+Q5hb6iALKdBAXXwURwMgIyk2Cgmy9KRfSBKwhb2yYXwmUyz5tsLya
T7lX7wFZCzcZc9AGH5pHS3djvb/TSJnkHffs6ydh5lEE8BZEZUZy5mGTLkwbwD/E
eEN4+d/U7fHF3L7Bni4eyo/Ed+19iHs8oMv0Ihl/o3t0TkK+IhaPUTQWjMKPWd6f
qddNjqWmzasoJK1bwOfwqWM86M5OXwISfo7CRIPmZFJPU7xTlMJ7vzcdkM9oLlTU
uGgxoFSP9RmAprvYBup8fkBzqWwk1heGqoaXzhHCpUh+UBs4HnpwmCIMffA97Uom
1kOjE22bv3yfHx7X6Mgb+i3S/v8X4FSLKwT2msPLB3TQZsgj1hbwF8cg/4c9+GDf
YLBWkRME+7HH/2OIQofT/DY4LM04ryM46qGm157S+Pw/czx8vQslZrccod1Zd0t4
FQHB7QvpBik3YYKmpFmo799N2gZY7SJAIlz0rRrX/D9MbXz+7QREcyJcDiApfhtz
WK2sVxVnWnLG5hQjjzGYUT0YIXKDLPxUeLCkZc/LPpJ2FfUy0NaQ6VJ07Y/c5mbw
OP/WjK92TABDp/kgLchDW9gtUe8mQ0TOtREaEYJWGBRmTjBm8vwrdFaq4mgRr7ap
UjUby8G80hnqqo/6UWvCsQ5q63dY8Pn6qd1RZY+ul/KKQlp0f9M5gU/xD42sgd8b
zjK65z5CzvxKDwvygtQCZA6T7B4NPfC6ZBt1jZapDC55SMtGRYHWFXfb5GO9Dwh3
vVOaOqFO8/I8c8NPS57FRFMU73tmMGjysg3WQLjHJxH5+dvE3HNlZwtezsxVSoPB
rtOOwoyJOREaEb+QYqKjjyUhk1GALKAjh4qG1dTliFm8snEiuHU8s6r4zxVyE8lC
5t/iWwlnkfp+XLQ6rh7emMgsamgOkJe3TTqoJVAeKQXnOUjQ5iuplMLJ/5c1AU8k
8u49cXcxpjbSByGNQRGD8DhkH1ZAxtAuZjj4EnLqTR3FN5CpeKFJ8DxMndYig5fk
V5mTyz3trgdEgVLD3DCH+GxyFwj3R7byJQO7cOg1eO+vP8f5LptbVZmXAhohbVje
toxprhog3FNejiw8Blm7lsX7MiWOg5sX6RlQgYfeE69CBJd9amJThzJC5WguVZ88
fu2XPMUZfGqn5kMBeMlADr8caYSnU8cRAws804zVGOQczBd3DmTq39IXD6yt1d3T
AjfkS8d/0941t50ArplbHyg5TpsQeuwe/O9DCptl4e3W9MKd9gUfdM5heD1MarOg
F1fgSO1pPyx0GwVteOJD6Yb0e0LW137e8Qz6/8mo028bPK00cNFeKpJ1JU3Jb1Lv
oRLsP1vw5Ikm7MQ2yjKJBFD5rpv0ZjvFpPhy+4XD0lHdHVgWmoXnPYS+TXl73uzW
bjFhdheJ0vxaRnAvIBqctGuWwZokvp8TFUwKPv6GAjHY1DCOmAi33gePwqayvxHr
7yV9OKP3cxY6enfBdXKleIPhewi3rWuxUQc1CCQ5cva7Y1mlLYAkHR+vGxLHSCRI
smjtzUOVG45xKuVWyTK5kUsk9WQLcdoTANBE+4EOOgGNJ1/ipMbRmS82pX5TJ4J6
OIhn/v4JOPK8CF1iaiMoBal4+xSfe4fq9X4/r8QfPhLHbPXq9dONXqHFcry6I3++
PgS17w10/O5HNJzVE0p+wtpSsmTh7MuDy11JHUZzNBAwbBeKK7W+LsckCA+MGeYx
oZUuNIVl9dVL7aw3dyujXbTjLm1hDsLszmK1QJ5bRrYPKKDQ3wtZKtNKC8Uu3pWm
BK0s3Xbjjfw5P2pIfGqOPljg9nf/sQuHIX5Xr70lqH5b5eZLtYnkN3c1PisnQofF
PYsu12C8m/06haUs3drDBYaWx3iWWx4PbCYm42jzucoS4FZ5qHV2Zew4g6JjClOB
r2axLg42IbBOohEG1SHKGM44wva7QV4J/yXg3mQ/Egv0Mf/biTvaDOCNPfbd/gTi
SmMt3+OllKqdr6DRyyROBZyQnASgQ+EvopgytcV5EP0vOE2KIlrXfuiKXe9Cm1Su
dRL4v/mN3Yaflz4lnSG4FAYUfmRu9igx9u1vsHmZr+WM8ueXUxkFfZapQgTYWLpB
5R2oZEoVAt1xFIn/+V9/l+1P3hTaPAoT+W/hkqY4KNS26oJ7x0NjuBGw8eGpCCkN
7oEmEbKIIbDYbUTEpvQDHs/XI3QlK7FCONpsuTqhJeBFg8jgTB228G5B5WB2QWcl
3VnKatvbBdiItorCvodHHjMe9M3iC54hFfO6rBiyNGcDpIwPVElra1v73m0HjwWa
g0meuHFlq+2w0CMLyoRm0dWRFI+zD7z9cjB12HtHvKdpavWlmNGYWNq7ZWIa3vgO
tddqywc1Klg2R91hWseXxBPTJfmpwwpz9o6cIiTi3pzxrNMJ7pkwio50+FHdPUpM
t1p11Yrtj6zQUI1RedqXwBngKTCKyl4Z8xeqoN5KIKiN1dMMlyUeYOihCdvUrQY2
/FEHcWdOIgCx98QVEwMOfuCZQ/4wx/hApoQd65f0ANcL4dmejRZ2PDpzhUTGVk7Q
29YB7EhtmXWrf6Doeo9GcLIQb8pgyJu+byy8xtVsA4u/fuZq7Cztgj6TljZxsLRe
2DQ3BHYOw+J6smoE3QhVXFx/5DqTFlgEYbHlTyLv20ACkxOG5lqAzA5rs3zIf5oW
PZt5MZAJ7e5pD5sy8cZ3U30EwUnbYW3wfxaiW3+FHMZdvj0c4ir98A/uUFoCae0C
HeFSATdRlfAORzNWz+XCKQQK/E9JMCPDNDxk8QJ83AcRDglyE6APf4BaXKTNdeNu
w8844vngqwfpyzmjDRK09WrEr2aTvpUSv4TTzekBn0zmGY8y3VWjF/f32CZJnKKT
Y/EW9o8lhUp8IhCSJBxsL9WbE+RYomhbTvdx9lUSBh1ocMCML3maxZr62IOXpgYF
1kf1x/1D381kv+Ckkr/n9cC3kyylf91Bz8PrJaQfHCiWl3FeH0SiSIUl/lYWUX8b
vnVizWpIt0M/yPBju3dzS5iBSHVhr5rVft12Zi6P3Qt1F7d43y5Ol3yTeb4FqziL
VOX48RMB2HMCF+oUD2Uu1k3YHHC43Toj58A+415AonyllOlPXkcINiXoW8R+VVhf
YsXNU+AW36/027nfEHkuKrxb+QPCzs0mW1Icx0/mNIL22X513STEziPnnBc/b7mq
pEFa0pi3oOiRhM0lawtneF9QX3NyfX3t5w82OIA7CXl68cYiLcv5oIpELV+KnTxV
5nZLk7AcbiOXAw959xNR30DFE7N3WkKABzPVOPRqnb1HBzCmTkglEJsB9TIg1FR+
KF9T6hU/cLmvkLU1sivfVRKRgwb23tLIWEtP5FsiglmbYx6OaCUP3r0pMOF43p5w
W3DCjj8Ivxda/OLbqctbgO49ohgfhdHtxe7kZ1jr6/cFZYXASqf81zHsy/FWhtWr
BnEtp8zf/7k0kIhz9F5DAhWAnpcwU6pstKY+hGckn5nhOaliqemjnMAkvNZVWavP
XprJE/Vs+OV4cjb57LZU+/wq3qtdYLfQcb4A3ITyrXMJN+kL7Uu5t85q7LGuY4mB
s+rOAQH5QTb4enar4B0AsGS3d9W4cMLchZNrQEi0ZFpItK69I+OH41563YFS8inr
etfUdxXoLklwX4b2qcHxUx7YfeDoJ5uYfx8oVeMIGJdsSRr4hoCGndf2ozrH58Pp
FfF2Ga5mP8GmvwXvGJ2p25+f0CkC3jP2U4wZnCa4fiQ6f0P3Z8+VPzXNTf0ubn7+
IHs3mpQ7cKt+5R/0r2nDrBu5JfFlahzd4cTo7yQ21hwLuuKsf3oq5LDzM+bjeHm2
1V27HtrtnDZOVCafXqLQE2MNMYy5mZiGuWeVfLwX9mKMTEz0WH6RvuaEpg6kO4Q/
4Rw3a3hin2L+lV2JxpFCiU0+9ZCDJ66nO4OcoF0dWwIpVGjDmjwKYD2tzLlUgUXD
i+sKoTMdKaP0h7Q682lcLvt1KHv/ysdPbfm1OeqD2cXdmKyjI1z0jXOuRus44dDt
ykcTW5e7QlhujZPGEcBeqx3DbcRugFybBKyY7z/LjN/Jg7N/LDCB1tCkfCQTzbtx
u3tw48tAOb/4/px2bup4kLASOlgJw2qFTTY5lcduaNtqXIwsMjvyfHkgPSVysieU
hMnig97qAZWKrg7BWXnJ40l1kS6gQ3PFWS+wsXLdMpW1mBYrOzcngHkjDMIfKxGY
vxvoVT3xhJspTjsIFmNYZ7M98uUJi2DnCzMb3+hskDgorfmLiWRNAOgk06oZQfkq
ZCbJwQ4Wg+VfIYblwDLkchdgwfVq9QRtVvpdTlxTK132VrWCRjq5zWXDTUHHKSBs
CGE2Za+vbauK2ZWd8C+BYXeb6i7aQ2qYNNbah/DdfhdnDgqF7ACJXOOWLhQ6NU5J
nel7kRW1JZZ6E6BtNuyAdfkDpI5GDi3JXdhSdZNc3cy+Aa/pTafwmIgcfiC8Goaq
PExtpGtKNMvdWCxuKOQ2Agq9L9OnbB+AlKWAbXzwj6fqYjlvpzqS7S2O4gPRTDWk
D+z7GrJR3qyKFEWJdmUKGDc8ahFgNhr46tnELbelvyA7HyPu2V7kFWtM42lcLnzr
aFcqOpuSnjw4++m2t4OqxHLqicXw7ckc5cTbR5K8ovDDtp1LrKQlBWi2GJG1F5SA
kX5pDbaH2KHYW/6YUkfrxOFbY7eBEDJtEHlK5d5ZggdS1uTUqU9IeP9PVPsaVt2o
M8DQvB1ktrSMGcbsL3pIbU6/MgJ0itKzv6tOLnXxrELswy+6uzjpZQH7UWJAjLfD
oigRcJDSiyqvZiiwpNN20dI9ivlKqD9Nx7nXg5icy95lcd1QdGlkdnSbKQc5f2y+
76ax+l7q7klf0s8xFdSXuxOdFnuure73MnwYHk8qdCIu1hEWb3csFGQuIejfZ14/
iaN/WTxbuotxcJQK3ZM1gvk4QzS1R0aj2GyqmaVzdpWUrXIhgRsnbklF54rggK4C
zVIC8qnQkhPOZeElS76JCu5ZWqBVXTnruaaKvFJSrZCmZJLEVEg7Um8RHjz0Dcn9
feWGbhPzwhA4gID1vrESuqfvb2qIiiLHStK6PlSTe2gxu5eoe6PT4H/xjkW+LdrU
sIdcnSP2v83H0OiByD/d77D5eVLf1sNpY9MY2C1+ZS7dXpO02KP09a0q6Wvd0P/p
3dLRUpEXY/oHC8tXPrM6PD1rXUdVM3P2dyX3VETlL+UfbamRxygBUdjRNMNDVDhN
pEqA/JS+mXvtk26LbGwLrSESvhVI4liXWQlOo3cWHyZWyC0duBUEcteQuvEHZeTN
DidozgOhBhlJtmtslOZfWsU8FU+emQ2OwXS7Nf5gdDbV5FZYL2JQeWPXCXcCiZEt
x59Qd4K88mqyz+GGL/FEpkAS+opbryv6DQRuY9Gj7yntx45WfM9rpx6WgXWLSmYp
Dr7uPWojKSrLElwChmqUomKT/KBEg9qtHGmBAVaTAsgGAiFF97IKFdBgY5Zxatvr
1vXQ3k+V+5tSVToUUhmLpuuR/Gz13P4pD4rU2U4yCiSTgb8hZbVjhj2Q51E0oBBs
txqciC1B2eH8lIf4Q0krwwIn+bkU9sxOLor83mV7zwEbJN9AigxEPjIRpMCqFh83
oVl/ZdPUMXoYf1um1SLqsLNnNfx1/s9SxJZUW1usSptQO9QZtW9h30BGOsrTE/su
QbxdO6YtbxprMuP2l0K2uX+SzfW+27GW241VKvo3pQcQA/huV41hJzK779bfTHVs
g2D5w/WhW7Gr3JcfX68ePyQ5+Ad4svsdeJtSZWnqefUfcnX8TJt+XufD9a2wqC1B
e84VsQXp6C4j1sU4aHa7nFI5/y42AbQLEYLv4FdH0LMqiLvC3kVsr3uFHjKp0pMy
aWiOf2NVG7gBSsQXcZQ0u7u9aR6UlO1EThsOB7gKNh7j9V1PHFaqjRm0hZG0ETVy
s1Yvq8zTh8PuWDloTpaz0RjFZI0dh3jWiP0dEVieVMNYZTBaJpsYRjJyQUYIhCjR
G1YXKBE/525+YBAubNBc2EbRiB41Eb8GKK9JNqzZ3fNOXsC8Juh1a4myCp6rH3RS
LWfuL4QX18gwwlCidMnYaKKR3kkRaK60oDNOtL5A7lH8PF3E16yTqPg6OZiUcWI2
O6zL4R9Nd5c5emIf0AA0psTjHmZRYfF8ONSDquklkr1nXJtZ9ozOVPI1ng34k1dC
Jn6GdkUJ8FtPP+yMxIJxW8fvlYyO2DrWmWdiqtcrBmEPbZn0+pprG8324Vnrr84t
eNSGy+DWNxcKPS0db4E8qb6UaYRPJdkFSnTQlWK2J6zxFlJlfQVG3zho49gYER4g
8J0uyESe3KKKy5l5A+JoU3ZPwffyWF7xlOFbfZ0Il6VcQBD48aU2qJveVSY5kC8l
Z3GucxM0aMSW7Y9OqPxnVnFGnb70YMVQ3b7iTBKIFg5PaZt3ldESAofNdjEuqNSo
lhfnPSVMwUHhIxffiZbzePRMB/UrQnxPp7fNkqfzdxl2Asvh5RmcRMVUBziUgRvQ
oBXdvkHnIjjTxIQ18daajqp7Y4+SUHnfrnHY0LXXUDyuiYyxPMVsfK9WxyuqJpMQ
JPuTVxRkf3hAh7QTzpLd7bjM3FcUQQpP4bf8UWxaNyvkq1R26FAExp5y9mcT37fW
iWtcAu0+66Bbdr+dwbIqiQPipaLXIqLvOEkJklo+N2RygXF4nrMzvd54iGgY3ZOw
bIb88RmcwYW08DGz8kPCI1R/Zy07I7+7Gv+/6FK9DGDzxwAjFp7kfwTkfzcUrRBL
i1gV3x2NW9Q0WYiu1vppbRga5DfR6Mp0nEvUfBxewKe94WpVxl2HDBkzrsiugS0/
QblFcKUCbmtFPm+C/6qs/3Gv9zKlRXWvxF4MCFDoaj6LMB24GKdC/Dsx2alUSgjE
gxpoh0IL6We4hCiQfxIxQgpSKVty/GpV9pUgbTiHz/84Uc9mLy107F36OwNxGYQQ
NI8GG8n9FTK1UZ/gZn0i/3xXvbMGN1alyD+P6101Q961WKVhDf1GTFJkI2WBvVl6
eFHVRbgKm9u9e3NTKGQiKJKEu46uVbA+3lJyEo5EJvGx+LmQza2QkvqHVmQPts4k
w7dYiAsWvyAJkZ5jeRkCesZbPuqs/prpZWLmJvAoHBNDraEZK9HG/YqxjtWqRkhM
hpAbq280vNmhV/oswY5Umv3nAZpk7QSNWmVO+/vUKocYRZV2cJsj6GcJN+KfIjx2
KdmwQ39m6yVZQzg5P4cQZjbLRSg0Bnwyn/HYDERDWFqdykNKOQXcM3hSXCeV44cf
cIfQbyaISyXikvwfBsGL8f8K19I0nh878A7tHT2hvXoLNOXWw60ceY10lmJPk2Hp
6m2GdZBsJY/JWE2k7XDpBSc1MhgR24IOqrBlQZPUu7s5RBVOTkc2o+8k/xbHl4iM
TCrLijV9soClfYCYsmxDYBPDSlolMzXP+8l9Mxdp5xwwQvP6612iin/NZvrJM6PN
8BWRb5uKOi2dxOzSXxVT8OAjBafNRZBv0OdH5j4CSqlGP6Cx0QJexRwFuKH8oekk
GPhStvLZlCPwSoKv2CO2rC9Igq1mCSBNAIHI3xTZ22a5jH52IQ0KKj4B/+STk/Pt
u3pEzI3oB4SD4+7yxCsr6x4o1GEetICRwKeHMkS75p8MoDGR4/fMK75l2MIvWmq+
`protect end_protected