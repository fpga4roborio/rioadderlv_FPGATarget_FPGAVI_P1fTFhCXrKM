`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
ddtXksX2+yylW5zu6QL2Lhnb2d1sD00763mmSITNX595NcHTEkwn0zB1Dry37fOW
FufOhVzEJp80NC5qZ/+F0Vk7Ik02dIR0elf3clrjeJRK85K4e3Hoo4xn7YbFUIms
l/8VZSb14+JVGURjfswrIyCUotIzlzVYZ6gzoZwDXIi5gQIBf/gI+KxNXPaKV+PQ
Ufys/12rjO6aI/pPlqSm0hCvftmBcnezN2hk1UeXgOIuKZnogjOsf0iJVX2aOOWE
6pD/psybjbnsNB6kH5uFTA5frkzIzkzl5d9+YDm9OyC+k84E83I/7/j+rk4L2dah
QJOvksSIzN867/4Qt8qYTQ==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="MvBXkzurAa5VTw+1JJ70nePUfoQXBvZOku/SMmg4TwQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
oRtzZL4VJ4iwysPsC8SXYCzXS8Fw2gtZTOskLcDV+1B9Nzn1zTyNtlo6lNICRmmK
ZRVu2BmCc2G+fmzynYlNTnSa7C0Cuel6FYpxCBlOuk3OF2tzAmLAuDyOH3Z1Yjzk
a0aHuoCdIRKv7BrZCdALt03JeUmXKPdOmIlkVGFl8yw=
`protect rights_digest_method = "sha256"
`protect end_toolblock="Jn9CQpRhJt4rnzZPRk+dOpzAubz7omckX1MrFd4p81o="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 12960 )
`protect data_block
gD6l00tciPUa6pDNTk/+t0OO0nC/UTtBwLB41d4inuAUA3i/ALrNyoJVcBnAmEQW
ptbcNp5fxEUJjnOxnedyZEuEBxWRieZFQnkRdF269oMrXuZ8tuScbvC9iK4dGf7c
0wLe/JVzMm6lNfE2cY5vcLv2LeqYMpF80YVXi/I6Ud4Jb+I0EAwumlkpoi+UFwYE
1umTq8DjOQwWh7AKPKvBptUxLqCk0vcaCajuRFCBT9fmDsB8tOIilxl7/kyZJFEy
wY1RRFOK5C3vxqNHQVq+KpYKTrz4pHm4iWCUOPCziIk3BIEEDGVxAMhGMwDyNOt4
dF/kAEzpxf6Jc8XDPFN9BKt7cvEH1k9cULFNNLeZUN7cYb1iGKmVhL3co8gMQHGc
Mz/qYYD3IZRv95kB9yrxEsDxuZfUDkgwv1VosWrfkC47UlK9uQaPf5SFFcii1+a7
GN3gb/HX3363zRQTbx8GFBgNk9lWeaa8Th/K2SZgfwYu05s5b6yYuqCAAHs5zNrC
6sn9VfNEf9MI2YFIl8YOWz6iy3Mu4cvVE7wl9GY5SDM3RLFL1KsfMROa8PYZl8Ta
SJ9VCyYjWOPNLbJXeRa25t6uNxFWtr48mME2/SER3ULXcS5w31DqUN0XGGtLKBfJ
j8hm9/bTWTKxP58QEfgQUm90cG3FP8v4MCr2t8RdGgP7B4IseJLdkkudurY1FX/D
jmbw8G5fKdgS3ktVNxnw882VetbjchmkAQTiQwWohU64aBfq7Mg+wJv7cNRP2FTV
HsVbVNAnATv2Al+d8sRX8GpUZojXqjfQueJGqiwzDOjVn135RoQddNID3O8X0vmg
L8tE5GYQhkD8gy4aNMTAzFEz3ZNr7aTyhF6QUeLhnOWXZeUjHKG7w3tGM+r3pwzW
iTE2TPbQ+KsjhvYsAuDnqoo35bDNSdbsdBPrEDoAj6HURm8ssbrFUERyeidimqid
rv2Jd7tZjtbY5/9ruAB6vy/NLNtfknKzrun5ajtV9UATS8PCFgDdyUoFa4US/Vln
vtsfKPXchb9c0AA16wdPg7BIqF2AUfPChR0wv4pVdk7QuQdx/fEMVOhbGQ9040lZ
OC5C4WZqQSJagZQsf/YDpG8t1/InepW6XIKUSViCXtHl/KLPzrpqKaJlApLvqsGl
FOLfdAXryTVegTUE8Nu5DYaZkGYoZ692h3JHp+CSmCYa6TqG9mhZ7RZXxisU5NXS
mwQaGWnripzaRLgKQ5mkbyV5ycD4sMCh/5klOuTAR1bkbzlZaOZ7LwZVO1+Vf3yj
atjxbeMbtdwQ5g+mxWHsRLUCto1KB7YoxfV7c2cWA97tPtbAIK/t6ftiwnRQgO1j
jxRmb93b+TbdCCQd25cZs2JleNFlHzcmX/77c1Kh5+6yL/v+xOqRb5Fwd3EHu0nD
G/mdwECbHbEIyiUE0WZ63whtd70Ki54UkOUwCZ/VHw9VnQn2+CONBNw/ErryKOJM
BWUmk+IuDnWbypefOfLx5MkQUOXl8GOsAbaSOtUHp+QsPojKcuT+ulSMk1qCeTf9
h8YKeEJ0Xx+YeX9dng3NQyBmJ86cljoFlCf0oCPJ6o0AGOEWVUi91gy2dMktOjgo
HOiVbEvL0119sbBdUHDDKfk5WRl6WOr3H/W14LKVrsXzn9MxRhF4xBEH8DRRGQ6r
7e5pxRk+uTDNgu7QJw/V+FUZSKdGhyvtVUd8DYujGf4812WdaaPivPZXZINq36ME
JOSJr+WTQ8SuGG9kmi/ECF+RNuYs5s3xe1b74mzqZhK3C+n2DMGzwSF/87yAiDH9
G8QGK5Kka6+lLLTaE51mYrFUGvAVEjOWSi4k8KeOUNS1FDzFXZG00tpa3r+rxxxY
VPWEmVqiZossZUNvQx09YgJfgS1zDQBfD5KkFs8CCKxSVPLfkJ6cEeNuK0uh7uUy
oI2KdX4TrXDyDXs+akAcv3xN3pcR7iqEHUeEX/nqZxHDifguD/owQOb4s2VR0lja
xN1LeJMVFHH7qAc5Tr9PF/muPAbjvaPqujQKNun245gMn+3W/3HcSjOxdukYpmoQ
WJWPqBYEa4Ceqho9J5F8IuRcK/bTf1EzDqS031twUkkDJ+DVeSV7813ILhDUdH16
vqugv3n0XHnjwuHHON2/to71Jf+4Zda6mCJNudY30S36jHJY0Q19Gk8RCDy0OYyN
W4mVqDDk20cbj6SPgF3vkaQsZMiax8M/NC1XImPpcspmLzxb3hmRIoPP7r0GZ5rn
kd5bKA1sS8CNC8B/5+I6yDebtkx8Dw+hamcJP+X+v5el3wXT4WnOPiPRQoiMnLVd
B+qi4PWgwHZ252+6n2FLlcAOVJvJuk4YkPu5SSm70tDNKD/xuc1Iv1ok+VD9I66u
Wfms8jISKqplwAMViHm7fxsnDGpc5SWlfbufDpFmkRHQhgsgWkRHxaRtUXHDqq0f
ItEh2ovBKYb1pDKyPXqHQo+ErT4htdpTtsBAqS7UImnQ+9/X9uHFa2fBVQtCQZqa
n2ea1Q6675a9mIpnnCEg1+bI57Qj0TyX7x5p3Oahsa5lMZGnNPykjUoIM0VZr2vx
UOhnlIxu1TM8gG+SGnpzpfO0RwF/JQuIgBqZ4R8pq55veA7v6Rm7m+s+eOhKDTtq
pjcAOsDEW4ODWPbwGAYNkxazjffY2LtFPFFiMWavM2/Q7EO7BCYjKv7cSC2N3V2D
JAMxWVyEaLRK84ptn/C1Zejuux3NVa5G22fraJzVppqUR3SDHvSselEMOzqTXdu9
JKPde/9UjbPb5GBSucsdfIPpSuP4W9J9lRcRzlC9qO6vPBH5wF3bXItqculiD3tD
dxWg/B+up1/MWy33YBNM/CwAaDL4jqbl5ANR+K2Zt9u87GtVEJSdZ2rAkL5bSN4r
xdv7dnfgMQmqki2P9RJMQPhIf0RR1u3Kxn8Nx9l2CQbquTNP8D8/cMVoLL6z4QUa
P8ctCjRicHPd0kIt8It04aaeFDIWtZ7lWMBdGDicMP5CVP+AijYfyK6oQNWY7ggS
plxMhmV71/7/zu+jameZqiTEa5jif+oHSm5yoSAUhz3t1/n6erzBLo2azyafZO/2
Az1g3PYlUPXNS5M4yNnlMBakmDRggLxbrqZ+cV9U3njTBa/8Zv1w/rawKj+/Tt+z
HTYTn7VOWobw1ciL8n4I8KXqJNbCfQebmn9XoYs96K7Ct5fKlmpzwr+F5IPfIO+4
Ucsr5r02nv4/1W+NgTCFwj6Z9sCFP9TxeMzP1NvBcXXHJoORmzT6t/a9XT8gPjPi
TeyKsqA/9lVOtuVwvAo3oLyt5AUyz1a/DyTnoFF/vGf0IZ2+zAwIBiYAxPK2OENi
vBh0TzhutgQEcgZjvhY3Sbo5+P+LoAJqfrkgetQzH86W3XXBs1lQOL2awUxFktIo
zb3pBPleLRsKJMdNqsmptIgsgkqpxqNnIBhr4jdYomBppDi4RpKBrWwomsQYQhRw
E2KPHGKubbKPhvIbIylsI+BfX795AU+bq/IdBmTZ541LlZfZ9oBQywR6FodGMnBw
RHyejSd1qF0UyrApLHpze8tHs7RZSKsvBDuk4ERLP9gH2wwRbx//Xyb5rcpgehzc
/BuEqfEdulG6cvJ5Tdaz1VW/WQ+eAnN1ErtTEb6jHeS+nRkFEqpHBHtA0+CnvwNu
tDlXGP9M3Aa4d0gx/WJXIGXRBYxlQIJbolVi5IfA5nI7QEjhBwVAi6Xzj3UXdZOH
Dc5zb00Y7O4QdkgyQt9V/jxWZ2GY3ykNJmzPzeDGNDo1/FXT3S2286HhyvsWkvEy
ZM2VpOLpMR32y/N9ne/2Ptxmj2vFWvxkcA8LzxYOCBfLxCkOGOqI/joETA9AdAUb
wSraPKcU26CQeNOwugdJXG+lOIhb2uZZq2ss8ZyUfLBX6RRk5o8CwEia5xpC2qpX
h/uxPaiF0gxJxJD055w3L28zoej5IpiYbK0UeqxaMyVkek8+Xh5rgYAvaH7jERjF
DyH6kKL2kPjpr5bbSebONp4yOaF/HuYn1T3/lygqoL816KxoEzgj8wQdo09HJ4de
6ypdc3t0lKJT5MRfHpSIp3pNyqY/YfyLyzbBqMiXGiYE3+w6jDGTqUl7rREH3EiN
TDw61u7hxnlfTXJuQ/uXlsMAkFkRqB4dBnBau3vmhk3A4U8pQjbSmBzxhfBPSqJb
33HzL0Ok+Hja9NUnob+hMf2OxmpmWOIOXzsBg0lqpzq8xz9LACYjk7M/XssKBby+
ZC5+u6i3r7yv1LotuXKKbuq4vvj8XUuqxulCIVbgyJn+NENoj4pbN6ceR9J/zUsE
/+VE/g5L6GHi2U8D26kM2kXpgP7ssOnELSkeN32B45Fjc0Y16NgLllyUD5NWSNVX
9CTAf/uYH3PbhQsHVhWg0tbUUeDCzYq5WRYL4w/m5C6DFBKbSBWTykK6ND5yPKTt
ACrMnLJ29AcOOpwxyjx0Ry1zhkUMjHWWbJtR3rS2KyQFUSVZNJAgBFx70lvqR+++
jY/X6Kc+kG4uHA+GqiVXGnBBDT5XEnewg0vuu2lYYkKSpjrFjzky4xyMGQ47JUJO
bXOJoF12VH1u3lyBBOMy9zZ7ocTnyeDxafiNkG19Fkd7mVLMtd9CXiDNnD0ctyi1
q+Nb5RAsnbtVyY9YbgpRF/bdzLK2XXMEM4oC6gDqRV3loQkxOuU79PjLOwVau7m1
7cHqJTTW586FT7RwQDRZQthdv3+HP+whBobsOLTfRI1GTUy+wNBVg91DpcdYK48p
H65wvo4AY/hTMcdR0dUdc7bAKqWEs/LMH9nH7w6BvRqi2653gb1fMvn90zW+Njka
774dPa5c7clAJis0u3AuMUptvDy271DHvGQZaS/vmvjXZuZKuAg91TabDl1P09WD
VGA9+BwL9QluFWh7wHsxWx5f9kIEWRs/SRue3V3FLaLeCva35Y9v92zcVzieexNq
b8Sm+JQn02tmHv2nFFip2iOPHIQM+tGGz6T9+GrrNqh78cRshY0U/soaAhOE21a8
ysow2+wj1BlyVTGoraFmjAHCfsrSD2fbLUdHu3wFjfkk2q+d6ifHeLHnEfxHei+F
+Rt03owqTtg53PgFgFkovGCsmHv0uTm4cOVXUSFTRhmal10drAVsqGvHNKO6GKoc
XLVn6Iob6o7YUH0v6LDNW5Jvdyy85vaLsQ4YGbe8/CVsChiWhZRrWDEAcJEBeLan
YuYzr3GnUpDsYX6KFDehNI0BcdpgjHwtKdzZKiO8aMihua1sryfyRdwX4uPhfV9Q
HXWfkqdmL1CLUN0l6WRMAO9VKcfxZcwOPqEKQ+s+siSv29O9WwSJsPK1bMQmqdRn
nlKvHHQhpg72C5wooD5aYMmSHGVNrCQCrJq1Jh2KQKmqdWpkjNact/rCT0q4eiio
bnGoM4/lWvyavfBrujfjiFDJ04ZUtP8ZwH2cQk1Y5ESXktj5v42pjvH34fmJo+hT
d9XJJZ/j4NoJ2vQsLAlhBXEsHsExEl84vU5yCZV/6EP0A8YhaHtKCIR6+Hlsu/9j
Z33Rj3JfEIuAspbYrRmhsoAMUL0+ZrOoOiOIBl3KWuGuJ4MIAqvDxVZKiYGd+GG9
5kuwU5XHxawuwn+DnsbQ+ayJZEWVBXU/MZC7zGxpDHcVPJgi0vLl8eMr8VxnkTc3
jTm5AUfB7ZwFokZV/2Hi7UuqcDf89TcBGRm539uYXy0OlOt8Gi02WEX2WhHXYrx1
ZL0SN4iqavIaRNHkahJZlO4gjnrI01dJEE5G78qofKdMZqABVUfCsr8Cr5t4HDiW
BOZKjCbmHyr8wGL5Oz85xkqDN6ZQFrRBO2pZC99Wu2S3Ul0M00IzFG6gQzZqSH8s
wsDVkvClGzENHWUP2+CIUsxX2Kc+9rBnyHFr4fDs9u6qU023lelJf6J11hFpgAov
1ppIKyOAAyLnF3dsLkoN8IPFiB9w3fjLc2rW/b3oweVimwBBCQP7PjLgy7lSEisU
cFRde2dKNRhKBEeZqfKmmpw+pEAqA/dPkeFpp2os/+A99UHe4SIAGccXOP3sSUyH
OymLCCfooy2+X8G/Slc5u3i8TwXwsAUMFjZLM92vNlcVGnDsSb9neGwmS1AFMBGM
u3bko/C46nJZVt729XJJjHE9pA10GjUYwDBiCYrcX6wFFBIqVp0JwmlqiyYdjRvG
OK4Y8M/FoK2jfF5D+99KAmKe/JENs2jaAxytmM/Wzl8GA9HIQaAG1zsGbAHb9inl
vZeB6xHpHd5H/E8SKp16tyDRD43msDu0ek6pXDJMIzymZ1dSl4m4JftZTIMMLQtw
qblSMEN290jElcClvI8Pg1eqbtcFRQ2JdH39fmKruMp5Kak1ATorw1YWZpi6UfZS
uh1d+4RucBL3UUCvVhXDoy679wqCKNW2kpXgkpz+NK/3Z2SabXc3pecdx04r61CX
SHh2hsL3+FeWZF7ro1jDCmYy8qGxf0zoiohaXgaCl2MEKtmt+K7zJQDeW36Tqgrp
bKqg3zN6gV7KgI+kpIPvzzmcdGr2w3mS7yVuU9D4EB287UpLE53E0Vv8NWVU4GfA
oQBSEKmTMZFndQ1AJFckqSHwif0Pt5Lbueyb+lWYW1dMKXYP6TJMc3YAV1zM/R7d
Sko5eZefYy6hw9bbfURbhZELy0//DMyln76OV80qHQAeyG7Lod0gBwLiidwa9pv4
EVq9CC7faeFsSE6i+FY+Ipf3a/gQjBjefV1efe5ZtJqE4jYK0Q7fFM4cO4dab8ys
yxmwzGp4jhElxY10Yarqu+HhSN0kCXM6icdcGiUXw2eWYWeQDvIWACxNlfJqsvxA
MG1mCqFiKPzLhhGnt2nBzDyzeTEA9z1Lqu9Qxi0QYuaFqgTXQ2Q8lQAROtGsdKzl
fSRYj1c4WVVqAHkiLAcZBuUqqrO6E1WA/I3lwKneEcfCp6OS1Iyp3u6oCvqdbQaI
Kul7hD2saGDEkD3u8/tZWiqQqZcuLQ1TMAIjV92AIvhehs+PDVwlm4k1Dy++GBVV
jZPy4Ye25yndz0OBgEyJTzPb7CK5Zs/lkxC2EsDwYzbXeUWFodEdVT+iy7ridFQB
UNTMj+DJgMVwpRbF2j6DLHG9BC4amIiZARvbzYIzt1Ky5/2UL/bd/gKc+RYCjEe3
KUODlSp8woW+R+19rGIGjEvUZ7OZUWtvBcK223vzMxnMtxrifhTfvNYRoycV5LSV
qOoTuZNNIk6DELYuPQwmxoQBsLfZeuIaCAV0Aksj3fDU/XInAabvIs0GgQnQEuX7
V0A7/Ce0s3DkX+dMnXYd42UvupOTWxkf90y0Rzf6POi//yghGnKSSigV50hDCVu3
anYOAZQbFLjMZREmiAc2+0KVnYCcya5z/H7TZKmvX2k3IDDFzA/8gp4QP1U4OY8Y
swZqf/fPJ2q7rNtO+L+hXZxQ/plc3plqKrc/fDpRRZc9V2IRCR61OPxBvsYannkr
JOLq2FW33ElbC3RnnnoMKzfQLQlF1wVaREYGJQmPmq8wYRRnRyEo0fefHE9bwa26
i6fbWcI7qfoG6pZI4rK+hiAvENaadI1aPeNzmQ5Jb/BoG6j0jLRbeXT2z1SMveQ3
h+hcsnvOotTtLtaRM1+3uob31vk1pzyC+PZ1xqzQbaN+chAJubOkbAzMmAnSZKvF
Wea5wR5BoIsJpJZbb9jG+DH5K6IfAlRj2QQ4ftoBWikdgmUWVMtW9oYYtcm52vGd
W++8ClwVzzlWphbyslGKaKKvos8rvlYS7lr+pFtqhe34cBh6k76fuEjzt2nKJbEG
WJ4E/oNsV/IsKWvCcb5+f2AJRs6ab0PiMp82LjdLdyNZI/rOwcmBKmmL7+0AEsto
7/FVSHqdqbrkyr3+jQSnAeFGNo+JR2rvX7X9GSUrxeUvIuOUkhFbJM5la63GVICT
Z0kf5jEVj4tJzg3CUgkLXoTdUt96lTFERg5A6jX+eaGfFy+hLeVH28cAik1CsiLh
EOlfi43NaKb2sZaQQJm3+kUyDLW5i54I4jv3miFHNb/oq7w92p4VIc4W1gLiQBrN
xlLeUuWjRVPtRJCjsNryoVJA9JGYZxKcsawkL2c+FVqugEyU5wOqP9VdSd34ACzU
azUkXqPoMTj1pVsfoQ4e8V2V1e4CR2GdjrZYoeaRXjFMpbncjLKh+lnA0ILlY4nt
e23FVexq2+/JlPBwNzKwJLu400D2Gv3xt90cUGJ9XtEIQC3ygWc8ytDG0KI7ZRdU
pLYu0b9pB5j0jUWXUoBh92/Lg3ZbqdQ1x0mHXkq87EQxSpDAnswhBjK31Qomj+k3
0jRTuFW/rnDfBlY0cRAMencSH4q/7Gf0tdpUP4bGhSJn2soc/BNIH6LE68nmEUIw
FK6ICuD4Odh4X2t3YG7LMeXlnJoowRLIqsPfs/SI2jc95cBOMiMft2ZTTp3jOn5G
TGU75Eb1yzqC9qaRLECoaDvnZEIkivzZSWCP/YXNmIqrblwvqO5HgCBVS3HpC80+
nvjXRubym+0XctMibI3QyKT/zNmYW4+lDuGkBvPi7eWkKVuR5Cdb76yVjY8YqJzy
dV+wqAVdWt/bdIuJ49dYg+vHoMpeWbl/Xkf/ypQRt67dud4UeQTNSDSttiS3Zm4j
IkBd7OuDVD0jYkPNn3uHoML12fsKUEFdyLTq5q5eYzHZkioEZdmPz4vEW1YIkrFl
yrWEWcJ058DCeVca6lStgVbctDGoAi/1iM0pD3LQRm3XWmEDwJVoTIsQ3kpYZzBJ
Gs9V4u/uwP+w2H7qm3vCKjQbcKNttrfHDuYBsgT+zsp/Ec934qChH3sEDS3sLPpA
/bLGDRBm/UY47qPL4lGJIohjDQ5p9wOSBq6dbEot4Vsrofu7sqsTqDZwnjM9Oanz
TnMXMIWUC6QL9bge0S5r/a48p6MV/LTGCe522GMNpLXsuGvoUF8SG/7k530AYon7
jx9/X7MrTk5tiM6xDjyD+dyjVc+dbqlAEUc2h64c9pnZIGew8sqrBJuL8k84g++Z
5/CXxjb/HyE9zNuWuEBp4vuol/9uHd9E89Fm84G0lyHvrXw9A2Tqo3M/mOmeYUN6
1j92VSD57NwQmqVbtdd3jfCMZNy6fXMlvRSqIpfB9nvGRz+5K12rZHOBdJCsU2ZW
zt/FZveUSzb3Mi7cybTNXeQpvPZjDyj/IiulecQXaz/GsAnAJmuh60bfGjy1YKwL
kxKIzkWE351FCG0jOnyjqMEe8FVzCf/q39q3CQUBwvG/xCcJ5tBdsZcWxjj1eqy5
cOyA2Wkdy4FNSfdQHfyXPm3P3Dl5y/q7PCY3YmkKjdEyg0aDqlvMu4k92rYp4AtV
TupEInGcStlrFW7FJhGjtbFne385IkV4vIanjcHpbZlpefZs2HdbZnuElzh0VcLH
8QzdOTeMrZR7mMyuDOMA3BHW9qOOvIHBILDws/RYO8MN402lmgHlYH3mSGaqu/JL
TrkLxwJU3yRtwx+NPneCudoTwopVg+BzwVCkG2ZtiN0lfeDhD8v9uAkWaBo2QcG4
PmiwM2R/bBg+fUWvmXzOl342pIVCXoHcCCjvBI/PqJbtCcEQQlgNqU04rfiF3/C9
NRkorpYMvD4j89+qV+vRT/Qox4tQpwq89Ru9TQOceFpN8W1XADpw1uBr9vpLcRZj
LaqihnvRCNl4pvMgnfxARHGQ5WvDEDUbYzeUaS1RFwTIQwcaKIMwejQtH+siULNg
XflRlVTihzy2hoM5z1SUNCIOnxyIxNlHZ6+8IxnM2rm/b5iCVsPy45YmMHO5K8kh
G13HjYNsH1K9O5Y+q32i1OzmgTOcTvIwz0wcCjvNPvxX3gS34QybhXLc8v539RZZ
xFsLINRqQk4D1QPLDm4BL7cEwX0EDM5oj3cbntBbd2RseRS/67urPTGfHkl5Gcw4
doWZo5F481UlhgEMqxs3dWgaXggzypeoxCV0X9QNyb+ziuAo/zHq87v9KjbWj1Qx
P0b4j7owhXuEeoCgFJvb9s5f/+VBN+aUsL4p5NDFT++yN34DX5i5Lu6YJV3dL/Gr
+ypi7k8xmKAkoge64G4hNMahq8BsJKWFHj57rv87KbND3dF11g1GPwCn+0tKGiK/
sYpE1/2Gvsu7aMIQZea1RlvGwpNMsqRYgvg7czU1bA0TAWYJ7cUHz079oAAzaJce
dlnuYLSCF6CJDTl8U0jD5xTxiz5kf7EnbSHjTHTEZqiHmeJYfUXrdRysy8hLRVoH
sFAl+vgRlIkkZgYcEpb5xEEIqHStFqJLbTzw8cxw4z9tqF+qD6wsT9po4D7J+EwJ
uw3kqtwy04PEWn2cwEZXV+UAjL0FYVrR5hznVtX9VbNZmtsW97Y6vb89Ef7WiQ42
41u0xtmBhDKZpJh57SSB6qdBE2atXcnOUtp6Lkpzl94aCeXCuDsecsXFZfdBjnCb
YiYO+vuRw2T+Pes7IuVwG/jZwpNPtCwCqPqCW7/eANeHKXKhmkyf7k+6W9UW8ML2
31mp8aUHDnar2wlS2GrbGp+hv+GvXdWx+WtTG/74cTkwB6ozB/FUF6rLTayfI+v8
lFfMK9ahsC4fiq1R3sCS7H5OGh4A9DxfbchSC3AcKvE7/6Ap8AT0BnP4BLXIlnsr
gstToX6EmodWxwEqdoPHAZ6WPFdRdrCUcNiJjP4TD3SKbBU9IZq3br/IMWNT+O3V
lJm8ginlMqdGNgFweNWxMs0TOX387CuQgU4OQWH7FKNg4Y7VlTH0Au8YCsVykHQY
tO6MM8apo42eUZSg6CSopb/U3SIYa11wrS+/nCitAWkzFXOM4oOyDMWYB+bgfAtD
IpBDUycr5LZfUg//T9wanL2X7TAoZFnFbVTxx9mTwBUjGwb+3Bz79R18w0cTiiMP
dLIjYJM1mECtV+sat2TMuXqL+dI6pufLMeG0O6HXBqOb18PGH2KYEd0P5FD2/28c
JgeLHlFmfdypWyZ72M+zc7UFbwOezbhhBfNeSTABrAXvZzvMjhkM26yhXsqlsSql
b52lUznDlYeAClRRKhNAtJi2B8ZSuwYVHwAwAPauv8yvBgz6vs64SuC8216sfNE1
qYIvOnNm1BJpSFt/Y1nOjW+J5ASR2DDDnbVHVL5M9zeE2swAGwp0GXSbh0UskWaH
TR6Fx6/PQiCySsFJlj+GZUsQY9SCPhNSuzN8WNvnXWD2w9VS6Dkmv90/SQzohPl+
3uDkNDFm2Zw9h5iNA7fHcZDc/z50hun+McUcz3VDYcwfEQj6+LQjsn6PT7KtUb+v
AzpBQSAWAst2GmLiq6/ArujAWCApOhBuGuzZw7NMUDo0I7uWEOT6YSBnCcpr4dYi
Vq+RqwoMtEHLzN+/ltRK1veHhmnj/xabJOEum+AXneJA+u8hC6C8kaXQzwb6Acz1
LeocuX+7XXlBd4M76DxfGhAGj+vNtAmALJIogUD0slHV3LCK2EYWJVkkmcwi5sVs
4lg83ZHTot0eV8Wn5gMjdkpaqpI7YaQ8Cq+E5OlxXLdnmSUR1Fa0+eTUbLRGg2sJ
OVJMtQfd5eRl69Iw4ecS8EDcPgDR3W+PyUt9qfNtk17w9Iko2kppEu/viJf4o/R8
sauqd08D/aDkjh1lpSNYJruahW5S0gKQmV/pjCa2n3Kj5UUJ6dS6I4hpSM8ftQXt
n5CPLB0njdz1nJKIguqqRPqzAJGOuAt/8uIHnJ5c4jJqTLjv0kQivGbA28yiHWUN
a5hRntQQdsY7l7jIcNR16hWFmzGeStJQejSzR9uOUDVQwItcuvBeXUygzA315J85
tF7rH7ajTxwOvivGDgt5QTLkkTocjVDGgoe5hhVxhc1dwm6nDV9rzhKcLHyQIO32
ayrmj5dZCBzZPSBpxcBLS3roVRCvwz3T1BNb43e4kxbM4iDidCo+cYQHo+P/tfIb
5H8KTFgkztsnW1p74f7j2fSSIUjT9ygHq3sDXMrog6wLgbPOQSYtbiw3QTckZn8q
ZRY6FrCWMhQdeNP1vc9pH+SFqyez+q52XMvK2E0ggZKyo68qWoJHxDUDlaYmLt2/
tPBk3ui2IlVXqXEeYMljQ0XpG2WOmrw7KIlL4CYN1I05+kiMWUX4qh/o0NeXLWUS
L1+NIAcmAW+dH/RXkq78Y31rJC6tDKnmQl/O4mBNzqCHh3h/2f3DupHUC8LMPgZi
fmWOi8YuDsOtuSSEXovIOTWPDFHf5Rbfv5vNAcAT547tpS/6ONVG1wUAiY3Q58q+
WgDv/Ciw+LKuTOWdsZlg7RZT/UzGaSXwLPLl+lVzerVVuOlNIrHYfYT8cd9vN8xa
nkkKmGHqrtjgKVETEIjNNmKO4pSldFACvAco7q6sb81VVRo8Kn6HOzLnO7bYJRjA
fIUrn7wMfmkMaZDWWyamCPo2tL2XoP4NSN3S5EBgb1sqPM602prgVGoRLZ7Dxg5D
m3e68B3UJ49VIDaN0pJ/NWWuW1u7WY6YbKmcF1jD3lTzlg8hPZZXH0dGiAxxLfBn
8VCQo65fHJnNF3qM+Ynam2t1BzNSCSVBQFYjeCwlwN07rqGqDocQbW9al4lupGy3
82zfTlRxEIhykE5vRt2iwjCBB9kB69sW92gzp4WvSnoU584l/SiLsXQhhNQz0k9e
VwDn1z/RyCP51ldB0zw+Dd28ZvvfMATTdfptPdi+PR6DZvHw1/KcE4yQC6hJmWxs
3FJ+WE9lDQotESdDX24y+sEFqWDMu59GWDf/hVEMgzrd8zjr1wJ2gjBFKUjb3H+9
iwsh9Fn/b5+JYmxpEpCHoBFCft7Yj4dlMvPtHE6x281ElCHbDS/JUjbv3g/EdS+5
lfgArBl+yX4G6EpteJ+nawHizh41fqoDBp/LzHcD/A9wuBhmZ5h3jX3po5y0hncg
MrkfD7DS4Uwshn1rovKeF+ae6x3kha5XXYR+yY7qTUaAeuWMbKlr4WGNbPZ4ce11
qMybBdc6PB8b6tpHHoYW78TBxqIYlgvK0Aj3tkP0HAOQeNKfpFv4fDKJxXDtZB0f
LRiGHxBwfsN+othBio0DkthArEGRBzH1PZ7jLr0QD0K5jASGvsNHn/u6U6xpRvf0
GQWDWVQXCijhZagqy08A1E3j5QCx9s1tmDme1TzUnEQPClMZ0ZeRYxsaHTqhuJhW
b53Us3dnrtujZSf9V5Nf2BUAmBbbHZemKXTOh0iq5usuPBJ7rJPJ0ZNqaaa5OlbX
LxObkf7a/+qKAm8WiWYpXr3sJwByj4mW2sriwu0qEv+z6VrHc0PEvtI2bUQaX0Y4
4tyjZGZtUT7+pSBlH4KodIZxXt6tXiC6mS6DteZbJ6H+uDmkvJpetLXKk53x4iB9
INwm1qjVFwVG54zl3LbTFgrCvwlwEH0/d32IjIMl9y6H2l9vThhrfSZS4af4CRKP
0qUPSMzX8kiMMMZ5rQkl7ujagLQ4iGXZRtEQpMApwHjNu4coXOeg4xyIZXsYRjd0
EEcON65CDO+dtD73OMRWQwHb8gSb58EV1Y3pwy+DTB+EZXFywvDdaHC/SZKevmTG
V8Xrd5vc6X1cMmiBXeaX29uV6xukCQTSPQMUqiBJ+Ix0Jujsqj7S9Yl71wWiyELe
NLmIpEgcIfmzWw4f8vyKWyhBPauqTb1b4wVP0IwqbR7IOuZcELIPcJl0xt7rhWH4
WurtZ5GRFnePBl4o//O+D7E1xwjBt5KVowjqksKmtOQWWLL2Ml39vOCAw135+aOe
YL/OCbxmJcfX/zsXqkMm00wDu4lQt7KV+/Xk6h/EloCp5qJo+m2dIoAMuXp2bbYO
q0RmDCjTgvtIdQzv+ob1BDTLIJizhxnxblaX/f9CIqJ+F6Yy2DOjNiKl/h826A+v
U6/Jxmofwi6veyJMGsVIxAuNyzyLOk1JhaqOP/padUQ/iWWQTXwu3ZR6dRUtg9Yh
uqxOv9FJwnfdVP8gyE0YFoG51RAlDmgjlXZXQB6aGF+gJlAQi1Lc9FBkdL7SXr50
UiS58ZRF6PAzsW8PQJJhaXnfiwt4/C/ith8CL2286yq5VdHhfuKbKOMQ1O+p+0dZ
FJvo7xXFycaHCtLTyFJRNAYbI/6nzRf1gCd54sk/kAmQbkeQq6lH0vBpxJ8aMMEq
EOe48fT5KI1h2eiODgVHVg9DAjDpomR2QMLHuwtfIdA8ikzhLvW+rtVGu5Cbxr+z
2E6vgkz0FhwszqDgUDytMrLragnuPa99x69MIC6szxFS6yIv9HohvzTPV0fOaIIh
kZ9ONAGwJ5gROYswsD9gG4hyneesdGGGtbL6FuL+vpd2gvn6XRQ3mH64sOeiJigb
pR4nd+Xn6gBFt31oRpB0qqOKmmuvjoJRXGGXG3XdhqAWR4mwzKIPJ8Lad86F9T3w
LJDqjUStt1sHAGghHE4RSXJKF+mAKV11LH1kBiiJFC1aFQrmehbeLHG2bf2JZwbw
zBrxNL6G5+FKTCT/bgGLV0luMzF5uoCH7CD2HhzQk6XVlASbVI20OtbJkWc46cEo
LUqLx5mP5igRqKpUnnOvB9AV+FiGooF2QIG7h1vrDmhDuQeaPSvcNv6Yj5KNQrJZ
2mOdK+PwqcKjpZnhmwnOLuY28neemxCoEg7fyQAoSAHRvkcaqCIacFG5dqRfdOih
xx8OWsu99bhME3q8dkP61hMgswOm3l8N7nfhKVBAb/hD9pGYJ0hoW/bWBPAnhAIT
UpnowqhoaQmnC4DCgSg52J9W3nXw2pIPsuDdaSuLmD0w1U7qOE3J7ej1dSNP056q
LguDx7SZCOMwjtrUJQdVUVfO5V5TXSxx5pU3Rudoyz8UIdA7g/PXH+ZuIfx8fh24
cfLUzWnhP5gAWOcVwYwZCDvvdiLXmRzKDQf0cJZG3u1KTcjVUGjf3qVHvYUMpvEj
mui7RGWFQSqXhJhG56wY0Un7IFEQXlFKLfOkV5rZuMj8VhZqPB8KYXN10jO+CuR0
qVPW70HnOZhuR9+/7HGFSfkJ4UTCiCm3v5keitGoA2uWzBRxa41jylZVjveCxrO0
1VVoBLSeyeVfVmGhayxpuaqPuf1X++iWR22GBZCtuurGDl3W2bNaAg9AvLlLw5zK
ikR/vcvgRWUH0Cp6PtKQ9yDx0vlfYZhxoJaBycoNH24EDky7UVGSd8M47auEKpTe
802f80dri8jbupnjFAIfwIcKhccr+KWPe8HTKKTOX1g5baPjwbMkRjcbJwDsAE7w
aLZ+E941JzBChdUI4p6MeVv9zzlBBWRL+pYlJ55snVjxy1jmJqx7jFZCgBWQeRQQ
IcZ3pWiyNk3YqTKhaykL6xVZvC2/p8U4YHrXPh9w/mh+MapOkNhUSHdkwKHNhgwJ
od0MNfoN8Wnl4LZ4huUENCGjdgpdsnwS8OGwDga0hwRovp+SFyv26QPkyQ4QJLVN
mzb2LOIBTwbJfud5i1BCbkHSOH+PvzmYNVhx1DffAF1LNShxyNtRemUvQpf4p0ya
1rIFZO/C6wBlgcLBIz80iMEMTFMf2CYrPFB/3oNXC4Uk7DGI/aTT3v9ZAil7Bufs
4Hu6BdqW9nAN01nUK53ZOYC5EfoczqesAjTZJGQnsDUjT7wXxghTQmXOblNN9pRQ
RoV/lzVyf/BlYBYZY/0chv0seR2H+wzi7nQnxOMqkAUBhi2NVi6HmVZSJlSZWABn
A30NwUR4dwqI7s705I8xeQ1umiy/dvOIpwU2rmtupaLWu6FUt/YPdP/KxP4my7ai
j4wZIHX9DrhB7FfmJMf3JTmiOuT2sE3LbbbTQzV+/vxZ+iSYug/lk3uMsA2pd1K0
5q/O1zDVcZPGQN9J58w+OxNw04DYwxfxwNzkwKe7XtDHrPEERqNbz0zhgZvJ/xTx
OXjX4T+q9JqzRqN3nzTBd9S/XjNxnTx8Xpf1Znbux0OTI7qOBd9rCNHgxPj6Bs/g
aNBQ3Bkt2ra+hAcb1w5SQ0NRUc7HJdPI6S6Ix2CCo/RcIARNRInseTqfZ1nsa68/
CfbAPK/cqqC/ofMc8+HDGVU5CHEzY9yII31KXn/Ii9E4LUCYdCtn3mEufl6aoakD
uk0r9OfkdWU9LM3e2iX5u03tgyqQqp7503sb7t3psnAZceOTP3FwB8VFELvh1zA9
LxqkIdRkNU11J9SFMRv4pPigJyy/yF7sGdUz+3lFIDf2dtMLjITVU5zGNdF9/2YA
A3AMQ2KgRI63j+T8UIkF69NbZnZQnI6yMAZTjYB9+9PBgb/seC6kXxccXebmtnkC
fiqcttJX1LMqg2cOfncFoaSQ5zJxWFr/fOzbycnkT7Lj5915iiW00DX+2FajUmvb
VbSlQRl9ZJXJKRi7XyELWSWx2N+AYihvAmKXguep8tV2jWn+f309i84zMzViXsZQ
M5/Pw6BhdMDPvBqlbg5w/Gm4vec1x8Tw88i0ItO9PJvZsvMlYadsPAVbo3o1AJyE
ljNG3rE18pA5Ta9lcyuKYX7FiWo9CkZlzalK2mVrSvtAlKP6TMTPzZd6b6iMxmFj
XJ+MEYlTO/1KJz1zy760A1yZUsRBW4SDhVOuNJZw5vhfkiQPG4xvh2/96AVa4Pz4
4ZRVhOdcdm7u/EPV1t5UpGeiqg1xojQrFCGcX6FceeMpJk2d3f2CrPiFHVUUJ+M5
32ICmmnjeRv1OcCel0riVHSL5ZeU/mbRJb55LPR0anbjHjnrRHnfWuCsKeBqYzWX
6y/wtLvnHGVjp3/usML1WnHVkshOOIGSFAdd6jvvQsBdhpXmcVccv/UyQrrIVrXU
8eYG/2sB/hGsmolZ0cQLJ04B7Cw7wTJ3X3BIsx5z9c2P2Br315y+FiRS34E9DlYo
h+S42CCfVMUWwRCaZNgjeL23TDUZ6QqaqieeN9CU/OCZfs6yvBuhS2alVrwsawdb
ALSGsYHax1TZqn6eyxaKhKoWems9GjcJhUuzQN9QtWBkw1069WRL6WfhKXvtoqaC
sBJP+uXOFw6LFHTmk+7sUAVLwH8gtWcPu1PTf/JnwBaTt21HSMaSDy3JYUeE2nCy
70Ysw4gwo3atkT3wj3OnIAlUzcHp0KoWA3yM7YZ1NU/XmZKu25TY5XdMlUgZLpsD
80xDvhVe/Q5mfjg9HEtnQWDeIZZvyuC4SnKpUVwuDivbjLZMtjeZM6OGUmA5/rhU
8J+zS5ux8Nge54/yAVz8LppsLQA3NJnoF36OWPJObP1xsGbvsXoBh6LnjTqvOfzo
NSzgYR5/1N8/H73jpTOwEFLtDQ3NoAk2LlbHv48sFp6O06QX8RiHTe5iRDHJ6Ql1
BSIVlhDMfjfPPL6Qsiw7BJNagQ/H7i7vVLAVigwcydXUrvFLz1OsSdaLvzhIhR3V
7deDBxjlMBHLcbrJgrLoxCxE1XJHfKkI5lbUO3MltfOxQAxi1lGXmDWPbGYJcIGN
`protect end_protected