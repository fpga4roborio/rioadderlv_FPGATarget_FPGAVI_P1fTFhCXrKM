`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
ddtXksX2+yylW5zu6QL2Lhnb2d1sD00763mmSITNX595NcHTEkwn0zB1Dry37fOW
FufOhVzEJp80NC5qZ/+F0Vk7Ik02dIR0elf3clrjeJRK85K4e3Hoo4xn7YbFUIms
l/8VZSb14+JVGURjfswrIyCUotIzlzVYZ6gzoZwDXIi5gQIBf/gI+KxNXPaKV+PQ
Ufys/12rjO6aI/pPlqSm0hCvftmBcnezN2hk1UeXgOIuKZnogjOsf0iJVX2aOOWE
6pD/psybjbnsNB6kH5uFTA5frkzIzkzl5d9+YDm9OyC+k84E83I/7/j+rk4L2dah
QJOvksSIzN867/4Qt8qYTQ==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="MvBXkzurAa5VTw+1JJ70nePUfoQXBvZOku/SMmg4TwQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
oRtzZL4VJ4iwysPsC8SXYCzXS8Fw2gtZTOskLcDV+1B9Nzn1zTyNtlo6lNICRmmK
ZRVu2BmCc2G+fmzynYlNTnSa7C0Cuel6FYpxCBlOuk3OF2tzAmLAuDyOH3Z1Yjzk
a0aHuoCdIRKv7BrZCdALt03JeUmXKPdOmIlkVGFl8yw=
`protect rights_digest_method = "sha256"
`protect end_toolblock="Jn9CQpRhJt4rnzZPRk+dOpzAubz7omckX1MrFd4p81o="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 13968 )
`protect data_block
gD6l00tciPUa6pDNTk/+t0OO0nC/UTtBwLB41d4inuAUA3i/ALrNyoJVcBnAmEQW
ptbcNp5fxEUJjnOxnedyZEuEBxWRieZFQnkRdF269oOe5/yqdGFvYCEML7PlEOzx
lUCDRK+jQ9bSm62oEvELnqxhguR4lH1GEMFVONTCEe+b6rjG2sGopDgF0KoT4aJM
SiC7wQjREQEoskO97yfbCWuT4qHidOgZ9Tb6VQIPhXfw0K8V7PGTiUHcQA1kd4H+
B0M0XFG1RQLff0kiKUjx5n+hxVeXkhNyk2j3X34NtVvydrbgxcmckbRz1gCkGLqF
SfPxBooeRkPVf4zQJYzU8kvknla2d8OoEE+9qMxtOC8b09D0HPxz208k5UwM/WLe
0CacMAsYawxuep1oRIA2ATcAWRmxDB9tXZm3/mE/YZmYeKt0nhK+7uAd6lXY0CjZ
2xIQazjT4QunYsmxsJHHBsuv/1+ZZ/j/frGjWRDLF27hYC+vT6NhiE0hXmlB/3/x
liCaXEnjDAiTaR5KxhmklJUo7cRAbax5cRvzsQt3J+1Hdv6vA7NZaC0i1pvET4eK
JwndM1LL4H5SWEYZ2BpIQf1eNTcw6Ys2AstnMu9xambq6EM2/YXv21rkyMEdfxjf
BRBYt0MlrSniWTZs0IWi3JZ8XeFNcn1oxpxSwcD5wOeDyd0991lnOJOhdNucsHjH
87/2VTBkgXMzHOVOQpPWX6VbZ/8KQYU36/HxioKvkQrRYCUmp84wfbr4T3EuNUHj
q0JWS8r62NwVzkS9c45oLTRQljpGwbB1yzDBtuLCWtoyaGQ4+CQoRPtjl5tdOVSC
Byk0bW+yfPMlWNcpdkhTvMBo43mYkszpDPdYSy6IjR4SgMvpurYKh0dMcZ5jls9M
htyHM453WXS7H8kgN52KFOxI+BDS1jcoln31aH9sk6IEg6IBRSeZ8zy3p2Bzyuad
cfAUYn0ddPE52VuTBPS7r25jKIR7qbNYjjB3WsEilfzWsIULj0/ED91dymvlZ9Hp
oI6IiaFvyfzMYkRAZPDtUsrYo5PLutRy+exYHeMsnj68Ops/hBTjpb1p9RYrsIO+
gqaH2Z2oZDoGn3gymfqxnRbOwFTOMddGs4o6w9bdz6epQ73L+0AviOfo8LGltAE+
aBjAE+9lNJfYdGdLLY/IOKhUcxS6TlGpESLYCoxLVYgF811Y9InnuCftIXUo3n8k
BpQ0qZycUV6tCf/8GcxjhjtWbb6JyDPT5/vcM446aA8Y6iSsbkBYceN16w3bV7SN
xIHDsCHFf9wI8kNqunD5r+uurgk3CGGwE2j3DjUj/KUyHzfNYgPKmDzZZFC+b7Fm
Zbduk451vJLLMlnRCxYz1382CW56ssRJCcxi0TgfOl254q3GDGvsczXMvrfmyl1T
Wa9StwvZAVxZDQ8MnmYSH6A9FRqDeKcVa0ZcAYSZ5TplruttEP7EQsFAobm7sZaD
A8iDPLNGKRelwq9LrIws9zolpsKM2aifQu13/Nk0U3T19d3feSFIR7nXfUoYSYmP
iwXGTMVaZw+LgEXaerkCOvpiXnGSHPDosBPcxt304GZSyeMC+fodTQM65EQVjE5+
wGoYhT8x47Nly34x0hopYL3dfc+3a5p3XFhDf//MO6RBkY7XYYmUWQ+ma+0LYXqb
IsXir5jkY0/CQzO913vCo8otRpOkCcF71ggQMrGxpvpWqr8yy8FQHV5sgY09oGz3
avUwJ9gUG5zsr2eeMhGsL8TKIpqskFoaiNs318+MGtinRQuH7CE6DSL3VjvNrRXn
7BIwNYKDEEaMryqLl/EkrttnrGhlv799ULRDPsA8YBXWu/KDAgFwy29N6StUfISV
dE7ZXHaKY5Id7HXhHkMxM+PWjEp9qdcs6Jc8eLFgyIVR9bufUB2yCOblUdpRu9XH
/ir93Lr5v0qU3+6/U9ffu2a4Kbnjw0dlTv3rZ9Wim73Vym9OUT3BuGPkk4d481xM
jIRuE1XOPtZ0DwM8YyU/bICMyZ0IMV4RbW3i+teDfqwOYkeuuFfjQF87CvNNAjXs
e9vDjojMwQPzk4XZH4vA7dCvRt6Er7F6qJPJxO7bNxO0mV3ZbqvWgIwSD/xxzMjd
zDKyZJUlTJFff+SRh0+tgCeD2D0HTk9XxlPSthtTnBJlWFik04vZ1bJX4WA5ZOGR
+jG1w58DY3WPNd5VYtuYi4QXZs4QR+fC/s3mJjDBcdE8PoOlIcxRR53349NQ4/3t
yIsZqRztAI18/alHgl7XY1asNdWJi+5u9DiC/3WgjlKo05gZL/QP5iVbS4jwW6Ht
ebHnyojD5DZZw9MDUBGfyUt4YkPXWgB/9Dd6YF0C//EFgz4dvWipRsHX/4Kwf3UE
yNP4IydE0gX12SXmaWVbWf2w/4X5t6QEk8a88exJDEbRLB7lL5F8kW9RYJfsnHRt
OnOgXRzekugY+36B5cOBgZWy8JZdmOsmFdWYYBcxGXLnDUv675KenhJHpj+BMHAv
x8syXS327WAZztlk5tblrmUS29AXK27/lizhgMuEhQYK65nDxHmHftlHQJzfRfeb
JtylYRW6t6DZOGqtlE1t+aZvs0K2D8JLhN8slMEkQXAWYtTwOLG5CXYArYX3C1UI
Vb289tq+dZznmXM1T9/lapPXeXTMTmueMsLs/Na0nAyzxtW+FX7uVev141B7STP6
QJAvAGz5a69IodoOWfJ80IKLigDK4XoNyw+LudhWQTplIjxcAMt6NacV3J9/HO1E
FwCgNjRFu8LN1qedjSU8ebqhIdaSM0PKxTIaGuHISy9bX5j90KkuRXd09coqR4Fq
qr0DXLjKCYGVwOjUWtDbc8NaXPKhOuYfrFq/f3HOs9nfAdx/WnyMK8SrJMcp6UAk
mGwWHTWa9eb5DTuTxzRTGJQOBNwmHlGqhb+lVoXFl+HakenZ/u/nNkITClcKLObp
EyuAsoYdd0qJy5uzGSUgpNwWUHZRJ6XW4CPeWgjSGtTisoxEH1hDVhziJ05z7Mgv
TDN/MbL7eXvqJzoxKpqDUxqdCQ8kT3vgbHHxntca0c8MMHU7PKywHUFjRt3hZYta
RDYDE2BIUJXeWgX7R9sqfLcrTOOVUcTyBJZ/mSwHYOD5Nfyr5yCMQ7GGqVbKpka8
iFFi2ztLLW1X9OUheZvdEXNexCWFCZvalCGIpphJWEDWR7owe0JE6sXL3E6Ica13
bD0LTxAooATaRTq46yQfAilrDaiy6GqwOjni4C3zbSJUEvfeIZew+Q0ZZbGd5GEF
CmzEfu6hMvP+KwVtOoexdKQmbxPXPHkiB0UVxcuF+FA7t84vk+rO0VpP87FRBcMw
50LhIhpJ8zXduXHbrJedw76CtuA/DNg7RhcELtotQbQLnJ4q2I7a3rcQfnskFiid
yJfc2rJGsoN9GpL27IUbLVdJSoFyvvtt36oUE+P4+BrNopeX44jr/fo4GNpp0dRO
eiVVtqETYjSdoVd0P2KPFFjqeXTTsQBTok2uPKuTB8aHsB1awHNcA9N8BfeDQCcm
9TjZiKcwngCiWJjCMjiEnyUX/e4M5XTOHAQYvfCpf6+YeA3fcE/lGpTJF/m+qe/0
tP2gqhoCRwv0FQJRrnFl8JJ5CSb/mo+L9ON6rhjtTJQI8jfwQn2DPZ98lsxyJbiG
EyMVdTb2nUY56yRDbzxUv7SoEV/PWFMIW/7r34H546cnMAIhdE1mMtg3OdfdLhoa
8M4L2Xp0BBAt1ECn/HzNqqDwrmCTzENeIhvRzrT9/u7Pz2olo1+Z2A9zwZe4TiFV
ih3RN+qzFVVd1VudTNDmged2XNCOSVUmBr+HTfnhmHgwCMngQHqr9r9h5xq38cO8
nNlwFcZtyMojBAmR/eSPWTaFSms5aI+7h5tttMMDU9ZycA7IfDnGVq+gzUV92VPA
JsX0DFXuErya3M69Nlu0nxEEwt15vZ2kwhpevDgqafF3FalO+N+Vw0pgmRxKgCLM
SzVH/N+drjGb26WOXV+ylzxuzwCloioIrHkuAbN+uGltGrH32voanrh/gHNOfGdl
Q3OwgECExDTi2pMjU7HrcwgrB1pDHpjfyrc4BDtAMcz/T3ISgXjxhbp6TCi0ENA+
pe6Eg1lQP1p7Qub98QQZ4jpxyqweCKZyGWC2ykr0iPdyWlQFQR1RZSGkYUrjKGdY
rr/8anfD4G35S39QwHmDoUgVjM8pMdQ4dEFYOxyPNPA5FBcjE860w2cWWKfekbA8
fMAUkLTsWFz7gRK5F8fMiXEflv2AF5DTwXT95w29x2qbwal7kMm97sLuxSCxwAMo
ou5PoSylfNuc87AEQgucFWJVjDfeJYTe63p2AzfaQPENFBG2VRqZrkCUGDmVVCB0
kI1ZerPcDOwyKOEbq/cg9d2mJsXjZZEi0GHZTEsi/M7aoEvnHE32LOo/8WATfLh7
nwJVTi/nqBaQU8JPPZPYTROXWOgpQngYJbfNZKQWbcEUN3Vpc0rfPA2RoDFKk7oD
iZrQB2NJvJ/KPayJLnQOl4klPqeDxgrSRLyrPOp0gMA4jYEwJgTtt35dtt0vTNU7
dzNrmgJyGsaPO0XavkCCpMW4SIIk79gly4FmyDjAREtfdSIl+iBvq15+EWUg/d5P
oDIblJvL4vMkQDntVKtVUfuGFypggJNMYURj/1HFM80RjbbBgb0H3e7fF6l4uzy+
HQJvC1sZPcS73LiDQTPkdF6Y+Gq4dx7ZctXJfsXLCU1KWhmT+hQbCkLgWRufawfr
RwYUbh7i8z8PZLvVK+jA7/qiZN82hFs88N+nAK8VconKekniS7RsY/mSQ9wht9bt
dxh1cBWVFKHRJOveMMr21yeUlrgZijaueWR5jBhPIAyG/ZOqKrkQbD9nt1m72FGM
pV9vi9h0Jut7aCumyns3dJA+xyWyTbiNZ/2GFwggbrVkBZxdfo0rfkY26XrlDvsV
ra4IYyze9Ejf3iJLcxqichFMNc6NdR1KmdUUfodLqnE3O+7ycQC7QNR3xjVJXBv3
qckC4TcQxEoMKVoqDHz9buZ6uxF9g9KbQdCVCcfm4+LRTqwrY5+ABRCuRL9eJeFX
gyvXI9qWqXtw0j4l10BdxBFdTc8Tm/Z3Zdw2riotrYq5KU4q+kZ6C6g87wcZWKwN
EfEUKbcdpVP4eQQemuMxHWyuEx/ZN6KrLKlV5bHAUfZ+KvU/+GZZ2yzwSnE25CNU
lMPksT0d9M2QyzmGs5qmA+sOBw2zwo71ntq+95/+GV9E45yfA2o6GKELuVYG8/n7
MN4stixv7W6pjXmyi0oZlQpzJV1SY8pk7n0+o071Q8dBaSHaw7tewXrUip6KAAb0
iymnWItZNDV86riHHbXF2f7LXEWo4L4YMv1f3UaFSyYoWh2ycdkH0YXC0v/XhHJ0
SFHL+IyaxsCPtfUWZujcaQxFYU5g5iNiJps63et8/TiT87igU9CgiRY5wBLpuMVh
vf8QqMmmfNCdn4reXMyvyOTjGNKgBtkEPhqo8Eiq2lwmHRGVvK+NWTH6r3CsT270
i3TvXCVOPcXBXfI0ENMcsuLFJFEwcaQeI+tNOkzkr4goc3YktYbM+zMwnSlwfmf/
9ssWw1Asy86SIl1amHpNamt7fWGwbUxV/hKbS3/qsXb3fWMDfavgee3NavwcwzLl
0368LVkme+c9gXZYBT3BWEa4AFZppxqZ/eCSzvNxGUcySgq4FXllnFn4SsfQr1Wg
5QYCkJu1zkfsO3RKnY9IjA5owRZgyoJvEyvxTd6YzMnfUbRlIK4uWuyyTifATgGb
pypOci/ZjTSJ3Kpu6J4sUPigrsVtVDIVqogT6VwY/RCLTLnUuqbbC2DhO5OTXZCR
IzCYjnKxasR01dDlakb1fMRDDAXccU/oUD/u+sjW98Cp6DrJaZZnSVr+ta61sYeh
X/yDxsb2MjUg1/Q2LNP4Gg33X0ND+3sQNWx0tWA3Yz8Q6tkJ7hRtrdPTYTT6Qbqo
dMhQAfvNDmlhNQ7HSswMWlDM/DdUhf5rizxsNcEl9Ne/6iywpMnWptxn3R0AdyD0
7vOAmsRvRwlfFMU9PeQTGEpDXwevsPRhc/ga2ISJH8OaUv8FTIIWdA3PsioDZDOS
SuIBwUJ0Y/KH7+c21/5881kfa3Mc6JerkEu2cdjACj4LAJrwXQanPf7OqKr9pdPN
y+x5TOpw2YZBd1aFOjXCOi3vEhUT21il3W8Yj8VICny9n6zE4W1C7d7FX1vc+XkP
YXDuKULdXtmI/8ooRMrnrZGmEdP0QDYilVwp2Egf2qLY+7QcFncguTWY8nz98yt9
/Xiu8SFbrCHlomkqjo92grMlKOF43pC02gbR2ausBlECkSLPzdq/SKPtcV0YBeDx
CyZZkMn8oHlKYnzthyg5jwOJiM/MRO7eqAXpH0w0borO1ggljCorHu09YKIKrGTi
A5BMIe3ZvhhB8grC3IDT0rjjACbyQ5aICDWBKlPQWjBsQV2XFAle3w3PkBYHwKs9
9NLEqrk9WmAlmdvmcwQ7ibU1gH7D5SpdOTwUArLuTelZjdQYl5jIw0H8el0fE5Uj
t5TRKteMYy7VrF3Qh86aDBFEFDufgiWXoM0tmvMkOD/Pcu301GVvCKjAjL0/tMZY
9wwS9jZgF+0AOLUoW4UyrKpH7wRj7LfKozIuPVfHPVapiNyzn8e7yRsgzri/0Hv5
aLgJ9ALHVdbihieZ0mIDgxuf5qiq0Wjv2xukkNZWM3aUGksEodJxRCOPuUcPxgQG
CPKn5HOfnuhvgPStkKCNQP1HNvEf7a/HxiqBIpVCVFsQEaAMgdHfSpmlvr/hBAEg
IozD6YQEZDQfQevoLZ6dtznUKDQKLmDvJHyejb8QYnXlTUP/mnGMp9X0muG1LskD
3I6y3zBVMG/kWD+0suWLpxOfLisbFkSWZrfP8fCurnZWlpvBPhBovJcJe6mKZpe/
7VD+Rc0H1G7O3nQZlqzNtxlkVJ25AQod6m5UKDTu7Q7Zq28HT80Dt3ZD6Q1HqQSp
dJpYNHKPYjay+nt5WY63j279/aDEr+Mrv8iB+MEv4kidpz4OpBDfgu21Zi6EF0xt
dvRZu0AOW3xw+qoKlL0fhRTIYWDfzIAnR/FdFO70tg/fzR2czgMZYecewaKGO1dL
I4HPW1tw4L5Uw/Q9PmxTxpnm4ifuejQd2ol+/IpghxX/J3NXn05autpVhdleTqp2
sm2QQyaTWpqsNPkh6XFwuh4XGGtokl+gwEAwruw1dhcvOn11gS2VTZMYQ23C7Xla
DEiccgiCctCOJ5BrSFcR56dcSh0dCun6zXMZymxSWZ4pt3nzXjgXV6aEWlJaTmgR
7kKxzMoRmZNaCarJdY33t7GQkhlwfwn4/LEG+rsmPqCP/JwzcOhGcOaaa+N3fAc+
hZ7weZG4eB7rxXNAOXWUFQ/+SJUh4bVcMPKr6oAcKmE3cw0s3JYtnPJwolZ3lUHY
H5Z8DuSyQCqW9Lo43lM54yrFIfT62C6m/4O74JvfrjdEo0ph4vOZ2tBMC7N8I4Y9
jA78OGgGnoy/zJjc7uObLd3g1s+OhchrqULV9CnDDPKCweWNHycomLCjdf0ZH1Qc
ERzR9y4b34Y0jAkQh15IAxvgUtoFAGaRKrxNN2zIIITfcaTHc+1scDUfeMLA5HO9
3vL6k2JfWLe1E0sARxqzBWh/jJKDYsuiZzGn35YltDwtlpTNPK0Tkvvp0xMwXf/4
iqVJqdl4XYpquHx+0ZIlaijOc/YRjiT7nklquZQmNX47I3w9isAO/J1XRHPbwvrq
5KyLAhC4Jde0JeQYB6UZpBmVaDUwmIra2CyL7gzY4S7Y5zauuyDFqy8usZQ68NFo
9cBUJVrrEchxnRjDie/NgyGYFkIEN/PlskfZ0mgFsYzTNUOWZljj6YViuDDjgZqV
zm5IrumFju9cU7J1d1qqxghjAV3pO9KoJnpehnHgRXstoTLYHDzJIFP3qW5Xowxp
rrBHV7qMpJhu/HdJOITUWyYXYELXcC+6+atrf7QGNRQIxCQROEeGAN9mbBo2+j+u
WjQkTAVAVOW8xK8pzCieKKi580hs8izEB71H4xDQO4+l8DCcYl2Ac0bVefxNwK4h
H9Tw6R+9ZgVFGB6plArCoe00z7pqykX8T5SbyHANhYb/3PPHJNP1uILsBfV30kIg
2CoqkCtzVIzPxI21P6Xoykg9KcshkKjdqeQAxMaUMy7QskgxUpPz+Z92dbEvzsLW
d0gqHDuvvdX2PAS8kqzh4k1jvok2QwKp9P/NNjtra1PRWO8ciBKSk+p/SK49PPgW
TSiswIYXpWzSyjjiuZrVk20jLkjv6nyeBdOCcdMOSJISgDIdYJ32BnJOF4166CK5
SMTBR8t1CchG0IgVGjTg3qqAToEH6VbjPG49zOp8Q/w49pAL2EoExnO6Sg5F4jWU
GbIjQBrmyIp9fDisWm7CHbOkIOyUALFzdKvXu6TN9VpJQ90ugbDciPO4bm4sHNCv
usKzaWXGXJcDCl+VeWZUitGvAM7QJcs10HCkPyljr0LS6/1EDOdDSCf5B9cNuqar
QWGAl+YuiBnafxUUQNfgpfpkoHD7NxGDyPjOR5MnKRfvmJtXBVsGK8NTfPjC+Gl9
sbF+JQt1ZYwNlcLyUnOF2ubpfvVVJAshnZmcz8JH99MH2VhTxAlMCzfGbR8si8h7
NH785Eja9y4zUgQVgYAxM5WuJIhjgtiZWBj1DntiuEDu7d3fJ2fx/uDST3pVxkS0
QDvOCdaKauWif3BVdIehHsrcsIsPasl3wouwv9FPvG06NHmr1/whswmcJB1XpBac
AWv9sIBNEYXjPsWhsZPYL38fO/nMnuexLpNgN6EIomxMlVjWeUvnBrdJONxgp44h
Pwp1ftH0T7r62n6fheUsvFYSOsgCtmu+ghzA4mc9QgfxKV973ZQDAX9NsTW2lpRH
qwg7Rksl2hX4zu8cl++361KtTKAJyAp597CFUmFTMK1kjpUSRFAPW4cCdgCfPAbG
P5echIoS/9O0pbshAekiBIFHRLl+ohVBw1APIScAMmmTmxowA076mBse75CuS8nH
tSVZ0rMj4Wd3/7mu8FrnTokbQiTryHy8YimNzye1q+Fh69HjR5ZtY7uUIzjwuPf7
0Un2zojCo90U5AlJBFe4FT1SgOrhB1OI1FqNS4c13a5q9c388XLYF6TJDa0cZ6E9
2WseSu+6uHS6/iwRtZ/uV9N3wW8PAq5yOBDi7w3cw9TWgQoLqewCLT5MxwPcDnzq
VaaTqs644DNtMeMoS01ncsfFZgaEYbVzphB7yU1sFJWUhtbfmknVs1Yq2ITI3Iqq
t+jKkt5vvMk8MdpZRyl6jFjd22zFqu4KfotA4VLyb1cHTcy5fDbr7Q1eXtMhJ87e
FEzBXs8tFE87frYb9/iIYr19MMsELnj/g4PP5hGW+Eegu8SI85QDErhFvwsJKQIL
/MwcHuRwwVuQO1GiIRBMgVorRn9QqeeqCxrxgijg4saqVSZMPITr50ebtQDJNhzp
3A8oX+wNwyGQDqyftPeoXjsS0B+a4ZUJOhZHwW6cZjpn33SfNJbzdg4AIyslY6DJ
+HiduYzyhdmr7NnVna6kKZTl44UmvnqqPcBG+0Ogr93ZuYbUOF+/wqL5ZtlLUMiD
deYI8RJub0lDKIO4wWDcZ5lgi6WAYMOZvMbm+/fgPVOrnIrvaLGSWI95GNPGHDNc
5GZ0bvqFNtJtdb8cCV/RPAUg1ZdfNdBOqrLDt+gJh7HBK/HFk6abyCWw5J8M5GH2
WwuhwDRErfNIFpQITrWiIQLdk5VXsanKuMBFPbboH5d4EKcGVJoUawBkBcJn/IZH
abvu0iYMKxAlrcfolJlYrlAtZgCM/bbMSISRorCcJi1+TEVRWLj9gXCDns5ejx24
2c+1KcVY78nLtlBlGxcy2eV730urFMy3Qy7o0PrfQ+wWeLK/2hK8elmbuLQf6UJl
N0rjD589IoTsmVQUyGxC1z2Zk1ZHdvSONrC79Y/6ahYD3TGdMN3r1P12VekANfTh
hufWnqydIL/IUsNUh/GorWKLUvVLasxFeEsfW5uzd2NDb4MGu56zA9OvTnfNKrdv
YzFgm9pWLQLSQHTIK8qKQug+N3zvxWUylttHex+RWa0fBjUjK841+j5KSNSG6GDZ
y35CVOOTzPbXhJJLO0n1eJInQHql9UWePVuVa9DhnZJGkfY7LJ2kJlYRWUBSdj1k
6iBZqKGouJ2iAVI0nWwsFK460X7oJ8FDxQVuOEmT0OpdLsAZR1nkoKP5OdxHZPPC
n2LMhNRwR7Lnc/J5ng9bb1mKxqKNB/VrXQkQqvYsooqC0lPyakb5kK2wu1hmV6BU
PhfcxFcqfESNQqFeQUNqVAjcODumHlAC964RYYb+O1dLxvSksStCFfKd86BTPInK
aNpZqlg8iviKMW9PGJVv7ST1riTPKtbN+UwS6SMWJHGyFDtXMxy7Zmvw8mz6CQSP
ac5D/CJUL92e0T75vEe0vo0bYzjERuNDJghxojLNWho4qGTyb95Wr/7R1XowvNJT
oAe3K2Eglz6RnW37xOHxELWWhySnVSSWiGxxejY2d4Z6jm8HbRlIA9CtLhmMO5i7
UlLo5H3w44982vdoJ92YR07Sp7yytfiGtp3hCwSTimYptk80WolFDeL5httVA6rT
RTl0P98P7KkREzH7GhPHAiwePlQVB5xz6F1GqZh8j1wcPSYtC0bPnyIZC1zaSpuA
mdFlF9FVIGEI9LRErsMnU0E5pG/xVwuGPmILQxpianWhHIVhAN6ixIR+ld6zPssd
2LzY4KkkP+MtLDJfjPWOkSgTlQFco4IYmikvLAQrNrSKumAwpAlBGpcYBd/fc1eF
yChUIluqxEgByZJyTQQ7RuXBU1eTUmr/aqYTbcGq+Tbcf51qQlSe8ZkvK9oGFExO
fbqubRdP6iDrFxhZMK/P0IULS+amJgCFbvL/F4jLT4eUaC8ibOH5n5XgY4JuVhrS
R9Cx+jLRl7tS062iunkuVFbGIUKwSVUjkNIGK7ZkaewvCnLVTRtZ8xjI2JOxZAEK
NCRp0iw5rRB8R0ArUDbJPFqbvfJpmxMo5Q5cla4QO3FpqnvAezj/UOfrASkLyPzm
f4xpESNqhBJzFmhHUcf9qE658X1vagGimR+vexrcRkc55iDduyswvhLFD4q8HUGE
gm1n/OsnZ8nv2SuBM+e+bLRxuetnWSrCJ+LYA/9nEP8M5FTByGM+d2x1WhL5woED
aGxFGe2bEXulVOV0anNrGxAEm34CYgkpi+bEp3ytrCm0r8i2xoDFYiUTrUQZMoty
Mvohs2s1/17Le7Krrkrr8ugkM8ERQ4sKRABIqOIBvR3pCnsWTZH7HTAV8YmHuF5W
oeh4h0CJ2Btk9ZTc2Sd0Bo0qskMo9elnP1KiQiD1ZCvl7FhRZXtV90Nt6zOlyQ9Q
LM58Pk2LCwNclTBOMMSRiU4cPizkqzR9cEvlIT2kmxaziJmZHjFCInczSfzloPe3
DHylN2LT3W7jBllBniX5xGVk55yx/Nv5jPWT1OwoGfYwZ4RS1e2L13g05EpKAstP
39Yrx7pmiTBHV4iWzEICAjo8jLe931FxlYrWCi+js4Jj2h3LjvDCjb0pOJRAKeFv
DKUMMF/o1yLWrCpFHCdeMF/NPFSkaPt5jS2KJUSxqEOg9tbFqiRwwRyjqPASekpw
dElDM5+u1GjNlOfxubtRTIKVnENCenlLknI5CDwd2pHi0jVPKRPSNO4w6TacKfHf
kRlOPs/Mw3zj68Zl+cvWfimSpcvKpD8xS+zZ8IKNBMKwrjSo75zyumfNGXtxZvwQ
+ug9YcWhgb5X+2hIo3bq6BcsFwADD+lN5d4uUndd3fOvRi5I6DKwLNVzn+KtNnu0
Mnq2ow61ziQnzURcnmJYfkLK7CUwGgBU9yJzA1Wm8mRHlAj2nzlUBljGXdMjRNnr
ZHUl3c25drl06yM5O8rtXmtuAu6CKl+OaH8ZS8wtAW5S0QVsUVMAfx7jEURH9ZwD
A8MQ6Ilpxw9ST2NSFN7ApgDr8bnISS2dTcoD9YgfK5BceiLjK00CsqUxLzp0a/wu
rNY65edJvqWDhR6mr+USiQ0LQcVDCz92cJFOgvS8b03/ts4DtW4gZlTevxiotRAU
4wFTGfAQTRbKeHATIFLHSbZ3tExChXF3hlxCOihLozba8UKgR4QxzeIUZDq8Jxoe
RO5LNVjCNoct3hn3lXF7KLXJ7CzIfkdce4FqnkFqmKHAt/4UNzJ+wAWREjkEP+6p
cdY7E66tMSBysre5CvfR32MR+K/LaxXzmbDaQ2McY92XRfVsXibkKDr+pyJz+pVi
qJT1PyKfFdzEfUx0OLvpMiMotX2x8Ce3VU5vTg8hViP1jvGUjWk4FYeqYlWi4R/e
u3YcbKAd1ZdIOCj/rDMKRI7xVzEzpd35WjhtKX/9tJcOK+zK+uolEH2pJhqiq7s3
ILgC/ZKRYp/kY9XdK3/wnlVzVDMfujoHAC6SMcDDIqmL5+aQ0V1DWtQvPRv3/0ku
72TuVzi4o11KhsDUKV66Bj8l3ZbAQQhZ227m3s/IKM8okB5bte8dVD2og6asRGld
qNKtcXN1VHswsYVo0s5byfZh/Z/VdLswb+SKyyIiyiP/F27h5bqa71G94j3vN5Wg
8x0Wa9WN+nl5UxklA6NV2uo6GtNXACljt9LeIxTVbYdJR9GBk3HMeSXVjP7k+guO
PeiPoK/2jdDt2z2BxRokItUPOfbf1TQCn0DOWU0ASWhrwnY08NULyYBS8u+y7Mgl
L+NXyV08ruFomYyt0lQEWYcdgtv/3t1LgpNutMAczW0puJION97hukkVmTOncAnk
EHcY5DNHMK1Kx9uScRyND7TMzj9woDfYhnlbIEVRdZNt50ei/SI5W2Ru5IUmSvdP
M6x9gz7mQwSSrpUY4Ph/wEJFaN8M7RDj90Q2yoOt/R0jmSx6z2xaWSRSHAgQnD+S
WLjlM2L1AsG0w0PkTsAp2EnHv/5MRaJDMD7UrUNlGxfNbLn9uoDobEf2SMr9sw9+
Rgss25Rn0uRLDaQbWBRNr2eepGoeR9V8cx7SoHCzOYdzG+u4AY5GPUXsf02+coUZ
pAyOJgVcos9ttT3fXg9329xEX05VH/o9r1i/nobBzm7peCtJa9lRRxOiqbm1r+dz
mVED3uX8Ap5R1wTMR+G642HGSxZbjopmCOkJQxlmidmiqNA6+kZMRJYMpXlr377h
2Bdw047pEkP28HyoQwRYtFvIla8L9Fs724CmI4MC1HtqG3DbALpesQnANNYmkeXF
lcMzPi594aYNEIJ/Nf6mEGX3H6vcUro75Nnlbdi7rx4FWqx/d1PHvoZpA9SwCeDk
Qzx7ysHocap5CpPSjw0Mrau9Qmc0tG4HIjP2VZ891mESKmCL/WsAPEpcOG6tJhjT
2+MaKhOBhEBpr6y2NQAOgY4nXUaUjTK32njfH9H9FDjlKwXBs2kAG9PxwAhk77Gj
nLkPvWqIAp6NewoU2RW617zXJ6OXMTVU0ya+ePtrLM22Gg1SPAPzy3cHTNNvIOen
IQs7s5RzpwwpZxYPJfFU+P1kBfhiyF4k4zg31DxgjTuxOqDbRZejVnCZLQHQHn4G
graIPWztnnai6YFDllQbmxm02AvkB7XHfNqJwtha+SHgmxva52YeLOTWLN83jaQn
6dpzd2B/jXpPhCiKYueJqCq048NvEAmcBGU4KrbbGWNlxL4plaahxCodO+eIP+eF
qeTATnjyQJEzkh0qOvRsmYeqcjkWcN5ZM24Qmhc8wWycMLIIH0m69vDlwzOzLp0j
TsJ/r4o5/uE2YtUVtxW9IKLmp8InjB3SlsvkIy2PL0hRFoGXQ+zMlR4w8B586Ocp
4glAh7y7OAJg9prbG85NopWXzFHu+fHavoM6b1urbLEO8fuE+inesvGH1+MtDDC5
H/7b0MjETxdZxZ/7tSAt2ZS+VkCOdgcmoKOqjiWyun7QWmu68OMkVlwcSJnYa1fP
0P91/wHtVWdhAf1WW5A39B700T15kYWM9eVcGPsWUi21oAZuKl/kck8HaaeIoc92
NxS6qt1Mk6hoNM9l/V+jOJOOJzROWqKeZMnTaRnGxpGCWBPNxGX6/UWntHVIA/O9
84c6OV7SV2H3DlqumEGBZ2TsT/xVoMRWpsHEcUZdZIaQUC4XZJ3xIxGAFd1D2hL9
yml2JgKP2qTQ4S1zIID2quQLh5bcivM06BAJ8r/GhZIpNO2L+PE08plHqsYo6Std
3oW5vyd4XXESCQhElMqyGr3MwKFRn2UPEBMz2y6twS+VZh89A2oTelbcsA9c4zfH
7vD3JtPUmaFUj71APmffVlZyHb4GU5IT4SKjk09V4xkS9WP7PymYjw4BQvLf6qDU
op4kRRX5z108WCkjhDrYjtLlgmzY2JaSTdQAJTBYWU4KlaQRfpDcRnWATOOvTqC+
Vgtb7ssad/BZdgOcYSyccCUCePU1yQlhc0NmnmgYf2D7V3ybS13yMUO5gk9YhDSr
CsD77PodTMagbrcWwXKiNFdAibf/28uS5d3G2/5Tr6N6LM1AFzbabnepIwclMwiM
ih+Qqed98rbItVG9tW0vDGxF17MFPRNNKAIevxG+3AV9xi8uTrbk4VstZoIgT1dj
YuDIYLIj/gzPAYtsoqBb7m2Z6J+z6JMTde3HuaTq5s3R8yDoTvVYx3OtVCDe3C5t
2xItbZY2nZeCdCqtzED8n4e2CuANuKV2ODQFreyFFh1B9BGSx7I/o1vAEdMVWnCv
9dCwHxPchO/8E82v/QxyMo8j3FLn16SaL5VlfRYlT/3Yfjt2unnHDX2W8ClArQTG
v2djs2HvcnzanQEabcVoXq1soYe479x2kHJAGvqGK9x0VPsigLIkTrMfPzZXl8QR
FYPaFlFs0NAAkUE4CmWKjRcbtrjjRSGg8LvoW1uN9wuKN8zSVi1q0Ht7UGJ2XaBq
sfJrMKq2Q77RvD1frd7TP0N4o+jBSS7+TjBjhDy3w+kx2Jfyx1ZkHlnVzXW31k/2
6+3KH6PiIj+L4URSNvzJeAVPJEfRmVLBO/a0rxAZhFAeea8BMm1oAve5Lxv81fmG
/CnkdSepsOfc8/M/bTljAFr/sJnWLirlZhnXlq04JIs0ynVlSbJ0I3VD9BOaqi2b
PX2Mnh8CVSBA0Gwd+RermdhelIsXW0H4pQGITc5xnl0Bq3R9kDP8Sdm45glmlEgk
oXNZ0DwflTF17CIT52R5O8c05XVil+4tUKxtA3jpD8IjepqPbl9rbkQo7KmJflTs
VVVLgvyuwV8QqRaVfOQHQRoQ5LfYiGuZyFVPEPI3wBe9eOkobTLpBSXfh9Lm2qZk
4GKCG39wB8ScqmbVAuoyYB9q3C2rGYsDuNzYViWZ6C+LxgNd11HFE/Zl2aqWL7v9
XamZAb/wVl9j1Jlp0YYI9sMFJ2sU1C/8oIvjOqZ5QQykyfcjQpFJ17G31wcbaiIy
8DncS6PVpICG48G3anM4UaR4O1X7GkiISZ7HU56176kydtQaf3BXnusbY2/CK5fW
4slVLqSWSikMawtFFWmf+ywxlPOQVYqnHSS4xfAgba/VPcJY/425wGqH7LfBoAuP
6c2ldCLhyoueFo3glqeWwS/Ota+FEYlsTVg2MHLKTJG402uI4Dh+mE7BTMTyliZu
s+UPBfDOVjaW7cZZb7aECr2V6y5IPyKQQlS58HBQ+IJe4Xg3QUj3uyGaLEtkvuBW
dXqHzPtx3nVFnpVq/k0793QgPI5uNb1pB0/p2g5xR8eCjbxUqiZs8+PH7f+UkPk4
lX0Mw6ALEGIQH6wPLBxqxyErxBUslXnkNJxLa4T/anzpnmMX+/xjRNzT731umUJS
yHqaVqfSWB7eKQzrDmheMlepAeXGrk12r9DBguluUcW7UVLFR7ER4O3yjURR/t/t
Ch+tiCdvmNVmbwcDaoceu/inpsVHuPENbUSyg/zbXgm3bceWbgFLYVv2+24cDhzq
LmAqgZFzQeND7UdZeHdSx+z18rqgrZ4crbK9YSjUrd95UVvr8wpyyedXbTNByo9h
7CpIhZPDNJORVpSlnkfMWIy9QDwkMXuYhLCvvDOy+h/b3Y1UHRfVJXhLma9vQeOc
9MVNMXE1WoV/gzfXaCd08RPD9s/hFiF1IpnFPGSKL/W4k0ti4RUvKwEeftYD9o5M
7lOA94u9lK8bgs4x0ILLNXu+HziwYxVm66vlTCYOBlIL+9q5b5nZMk5CEQl6KviT
cemxadtFwslhmeMUVcXi5iJnWbMkNezS28uSf7NSHPTLL96HuP9Jrn6dTfOjLdqP
4Mj8UOacWyWX5R98EwjbRjXtRuk/lWo5ZEeSxYqjxskeLyzH2bfRgzRKPeG2bpPD
wLoNMgAXRNNLVFpGQwdnV8q3lnLOo5/Vik/GL+ljZmqs9MTS29isEMbWeZtQxqd1
xzx9MW8U26GEpU2uPoJuuG7AdqkFgXkWbgIWVvjfgeM8DC33jV2CmTgtgoMAQP+o
ZB72r7lJYFFX7+tzzJMvuOHfZ2oRSv5pnUsuCwRlxMGYoRFJDjRDAGiQiH5C64no
N1g1SEALePTkJJ6FAz3k99z1nof+2IyqGe3p5MIfTprMWLMKB5QHSZryMtuaOk7P
kdfsEgh2u5GzG44D/bGrHjmAEUQ/KEjgGdUtIB9WIMFcZ76YEnagt8b9b62Nsuni
HpTak3omKEGrzKEcRcQJC4Yql8Q/iaLJQlUE3dMRh02ui4zohlTyN7QQeAcHJurF
9TuIVQPbdMFf+obItZrxB4Ui5EAmIvzJ0Q/U7Xi/+T06Z/ZO5Vxky5lua8IoCe5t
ZbAYNxgst9zNKYlZYCkxOx8Ckl5RHWzFMYnBx9BM3q8JL40FpOV4aSnhriRNY9/I
d2+PZlUNy09U30BvMADRktQR2VwY0qItRDygjh4IdrbzL6xsAao6az5i/M6yko4K
wAXjBZof4GaArPvOk+iqVSacqe36ASQ1qWLkjsVqPcdJ8JxhcX9FxRZ6YlGRPsgO
Gd6uMdzvZsi1+T20kxNsAAlbdC5qWZTzXIXZVJ4sCOYFp7S3Hc5QcAs0nc8kdRHR
Dezosx4eECZ63oCPgg9fZzfwrYK5NwLkjki1azJmSeB61mDSvQRYhxtnM2v1H0X2
tzwXsje5lrtiy6UC4gUQ5kqTOQ8/q4ZLzaUcPQ6LcJTDc7HEDnhhQE9JvTKrkjYF
NZpJkFQVLs0IBCGhHAoU2g3ctenRkXD4PttNM2cp+5dpgE2IBAFX3PuNtdzPEM3c
/5NGk7O9qm8NKuCryEjuUQKNwG7+iErj2LXFE6m+3Nv7GZ3oTm/DUWNiygLzyNZq
TmXVUAwwvm9RmKjeSlZkDTLSG6/BHTjwfO2XdVyx5VC/6EcOxs1RZYWWvtRS/QlO
lYrAfQMLV9NaMN1PXoMNDko2a3iTeuwEm8KS4ldrYMVQyaAnJXD++aesvQGvGFfR
8pp8UiLjM39flC710JLw9E2Qju3iUfzZ25tMr7OHrbraNO+7/hnYiItwHhUvKOBL
DFIqWEg5oPYSR51Dd/bQjSnjHDYikqzXJ/y44rmxwVjcGmnz8DgBJAx+f/+mvAf4
0HVU5KCWc7qShPqaT1SgDinNQFxuBx5ojQqhiiH8PzlhfsZBOjMlCW6ip8sFzCU+
U0FAX006hFmk/p+dIItc0mFLZb5ZZ+WV/hGTVGC1wy08w2xwIcLpv92g1lMDMgWq
ERcsu7TJwhEv6hSZ2UT9I9OrLf/WTVz9kTYUE9kFHrJOOkQbvtqSyFJrOrjTDmIk
pxaIO5cMbknYbow7RTvto940JSj5as/XMlXwM2FUdVEttHFE9dbutZHF3poLrg6O
1v62frYR8lDMxKfkurMUKo33r9LsfdNTNgzImZZ95SLJmPZW4vpxJnGHHf5FhciJ
n1qIrD8SPv04l5KsmIw2JTrnoRMb7HODy5hcAwo6+cvUc3PcVwrcCrzVxrS9UEWa
uypbJDypmRjkTlf1B3DrErmnrVIgKvkkV8xkFBmJBxFXDMxRaoV0zUe9/IYrbiqT
u28VgyK5DZiGL/kQMVdzlSr607WcOooFe8QNyg+4WRe52UtrQAwmCJxgR6s21pGk
uXE4bgJwrNJgbVB9zOaGkRVAzh2sUZv/bOwKrcFz7peshj2PCBMd5kO95r+ZsHEs
E9TBoyB/rGrph5UAx6Q1w1OofLbLtrzGAPmn0Si0ClGGs0E8D3DbskqSop+Gi1id
/4C3uZMrR2I51+V04LibOxvInJXtEvzVjof7B4JODK2TVKzkd9v22JESEl78to05
u8jjuhSMGZSkXCcIC1rFWbkrWpbM58bPJdaUfDJZbo5NllH/IEJGfzWjGoGS5EwU
wspB0QX9lfFiTeUimtmPzr38U475UP0trdoiV+4V+C1pzvjSh0S6wv5X89eQlG5Q
GDlMjCEnP6Kj/pViQ0OrBPwwoO2aaquUcYiYjoRu9U8ABjepRn3cF6LvYOQOIjRx
o2DJx8Fra7xK8B+5cNutHVSHbm1sNm4SVr2Vgv1Z+Sw3QHlQiQYBvmK/TYRm0jv7
PzJ820b5PcZ432yHEx7CKnH9K1z+RboUBhVz/HPSAkRbDhUl1Xq0l2nLxcJ1qo3B
YcS6dIhIGenVXHOvBooHEi4PwCDrcdngFo5urb30HFBqdOnP+et/Nc4B5Jke77iU
`protect end_protected