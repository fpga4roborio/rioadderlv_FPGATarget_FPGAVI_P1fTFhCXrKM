`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
ddtXksX2+yylW5zu6QL2Lhnb2d1sD00763mmSITNX595NcHTEkwn0zB1Dry37fOW
FufOhVzEJp80NC5qZ/+F0Vk7Ik02dIR0elf3clrjeJRK85K4e3Hoo4xn7YbFUIms
l/8VZSb14+JVGURjfswrIyCUotIzlzVYZ6gzoZwDXIi5gQIBf/gI+KxNXPaKV+PQ
Ufys/12rjO6aI/pPlqSm0hCvftmBcnezN2hk1UeXgOIuKZnogjOsf0iJVX2aOOWE
6pD/psybjbnsNB6kH5uFTA5frkzIzkzl5d9+YDm9OyC+k84E83I/7/j+rk4L2dah
QJOvksSIzN867/4Qt8qYTQ==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="MvBXkzurAa5VTw+1JJ70nePUfoQXBvZOku/SMmg4TwQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
oRtzZL4VJ4iwysPsC8SXYCzXS8Fw2gtZTOskLcDV+1B9Nzn1zTyNtlo6lNICRmmK
ZRVu2BmCc2G+fmzynYlNTnSa7C0Cuel6FYpxCBlOuk3OF2tzAmLAuDyOH3Z1Yjzk
a0aHuoCdIRKv7BrZCdALt03JeUmXKPdOmIlkVGFl8yw=
`protect rights_digest_method = "sha256"
`protect end_toolblock="Jn9CQpRhJt4rnzZPRk+dOpzAubz7omckX1MrFd4p81o="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 2992 )
`protect data_block
gD6l00tciPUa6pDNTk/+t0OO0nC/UTtBwLB41d4inuAUA3i/ALrNyoJVcBnAmEQW
ptbcNp5fxEUJjnOxnedyZEuEBxWRieZFQnkRdF269oMWeBCI9CVxHkNwRU5e3e8n
3APDura+qyAaSZEnkLXXgggy81t+MqkUYSRZ+QEkqCIw5QibLw0qlzmqcla2pzcs
GI63R93w0tWdKOfXtRx0+sV9yFBgopOhptf8PwVQG1Aiqow6i1C+1pgodA/PFrAK
mIc5XDexfosw9LLfl7aM2StQ5ggMJcYjtP++jDxVkHmYcEISesVEYOEJA/E99NBt
tuBCqX+T2JxNJmSRi1CVsYhCavcVXWH0TAZxXy83oLvzW853KBOIc9sp46XHXM7c
3tAx2J3onY4AU7nTICQWLAoMeMnve5+O4LCA1sUf5BietngHiC0cfgxZPL0nm7Ln
Bfhb/h9FAAqHLlImRLn2SCwK6f57vXAO7HhDnesbMLP2GyMHuLIplsYDYljTAJJf
m/ExBVomIVBq5C+aXPB+AL81+oLBjbHqWgpIbMLGYm8pkut/GnexIoohGBjsNi5L
X9aFIi65kgOsMhouy+202sBEwgIE4T9QtCqNYFUdmeJiFoC6FoFbjIFZxzu760rA
9FQDRpu2FDQMLSwxCiGb5faxntb5qpHRekryt94GPUeLthxybylPvhE/1xKDAnTq
7tUKrQizdTpqB22/tob2GLAcXO8+Z47MxJc9//yLulLxhju+4ryvQqNAP8S4o9T7
Kt536MNBZXhmHi3/gvGiPRdWF8O5PcmKkC2QqshhwYR2XIZoj0hB3kWG4AnKnU0p
B6qYb2zEYsOBDZH8671O1v/7Cb53yrbyVuAb5uE5FqP90Qud5l5gMP4rBgzkm9mc
60RUb27/Dkw2ri79UGGICnAX1iRznnw4yk/iWkAXfMg9B1KUWHJrVIxHpnsAp0PI
gkxCTVf/pS+fq147rnv1NjYqT0EdtKs8kcV56JDOo/Ta/NIsDtFRvs0tjAg5U4Bx
qHvp86jh+1SQGqFwqAu5CmCs+PXYc+1iu3RPuBVt8/A5jfo9wT+y2imAfWNUXZmi
LpiWd87Edhy15Fo34bgfBt3jB6qMfOvcF9n/0dz3SM2g2uTfOxLLH+jzxYtnQy/K
hJT2NE9B6jpG9gBahSDRgtgpRig1Yjya0aV5cVmUxAj6R9ec56+mH2Z3BvwkSe4q
eQdK60Ve6oOr8O8JJHpo5fNgr36an4q1t28H7obNT1MTymxw4DgaCImQq2M0SQw9
QI71yEfylY2tah/ZyXrXxVvmwfibiTHDz6XDW3Fzi3exOrXUJ00j1tWIVg/MHkRA
3TSKmBPKeONdVUV+E3xqe5iYKhpUhl3D8511GKVO+75qgDfZTekEloxdBho+n55i
RwlLUQUWDrMkNRthTDRqvF2A3ExEh1bZ8sdXhMb9XWbgmhbWFyF/63C0nLfL94HE
6MBY2s1DLf+GV5sgdinl/CKWfZ6LKPInmQbG8+DhMiJxZCIXkXcPdhSBY/dQFq7i
/9qgOrZbQPsiKPkRiB9SM4koG5q30hCRMjVfmI+00phAxj3ESSXi1YWb9CfUscqk
H0wu/UkpcIXhMtTgWc7IrWmafv2vXhQkIsTkoijc9eAwLbtNVq2mU+Hx65y+EEZ+
9uDb1nZre9XnWQlt5hsu/U8VQFA5/YLL5pT2whEEvxmKivkjJMyQOQ47BXEJE/pM
OGFJNVR2alknJ+A+IWHyYnJXKRjjPo/eNLIvVKTPYJIK/SgVi6cO3+YUXw9kkvAA
hG71nvTU2kg2Yv2lIf17KuxS5L8pwc5wMRB7+EDs8bWkSRk5qPXdq18loNL72RUn
61OreDdZsyBSW544HAqAg/kTgFlD38YYrt51Ve3GxUoTiNvqP/9BS5YVtxIw1hwa
o5KphOEqyUp7bpC7JSWIFmN1Lz70U11m1Xs6raIwBsB8j86dDrhQQb5llWAPEZmG
mT29rqXfeUVVFlRA78dJKJlA63+KIMTfDhPaiRNqzSDzYsn/hHW51q6bCYFE18Rz
kPjCyJmBuzy3pVRRcq2eyye6IMStwsAnJPvEycp58xfTnsyyzvl7XP/gbBofVKdt
QF+DZoJs6IGTuiKc6VgN2OCYPSIRe2v/Tz4AljsU3f0oyA2DoxiHYUw/gaNDVTV0
2iEaTnfdBw1nv3jN0nkNZIBnLTkFZnC5r0j9LChl9jNJ6LO1Cp7bKEacSA4qpl20
R9DkKutMuJN4DzVOniMzN0agsKWvnjyGAttyglR/hJVm1+IAbnvX57hJ/s1vBYUD
1DsrS5XqqpS4q6Qs20E9ewn261in4B7tBnTOy2yxf3NBJbDwdZjYAqwg5Vwq6OhJ
hq+zztWbf/xabLfENRYf7gILIwWB5Kw7CUk6Zd0BvjbWM50WK5Aswsnq3ihPQJmw
nnLsKBd6V/U6omp6CUS/R7EHzaV1uIDjx6FEl6N7DGboSUM8U4FvFe+ZSDJ5pSwK
H11PlLbaGEIWZM4oEOmbJOLMwueKVIeczWFscTHatD1+TszQbUAz2LWL/O2NZ2ek
MU526+p0hvDpauMjGGR9YnMmr/1NXK0DUDuq3hSq0LrgCywzV5W10+37eyyrr6y2
Jx5YVBr1duPimM8fUM0kq9SDLcTu0ItaGCNLSUPbUpGiUex8R91YLJ03BXNsL7lo
iI6G/rqbyd4kqG7T8HESI5Vs9ZYbgqMNpq/2mGrLh4SP9c1yXeNIzzYS8pBifar6
mvL0b4Y7vRqmw3nyLSpa68XBl4TSSlvdM1/itHCqCkpgfC05Bm+psaf/Z9/u2Mly
xI3t+UB78CGd0tTT5rmugh9Bab/2luqW2cY6gnU/XTs8WDwKy6PTb8g3hT1T3iYA
lI9a6IsZLpycFRLILy9eJUUXK6V0jvQHlkC7HPHpAkdbUEEnZTVBZWX5rUyK9CRM
znn1TcdGkSSaEPQdOVSLsZhQVGMlMpMb7WkSYAxRuoJUQ5tyFrVDV4e7cUvEbDxb
IQUURITm4JFFHyb/X5kBKUJOuDH95djcDHl5J/0BR9mQAJyH8BEUj32j/81KjncJ
91P8+pc6xyX3SeTyIVYgrTBtQmE41CrZ3MUByr56Ki+YWvjbkhWXlijjSVSfEsuu
U6UUV8m9KeSmFf24emjbx6mYi7utR9dsS0hw5iYy4HtHSKUrvx6T7JjKNJJEOorS
ijrK2UaxpziKjs0Sh5r4Of+vGs9C6cIMBIH26QHOw3m0zv075jTp5lhwfGmN+mYV
FYlnb3SmFeVQQJGmIu3wzP3SAW/q3PFIxiranyXurlIrdnO/G68sFTfezXMCifeF
GX3htzQgX4xx9AtVCPeyuCOEY+Dgp4zdXVao7By1kFFJpplssdiPacTFnpSS4cdG
HRTLAAlpEONkWSfr3hkJPMsUoR8IBhUPPfcjd/RlCWXVcyBuOcxiyBZPxWrvimUz
gQE6JvmEykX/3mY1jVEcbhmd3kRWpnlxAOyMvS0jspMwLYDTvDsCGfQQmmBizktY
IcjrEy4K5BLO7RI9aq1t1Z699HR7gaHAinJQU8oYLEIaPvDhwZEaal3kj063HAtA
sXVeltWGvI6yjbZt+TLKPy3JaBDjyP4QayM6VaC/42qdaSeopHUFoUVsTLwvH6/R
cdfj19n1XziLRI/lMriqMMlEaaEk7MEcM/gwM/FwW1mfkHlPQtYH/Ht6QKwMwYe5
I8YLTTxmiMd9ZUc7rYlNu29/iuYvKmhE43nOfMrzxffTgWsnl9VkaJQ17GloTz1q
KC0fjk27RSmZJIzHz7iXcC16kV/n6takK/agXJAte+UBt44dWcfbaeUNM8qfalJo
p5QCEon26zxK3jWxQlYaoZ7L/0jRCA74VlccBshOIIW2/aw9SATax+Mkcy9ckNOu
qietpqtr9BcnzX7/E5pDnLLmGlmSRsdFCTEJWok8PcCWNu+7moAdZsl22YSWeJA0
RrftZ0UPy05qN4ALVSIx8Q==
`protect end_protected