`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
ddtXksX2+yylW5zu6QL2Lhnb2d1sD00763mmSITNX595NcHTEkwn0zB1Dry37fOW
FufOhVzEJp80NC5qZ/+F0Vk7Ik02dIR0elf3clrjeJRK85K4e3Hoo4xn7YbFUIms
l/8VZSb14+JVGURjfswrIyCUotIzlzVYZ6gzoZwDXIi5gQIBf/gI+KxNXPaKV+PQ
Ufys/12rjO6aI/pPlqSm0hCvftmBcnezN2hk1UeXgOIuKZnogjOsf0iJVX2aOOWE
6pD/psybjbnsNB6kH5uFTA5frkzIzkzl5d9+YDm9OyC+k84E83I/7/j+rk4L2dah
QJOvksSIzN867/4Qt8qYTQ==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="MvBXkzurAa5VTw+1JJ70nePUfoQXBvZOku/SMmg4TwQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
oRtzZL4VJ4iwysPsC8SXYCzXS8Fw2gtZTOskLcDV+1B9Nzn1zTyNtlo6lNICRmmK
ZRVu2BmCc2G+fmzynYlNTnSa7C0Cuel6FYpxCBlOuk3OF2tzAmLAuDyOH3Z1Yjzk
a0aHuoCdIRKv7BrZCdALt03JeUmXKPdOmIlkVGFl8yw=
`protect rights_digest_method = "sha256"
`protect end_toolblock="Jn9CQpRhJt4rnzZPRk+dOpzAubz7omckX1MrFd4p81o="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 13904 )
`protect data_block
gD6l00tciPUa6pDNTk/+t0OO0nC/UTtBwLB41d4inuAUA3i/ALrNyoJVcBnAmEQW
ptbcNp5fxEUJjnOxnedyZEuEBxWRieZFQnkRdF269oNomtS3jDF6BIQ8Rjo+yOPA
kP0pBKcek34xcc7uuMQatffRPVzTdr0j1w77GoVXV2HSQQ7yIntkeMtHyKj2pN6W
KtbD4XH/mgHIAosuS66FV87/8ZSqQ3/N/EHWIvzfEEKK4sNvX+axDiWz2XQpOnEl
HOqkfISqUbUxawL6Eea98KIpAtpxIxC5q3Ee8801Vz13OCBFpCJ8OqGOr+Bf+9J9
SEJNDsK8oyxwIoerOA/wvUahr3xv80H40btsigy8jZsXzZrCF8XrfKHwKfShxjLn
oJVNryD7PGGvVrLCajA/nMuHBide9hLOOP3v+1Al7fwM8R7Tpos8tFE8fL+PK+e5
+A4sasCHAfxBUmo8ikm57FXmKb9rEdPxPPSzUO0a+K3QN9DZ/Reny5z/IX0TsJn5
QoXVq7fNNMp1HTAbm2C1C5AtyVQSzCoXHoMPcmodhnn3M5M/p5A/pj5UnmDPZfj/
4CfisVJK8nBg+RlhrKyipAngqLGgQAVrXsFOJls6QUHHWQvt9YXNsAWWmEYkbQoS
5Kgvu2IjPgif2YOxljfIvBfVd29nfUvs81OuzCmeg+OW1nH1ZWuMaWPfs4zD/ZxA
7ZK46ugfHad9Ky6woGF9Sfh3YE9vfezJqOLKYRj6l5P7rvn/N3he1sovJdOFgLgp
Ju70KdXcx2pRPBtJpIkH9CDla84ryzCqe/KcAgvDswaiMOA3tm3HSG/KvvsT0HRC
prvAqfYCcz51R4EuCGZr34DpswFUTPg2JeD8wNp05cWkRkg4dwUawfrW8XaRpYAy
aDS2FVvhsp+Jx5Efpy/Cc5OJvZgVJIDwg1yMW+FOgAXmuGhArf1OzlZLTH7ZGF8C
x2BeIE78B7wp5X+W1FCgJu2lCp8JbNzjLxr7L72vh6TZX8Bi8TezZsbQKmaCEFlr
JNyNnFCzo0qw7yPKhpCpk9vq2dXn4S3ilSh1KCyAIzHwH/kSNimW/g8uKpjdXfMp
sAe19g6XROxBa33GFjJJ1fcfl3gZDceI2cNWCRnrQ3I2otQGFgPFp1ghPfeh0ipW
eeC0B7aOr0cf9DanMHQa4JEsgOHlKK/2Amwbc9e8wcEgnpFWEQ/6H/pEhNJS1RPe
r8+5xx7B4Fnv72LW7fe36Xnd3goWa41fmA2HJPiNLSlF2nkMKGF0tuzXuRCfglH+
7b4LuCpyLf6JkIQC5u7EOXzCA2UzU5GkI1m+SQizdKf6/HOE02IoQq9GqbI0O6aG
9VsP4bOBOeSXz5C1L44yVBUHSckxcBZf9P466ck+kNQBPpNHY9HylRh8NjZHd6hz
gugsAMMxV1UpthgtUW65XNc/ebcYVHsPq4Q00YlPL+Qa0rDL9dQ6GiYNTXlrVf5E
s+4yZA0tSzMpCXRcqYUGmv/Ca49pSJnEKcFLmkHR8pgSbV1ogEg0zjzOYslcXT8r
SHZ3D0eSHNguSdQ8FPYOZw8/SQNb8AA+scqzeoo/uo3qehxU7DGK8Hy5OARgeqqa
CyUOLUKkcYBfD06cWfU/cdZuu96f5+TeJ6aSKJ8F1LXZKJmZMkAJazHKtzZMteTN
0uk75BA7pc5Y4D8piPEY8Or3BjhKxmcOUGox5rZKY7KtYvKPyWYob85uo0d50zTU
/OYYvjDYlYYGaXaRPFR4q+HFJiBeoMsXKYqzxkO03mIX8hA5tfVq5mehGmHgD+0I
+iMtbKj4p4IOn3exBvX/9PxjG46rlSyk58sHMzPnkoFsjTe1eduCUEW/II2FQCpJ
uVDLfJlQXpjgtos+e8e2y4zof0oUMduJQ4EvLmyoRJdiBlH0liMjQykXAPCB8KRs
B6ZBQSZdhzJ10u0QMRH6osHgPk0AqPRAOx9K3fdBUM6QE3o5du28UICOrO4VYcMM
VrOI2vxg15ym/2wud7fYg6WrXtPDLIx8PXtkcbxs7nJhWMRRhw2nM7Y7adZZbmdo
BswKGAq9LtlL+jC807FnzlA2VDNSNQ4/pDLPRWSkD4snRrotckrttP8ehWj4quDb
vZ9dq/cR376f7jkbSRp9NAhYXNYZ9aAy4dJGvRkcgVELrH/OBT7YLWbJfedVN40p
IOCDPtv7qR7QU6CsVWrKJtaUSmf/WaKgXi9ANUMyfzpU7HFfGlyuBuO90nmq8D7i
izxAoBgmcxJTjdqotq50JBhQmi9egbZQ8c+/MtH9jAfO0yoIJ611Pxh3VhRcx6NI
HRZe2etQbZR2BIqiN0Vzsf17QUPifeslY71VXufkrqi0iPZrueO2nCruYsoCqS7f
a4ttYsAHibKuMAkp0fl7Et65TRom2kOyUow/4Np193Js4F9NxHSIMS5qyb7nJPsw
QIbxXCXvcQ8cqI39NeFPuUHMg2jGbyWqWA9c2USXqt9joqf9alvf1nIXxc3Y/dHZ
PafOG+aNDI3AuKXpMHmCDh8o0brrUF1nPVnfn3qEsmkgmB14WRomrgL2SZQm5UtC
iJ9i0vUG1TeWNk4qJiq4xUqMiYhci6pkjguQehKyyyAk36Z4fNQxJiHDVH2SOmNY
7HQJJkmZZR/DZGmlRxPaGloDh0JYQ0VHMRF/URAEF24IjHAsQI2E2r/M5OKKguAj
c482iztco1YuJ/EfM09gc4ytNoNFIA8oL7f1M6ii4UGc4EiAccmb/nbO2UYyeGCz
DoocdPt8kogqNJ1dxReO0r4ZMmlv24bqWbUsG0jjNNAQa6KyzK7iqW99BzBe/DqJ
25lF3eOp/DGCVsyPnA1PFFKBLz6bFF1YllUklmUPa59nesVtaHX/uVuc7er/10eJ
p8y5aZ6aAaKcii86wrIXXuukibFFe1F2MhZmiQZhy5mbAlWz2YJFa3VM70ok7hva
Ewy57jmys+PGoiQxVkDLRFm/p+62mehu380fVzmrV2ZLVw753klUUdI/W/tCjQzH
JvZJzmToVgngdKZ3ZYYjmMNR+CgV+uG1gZjlyYQmk7yTiCNBEBU9YLFCv6gRlWkZ
RY7sE2jjFSpA2VNA6NKvUuhFrmZhbh/GAM2Q11HORCV7XY2ZfYUWyAVUdTWbt6MF
EIMElaGJQBMKuAlNlydY89d3GhiKYinmT04RI8orkunN+bvv+xT0kbsJ/Xbhlypy
QrsN8ltJxSQiF2XpWUX7sMPUbvTUYmKt2kz4juyvUNxiMY6jA5KVky5ihDDFcyVx
4Gq/oaUHo7HPBEgIr4FbJ/3ZGZZQJaxK6r7/Zgg6cfK5XKAfjyrNib8jSRjcadOs
FICAPkKUGd4O0aaWvSHoumbPKxxC+iH5v1lulkqO8hY/Xrrz7+KsD4Lj7I1tiqRd
IEL2RFGwiZn79GMw5MF4N23vUtu8ZIXtidadhpfQ5gu9NbzzTuULORxzw7QgInFJ
MCTnXrFfw3IxfMHn6Hmt20o1hY6kJmKdP1J1BAPxtgFK1LTe8Dd3k1xhEWa4lGzS
E4z3X/GgjczXkkIEvaeqrTKOblIk9JO9DD1DoLiLrT1YUIY69pWAJLxYJEkrtkX4
6u6bqYWMD7teZtOEvFifTJJiyw/jAjYOSGsjNx2XHcKSQ3DVGx4oYpfX4MUZsnEf
nZCsrJYwxyRxuIAVhwtljmxGKfVFgu7uoGBnfCpmJgnEQkNF4Wn004TNsCCxyz+/
+9WBIojJad1vAafPst5Noj+eZLzUlkyFCKBV+kCnrpaBgaZjq9p950Sp/th3w0xS
v9vUumju3QLZSX2nYdIgK7DPnWdDtfS3h8clBDVE/Akz9wxeSVVaMjTM+as3eSak
VufbHuKGZWcoTpVr2WHTrIII3HyrXyNzQ8iyIKCFXv+Ms0XOTcWkKxJkqQ75qyM0
68z3rWCjZWILZolgoyBi18lClAzguxl1wesf2AJN0kTdReQSDTKXCTO82hVMu/T3
wPMVxyuzSvS7LEfRBU2Ko8oiIVzJFqCHwPV5WTWo5UYAAvgpG+mEWp1FV/fFUXFn
mlKLROrYsnwrGw1ySgajVCTP4jwmXfv5a2Y3vA4j/47dVQTpXtDSD9SyI0XL0IQz
pmNisu9jKvZcudvPj6xyCMyUWVVJSx98Gs4tT47KIDVif6GXN0VKpqfjk49y/HDv
VMgJt9awdKF6EPs3+nahBE2QzOfHyWj0+l+YTSQMV7iwjUiUC9AA6z83PU2sNG+i
KNvfdBu9vkg4GG+HdQyUDJylO1phwyc4OD/U7Hmr5O8ApU1TeyxRXz6qilCgiTmq
6zOYM8LfN2b9ArqSTKynQngKZ7bmmujQOkyB26R4/5QqkYzN/pnh6+KwbA+SJcRs
1LPrD4iIToFNU1bQiR30ygMkSMXUZ0BOvJ2tcBbVZTalSxJ245mXxQDtmlwCLYvJ
oj16vi7HdGyZ1P7ACKIIe9uiwTqQQsfFxpRjNXoem8XJ76QHj/5uMKHd/nERx250
pU6WVnwRC4iJKu0M75yiUlmwKMS6rr1mNPKgyXxOiQ6wudNODxLRZ9CX6/T4YTZo
oCozkh7wLGPLGJmMeFr5541kIpableFSaGOe6Ee/h3LYyGQkTRAozgMywEWHtMAN
CTXEsmho/Znrlis1Ff+RBAX2tzY9ydAN3Vujix0kLlxS7fQINQ8X7v49H0Iu0FVW
QxDSLpkfaxBMXuGWap7/6xxsGdu4fHyv2FSOlDPi5YbLN5YzT0ii5Wp04ujv+Z9c
DBGRuRdzn/9GoY74rCw9McL62pEmqtvZNWlnpCp9YR2eSfp3RlcApiUUtFNcd31j
Y6LCxBVpw8sl34hVSC8mjFSu1/OEeec7503bY36vA2C9vsC1vf5fdEOc2wVjhfah
WcYRnjnmNh3aVSH/tgO8h65lsVXDB3OI68wv9Y8AND1qs2y/jWOaZIlKy8oJMkBG
G/qFjkq/YUzpqf/jQPItiiaxA8MT0SNujrPzszOzTELP28OVVWCNXX7Xx0qQa/mJ
oCrczqZb3VDSO0DZEyFdVtHm7uqPeeV2eMJL69hwVUMSmQX2V9EezjAvkSMGY24A
F4oMxXfG+T5S99vaXKDEOnGK8RL8Psg8jOgg68FKR4db8lK3MWQ+paUqES9JuaiR
pliq/8QWLpttIvRd7At6KUSmm8t+YeskRs7T3l4Y39MA75ibEMFvA3ilKFKEkGfp
hkrE8ZX17yvYvw6qFBxGvQo/le3qe2aGMMbS0Skbd6tnzxUNZQEUCRoIl0kXV2wK
X1b0VOOsEWbKn7IBNrq4kTuOvxaWz0520zKzMOXVooE6ZnqORQuRr3AdGPckteCr
bNXpoPTQlyygo+proeCT1If4WMBvHVxMSWMB6NKOX6v/0MeQJyqBBmxCb2CWS8xE
Sx28gwtszhiWYdRa4qrjVQucYI+KMVDtGshIdQwVawJO2L/jbFKPgN/6aifKTdQN
LgaQZwx/AttkfrONzSoEteAmPbQ9C4Pm/0UNYayWQf30m6idn//DxjFf8FBLM9Kt
UdkzW8nKzNZb6k6AX27ATrFgdmc/1OD2t+KtkQ4Kk5C+aJx49vQ74WWqGBIjSL89
0FXATBfKC+JeTudVuiET0znz/FQLLB+dVC1ZAQHsBR0/9ye5WDhoVOf91v5fJJuF
k0d0IBMH3+CdeR6QR65HZK1fpzEJ8J7KZuZqWCjwPeEl0qnflLhnD978nGsUQ2jy
rnNrUYbpZBeT1ugPDSxyegEC8D+stneIl3FAwOM33faJUiR+mrOm2sZlwgVBwbYL
PXD0+zqQFu88uao0Lx8JFYHTJ24v65eaPIk0Z7TqtwGYbhTfx/5aozYE8OwH5Qt8
aG0KVQ8FFGGMXuz07f+QYUjvRQgpOhcf0aKXH62fhbWO1RvDX83xumrO1eXtopGd
iNcBWle1jf4Zj8nHqCiOdEligfV4F6BPtJMEyaxI2b+C+VJ4h6/uhh41ZPNHFNL0
Tja0IjOzm+f+skmfd4dVn4TJTNIEwKdYhI5MLVKLK3EBOygpYRgTmiH7Innc9lsj
zJA4SDZ3F/SJ6vQCUKVnSFdg+0DNIJbgO0IN5jUWBUC9dUCJGmr5V3QGcyCCYrGs
bG0nTQOm+9wciX9wfMZAmoiZ7/bkb9oRe3ThaF96c8UPlo979p3/j4JUphHMhRI4
8gyGk5IH3gXAM6piH51S3QYbElIRgpyGXN7b9SvowuU1ODlykkm1jK9WP1OHkToo
SaSGI2P1xZRzjIWIG5rtz54XElOEDUQQXg0etFoVoH82lmJ3mhLAnRnvPLuFVj+Z
dcg/T9JB4l3whUeHyn/76iw1tWdg2uiArSLI6++OiPlCQDrB2n/MBinYw9qw6Jci
R/hNrAT5Beb+ULhSpKJjirzf7bAsQa0w28BOVl1doT0vzX4tD4nToXSow2Pnz04S
GykIR0+dcwkpJw5jVGAHnMyFLKfhbfbUbmFeUna1YhrsPeTTnveUsDirQg6XnVEL
QPz/UlJEbx5HIR+oOvg7QS4/wCC8mOPZ9bbyM61y/FA4D5woE0DOK2nx9uwRXyXq
qkOSuWUntrEKAuz1E+trdQATtKPgo+2YaamU64f6qsMhLyTcqMpiDFqXXt2vq2Bq
itUMiJPbG8GUA4FzLhGa81otePi0r5a/oa6aMMHRmW4eDpG/qz55n8nDfub4gulD
Y01qwo2iHm98vO06Tgcf4jbAu+6zHs3hCsBCB8hh6USnR2BPARmGXvlfGSAsgUYA
3rzv7ZLksdIF9vUAfb0vHQ6K7SQpLeWis43NvhigMRruiRHYtnNLyBShxO9DW9eW
M3S+xuCCZutXAFtW2JH1wSAUieKvz7o3kc0iygmHa05dsM9+nCfptLhnjNXX0ahl
YgioFKnneoJTUGZApEMEuPx3Xetu2WoQnyJDdEdFt1wYxAUR7g6I8yU37dx0W6mf
nGsCmG/oJ/qeywtpMjsWohCEN07Kc4w25VUxcchhwLnin3pczwqIU/3WP74XztVm
Q2Peo9gBPxsdapMvKFanKw63Rwxj4z4zZCdnAVv/p6FKlnZPEZVge+9rloNn4wRR
zf1AAD3v8e55diGscPg6JosvHOl0zewckTJJSrFpsW+7dKImiVMk56GrHxSv6XHQ
cqEHgG3zW66khujTtNUa4DL/3or/Yfmo/5F9EUXKbNOEwmvQHgM/LED3O0fkxJak
pCCaLPIIMbQBHVCF0ThqErTD7Q4KPdYEUmaVjwvjoG+e8jAHn2m2uypPvLdVYfmF
LuURusA4T44vePDM7PCsm1MvYwbPdeoOjhxl+3vXPV0XnW+O7Yij/cq7WVt5yZvU
9Mr+Fi2xs/OdTkstl3tjZ/VREDC+LY6fpjfWJyJOTrBJf0TX87SP9+JDDSIIroqe
7jkG6Al/f5dAtrXhpZqsfdDxRf4aOu2dUxMCo/59IFt9Av4sZpLUvP/ASmEr2zwf
jm0zUqIDI/kX6nwxZRxSpScZgZ41P0RCVvY5tWRWbyL7zhyFOQZWHZ2vzUabz8TC
o7PJ5TpKArzRQmb1tvwOB0SCuKUde0JcXrVvN051b/icb2PyciXgRBF/3x02qOZo
ev1Z9iJ1CJhMoBfJ92T8W3NZ2RGUXykt5fML3CL9y3t0hJqDk2A1lNJUT+fvVkiM
X4vHcrG7RHiD0xzyt7d/KVxIlGaY9jCxfqJMdaIQ8v9l2cxXjp5xG5n/STD1g3NO
oPHs688sLiZYRVQwhI+QRJX9IZHZ+w8ARPE+wUQ+kCiaf/1ESAtYXKQaHwrajgXW
j62HMjjt1aTRbBz09gWBkrHSj3AIBayO3Rofx7jcE+BKjugxMhBqan55Ws9tYLN6
MeH0OK6mM6aIskXm7iZQRvVUxQPU2+YDMK3/VCeu+vKjq5MwPdDjzuvkUBbGiJbs
xl8Lcht93lKvljQ1rM9eTNeMn/AXBCyHmDecBDNaO8TyCG1q2xFClRk5TUU6t77D
Q88II8UsXjY+2tVE7u5cgS7zg/0WNWWErc/Kxv3F13z23dh9btFNXqjzk0jr4YZt
t+FJaMIEjIa+VYzga6vKlZV0RSAmHBqnFm8UQQkw1VA0y7E8uh6lZ58znnZtVi1a
+yuVdOB5T2S2+Nf5EgvI8mteO+2trQL6r+skSxztpS7ZjtN+sseMvZq+wNdFIYj6
rXdDHY7KFA+sYBp1kXq2m1GxOeDI653pBCUBY58gXuWrOK165nR0AiaVi5cNAOuo
tHKWKiV+RoFZp159bDHMR3+Xuh1cRjqAKmLWu5ezPhHJdFjZ4sokUZu3kNRmwOQ6
U41maZkbyc6Lir6kMGHYn9iS9D5CZA9FhSIlWSMXUsEQVLsMLDDVnbdnZc5l73Bc
2Nmun8Y7R9qsqUoIoF5SFZ5Is18GTtt+K2PBUDfjSFRfnOPNQDFJcHu1PWXs0uw+
2zrNOOx3CiHMMtqjSDStQZOQdSTptzdPFwjJ/lZ4qGw38eRyMXZwP2LgUBFnhUs9
qXgXqx6EDPzZBGuJmRcWS4av3yvvmSVvK882XMJZV09wNLFr3MUt2d7XneINdz8J
mOwh8bOKbX1PXvSZbTIxlcqzuhfeYmfOBdwWWf4nnA6ptplNpbzvMCjrlUveE4sH
RXiVNwNHHctOozq35lLtEW0lVs/VbwXuJkJIWG4kScwaM5u1Vt/KYnP9iw3W9Xt/
SDa8MZGGa46U43DOQhUVb3+dBJvOM+etypjezYxDJUN/TMTts2ms7dqFOB2muVTA
QrZ43w1lcP7KXybUdGgEAQmhPWNIH3/C9Q4KQmMAIHGYo+ULraNKYamWMc7A3q2M
IY+iiZLaLXZFZqshvGE7rnWfRvHRmibwPS6m5JmpC2QxUXeF+Gm1fGTyN9Yl0XM+
on4FNORGYCsuLtDSdXieHoHkBeu30rns24qMI68tyRoeKhZMZkValEpNorL1eeUh
IU/MjxCcIpWvxQJd3bDQgGOj1wVcbNr8kyTsGy73a6KnYBh/DcleodkMzgSfvGjM
9NKOpMxGeqQrVL6RMLgjfUjB0AU7U0ljTdgkWBR4tH846DSWnQ7Xl19JMLXknOGJ
n1KdOJE8zeBpni4c2ut9DF/pItml3FmvLKWnqr2nHUa1On6tpv8iP2qv6BP8lcVg
CLOfiG6JMcD3Ikq9dLxlX7ixzIzPJ6+m/80aVLTYDIteKTVU1OHTRpoRuK894RmQ
b7mL59zjuGkCVU0utrKmrf60TI3k07So68PWowmt6IpNjGdJZoUTZfHHWIl/b4Nt
sDeXKRHlIp2rFLfTg25jSoJ/gzRCeRAkbRbD99GdqVIkEeHdgKQt/hRb5fd18ZhE
EIp6UN7Ip3hpgnO9tFIOVVUXpPAjPtWMz1hUHwIaxiEMo6Hgc/yDyTlF+hqYSuKQ
4xrHSeQM4pTBOPndo79y8a+SekyN60Mlh0XDIYSaFxSfzXaZ99KND29CAH1x1/mP
C8t/NVZsKwaupJ3Lfv1L44eEw7gIcQ8gQeYCG+VQMp2x+MHoDH3E+hiFn3Kucw6D
oBBoEsnWVffN5LFwUy7eflCpWcFLG9wNdOZ0h60iDYaGFXJcgVpr9ZLIz1BT5J4+
iawHBkQt7kSMRG7wjr4ha2sNuqYU+oG8qHoswwBT7MizFeIDPLU9GoQ/T3/P6Uex
R/vRQQZvw5zT6FpeAjHxub8WEILAptv8hTIB91OJznizM3HYv7xPh2zEMdum144G
9gMVt3SAUaHjIs8xOPgQTbxpWAGxhpO/JDFeg8hAMNDJpsaKty/IfgWOZPT5NxE9
SZl5P8KK8AasE10YU43EmdVeIa1u+DYxcXQI3WbMHr/0SI+c1RqsWkWw9pvMDySY
pKZH7VJjHZTRmbxBd+rN3oq5HOpvWrlpXFruq4q1tqbbbzm3TsMtGa/7jJ3Yi2zs
8hJXayrcW+7/Nc4UUW5L0Z7TpQ4bQSh1vLLOnZa+dijLxlMbqSPfL72KeHBPz27a
RP+aNqHsYE1d32DKOmc30GhT8knmzRvBVD0nhv+VF0NVsAT3p2WYmxtD0y7Z4357
kQFfij8X55SmPR/3vTSTKKhfMDXV8ATyOnV+mpcZWWpxHb43T8729cgdEpYoinZW
fnynPwFdCj4ZCcyPPCSASYvmRUgMfhXQoQL5kes//yD6n28T03jEllf7zvk7U1Y4
0z/uXJ40ZyXEVjgyPGalCnKtxA1QNrNpRZoBTmY6/wHw8YFU48BR42G2wXIsOZM5
uxaLo7Pea/oSMasB6Qv0JOms9/T7PmjHgoTvf0yi4WJSXzBJl4xYpE2APzToupms
WvuqbyxeEeraOXpWDJSh0Gk25sMDdzL9xWvnqtsm3hqX6dRtxuCMbaD38ZvBkTrS
XcktbubLYmlKRs3DvuirGLMtBiWFVHt2Gtqt6d0nszeJ5zIwZ1TT151VTPPlfK3u
6x1IfNDraqLiSZIGaxn3Tf0A/rKTM+Im0XaQU808jftL7siALckUg0ORBjOVe78a
NnUBeg+YQ18UywUsGql+2YZTyfZ5NTDftP74JImbMOQmURZVY0cxB/tODSUekxEQ
3PuHkUfIH6hQbF/UIb9ENOjpTTcvii6hfJqkVfZnCE+cCOjkMpB/2XS2PJTux7Ky
IhVq2sgegXLOR6r0DzL/j1AMk2S4KixA4zFromF+lwxqsaqub08OZa/POaF5qdng
TWyVUcTrdB9vTmUoz8MAsbTES1OchPAvB1V7uhL4VTkF9MQ7L+Im1haP4v8MFIc/
SWqiP7pzUeVHDmjB5C7hWtbxxyj1n2QLCaM5CYXOt4Q8KNsvhkQvJ0ak2wLrAjXT
9I/rlvsrlIbqiJuFrpB9LmGnHm5DnyweQNHOGw17FvoyTObDMi6u5s6Vbqljare+
IdN586nxlnDzNR3xW4taPwRdnRBIOkpMduiV/2SUZ+pKb2fNQbgNmghmRDnae9YR
eE8kO+hXvtUAoybuhpT3f6sbN5WVG556gK4NEBcLP2xlxZgQwhp0kRE9ddoBBoAL
gMJQcKLISjv+MPSt9Tv7w8khht+G/T0h45IienBwfiR6fe+ep2h4b+FDtu1Pj4cp
QbqkTFYJHFjTQcrt/0mF6EYJXIQasE5wkamUYyPings4qxoXKnH0iU0m33aercBW
nslUhrt/4AUphY0lX+8jx7zcBpS/r7InVFfQsOY0//6o1khd3/JtYh9DZMFFB5TF
J0ev6SHPexiE+UGC5q5rwVe8SWdmcEGW7Sz3k7Hhq52JhzXGLWBn7E0BVjmxbiJj
cRpyDbxM3C/3ApeaaS5/QGQEdsLL87ySMgSF43BnWivFHVO4wzPTLwUkE/Ye+Cpm
W/D9hks4tNGGCiVkYLb7LOLi4OUPGCybM2DEN8IkL3X4PRIv5/kC+0YxAUBnAB3a
iCs2TSCz0HrCuruqe8sostLekFkMHmV9+YDUrdlsgfyjyj9fYQweDH025H/2Q/fu
DhHZGYGmjXXLUd5HyR/e3aDJMBbVIGtCH7elYOALyPu322rw3JgWFAqseNOCx17N
ULeY3XhZEBeoE9infxC7XmDA87M4WcrwsZnI7Xqn5N/GuPtwCF/7gt+T+zt96y85
bkJM2M09Znk4c8lgm1jQCIkq6q8WQWzpRREhrmombV+VFAWmA+cMFJs9TjR1eLX0
Sgk4PuDwUSyyvHtM5eeloGkwgYLgNVmxfh/52FpHxuMmZcK9Fno4C/Nkk0dDA5kO
1YrHlPyWv23BjijHy+apBtOrLdnI2HjKPxt3t2MeZByqwIjv2NONXxagxQnXgdqM
rgJVjVrt8xgTHegdlY9fHfrH+q/8HL8kBAyTqPD6mdlUhbbJgqN6CJv1E2960nWT
HtVs9Edw/Z/Wv+gz18DIThi66HSYABJZ9OeGc0EkC5/NhJWf7UgUDV5M942BvvRm
Vz0EZouVBwWcGwVvF1biGHqDj2KWEZvOUPaIOSFPk/ighpfLlApPa2DkLdTorhMR
xuLbYA0VNNAD6e/1eTlOA1BKMTV2P8o75vIbYNOMi/l6/qddCrD5bb+pdLw5ccnv
BvXi0bFyzBOsOmwGqd+mcvi8RNk1EUTKsqDIFdH+1eoAu4h2OoAFTQGgT73RQGwN
p2E9ko/BXtesPwLjgEAMDmoiXIBtjOYUZY8DA1GwulcHsR18to7M+O+gYX+nyOeU
lfPuGt/Hy3ZE6DmLJt4V5VDY22buX95f1b2XYFJIQq1KlEYWg33Bn8Zf4zKgKzQu
KfCq8k6pfd5OPFx06GgPgKKopE5CjtYNBhjHof4BavnNgYD4WmvDUgAVRSBeLiel
ctgS0tCYyJyCoE34TBtvDGCzSKa1rkTel+UsrzNPDd3084PrWYcnf7JIPMpBphTT
puWS8WsbeSKbh5OrtqZgLgIJXcW07MACrG+0OATbRWeS++nQiS/Hr8SV7BczcJiK
rHhMVvVvsyhzqjSASvtyut18NvP5SFzBHKvLPQentliCIH866jzVv6Xk6x0RXBZS
gRBSVUHvGUAK8TDpsfUiNSEo+P1Ku7JmgtnevF4LvZ72Bf2+CbISH6+HPZ2ypPRU
DG6T7xrIhf6xiJvyTzp77IPQp3Se+vx+3EU3lh/3F9+hgvbs67UYQtkH41uI8UY3
7YxgGkHmmWGjaIpBHLDpbmwwxeZovzih8anwb1+3/YgcY3af3g593jo7GEd1iLAO
qZJmcl8aE7n9Q0ysHrc8WLn9IPz5VeXjImeyjBpCTmiZStFxGHXScq0BNT4073+v
IbrG0/cYbUJA2cOXbpQKZl3zdl3s7ihOfqIN9Gn5Fl5O7d8t4G487bJwQHXHEj6p
pWKv219/Fllq0R/1wH/7vytSts1U5oc9F2ZVZPH2EF4v/2k+VzWoDclermJJE4Eo
U5DdQBS/8Xz4o+Ss+BXTfSI77Aj7S2aVPq/vEBDinf1QhAt3FhQ3BBCtrAlNNaa4
ycH0K2fWKs1zTFLMLQDKAm/zkO5jUyB8KCIX4E2r9nmg8eW/Ntwa2hy8TV1T2sXJ
si9wwN2eSwtFlgcBOzxp+FaCkHmQlZHqTqIwePEFwmQQUk8GM9Wk413GjK1BjGqq
+rwZTKRdzVqLyQOo5hE2KrGxFKQnF/42B2+DmhDGcQhn5ZKcW9OCO+Xew8yIsUs8
+dYFqqwOqyO5BDr2sF57GZQRhGVwRgZnynbb/JFlgT6S0x6lFHlYFlT/R//0UAHs
4J71TC68eL8LYjByCDpwWNcAFyt6Ay+1MMUG0xcUvVlVo3hpqYNWgVIKFFtQ1Wyv
UP03xz6e9H/w7kLiTowpOHgyp0Dcbn68fD/Bq0fJ6hudpcqd2VZnyHz5FAlh5NJJ
pSHZJGZ++n+eL46I1uy7e61Kn1SWVVBYlOBiNJLmFwVgGq4MjdAfzvVvCLjQsi1j
RVUPKD8OQ4iRW66VdUh15s2+O9G4zkCz6xhdkFQEWCJBeahyGxfmZ44c8SBj10c8
6GDMl4yPRNiVRF7R2D8rY5Ane+88a21s6IpwED9C4USOiXulCNo4YiMdhnTnlrZV
m19M4TgP3Xwj2U/fWDJzxYqTBl4GNtIPNeFysuKNUPjWhb/Yhrw4GeJEo7Bc8dfT
Rgm60GnXnOCT8VOArWAk9PvIGwjIgzFER7BG1DxN12epcEE1V6qFGPLUKpWyjYRN
UNNSpfVYFNmNLxisMibbqZ4hDZetJhUmuyigKeiZHH8mmJ5KlGXY2IjAtMim+Y8y
RddxFq7gZQoXjPBVDnmekhu7Jg2EmULlL+SUhojHmXQDkCozpm4qCxaXlqOSg4lm
sIofbOaKh4m86ArSKadQL89BeiPeIhvbgzwcnSPDgnLFUHFh/KvlQn8b+bCV+BtE
Jj3iiKMXbldCiM1gv/yCmbSg9L472yWycXQDoV4nX/9wLgJmk1nENBpHy4kzjjd6
AaMh42BeSgGSVME/TEzcR6eUY/Wt0qykzeh4OL56j95Y9Qi0BMZA7cWXGa0blq0P
I3UtqqmBp3U7Cs+S6oEOVUqt+OfJWYlniwPpfR7IQFpJvGTq4jAfS+EtIEf+/HmJ
F6iIHQEiK8pcdIYxdCLCuB6hQgYdC+M8C8abWij8lkFO1tcL+ExhAnpnGuzLTEvj
OMDqzwx+MCxqSN+g6piSW8WXMbYHPTbA4AemszvDrh9sPbDyL8j3YsYRCTlswUKO
TTHA7RSyz0ovj0SI9kOd2D5KgCLoKpe2CGgghfFH5EPZFWuSYRc4JyJmAvyUS4+p
6g8RgF6bvxH4Cl9Xd3CKXoyvNaaOczm+ira2IfOhytXONf4nVmh9x/qlkpVl57ql
8DElRDhYpmkvFf3Z98NNyJVquKaHkB7Qvzhyo6UZU1W5qLa7MQSRvQMF8aT64fxK
pRQxfaLQGDfSvM+hZ8WA0Tvf9U9Bh6FQLpbjyy/VnWUFpJ5FVrr1YIJC0ethUCaQ
P2ck2JX3fqCU/+tvaHlyfP1uUNCSo94+dc+em27QxEZsjmQM1+g8u1AQ6qan9SZ5
REIjH1OYoIiDLhsHtQKhZhr3SOXgQN73Tzs4iATN4UlD6DEYoiVqWRR4Fbtowg1v
w4LLUuFYRzcP1F/8iTmBeAIEgW/bZGC5LdHpqMKX9k3Wz487jMMf04ku24n5sP7u
UTe+k74S/xaRMaFMZKyQkTyK63tU7JV6s859ZIxfBusliQXKoX4iiBlVNLTEGSIy
bHbEWkAy+fuh4h7S+XPeNNqZN1e6ntfYCrerixTyPeuP0ohN0PRuPk1FNeXLFDbY
DagkYsIVFeSfM8h5IRiJ4PJAEjMFfp7bBFVbQwhGjAClXvIAMgQhBfez5VjxsEB1
jj/iQ2lEQlmkoSoLSNW8amdEzaqVWJp1spPR+b+u0WvZrgkmk6xzmvV7inOvNI6S
KxB6iid9fhTIF78BHdjDn4fLuo+M/5jWmBvUPdzHKLUCtf4g/7k1XWuT4v9SsY3Z
QTLZSa8DcpdkHr5yAq8FbO5vTopc/S8lVb6YNYH79eRnFBjHAXpsYo1OTrsT6nSx
a9WBX20+qcO1d+FmND5tdQQQaBV2oYSHComGvTyRF9TUkxxC7qDbXn88FMgPTE+5
pNb/XnQ/DPbltcuQkVCu3lblUpOs0EPZf59gKxvs0xj8NGn2uyxPkkl11PDW9Pvy
YUm+yj0ghUEEclABRRNJ11WkIdmpPTDEAXMDu/HcoYJpY1K+8TsOOIwXtBcBfSel
7fiwP69lMl89v115RKFewpzjQFSugI7IZ3frwQlDaaLqI8ZAdvxMAmJR0OiBlMsI
DMuxKUe1R8dMMd+m2VRCDEaY+ZyqBevqCMpYeWq0d5uzfV+NWRpjoNhaIQC7VSQk
JE4B2m0rewhryqBTnQGF8CoasRq327nExj6ydgxwkjZ/lNDBsoJ1GYOX8FLhWRsP
61BX+aQeoPZwbDP70XTQjgkP/o3AOL1bMx4EVgLVYs2T3MZJZBc19QuN6hwZGsrC
wd7WedqtSavvYX/CKYkAic6GQiqwnbFPV/1WWL55m+/tJbR0vJvHF2PsOJ8eHfJ8
1ZoZ9Z2nq2J2+qr9sgXmkBYsxxP9VUqqZKwUA7Dagk+oXtxB3J9A1e1eIA72NIHO
Loke7Pt6ZAT6qmBaU7VRBhUWOJ/zbbsTkRJD7tO2gIbUmRlpE6vpEsdMBUWb3x3c
OPPeOli6GNv4aqu6C08F97gI9/5DT8sbZJ0yC2Bi4T+sM0S+hqr+m2z+e2m0+7R+
+XlBmLyneTw42wA6ORsntd+iKRy2wcDsLRQSvopa9GGC8ohq6zArkBod41qvRdXe
0sAae4WE4S85vjs6yUET5t3paCskHVRADQPtGG/dWyat2sdQRtW5DTEQ1jPHzlFd
h48uWVek2rzBTwgWkVIlQsuFN7d400P5kcsLfa0F6JSyNcy6muFX1RzFLdTuaNzv
UqwVkU+zfyWt1OlcMFTodh93jtYRKDvrUkazCsG7eZC7Pl9HFLIVHBNzxoU2EFky
MvyD6y7NYE7QJO15IhpruFocH0GHswSzYYMm9MGvmE1ITdwlVyTXCEs2t6chJbk1
c/am6zETeHYudoHUU0HPFW1MRzyipBqm/ikmCI8ogaR8p8S3BsSDW6SDsdoRlHFy
ge0dl7DxAQPa9xm5VkKhmX4837OSY4QDpDHqovla4pcAlvHSgnTzeYQY8bMQcdHP
V5+HX8zlFsa6j1UHpmD2OQ6V89YOS9Oz4Cz+J5abhQnl/14UaMzFAPI6wm7zAQXF
kaF2P49JpWaRTvjpVm6jeqofuuoDyQ9FvvMXYTeauTFWIMX4j68wnp/il6+NygMT
MrRKNRFxvq/U2Cujj+CjmzWZ72S5rFGFKURkcdb7qNBqs8KMxZNnPz18b5iU5GIH
vbsiziNm71sYasv8XBbk6ih/PEu4rktsgRP2EwGPumgvVqO7DNeeszYiA+zZ1IcN
3LGvLeo4PEk63n7VeX1WXsnyMBo7gOpbnfkjfAnfyOoUL5NdPtUSbunOQoCWcrn4
qwmFGt6VyOfwtL7xUgYZrsJ6iwJAFMgwJ8aeqwvdlJHruxrMBAF8/6DIz7iTP+u+
t8lhl3w7OpNMHBV8NgALJrMOLNuiuZNepy+Tt/woAsO63JArYv/wnhIjul3bjXiy
Xs+V/0ddKZEgCD/AxrUkqZLLZEU/koL9Pu7XFfRoYr1Ps0zcWozvsEfkpdSNiHMf
TJUvz3h764kZ0g+vVlyTOKrHXD4itb0tS0KHWCKrvKzaIJ4iTYVBOEIE5sN//uzP
A2Kx87a24t/ei/vbPKI8yARzHieAf9/13Og7PTDreCohGoTqXrUJiB0twn2W0Vhb
4TtBzN9XIbvLwvjEUW4hRuiDkAWu18n4AMDYDLK7pAERbvBUJZUbTWbiHlJxA56C
t/qljK03sJy7ODSsEG3XNuMwq2LnTDNMSkVgC07dGIrN5EnGCjkjYt1nwpaTbbDv
yz/53BNOh/q9gfByalnD8nnrTVELHJjPRds/ZBhrg2TBiz1gXPDgfMcWBZdQlvRL
UkC0tYXXyjsIy5zIKrcfJHx/x15QkfR7UilYj7CyBj15FeRO9ttTa3zU/AmzWNtd
KpiUp36vUGppkN58EZdvaktFcNQ7pPtsQdLwXh7poieH7S09rZMhLyDSCXvkIJSd
FklkIZFGWvVT0g2id1WzZCjtviSrLzVzXFPCBfjtl5v7NGwLMAz4gxJi+of8ZWFy
xFAc8UrbrSIWtSv4d+JcSLlm8tPuXyhIaTPs7Z4eRZvW/qTa9MRjOg2d62j3sJyK
rAsA1dKAmv2n/hTS8213BgwLEeIhZcJ2Yb2Mn6a/s8fX+ML+f7WLPm7VvTIrAFKn
4xDH0uuidd8Q9TFD7KZnJeghogUqK1Q+w2h4Gcwa7q+QuWJmmVa+cbIN4LfgkL34
QrBfkW7//8Nz8C2SA1LWFuoh5eu4xQ2O+Wk74mLqe3CNEx5ZXaBb0MfhDGKpdsm7
160+uN9pzhM4LalN8cDEs344sDLoq5WEYYB9BQJ61GM/nVSPEbsSJ5dLassIo2Cm
Yd/welKeRjl4MCAYL8TFMYc+qaZTTUyO8ypzoqBJ2G+Fo/gV0BXRWiaw8M/Bqj00
dOkpPIcsBoVTbTCuNKYo/1liFRAUEAeCJOa6F8i8Q5SSLHHoFzNiC38kbAuWcYI9
AnlbGbPlNNfGznxJrIwPBlfB/3Cf6FvlVX/1ZK5z3d77QGfExHIAtiL41BaRckA1
RzsMd8yD2es/0nYXJC+j+ZgLHfBiC+gE+DlJwN2iTdpS3bH9zeX05JUE+Ig715je
ycqp9/kX4B6Um0pLSgi7EHv/EL7rghTXz+DdQxySVEIG5e/p2NQuof24I7hYuDYh
z4+Za+rKi7cicJc6Q6IF8lqnlz6FaFWlqYf6cDgvvQYEjsi8YfCSpw+7wt9930Lk
X1eoTUCyLnp34fLMnBsCks55FfqKGvQLRG+fuqjDrADpyVCjzIiFgF94w5oJLpkW
nXfCLEpDG8RfEU+QTZmx//NeQT4LTkfGoigzi43eG0Ppk7Fgw3AsRfn+d3UqtCp5
Pu5iml2xUZGehZM8zWeEWHwHeERELsOMpoHuOUXqIsklXj4qtIl4kxPuTt0RYMrK
xI9bGK1pBpuElZwW+wLpnSYZt/U3Tj+NlCwIx5XC416ZQDCDOe8DCkFywz8rm6IV
L5naG1BfHwHYbED0RcULchAHq9TQqva73rwfJp1cZohvM1jDg/rJ1hz4CN6FAxC8
db0pM8mIT5i4D9HKXTkdMub/hFFOn7T1Ek7ItlIKfYLzzh5OXpSr3e79mtpNDmDG
ohbZJThVO0LZcEN99IEwb5dvObW5CTwrq0Ca+P/LFvM9RE+bx3/5U8J36/y3jk9I
exz1gL4+YgsO30niEk+dJitB6ESDckhHgixoCKJRud/ai+BKNIY1RLIIJVSBNR59
5JY0uHMQ+PaKNT8hst0FyLeNgQnIoNu8udJ+UndiLK5nEnni+WGEn9NbV/3QI6ri
tfaO8/3cjmsMcGLp888C2UiklRMLn3AldKJIzg6xOWVzA56e+uajMmjkArTyT0j5
eS36VL9c5RA0n648n69gt3NrRM7I1PBuBRXW28neXE6J9ZVZfwyugDcQwWx40tSw
c02xmbGQU2oNKfuwZEnvWzvQk6qgvsDr+MLxqgaocEI=
`protect end_protected