`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
ddtXksX2+yylW5zu6QL2Lhnb2d1sD00763mmSITNX595NcHTEkwn0zB1Dry37fOW
FufOhVzEJp80NC5qZ/+F0Vk7Ik02dIR0elf3clrjeJRK85K4e3Hoo4xn7YbFUIms
l/8VZSb14+JVGURjfswrIyCUotIzlzVYZ6gzoZwDXIi5gQIBf/gI+KxNXPaKV+PQ
Ufys/12rjO6aI/pPlqSm0hCvftmBcnezN2hk1UeXgOIuKZnogjOsf0iJVX2aOOWE
6pD/psybjbnsNB6kH5uFTA5frkzIzkzl5d9+YDm9OyC+k84E83I/7/j+rk4L2dah
QJOvksSIzN867/4Qt8qYTQ==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="MvBXkzurAa5VTw+1JJ70nePUfoQXBvZOku/SMmg4TwQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
oRtzZL4VJ4iwysPsC8SXYCzXS8Fw2gtZTOskLcDV+1B9Nzn1zTyNtlo6lNICRmmK
ZRVu2BmCc2G+fmzynYlNTnSa7C0Cuel6FYpxCBlOuk3OF2tzAmLAuDyOH3Z1Yjzk
a0aHuoCdIRKv7BrZCdALt03JeUmXKPdOmIlkVGFl8yw=
`protect rights_digest_method = "sha256"
`protect end_toolblock="Jn9CQpRhJt4rnzZPRk+dOpzAubz7omckX1MrFd4p81o="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 960 )
`protect data_block
gD6l00tciPUa6pDNTk/+t1gcgy1iCdpjTkA/bOvU9JA+cpFEv5u/7dp25hHk7lLT
6tYtR8HgwcLXTcx68BnPlzdPHkVIv0lwXo6yhFVkYlDWBcqD9ubowgKij0UjlXmV
p4anbpVt/gKvAYRDYe8Q5F2CQ8AIsxOuOcJ2vhCPchS4QF3n7+oG0MKU5ZyzxTu6
XCtaTx4goSIs7c8jbVtrPcFgIsEEBe2ffISUgGCMjcEJVazNyzC9sGK8HCEpnYib
WQskulEiwfMACxTmU8vWyHRiVH4pbKZ0DfMf7Yv2TMhuefELTIM72FSc9VgdMBMa
izMbxVCnfUT8ikCG4t1OzLHdrezrlArJEJpklmcSlgFUsbqkt0xmQ+ky50SUZiK7
jzzWfwkHK6Jrdo5/qiPpvRprm8V/lr7rT0/F8VjahALlAssKsWhWCNg+7kixE7PV
BpWDoYzDrSerpLn0SidNGUv3EJx3Rh7tAST4EdUrR8srMBhfXvZ06HWlBcGFHuYh
OkC4EhDCXbvucI8FFSHsyN8WqsdUVz+6yc/99sXPD8ZCzDa3vZWW99CkMkDLGDH1
WJ5UIUMroZ+3x8Op/ol3t/eKtkB0NqJMDk5XK63cVrDBJaGaIbGcvLLrNCS76+/A
cXAJNNXSTQ/tHrO/4Ro2y966JnWqDbrkpqBm/+HY3Hv3AleHJZLpjpcsxuu0H2Vv
GXU+Qf8quqKdQnUEqs0McAyFjrXAm8JK0W5E6ZMOLN5ZwxCriM/am3dxjgz5riR/
pUVLt/lvcXz0DPlsFiht9Roi+cZDJiRPQ5d543dWR8ZYpfnl7JhkbWeKX+KUs3CH
ambWjiE8zVOYvrh9d4I2D3LUHxJk0DNKBcSlEr023lwlr1pXRV70Dc0pZ5o6RHMR
STWOv0Yddur6AQhEZE3yx1ZhH4b6QaVAseupJolAlom53P5uorSmzIAKoSvhNqAS
mdtmJXpEQUKrSDi0j7QAfKdZTlmf/eTdd1AG5kYZ57Z3ITi+uSLk1k/Q5ch1jWtM
nhdenjxhXOaXfCT8iQ4ASCE1FDhiSseVrBQ5TyTYYF8ysjdbXI4heSPFHp/A1RN2
eaL78zkXG2rY7/PAVJ3F1V1yCotv66uTX0HdTRrKhDKLtTtS1Nrwzwz7AEgKJEpi
HqkJpVb3T/o8cjDCRVPHvjc9SgIwyDFojnf4nuTmmyxRf9vjfcbvAawm86bV2O7j
TSj3BEdWhm0DvMN5xbMPlMbFXoLcZKG7Diq8Jj6ZC6IvflfpcKbX/bbtLK/Rh9Xn
`protect end_protected