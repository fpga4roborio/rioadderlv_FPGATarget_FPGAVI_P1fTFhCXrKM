`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
ddtXksX2+yylW5zu6QL2Lhnb2d1sD00763mmSITNX595NcHTEkwn0zB1Dry37fOW
FufOhVzEJp80NC5qZ/+F0Vk7Ik02dIR0elf3clrjeJRK85K4e3Hoo4xn7YbFUIms
l/8VZSb14+JVGURjfswrIyCUotIzlzVYZ6gzoZwDXIi5gQIBf/gI+KxNXPaKV+PQ
Ufys/12rjO6aI/pPlqSm0hCvftmBcnezN2hk1UeXgOIuKZnogjOsf0iJVX2aOOWE
6pD/psybjbnsNB6kH5uFTA5frkzIzkzl5d9+YDm9OyC+k84E83I/7/j+rk4L2dah
QJOvksSIzN867/4Qt8qYTQ==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="MvBXkzurAa5VTw+1JJ70nePUfoQXBvZOku/SMmg4TwQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
oRtzZL4VJ4iwysPsC8SXYCzXS8Fw2gtZTOskLcDV+1B9Nzn1zTyNtlo6lNICRmmK
ZRVu2BmCc2G+fmzynYlNTnSa7C0Cuel6FYpxCBlOuk3OF2tzAmLAuDyOH3Z1Yjzk
a0aHuoCdIRKv7BrZCdALt03JeUmXKPdOmIlkVGFl8yw=
`protect rights_digest_method = "sha256"
`protect end_toolblock="Jn9CQpRhJt4rnzZPRk+dOpzAubz7omckX1MrFd4p81o="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 15808 )
`protect data_block
gD6l00tciPUa6pDNTk/+t1gcgy1iCdpjTkA/bOvU9JA+cpFEv5u/7dp25hHk7lLT
6tYtR8HgwcLXTcx68BnPlzdPHkVIv0lwXo6yhFVkYlDWBcqD9ubowgKij0UjlXmV
p4anbpVt/gKvAYRDYe8Q5F2CQ8AIsxOuOcJ2vhCPchS4QF3n7+oG0MKU5ZyzxTu6
eP/7ob0Oeb3c+kpwe8dUpN4mwchX3h9mU/AvZ3soMbCFLMuV8u+MIwiBpRE53hD1
6q8Xac2L8CWEoWydM/NScH9gjx6Bf5uxZNFPjffyr8gQqsM9qQ2Jclpv4zf5bUdt
bZ90gfFHSxH3DM0sa2AYTjm+ofLopnDqtsUTYaWe9lix9BwXvTT+/qBdqSQOSgF+
RQrWPIq/9jsI3oCAm0XlW2lUsmgq5n8H1GORH5k0bnVm7ubSbBqzgyVegEEJEr//
9MfP90g1PZ8j/CRI87r5o5rXtrar6p+7kz7+JHrbPXOXAxypiU+dsyNnmtMsP7Ao
GDHgOWEhML6OfU42Txnvt/lIqttpHNVas9jgzaiHp+jyjvx3nFhrOxUQmPvDFekC
LIl7UmhG2zNGlzXL3tGUfDQsFfwoNof/ElbhOydyXvTGNgjDrdE5siJJmOppN10R
ZGJp+wdkXkUd1k4AeGiPB753fOlY6Q5GM7fuBGlBigrDyqafGKwOmDw44qPyi3Jj
YwA1/0PdimVTYq8alNSrKEXgxpOZsOvaG0dQnja2fFNvvVWYgThaQ82r4rVbFwVh
yqdMr8Q2gS3L9ysdw1K51UMyMX2j3v9zEoUeCr7TvKE9b+/FN7fBh85u07dTORr0
slr9wsnRUCbKLa+NSgcobEuLL4J1DtGhsv16MR1DVs/a6LU7dooXbPDJaI9A4++2
Pvh0+fN5A2BTn2q8HLVJ4Y4Vig2uJYbUgZriL3wk7IsCXGmPQC65GGbZh3zPf16Z
6XCj2ypGWrzVtb07EzaWFFnkJqyt/QEFr6Fo+LFg0YdhO7vgat6+/Istq/QbE98c
Cdn/09cJZWwQcyqOyxG6JDszxiGheqz5kpG9ctlw7tRnMkXgX70E4gMC57AB77PD
mCObgiyspayv8Fz3r248zhHSOnhGWrhdbWBgXrPl2t6dniS6gFLEDUIn7AT2JvaX
bTC3kKmmMTtudCatGwziEq/qqrlAjYyDdnfSwEEknb76eCzINAxzNRU84kEPL09g
UjaO4CJveLTQrQBjSTh7wMU8EkdBDie++CQsutPxXD7EnG4U/XZfBNU+t3MczEQu
C5Av4NWNK5p2FUI9Ac2RcdLn80Kky4ckMM0NTBjGF/eCFRQ2yCHo1PRuW9Qk2Un1
hSDu5KGaJkKVPjH4lIQlPvcpAi/UlUJwA/jaAyQJlC0jkQTXr3sG/we2zH/HC0Ub
dkqkGWMFsbkyWQ9C42X6N4uAEPyowhVPXca0gYBWLmNt3PQquIQJBR9/mc0+L9H2
CAroYCQMayqmhk81lA1IruvY94wMJL2CsmgTZUYdU0+w01GGaiUGZ1xlzV9MlIVm
PDMiXgEWkvnfpVa24x1BrPFlMDdivPSUkcBh9lM/oByNYmXfGvJxzWJjuPr76skh
7bXQipfcu0LgjiIgBn66H1bPfTp1JCHN7CeyTKwQypa+jrRVJCYqYb08i1XAeVBD
WFhVKTTF1kH54iSgkN7+b8ncUZDPfQICnaNBY3PyQprmpgjf1Xqlb9fyUWEFtYhp
3E1XcPudpRLuYzX9ob/Sn9PzL0NeVA3ry9shTn3XOkelhZgTBU9A4+QE9BLdS6DS
Ddop9vSoUCcRU6lskwecrE5clTsKgu0/qXk681Z1Q4Kl9k4r4dw+axSh3weQqaIh
CEtY4X+uyJv54eOns0pu0Ft3M0fAKvURm1ZZAh20cmK+e5BdFnXDY5EIDgFj4EzQ
EgZOEJkc3Xgm5ldEj1t1jI/qZefovdp/jF5rEN3aQZ6oIkb/sCYJw599R7r/NWJe
nQpVGrga5lpbS4aoCBBz1vquOteMpRtPiaFRcpkpzFnT377HLWhr1Nbhf7Rwec0W
S2UNlO52CI1WUN+Gvrf9482FoHeioQSRWxQeOzMiL1Y92jSBAPhpFHvu5pEooTKG
pqEvQX3AGcqm56G/ckBLqtIGEIkjMWu6tm08AFvhzXQVyG0gc33jY74AmsoyB16Z
eyLeiRR5hWyfcIuUInLnRnC/kZTvIqRCB0cta6WsQRKBLWb7n4R5dE1dq0wU7JRA
zpmT0vh5bSz4i/YhnQGh+isH1OAiP6/ppNAG0WCLaAao3GLqjuAjECWEE8QdWMoW
9Bp8QR+Uq+xEQx5gWkC63/1SsVpRXnznyUGQr3rCZVtPzv2GQHp3UCu2xTpBBwV9
JGlBNvuYATOm4vWIsNZ07DFVz5gSpxoX7F6EsRgCUgGTbcn1lA2tFTFKUeLl6Jx2
dfYG29kgxFciX2XQnUxmo8eonJKYhYhMjEerCcrvAaWr7ePlkZ7/VGNzEOkhJcE9
EpVEnHACzGzjeBeWtVTes32x6iFzdorIR7VjlCjPLcouLujySMAN60ycjtW0jaLl
UNwkfDL5HvoxlADhe7JwhvwNYpZ1Y7HMS1XEnVTT9cqvRczyBaNWrMgOtH11vN6Z
xTzpGZhRp/AgAtWy1FEPzxIVy6LFKN16pP13mNfqGn76zR/vbVNh6rRd5YaPmcbR
3WQ3SxymCFiNDf/i+oKS+MEtlF7CoWioYP5aup6ngw/9d1Zf+YsWJmFSu83oiw9w
oM2YXIp2snRY2bHVxqMm0Wo9qoYRa2unmVva5zdnRKNFectr4IVAptRiR2wXqCa4
VTokdu5i1roD+23mbTWbEm+sRkEMlk0sHdi1j7eYEKcuNPY03WpNGW/xfxYTg9NJ
QxPdIkj4tkRnXH59RJ/EFYflHL0G3kT6Hq4o6FO+QLTibCtlTSSePrmUNp4Hikpw
fTlHjGWSi12bg6tkBgDl6raCPHZuQWJJar8Hs/uUJZ6GNlY1Jnn56i6zoyzLfqoX
TxFfrFBt8/mQFRQB8S5uRSx3Txa55RQe8jVA1UscXGTkIg4aW6qKNMwmSkpYpYqI
t9rjuyP4ULSbs7HDDEiGXLdZegEFHXBTfFtIdBDAlk0TSgxdwQmM/ACuTm0rTTKv
cXwSgsnsWrTCl2IWSKEVjKYYVsAW4GDUDup3N9miz6tmKHJrz76P0q5Q7Yx+AahS
V+caCB7hL/KrFKOF4MkJzMhkByUCMNQftQbbA9HZR+VMFnGEICqKxatCY14kXycR
Yg7bhVe/zQraqR+lBZWVAUp/t4P2vXKDON2zzyh10TByiEVkHorzyjSM1qfIOsUr
V+GIcOdyz5HJ2OvS9wqESAU0DyngvPoIWficKSb1gH2NhUSiuVeO/NE27sSgYtfF
jZoUMoRK7gg54IVslStwAuYhY5OG6Cy/wJOQ8M1iu4u1CIGV8o+o+ZZ9EHukcEyJ
RqHOUqWR58YTjb/2zQdlyo+4QezUzm0OzfTw+rHktesSMt9SS5Tgh+gF/sy7J2uz
wHXJtNcvWX/Qg0b7Z6+9ZgLV3h2CCxOuxWatej5qTpkj0s1uc1e14xBMwBYA/Xro
QB/ek+N2yl0ZudGMdhmyB8/6gh3PDLybW0BjxhBCmGnQf2djnkrlMKczrguT02pf
h9+ereIaq4Vc46bdppbZzFXCZ0J5O2O8mgQiL8PqpctNR2vlLrL1zHTdX9iILXeE
KFTHS3V3pSjeVrOoH5V0zHMyUe8jvLr9rOO0WUNWFCLZpUV4/znvDIdcY+Qpp9hr
ApTT0SLFle9wMbgoYQcuCcEG65SlgqjcyuqjY2+l+I7FdSz8hXx2v6ItblU+TtQP
1R01je4T0IQxWwjQYH99Yz23veKOvuALaGvXVvktgBWltKrlp0n9DZKKl00qMp87
AjKKzgArJnKGJsikUqFzDpyWKUVxdex1D6FbGUdoyOCWIOcWG9PzfBw0BD6d+3xM
De4lyIOtt+9wG4Mu2lLxLzPh/slP7mduU8NJoTE/2V+pQNxH04YXlN9UCYsFI8Vr
j45GQYAnzvIgZFBI/2lwM9kMS1QxgE4uHo+QObB8c1jN+f7aW0/HFT4ZlhgQCRO2
VWdgUooIDQ/z5mRQy8DS3Ivr3ECr6s3G4AFoRcZBrfhxKBn4vE/miVCZJIb6wMzP
T9+yEl8JUD8B2WSI99kz0krgYBUV5CGhY0BUL/ENqaZ+m5P5zXacsHS9tsXmjH6w
RO8NkuJ0n0Wxk/aBVJscMsRMZnEHHO7D97vB2W0xJgvtmlwrwXwgWQzKnCoIw8/o
QWw4XLhAfjhUIQvaU3xMfx9cW+3Q10ru5AZyHqUUm2jb3yXKP4G+SiuhCMIpV+e1
pURwUzFPQuGhbdBrHcpv70PGmx3mDwGo15jhi4D3gOa6fi/UTXeE20gxgaS4W66C
hAUzjaeFG3Jz3wkhWNnOkQgNk5JB7bOWgBRViHwL8+ShFqNQc6BXmDH/bDq5qyl1
yOqtlZSt0IBiklowVejthJ3aCUHpPa46gr+xdM09AUKZOgCJoybtYl4xXp7IS7yW
cD5PPt/RVESd0xSyUE44yvpx+wUN/OWTQfpEPgoXirCYcJ6B4jyruHGPr6fQk2Gc
1n5gWKStqNrGm5vCJadXWhGhSkhvCGAXj+MRBX76bFV7Cwwg4jCx9/ZsHRO0mGkY
6eJCrchJYcfnfWlMmwfjYMYCUiaCNnQtglnxOojecODBjZ5XxLaN33oDfgxw7T+G
qIQ9k94wYYC60jQj9agwAbfer7RY2l5JNt0X7q7IhjSbz5tp9D0FkuwtnH6PIw4I
VOeWi8jSAtVKrA8JFxlMeHalicKl+48gWzbEN95f+9qYDXN3Inn4odFYsQblkpvS
qTlLQyFuYW64a2fH9QtO74dO9tt+j80SiILPOmasrJGiGjHuvKwDL8DF8RQ4P4Nf
S98YMlXOQPtwEsznRV93itmjnj2NB/T3q3FaEl7dDD/lenrDBNuI4Pq2mvS/LE8C
bxHxksxzWBuZ6hOENhRfR271WfIFohAdET21APcVcbxwzonU5XMiO1/BK/0mJ+a5
mCfIoHul0tHcArfzuyPAmAUKZrUpwli6rQ264tr1GE8u62p43STaTxZdt9icuIGO
dqLFdjTMdRoNxxTwTIq2zzMncVEP9MWWIW9K2E9Ziq5Z4HtF9R+eTircQTXgUe27
n2KsJYwFspyPFdDRX0abLHqkp9qT2OH9cLGy0rn7JriAt9aV4If+sJwhmSYWUrKY
BKMK9uQu97zXeEqBGsrKdWwDO7f56Lt2WZJ6E3N6aaFdy7/Uuzm00DQgLT/+oGQH
Vcv3ym23Tthd4OgZ4ZfIvMtXzhQMvEdcTCy30kxcCzGEqb7mlDVcB9T62DJIzNca
Klbl7grIbzpMATU/0YWx5XKoBULqgNVvxdG1DP9CsMShQMDvGKSUnVc1i0KC8/LQ
dDONJ1cbL6uTJnjcPTLN0QUgPiDqEAuQowom2TXCpwq4MWZjIcOGCYxDb2jJat/s
DRPEibFImhafY4aVbVQ5xQJ5+TcaDPZRLnepZYsk4G2w1J86tWKnk4MszIrvZnPF
LAG94/3EGR4pzR0Nh9P0hciZaxytrz+nMYgB+41E+VKxbb9ZxWPp6d9z5Ds0/d4y
ITVIVynRBqxFRk9Nx5oUZiWLOE5hqS69F2QLx6qq2rvv0mMwmq6nTaUIpb+yUkbj
PfczpzLafVfV0IRt26EmZs7oBPFAwcufBR4aIRA7rdyauZ9BwhVwBkmsSK3F2D3B
Lal8kn7UcIxFMm1ZaXQdUe5DPVB27R0uMcgm5/vVLPyZvh4VK7C4VpHSh+sF4X9+
/hl4OOnN743JE4AT6/SjgAo24vJlyF5oPGPZVDlKcrPdtLZ1IPz7chSkhoOA/5vj
zS0KgVCB9L9SCb1x65n1C1m3e8ssn6BcANRLVq1kzsvGfLaSClxfln83gAhzz4U3
Jx2PL0RZBUtFyroC76VrKtnhgKfCXTp2+LmOnJ3x0AwA1bS4wqjc2l56HP3l1eMa
+5LMNK+JqCSc86eHR6//H2VglUY9ohBY5s6i1HqmYfJUmBTd5OpMDWyF45tXini/
jfZVQQrMnkoTtkZfjI1p3cMb+Cl/dwj60VOv32NmHTf2y/WvZh6XBRrziRDY1bEt
sec/jdRRytHghz5xdXGuobBzq95X1wuM/iyYDUgFe/pzzY+zMu4QE7nlGiTyRO1l
PbHvYJNPIqKv5xYYF7/LMdUqNk82WOin+nWrDITV9wbob9520unDHR65UB+0HHPr
9SLqCJIt+0NhG8JikxrQXvNFVEexXoNIyk9CH+ZC7hZe0SoMvBBdf62qAbSOQxvk
G9usg65wlvBUHWanQ+mpTTsfRKgzfXUL/JssDfGUZ4AYZa4p/9vWbO5vftqbi8V2
Bpo5RwQQGqZ7ONJLF9EutDHzhRHvrlaqPCxunX8Y/lLftA0/MZeRd50MLHEEtGGz
S02LG4hvuhxPQ6A81iR/rR78rryeDAnByrBNYChKVGl/KClnkYnBbiUJybSaOvZu
iijB0eFrm2K44XeZwI37vjB/wpTW5XA7UAIeSx5eFheiQO8VJldbmTnz9SFM9ENg
Hfkq4snWz0xiF3jEpkZDc7HEUJqD2cWTWTDEA7Khi23BHf8hja8Lc3md8cqMYmz+
1QPnQMxxQU/lfNrnoO5yttB+pvRgjrRWuvGeVhIKpM7Iy8OgIL+6+wmZ/xHLGVt8
W1yHZ490LKkG+A6nvohVNVqCbD5CFHHuSveVsSqF7kQdVHcHLXKjSQE+uoHh3S1e
xxKrthf8/QtTS+rJ5MJME1+tDBkbCBL9IGbCI8ZiJTyrVJiHAq1qXtc2RLWDQAEC
3ZwxghhnwZ2TwL5kbiKtFOTMhpAlFApTYXdUpO2e8Yuu2wHUm2zmPGeMW1WVOHpV
wG8ikPO/TtAxuwWLQZZFW9HKFn+XGORFa7YLSFBSwmlfi1d5nE5G2IaeeeVHRFV6
+pTnhmL06U6WxRN7p2cTnHPXNl7BbZTJ65xwf5Y2u4B/OrwT7SK2cu2q7HrEc7ez
nVMCbsEun8BlAnKIW71dgj78b37sHeDiXtxIrzuSnOjcn5KPcZKtQvAjMCGsrvVU
CkEcuwUg1RIkeilI7EAenaxBO6E3AxZ7Z3eX+j6i/fmVhF7bvV7lmddnrUXethbT
2TCLdMsOAohUhPVULd3pm1tYuEJbvuhZMGwKyU2nnD+UiuGDyGn1FDoxsEqQZ0NF
KLPWiNG8jI17E7eT1HvRs3Zcb2tqYbluWUfI2Wb8eQNcoHSyWPkYoIS1JTPop4Yj
E8mUH+fQFhPemjaSZiGEQd91ilFQfLujSTu8AIrU8XynbhmoIHrjLgXbiybzqMMD
vZ+KqC6p6RKuCclTHgyZHrra6WIl65JsBJz4/G0brFEU/FmGe+FXErnpIgrs1Wsw
2yGrg41yKCPrhNoitHKDsRXJUcusLwQmyZmkCYRCpK+5K0w37b0Od/Lce6dXgtCC
jf6ncnFydqqhpUP0l+JS+FhMe6qJ8yKCFqL4/hEz6tQWB+JMlhHAV7WJeAPklsjy
LBjEjOPzw/ZXmwI0M/JLbA1r0lLSoW2CjddYp/N620k+4ktlYpV7WeeEkqHcsaF6
a2/WjQPcfWlFyud5mDN0Qn67dHYmkCB5PpB3fxFZM6d+Cf5AgaZmu7HDmah8LuyH
AXT4A56MwDoWHhpY4CxjRxzW3g9AOxh1s43zzGyj7j1DcSzImVr8IZ/ldIhAmrh3
voaR3dJYOWiyr9hVmVM5NK7LNigbfNIDuataupRjUSl+zf/Zoc4lroVdcdvyPDYJ
V+Pu3kAXAZl3Q0RhVndHjOlTi+6b6T5kUnOjMl3V31GYGTF/xa8hW4blltYtWlHX
YF8fZmH5N1qRZaP8i4SxlozS+3ZrT1df87MuJUmbVrO9fAIrUAXC29F8M8H4s1P3
GFgWae7OGJNE+HGsGC3SqQzgF6zzCP2PsS5nrh8dfeHD5pdpgLvBL5H/nADUCmEn
Rfg5dT72obz0QskQfP0pBgFipO8W4GAwCq5LiGJDXnWPuSR2fXKTXNrUgnvfbocA
pA7lg1kn+zupH//F83J0g1nKu6KQaAYDTjshS1lo8Yw9fOd7sLNfyQXeUwtJUR85
MDc6uvZV0Br2tFpY6UGD0Qpau6sueRP2mW4DmdA57kzdKyuXmdUFI3N0Rudw/oTE
GeOV/O+6nmsYzRpdUSYDEvgRHBRquwUGcyIjXRb4vurPJ1IO9xnS1cNXJyoR7xbI
GU7IsPjR3Y8Yog4POH0hyfTwirrl7k3f8Qu1W89fs4nV/ZXaqG9roYZJg2Poy5B/
8LMDjL+e1PMgMqAcsglPXzN0vPBIGRcVm2N0fBt7tQF2pWLoAFiezPoveNeDL783
EAPAKxTiYk4Hm/vT9HCFDYs9ruCzg7clwUu/dz6y0dL3VOPoC2LI8hrNEbKbOuSw
i/1yK8cVFp0SgSdxFm+QYuxJLyHprfUK1iuINYItm8oQ8dEDsVxP9+emFMY5t3Te
5+XmY7c8nKiY3yMN3tmFnV1I36IlFAaPLyZhng9EfpxZSTnC9cseAXRTkXo14yBT
pHk76v9LsFMzKBOrYCX8UcHiiA+RLCauj0jaFaMt5OvM0Ho7+Q1PVRK93cEkRSgN
Tm+rLvi2+Kk1AiOQwfcQrcnTIcIc/mwOi63WScinuAPuGOzskVE82Ks+q7bPGOCc
2EkUhrB1d6vBPYD+mysRgUin1aC+7q78S3/+uofo6y85l1VQgqzqTZHCS1fbzMj8
nqd0Lwuq0RA/UhntHzVwgoQBchNazBSEwlE9VlyW86QqVOYB0G0vIZQlbzqRVB7y
gj4q52uWD8AHV1vbTZfPFlLTOER+UeDLVU0CcACCHfP8uYUPR3ube79CPHsoS37W
Gh+AyZVaqhC+3P9q1r2p9uEaeJCL49SB3X+bWKFtAJVjKqfA+Z8ifVmmNEGfk6fu
4UOF80rfmIIRFAmO+QDkDsATav4d9WqM+SCKPnYgziK6NS5I1ehovAEKzeQo7cgo
XBpJq9PI4t0G6YdIZwizZBT/5nR9Y/4psr6D/U7Eek0OrkVLTz9OlAvum3zRiwLo
WbcLuk6xvE+yIIkYc+4sgOjuJNAVl4fVR3aof94i9FyYGfZd/mWl+Mi96oXtF3bo
6uTO/0WuYM+iLKAWLC2LsbW8n8798cNuU9h8LHnfxY6m9PojywMQB/TaI1HBQQjO
sG6RlDNn4or/sN2ZRSx+cstue0r7DiMfqde89g6aNsW/ED+HSiHF/TyhyWYSE7K8
Aw/J+EPWFOythrrznXQHKFjzOgtmLi2AQnvfWeBYJ1KoXvNROOXj07Z41hR3zf08
b69Y8r+R9EEErcIP+zMA+ghWKWV/5Ua1VsdtUESa+sbIPuE+IzyrY3MfPUE4/H18
/o/CxzOZ0obS+IyhGAk8qWHPgvfayJPxRUMMnrMXTcAKXLMK19aLLa0OjCh/jm7b
zxjK1bHA/4pb6JGGzFoT2H9/5Y24lw2AQJjiOgsyjO4lXP8CjUO+HsyWSp7hrN18
JEs+a9LyJz5/TSignV6CAyyMFYvV21LLkweBTD6zA8lkG4nukb3U709hSzIk8tkX
xTYT8LFv3DfYURS6x7dzzHEKoimp2Dpg6SnOlwFVupPEcaaV/DdPI0Mg5U27Lltx
kFEJRHGQz05p6XaeMaVklRnVDCVUAauuG186S7Al28fCc3XWzKTKGqXyjm2yTvni
OSxREGIHpAKIGBRw6cWftXPAWOwQ7YgL4ouxVLl5wfNTTkGST3rLIM5EopBnGaQ/
bhFqOJZLMEyv8ZYzrRPSwiOXvOyqXr0do1e4zCG644TjiPHq287YPio7v6/9MEkv
pucjPTmx/1JMXUCiyL2WZXRlyqf3TRutDBZKvmuWqZtAaW8564uORNRilknE5glP
qCF0eP4OYgke0Qt8aCcyDXqaaECdGTpNJihuS0IYpccRDQFjJ188+LrWaKBp5Md0
ZR0gnQnWLt+UmVEjjifBU9mvVvUOYUkWNjUNBgS0vyIpt92KWDYpIbaEgUimu0PX
/B8V05ZbKa3YjkR9StexpSpRVuKPLzWplw+rqRAhvHi7O68frO9rDCO4tmUr5gpI
AsfPl0fE8D/8Oafr0pfR2mz916AbEM1UmGA9xU3XU7I6D0t15Ea4tDXaNTYcSviG
qkjqd8YtgEc2kJx2WHuyDxGGytemtiG4VzOxLmwTxCmoJrtrAdaBLTxIJy2evcPW
xdk1RJPhoia/mFscAjF1nN5409DOjCnjPBaJFWf49snLs5T3iEN5CY7A1OA8GA6K
4mo+FkJw0A1ih1io6prSyGbRO6rGW8dGEmEcjY+6Qlv9LjvI3LvEUCsiVGJccoaW
SA08IgPaBF5RzgG7zG460yeqQPElTZg9twRtoBBqsjlRyXWG0K0a7lyt6Bo8WSVB
648f0fWGtcKPGxGQX8fWZ3oEGnda+eoMhV7leJW7WnQZXGYwfCmzfoTlUoEP+J3j
nlOgqC+vlGy10LSLu9rlGirh+2ZC6lYVPaoQMv+pb4+h+h5cht8lnv2BGlhBc8UK
jbsb9BPnC4XEcLlyuoforKzHEmGW4E5IRZxY4oy9nPqPMqszCb1UTvs1JSLe47Iv
RGzDuZ5LbXN373+Etq2ppK5prdUZuTGfRmoQpv/xdHssV210wf5z4nWEkRoEmZMf
cPgR+M7GyIvd5YS6elkrKFhpq4V8o47J5Ez81wBVR1Ezhy0ZYPlrESCb43IlsC5g
T0CG5zvkae8S1pysUZ+cytG5juf+G2v/NDZuFuMbAy7OVUfk3qgNW1DlV26lDZIS
k65v/fphbaXohUTVICT1gX2TQ+njFQ2wa6hmVglr4yb1Bjscfezfuff8fPsu3W3J
7dG1mhf9mDV7brDFl8hPgVvG+AysyYN0XED0diwXsXmE+ivpOO5Xju27o+Wo0TUq
ITdpYBGod+SOD/lvfzO/rHEu8QuwVisiCa97VEo1ld5ngzRC75Jrc9riQEKIuhzi
Yj/feOOL6+E/ISJMK7CA91hCEkiz0vEv+A/lh3E4jnePCQiRUL8wD9RbY4+k0oxQ
oEc9z/99DzhKD9p9vRs0QdHRoz1PNterE7O6nH/fKL5ZIuMWpHb6mhWHIo/VYpHo
WuDsUN8Ro90nvRrXINb9UYX8I74zE7c6NHnfHlDGRzlOgkxTPYMJRpz15l0mW6m5
HITYeI+HT6rYjV47MUA1Jq8n7+G8xQvjfsxq6Rjxz6eg4KpU+zxd5wSZI9mJ6nlW
zflEODyDTmjxcSflVPJS38pkRRXAtnlWa6ljvqqny5uIxrMGcj7irYkyhsnihxWr
db2N3WG6RBHFlrWAlH90qdFZojeNGooZRpk4+EBWi3fGz0am6zAJjhvX7/81GgcU
0cD09lC1z3Caj0S0c53Vl69XfR92rQ4Y2MScD9vL2bf0FEs6zoxiPqubkmZ7tAoy
6NNZmVDiM7NrpN0I/ymLt368RnsSs5mIJRGGtLi9FIMv5E5FfOA1kEXVgvMTXWcV
DpkYNX9jyIOrq2S30cDTmCb44pUV0RqkYWV25cqywGNP67cHECWE2cs3BuE1mCdM
rnNIgPGLn8FfWuSIdJY3WPnWt8tyyx/kJMyB3dSk5zwmdDk6tEQpfsYMmHluwQMz
3rCiKVUEYoSDlZ/LMtS5nlJ4xxP1V7nN33GUjq2a4tGmqfEHtBlh2sOBMCRBOBJx
jYlqnx41m5Ll4PMjq08+LtSEWI3FXbcafmbeeVC2HYBjnKJM7d6Ssd3odmUBgBqJ
0e1S30oPlpnnIN+79rSmlVuKlyorupmzB5VxBes7CP0COUZ5JB5KUITMQuHRRkFe
N6QPbAUc6eRfRYJ5D86Am9256GCFlbCzqW91Ub1w+UecsOjapWw3p6pteMYqeaxD
/cyI04sEFzq/PkRLcY8b6QkJmCGvqvYs1vUaOJhu2gjsNfjrE5QqLKSrH3WHASAf
gX1naNw7LI7FYUE30ZxGzxE00ycYWHOra0QAmwJBxxST3t+Nob6zsQg6ZCBnrP35
mPC6vnDJvAbwfnHs5DVioch4djvTj4jt+dg1Pvex+2uM61Hqh3Yoh0VMq8z5knnT
ytlMwPsLd02gPHsKvXnsjPTBXyLxV1itK/LmNfwGKLUckT9sfvMEN8onVAUe603m
ZG4H5i0y6/mSSWXGHuF/tIYFV8Ohmr+wEFubyXobBdgwRfZaBEasjdYKIFtthT1e
ItglRCExms3LoOZzbh1b/z4QzwXVCQTyKMIGfJAPPhhLV4ed8lwSnALyIacbQXeC
7TWLgiShRuo62MFvf00xd0XbBDmD8uObf2hhD09nt26Hq6/VtkDxbwhZ6whZccto
9qg25ewv/CvJaIjwZTNGK+Ok+V0XFka1JZZuDmjj6jiwJJTwH6d+e3+/m/ZMnPME
/xrs+i7BaWmKkDJwNiwX5AdXm/c2lVEZOMh2/Hrwa5W7p0XBSKGCzhooP4aoXGp/
PTPyNzi8N43PW/8F4qD442Gz2N1TQ/zq++++Kzs3KdYaw8rfYbKMZ+/YMkMHRLBJ
qqLHyO2lMGzF2yJ9cG2CWdqRbL7rujJ8vn1QFqYnYJwUwS3pID0ttbp1B528LvC+
e2IezlOtMg0CUcGLWyPQH2Pye3LxiDbkukF4jG23ECVmdh108Qe4Rz4qSLnAHrH/
Gs11Cjmm36xoM7x0wuBwrYYndFUQTNb4jXTPBni9zi7EpmAizODhxKgrwuEEUIAG
+IcvDoxkxdXjC1E9h4uKfa2Ma4SZpu1Fj9U6CN2TS40YGxlBvsharvzfE+ci5Sud
uga9dQ+rUey1uZv9cyADzTRoAmdsdilT0g1jyzbt1vvSsxdfVgc9+7pIwmHi72bF
fxqsVkIgmfMN0+QKVgRzv/p5SrJrP6YRdgUNO98XHrLrlh7Q/7xoj/zzd2dY7oUz
vwiTt2UVYyCEnXyo/DkYDUp8cOPxarvgaAH0xL/00PmrXF2r1wFe+RBRaZtSReH/
jtmxWvpAYrOlY5GQYJE8dyjC+W1KUL/uTnfRlZFuTZM8UhbqQ6mBjy3n80PFMTo8
8FIP3ZXbdSOhI0Sf44qEey7B2uBfLpOYDkoFUh5vrQPr4XFzapTHZpNttjJ/TakR
036aXbcAxdkYstiN5cl8XiG4dXflvY4zZJmDVPXvnDETrZwRfOJLzrpHReBIlzeV
mf5Xk+SnIAOIuf+8Y4tO+pAySsj8XPEnRDgKvFU66DGY/KNEgOvfVm47RFuGT5cB
S9teSrYbXvHrgRNJggK7IzMWOqQX8TH1mEckfrb17qzeZcVIduH1ABB5m3na06ZC
A7WM1pS8oZrs1lUWX5dS9iuUvsndc85r+ynMaH6guhe0SOqQ+3VHrE1yomPSeBxf
lqfrDxBrUVX61NbZt/QGtWANPbVMqgrMcgsHu05MWtHO2Zywoz2m3sYKXoUXF8hF
6HT2PdZWg1Pd6F6DCi+y/pWcorPURqepDZdZXslQPxRya0nSsApQZ0wI97/jRl+c
btafPf978WR4arxnk10XWfAfBi6R4JOrECljQgDfoYB3Q9t3oigq3bv7hSWzokFJ
dAmumP/J5QKvXGy8rHMNPtPoyuBtnCFBnTeAHsGz4/Glcy3bwx6dhXXcrP8nAUlq
vyGS9oPRTQizD1mYPkziKJLYjtC9tsZM0Vl8OyFdYKFHUiyy/C6Sc9oeF+Mu58x2
y7HKl4KQ+pw4OwXZvBAxRIb2rWke0SZoSp63o1jLkFsHsybacyWBl1a9zHlx2EiM
9A/dEKFNmLqm/oINgxSAcfq73lCjFm9q/R+0lsXrwYmiW/oCWSwaWLedQ5wwB9wM
KzTc84HEtHHAgktC79kMKeWZPiX9F12d46b31EZJUn6+QvBJuJB3sTwVlf88ogj9
egn/0dQXiBLy8BsNsbQ/F7cZUpV9vJIaSm7eEH58B06wQgvrGtKcvsBETM2PgCO3
YUPR60NMq0P6dK7Ps3//4iMPZihdXNudqMwa8/ZnX4tYLh2fJG+GqNzNZ552/Vaw
Add8rE4Z8IKCRvAmAIEvGBhqxJnN1+Nj/Z0y+w+PsF7BlXnuksAhxmCHhkO4JyG0
xqzVrG4X6neMqfBVmNIxLVtB8nnvTt6tyNAIOzmBO1H++c+Lb4P/m5AWPypE1xT0
RzN4Lrkc4R1o8o6ch2gWR1AyI1x+ZdnEmJSW7NCle0v6GPCDvgU6F/8liQ8tYQfS
HHbyMgy1QqGyZ+mGrhO+mjvYJUbsAOso+EmJ4UHAXs13587yRMBhwtLF/iMhb3qj
pegXpzKkEBnzZHo9BQvhBQKofxU/hLSjbAImH/Y6xViYcWCMxVSz0HMnY+FBlMKa
g1cqnV95+K0aI79s23esWJALD07TRcJ5FGVyCpdFoOvqodWeB5ZIGdO2pl1xODEg
52n93XqEL88UnTmJBNweeX/hCOfkxDgZKto/rzVo0sK6CjgnccYxbGZlof5t+uGt
Kugo0yxEY08vxqoveNn4LvyI88uSKSlE2ygmRxjPvzt/tftuG9s1zneJIYSWPzS2
6FRqoMq1HgNO/QW5AgKHMI5iyXfrZyxQy0flGYlSeW4CVGKw9+lSGiMZETTGQnth
ityxbVxlEh7STRTiPeN3NsqXxC2ggM7YGj9lVEc0lIaW59AAweJBqAV8KEUyZ0i1
njgVmqajJPi2Zrpo+lzKedHMJha0BYDyigtGm5zWvRD6GG1oPoL4+3ldVcMfF8g5
0RNcYE0iC5mBHZa9PgYDNMdEFF2djtz4FkGJn1tse+sgYbaQp84iOWoB5c8lJr7H
10CQnq9i8bjpOG8YPZ/LxO3GFLk3adn8RzqaFk5FrfGwqKz9dSFiXL0vcxYvty0Q
H8qseeKCwnGek7bIa/sVmgGqnPRf7FWK+d4vW8JHLMOfrTpoEINftnbstiZAnfXJ
XM0QTVdJTs1zN3h7LKitG0USSwptALnZQl7im0we87/tKYK/TWJMeOX1SaD0gmmz
iEklVGy7PwZALL1ySZjUImN0dKYyU7kv2NSUhTzG3aGReE9dRKVgWY0gmj4RmeiD
oAaHhBC9DDIej9/ml6NbTKcfojwuGIbD2Wt95T0joj4mHO2rDGEUbRXbE2b7gZN3
VAdUQhet4cn686t+8JfraKUu5G6EVkV9aHiTTlUHzTfwbX9nZOoAWGFIorw4/OJB
3mnKMUE2W/+2H32PorPW2RmVbE770jZYPrXmPthB1wkhdPNa2l/yDe7365CwM3gH
NQIPbxWYAM6StOudd553FUNvFinPtZ06K/6CJ9Qj5KM2qUhPBqK8RP//pfPZla3/
Wi69EKdKc2ZTxtJRcDY2Qjy0SMyaUebufOqhPmji/yi4U1gI4u4dB6V3grZ9Uhnb
iVM82+UI/2wyIRiWFapwQTOtKp0Cm0sikSVQGCfbUJLXqK9vsKpTT72laoiVBkhq
GuOSbnYrqIUbP91CZ23ZhGpk8UQeiKZBIWMGdBye65P0NrlJ70wfTEu7/tl2zgq6
qW+Z3dewoRlx1LT/kyGeHDi+GqjsII0YTxKvFT5wgCwkS0X669M5PzSsRNxujqln
2/PlLEZqxLFTysOCUgZ/x8qUDCBHceYwS5dOUkaGPMHwCzeGGVd0zJJF3ZkbvsJk
4ErC5W26GbQEokbLUQyJ8vA/Kzd6y/bZb0P5KNRf587Z/A3b/xWyTzY4B1qYsSw4
YlLZD5Hbivz8X521YVDaJF5m/eUPRMe5G0MiKESaWCQPqvVvFmxUCyCC5zxWPJ6N
FTYPYqyX+Bj2IyBpwf3nn8eh5v1NEjkWfpwqfg6N1f0eQiN6PecjMb8MbmraozmP
GSBB8F3Gxib8rBAVyPn7vywzPWPDqcohGrj5Pj9lOYWwu8qyys7AASwNPyoPKybQ
tKj+eV0Jye/zrmGUbBJknNd6udvVRW25CFZNNIznRpbxbLYAx6Dttwmpzc9ixoBK
3lsTnvf8dYypyevUsMxrGNW/uprFfmQRjd5kJcrr2SykG4vvyttRHJ+HjHy2iZnM
6JEdWYcBGtpYCJrZv+0OCqZW1P6HlqYJClV0k1H0zd014PCk9acstuixRslE0NuV
7JZP7mXKTGPvI7GGv54av0UXkFClw/cyde1vS+eq8SI48ckIb+FuwjR6I4D2W4mJ
dWG4B8weNijOxsEc2EEOjjFTZqxnk7txLoygdFt6Tfc+i2PjP5/f9FyXz6IBqex/
pYK1Cg4FEk7DiCkHnu36HzgE1Cq7Y5ygxXnGG899fPulIwlAkoT3YQqJMlqgHy5L
enLtixqeBPUJiKw/DIDL7YfkI1fhjz9NiwQxMqaXoMIit+fKmF2IvkQRSPMcbIJY
oAX9UfPpa5JgG9D3grTWYpq8Gg3OENIIGtYAYlHnoetPIsAbYr90gfgDSC2DEnDl
fn95LKkuGmWl50f6L4TAxrgoJGHx+Nm8u1zFVJ5In1lLIps44yA0W9kH+iIksx/D
q44U+Yqwi6VSy/peqAT4ItLCAXOpQ/E7XBLu0Qc/zaH7ta8EF3UzKi2oGhEaa/3C
MaeGSFSHi0x4/MyB2ZSiu1hGTUUUi0p+4TuoVYVSZDwimtpz02u3eprj/4r7XBGU
/PAZOIYbj3mShOgocGQlyxcJPFRqg+Ff5uJVQKqr+931QuUNxzMm65BICKci3BnJ
eeaUmr5FfS1Ozjoc9slYkWuT4Xln7O8kTeHislEjwV7h3eVXP2x32CY0/+Imy24Q
EDG83CHFOAbaw+/QW+Mgftf4EGyjFVxZ8PVqyn/APrXwGYK3hs5Sqk89LvAYXNGl
Od0xKUDUpAupWT7DE9lawYy+gXAoNtmoumy54Kj5rd6T6U4mAIl2VclQ43h5Dq8b
VDXC8FuEeyZ9DYjO2rRS5Mobq2Vb/sB/nvZyFbH1eXG9gLNg/W5e6Vgx6MNY9ScA
7gPH/4qDrlqPqj3jCeX9KlhN1Ag85wvnXSVmknfl/Plq7kEMEqRlxfYS8/8EAMY3
KQZAld7iTY13n4bJjq3LiReOUv2jDPtEYgGqLLX6xERIFV/RIJGHgII89dTeuXVs
NcHnoRpovMXruRdj9qAYCW2unkGc9v/rVdGxDdgYP60UmNwIOUAUyd1OLkOpYIf0
yD+0dWLjufQ1QlFslV3h+zWHgQgiBCI48XAF1vE0lTKNNTvW/e9R/52HKlubSq5Y
ryz5L6nqRb1La5naCcLiBUvkIv0HtCyOjpbFZzwZ6/TRBu+fNnH5MUvbmOKW68dO
jz19IVYxNiFTWNZhErBmGtaynfRG6xvNaL92r8+j0Dk/kq1jwEsmvvkLOUU1FlX3
EimCubX2n+8tCoqbJPbnl9OEB/zECNah/nR4hF7DxswwyV0SMpbjB7s3YbvUGj+H
vJAiDvwfIiMh7ql2sMT0b+DmsTVsyGj4YWPTg+9UuvUxCMFrp7CnOyuio2Oke+xa
OBTS4niV0Mgj8iyOWhupJEqnzGvIx3LUgEwt8jVokFbHIjWYyl37YXh5KSO0/+zp
JSV4ndgCa6XNYjJCJwREyZEoqD9FIc9que+85aSj7WNbYhyRsSapkYDnpI3L7SFx
/jePxZ8j5dJo0pYATP1lnxaIJ323W3h6ABMkbzRj3bLyIS9kk52GzZ6dXfO2FyBN
B+qEGBc5SOvOw6FnkZa6Kf0qX7g6KtGrXPninZkyEWj2IGeQpTcqRKJ3W+L0zVpn
ZKslcqC9hHtmg4Y9EiHSjGkrplIqJtIK2unTM6SjULR+EREqxBbAz8G0buvRqMJI
CwHotYNwxAf5dytMe3waDqHEFfhk5wnbJhjJ1qi3RURe9ZKu7SGklO3HefGr9x1k
oYpU83Nh8+t6JnFdmzVCs1SchL4votZMBDqWZPAbRxP8CL23zdRICTBO69pmM4D1
TN4SYf0yCkmCaXRXJk3Yoh8VhCbdAudWYVbzj8ySQuCPfNYBqiF01kIM8JD9Txhi
hE9dvNQMD35/WqpqdqjLMBI6S6jx+2oEaXeYDnow1Cvhcw3XlYoMOfTN5l4XsFXp
rtLJIPUIvylXX8JXnepocPj+UHGaKhHp3fEUWv+Hw1BbrJxIUKqtWs/XkfslZFYx
kNHyqTFgsDd9N5pRhP2lMVOefv5wxAXd0wJROxgOsi0A3BIJpEv5ZioHxJblQPZ3
RZbin6aUZZg9OH9G9joMYymrJbumovN9PxDLOfntYKIkFbIuy0/AzgYBh7hACvze
g7IeMk7g9ppjkFxZL35WSetzyyRxveglX27p0vWxUXvQqP1bNMF+XNoHyZnXkc6C
364WTaH1jhTQdOBCWY/Y+4t4c+BwO4/L/Itf9+psysIU2A9sIs72AhGYIzW5AzxJ
UMC2P5cH4g2xAD8bZT7i9Rk3R/ybplQYZxibWWp/MRG2aMLdDcah1iQRlVBPpXJp
LwCXs3x2/zn8rC0nH8bt/ury+20gqCH+osCWGFNOCdC9spDa6wHlIJKGY6AFkD90
HaY1MMCurLiwUvtcks8emE4/fKL/qA2ZaseVirBnOUwnF37wDb7VpfZtOZ4lKK1x
mrvyzgQj/rV1Ywrngj3iS6cIYKjr/hWsyr+I2iDdC3S63bseZPN2qAN6ei2MRt8P
Sp7gAHPQEI5LVCD47FyNi3NAUWIJBBNHFhOBk/RN0IzFPcgaULVnId9I1voK/dHm
yndyWlbdXWXdwhWjRPjlZx1yBAMpHjAxUkhJiOeN1Qya6Bg8A7/sx/mkf0oluWGB
hRbqhIzSLKjGGqVYi6CsCjjGwcGk6+qKJo92J9coIYqIup7b2AK/JpoTHFvNwcTy
Hz3jukjBxpLev3wofokpBhJ0NSCurld5MiUQ+ptdv5Dp2Anwl9kvrHmFRzsdhO3O
KyCkfJGYObA+Uu6RETzA55aKxblwYYG98Z+zxp7PENeL4cJN0jXt1EcY/dyyFY/R
3mPji2vj8JUr7DhHX4OPdZbks770hZihBIdq44Q0VTecQmmxG+7nLLKo2ruWhUo2
Mt05yoAq0swpCBR2dupoqQcWI2wRqlSMYk8OzOxNHlnI7K85psu80HEbVyXGBIfm
8D+8kj9bUH2EWuR5jsV+8AhZlz6dgscOQcjOdjftHTX2Z3hMjWZJ9YPNAz8gksmZ
J3i7Gmg9xaj4c19osE0K3ZG94qdD01K6ukX4b+LrJqspwVakMX0z8bMLJeROrvJV
ZiPW2c7kg+HtaK3mtttiYcmEx6bg2lxScHO9QdyUGJ5pmlPSb6WdE/KAjSYCkioo
f8Ka3FTX5MXla0DzhXyITafd1e5xx+lS3vQ1f6lT2i+4MQmEB2FP7i03ZaLkWdln
L01VS97a84f+13u73Pvca+8mf0fs2aNaUIo2tHPYoogaYibjs6Weq4ERCYl82+n1
26y9ZurZOwLq08dXch6OAtdTkkB3C26gpeqaFG0t8R6XEp2aJWKq3OhofBSnUFPx
Phvm/BgiuT9QcXAiZi2OE8nMmEYjGubZAF9cCV3T8MgB2VV7YGYBGO/T8M7Pu3jU
0Fnu//tLQtyDDK2aFVfKhSHBBzMOxWRE+7VOrNQgqu4E0nyvlQS5ZydtA7evCP5u
RxAdrMe4bnaTxFTGIrYwbZTGHrTUDQIvBy1tnx7n/hbpOsVINyIr+UXObQt/mWzG
RcieYpWio+Vx6nuxNLnkFfvjD9DdELkHWXdxvSAC1646bwCPe8+QNZbBKZlwBrrD
fgdBRIJutk8v+3nIFU5dRj+lKZAivrDF3sAscGEZRDKaNfxZe3v7bBN0U/NXrzlI
jMdlkLmT0L8CPwic1hmh2R5dz8wCB/1Mg4m+JNmOuuXqmPZpO+khKV24tEP0Kwbf
UoJsb4BD93f6GJlxcGscPfsjGW6wDJEDxz+ZNJnQI60GxxiKI5qDTCHB86eQMW+z
WrT5J+FNrX+QqiSwciMZtDdKG66DJlnKl/q2byY59vYOELFf2zC4WAiEbPZUmV5e
Md+TUtbN3Xgv/jlznXvHW5ZjeSY50hF5oALx566HuKRjSz5FNqtJGFtpomFK7ddk
kfwARRyZTsiWIjJ0ZZ63r8iAhkDEPwIc+4jwC7iqWH/45gb9X5GMWgDIWDF8QYql
oSL4n25+vubBoc2PN4MUBBkcTo4Sa8u/l02FJAWyGM+3PISqoRIp9cSRJV6u1eUA
s1oXzs51n7iKikn9URLtBWRrJUIjM0Ta4yPIbpCL3ppJdCSBNj/Z/aM+22LWo/UR
YVK3lvvtOXRcv5IASSPO/CVxy0n6KV6hDHztzf8m4VVxakUj44X+QdIwOhDrtjSQ
9wN4eKaBZzH5Ir9/P+zptcJrKazCTilk4Z74Ni33tWE/FlljOnYvGguAnyFlESDz
RwLi5AqCIOGUAVeM8QXUfp9K85/kOD045JdSTA5ATdmV8snUT8NjjB6RuoC8Qgpq
PElWTRTlINhaqJowTzRthWnjV7C+QNDxslK4xQD9YpEL0hFZy+GxLl7toGOaSHf9
3K+udgnDAlq8fP+2ELcNNtVtlGpDIwOY05Kdu2GPOrdhc3OkAC10DmY3fhrixYSu
RS1RcGkwFEASJakwI476p22k6VqNRdNgD+B6qGT+pxDfVA2+ijktoy9D2F5MSvQ4
fhyyYSBJrJlUV4BPmjFUJ8cFrU/g+6nBccxJXb/2U1BYkypqmLbxWNAiFTuPBlFM
sbJr7d2sHXwrz5omR1b98gtWi2HN34jBLiuP0MCC89ontLFgcGtmaNa+MCtQPio7
pxgnj0b7L8tOVyWoiN415WS7GN47MsfYxj69dYYoX0J9yuujPX7egOnM6AMSL7Hn
sdxdmfEslYFmwCqxHabI1rR52cK1rAkKWvoQZos95eSeqmd6Ugoyf6eOXtLsJqJf
DfuZx0ZmUfnaDAipy40ILjHcYxaqQzWM6FCe+XxZrAcvfLr11AgzNbWxgSiT9ncP
1HuudSDPvHdWUpvZFdBvTa6ZRNNjoVbSel1BWIQxY6U/0IA+BeV8EkLZi+mQF8Cx
OmMxkcbyZa23ZObq3AON2HouhJV4Q08wJW9+DwOZd/X37kaoaEpybsN1S9DOzUf3
zjV3fA6101pYAa+0A0eiiUqpIb8hVgjT/Y5tWnwcV6HS0NTmmU0ZxVQPnCDgazow
PaD6mBZU3f7dScEc7MPmBA==
`protect end_protected