`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
ddtXksX2+yylW5zu6QL2Lhnb2d1sD00763mmSITNX595NcHTEkwn0zB1Dry37fOW
FufOhVzEJp80NC5qZ/+F0Vk7Ik02dIR0elf3clrjeJRK85K4e3Hoo4xn7YbFUIms
l/8VZSb14+JVGURjfswrIyCUotIzlzVYZ6gzoZwDXIi5gQIBf/gI+KxNXPaKV+PQ
Ufys/12rjO6aI/pPlqSm0hCvftmBcnezN2hk1UeXgOIuKZnogjOsf0iJVX2aOOWE
6pD/psybjbnsNB6kH5uFTA5frkzIzkzl5d9+YDm9OyC+k84E83I/7/j+rk4L2dah
QJOvksSIzN867/4Qt8qYTQ==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="MvBXkzurAa5VTw+1JJ70nePUfoQXBvZOku/SMmg4TwQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
oRtzZL4VJ4iwysPsC8SXYCzXS8Fw2gtZTOskLcDV+1B9Nzn1zTyNtlo6lNICRmmK
ZRVu2BmCc2G+fmzynYlNTnSa7C0Cuel6FYpxCBlOuk3OF2tzAmLAuDyOH3Z1Yjzk
a0aHuoCdIRKv7BrZCdALt03JeUmXKPdOmIlkVGFl8yw=
`protect rights_digest_method = "sha256"
`protect end_toolblock="Jn9CQpRhJt4rnzZPRk+dOpzAubz7omckX1MrFd4p81o="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 55856 )
`protect data_block
gD6l00tciPUa6pDNTk/+t0OO0nC/UTtBwLB41d4inuAUA3i/ALrNyoJVcBnAmEQW
ptbcNp5fxEUJjnOxnedyZEuEBxWRieZFQnkRdF269oPwTuIT+eN4tcfQG6SZw8sZ
VGAG9FsoWO0jV6WBTf1ZseBZzjUArqKXVt6P8oeyJY/lxVyEYLB71uJi+SNepGX4
9GxBgGbrFyThAmHryrvKgNV4oBlIQzVFF+zglhm1lUKffkRRK3M6+nGpcKdvng3H
UUZZStRriTSs5Iy7Chdta/G3ikuiHEy/7ZTHS6G+VThA/WBNvCcwQJ1amiKNwMv5
FulC2dkVLhSlef46VNrZ1hDjifYJcqDsEQyFFwLuT+EAHNG94w2fykI14uWFrdP8
1rKUQttNVsolrQkNShxzmtJGNDBXF6L7G5U+CQGPzDKzE5GW1w2uGhQoVvPcUxlQ
2Z0VUIohP4o+YLM1FzLQdVR/zSOnY5seRF5rQ+NH5eZqP4RdiRSmA8PfeTRw/zj5
zvablnF0F7lRiZjZ9qNzsVga0k+o6sxg7PhJL/iWLsNWQgtBOo0otcGLGlaVim6h
BMbMBm57DNVKPR+kqxN/oZYANlRErcD0VDXCKDcN5hcms7Q5U+Us/RqdzomfdyAM
4Rvvr4rmvvojMT7E0oKTZiaYTedvG6RAomotaepnvRL+zoTihW1mTfayicgJzzzU
D3M9gg80hFVrre+vjU3e0aNl9wXIjsphlV8gPM0KtlEhfWoOxO1fLU91kVy7HEfQ
i00noAR9QrbYWYxLPDOCERlU7g8SGyK3AHzBESRyG0XxUziNop8I4J1vgcda2N55
5u4fOjzVRQm4iA+3AtjzwyueBWS1lFFmLleTbEDdC+5QgTAT+lEmEpNBDJYl6wqx
OS4tm88cHFbAFJscHMudXGOXomRAo3FQ+e54dRrTmF6FmDy1rqTv7gbkTMxD9IIR
+Jsg5xD9Dc//6vVosRK+xsyEm/PPOtBLRKJvf1zA6yQzy8zRmY7CMGgmyiBHLDlN
lagMNnzymbW+5EqSMj4EUnwIssfFcU0L3V4JKYQWyguUAPGhlXc0ulwldCh8ssFy
suukmUTD3WKcbKRsJ1atGg1VTbPg/zyrgAmHNMEVde8ltCTViR41MwtsoVKYpVka
xkPVz03dDPTO6MMCOwam8ow2Ziq1CDG3AL5h8YXoMlA3N1EJD4WJmX1BghGqShl8
Cv3RLErJhQKexchNlsPOPlzel3Q+IVp/E6HgjAX/Y0gja8tzc72ZsSssMCcyMWUV
u+X2kNJmIusywdELCJGP4AgJlYM5NZnJflHdgq8gohACtdNaIo0Vt33x1DDfT9FV
ESeysEVSh4PqVNq6/IIjY4kVP85TsSkz+ZhmAxpkuISmLqQjEP0C2KgAYkMRgDpN
a+lftMWY6rl1nA+Nl+Qb1NYnCNLZ1bxuAGs6Upd1KLCOI2QWu9iFlevflDEnrwb7
KTX3IZx4u9WETrnxwJig+YfXTC0a8HVjbdj9/6ZR9YTiIoZnTKj+cZUubcwNmlIL
9qbqUKekiyw8vVDrb4Uz8WUK01mi9u+glSoDXjn7xs/ZUJW0UXkXqjVmt+8CzP5k
O3+iTMFlug4SqHNQWyaQV2UOOYrjErAPS5z3LN3SjUAhgyfb6H1T8RbHUuife8Tu
2VL0f4I/5P90ZLmrPGwM0Mo3cvu97PeZC+wggHkR+GymifodrY/54JTcFGUVhp/S
kKIcQ504kdOa8iqYTfezYtqygTpU3HmhCaSG5jOhHoL2Ky/fsD1owi/DFzgxiXdi
lzlCOBOJTIheFLPLi3kocDdXrBnPU3Z/op9xTcZUitOAiWsVAJMWIfMHwLwdWxsm
AKu+hAYq1NIw6bVeUSStruAxuh11SGzscICswiMW6MiSnQmh0Mr+BDGY3WvoS6qc
aRh/Y6n2Z3dyPE7Z5bn3FSnPuhVvapNtJMZNw82jgWQ6yeomTSd6ctltJUlTkASW
1rJVCmF8spRqYImG9sqSolNwwkwCScPnjRDLd5xdS2Kj3uPousimY1a0QkeRburY
CE2p8Dy1UX8eiAb7aNjQjojCo5s5XU3NnE0uE9wslZOTkosdsC6k3fP+aRahzR5B
SwiTwCmXhiaFwfTGSk/4/C0Y6UjE4vmECsaT9TR1EbsMdYMR9W5ZRRGFkYxDisQQ
UVNM6bodKIR2ttLmSZ8qRyg4CXQAY85YNiM1zFZO+LLYuq3c2kcCXNFcEP7If/kr
m68ZAp0CmZGYYZLsSRgfRxqIcN0T2UYZgisRcZ/UCpGUotZgO4S6TI2raayY8TLK
RYVwoHit10DTP88ciPkiT/fG/Bxw6k5300yNFjifI6aOP2gr61jIKhoJuqU4IKtM
YdKOzzkr5sliNV3NO2SE+ZYYepFb1zReVlpbfpsSiZSSkM/rSsF1Tu4u8B8jEjst
xZO5WJopFh3IJPrg9KGvg3avu4KphX/HbraZYTym8QncTc1KakvyIxdB87h23xEh
Bqdt3ZSGsu7gkP9KhKVqUCIioPm9R4VvO5LN+azEpzVgLOXEVUOhxPUWTKiOWqWw
63tlLSbOtNtm4/U7krIMLmOnappSuXe7IX3j10Yreaz+NptorW4t67sjVOg07Yrm
0OYYTz5FDnuskoYZpbBA4B/faQ5BftXpu8jHVMZOUVYGQ+hiKyjQV6PKYVcfG1ze
KSu6zox7XyBfewLf+UZnMmHQgAASicGopuv1kyQfvDEk5kiWot/BycAaCw5iO3Gu
sZy0rpHaBnYrJaUat18BRmD0JuzpeL/RKIGBHnO2/WIl955ymM4cOrglvGYfDv95
qqW6Ftl1HKr/yyhwNeiaw5I1jNKaEmtJLDNO0mJIrn2zKJj7dCK9Ecj7KGiqHXBn
XPZoGBsc2CMx1br+ticNtDGV0tP8L+c1IJjjX4zW4YSa56YVT3f7eLT/xIS74LVz
XI49uvSBBd7JlEtihCoZ7IAlQkgwL69CAg98gq3uTdqTANxV1PwZDJK5wKTveJDh
0z4xassQnqX+DPea23njikHwuuWcaKOLi05Y6kCBSo82L1IYXsFVzUNNFWTZYN75
wTxW0Je3ED0049WxPRwbOvZonT00/5ppY+oP+zDemRhbWbwUYG82nKqeyLfaYy+G
83Sn5gc0JsqMTlqKvn5VC9idDxxf9Z9rRsG4olFe2IfRWd2SQqUbAL7l4+9LlUqf
5Mp0oXWHkp65KaxsrevWJ+wG5io/IlRySUp3QJbrM6BkVf1+TJFvam2yxe1olbdD
Xv3Y0c67o2lUXTHgUGA8CCx/exK1XdrDhsDmbaiMn9oknb7rP8czYEqTHTfDsM8/
titmiB0g7v+GvZ8e0tVHbI341ZMgqZfaQ+NXzmI1updupRIBb3BNqEEo2Vf8ewQP
JkdkrciS96VIg7RxGkiwDL57yvEYT3c6sWDI4EE9p9Q1F0IAE74629iyw/p+HVBD
h+UMNhhg1NI2FOPBfoZtlBdUdvl7TWaPOSmYrJhVUCEebeynwUQZ+XxhXA47GQEa
ypBsN8kbXLJ9i0s8QJhnqKp49y1h6DAUyG/yED1n4/TKH0NmfZijP7S3ss1wbOWH
dK/rflOpkqTYYJgdF0iI2rhUOekAiWq3j/tyUDhyQ4ExojIOuZp5KH2IbMq/CrvW
L71sinsghVIC4mnoYODmRW8s5UEuWoTxBR0UYx5fD0E+cuBUfO5TBkaBEHTblTvI
7YBz5IatKS2yJd5eEnc9bQleh155G7C5fMy5cBI8yJ3ggPyPf+pOfAeuMoivCkOP
4X7nW7X5O2JtNA4bEttT21lsggK2tzlIiXNMCIjHX29gfXK9K2/CjVkVk0CDE9RW
RA5v5sHijwH1td9JAEmWsKgucwLMgNdJcGLyggw7bRsFYiwBDByYjzy1L8lBwERc
7RfPYarZdlUAYVJQDAQPYlkRBEOTYnDtV0zNzrhaN0NcVUmUphtgDb/1jFVRsdYH
qLrRNSImj4P0yOmrErppeliCWMMH752gmBBRKCctaaUVNqnYIEdIrhQKIXJeRUnL
0VdDYK73ieQMSqIvJ9YvTMUEVnycO+QaMY4OiZLWuQlv8Rci7UbM+7zAjDgpRB6M
0cVfX0lY6WuhBAR2t16YNx9+6lSUrG9p/a17vSvCo/2vISWsP4VP3+9YhJ+/G7ux
oVIrvVZmrj4JOV4c1Yiiu4QctYh83CxUkbwlV3MsmSoG2a0lorHyB2c6bflwsPP4
3A0PHYD6JA8w4vtsLMpCcLwU/qiXBxed+ZkID0cHH3sCFj/35l8F1qGjOGPVDHZ6
jnuvNOR/iYEcwapy3tlo8iwJvU0uZSBchOy4N8YhWd8MvmM9k3JKV3nt8K2Q8JqD
95/3q4w8JC0WJFpkLuSBQj8aT7qjpMmU1+89gSGy0Dw5/LPcqDqgrlo3iEszFGza
pjZD+vX3QuHCsQYth9H/ZeYklYf5dVvdyA3g3iwR9ljmaQgL0xWTTE5NmuA+Z6dy
X0J3AlFEgHkKk+5oiRxLB3q12C9jKYTddUI3UuFrPciXJ+DVS7CBMQD1+NfxkYAj
AcJGUYinDwNER9Ovp6LQblPfzdaEvU0yREZFpN5vOkk2+AXTDt1DiSeSA0YKo7Xy
PzLdHBVlPNidFYhyfY2nlerZI6TzwHu+QV3tJhKbCPDx+NOV/5bv6G/AkaDCmvw5
/ukfO/9WOVNLLX8ZTBITcU4vHpKgrW2lphnktpjHka1VdiAgdMMn/+gI39b9ooPe
z/TvARNOxHGmNTp9D4Lxp6Gnt3Y3k9cvkIkBmqRlzQwRSK+SMQHO5AcfBxDvyxmm
4z0hOPcehDyDxqPfuRAJm0RVPvrJGwS+w3vYhmjRLN0ufOjq6tqUomVhk5Qj3F9f
2sBmUqm42ue6hSEbTAyQkpll9sZesMwHrsBir9imjdbLrC6DDVQwc+7TgXRenebn
TkNOtATqUjhVtQ6SwImvxzqgLtze8CiXoGEAkpdCr31sTtpd7+b3tpr0pA2quWDq
XoA2GnTrBnKEnogpwmLcoeuRNsAkTMF/1JhQxqnjq6odRmOPL9/40MR2UUPsYJ6l
COKpEJH9b+BT6OtoUjsqh/VIaiNtdI4eZdOyx+EansVkKGot7iOSJ+4SAdUEaxed
EkVaj+f/UKL+CtYpl0wTvRhKladEPViyVnlRoidC9IABI8o28uxYIPFv4N39VzMm
uzu5vixOO0K/5w1OrNT5Lq9Wn871zFjzc7Mm0wcN2CF4jXr4ZgM5F4BhB/IZuAug
ltLhBjZM8/N6sQo5IREwOF8Qmjh0za/Ric/PsxoYNSvvxZMdOXF9pmZeDgLgYPcl
Bsk4j6N+9lNliWDBhsXEer1yQvj5zECGjTxdwGvze6798J6Dm60ermM77r/xoNC9
CYsboZ1IsFPNRNtemvU3LHPIN4YEFXVxXCEASEYos8HyQ0JG6CbKz3jEXfjuSSm6
sKWFalMgKB17ADic+V4MC7YIal5H0z5k7kmr6Nc3sKiDQsWFlaTXPo+QPQwBPqyL
oodCOTiwDeBzArA7DqNDCuCGb2Pd1yRB2lzhh7WpquFS5O+C/GwAIObT6datwRu4
6CJ2wcf+WtZ9pskgkfYQWCfPD6RitsBXAt1iXE7qcu9RHnCF/vywxosyMlqlaP5C
Gb/JxoiKvn7/uPEktqLuO7qhyISjuzmtyfFJAve1TASpffRQuTObkQPepWMR4gwV
ZT0ehP86dyMxQxREr0JThRY07zT21SAkmv1NLho2r3YqvnkFnxg1UQXwsJp+HPze
yXb//pDa+EhJ0tDcvROFicbjxDPqDpBpYbBs30D18v6DHY3GKerBKzwDwQ2ft9h0
i3pDAxLkTYTKHSYI7QlHhnf+4J1Z+UKNZl0hJVazGMaulUHuneBgWBgfHv0CFes0
GxTE81tQwFCRNqTIP244sAJPV853SC5sD0qY/VQkQEpAzkKRyZj/Vie0dIbr+Wlr
Wq52lTGK8vcnjSfFHMfHiH3EjPDN8oSjP2ECGYt3O9sa2buMeUaUtAfmwpf6/YU+
H6HM0g2fN1JBdC52LIQrNWz2EfeeS/GICBbrTw1ThQ1X3/UIvAkXbmC1Z7/7Ixsg
jnBha8waBDyySRZupdRHwE1/bLKJlRZqebdn21oh77ypcUaRZV3411vVOhT1fsnf
Un60GFkpCK6+e9Xhcz4qboXydUH73owbh7UAwj4MCoqRgayqMXC82LVBbde4lzXN
oTPahE5EkO9Bcy2WaoyV3zI4pYubEfnb3LHIQcC5fgRehzplYE2wNY9HCWz4jINy
iIFSmQXuqpyyCMhBgvKBlGVLUJsIhWRKs6oJXBF+Pddd56aX/8MJ+O42KdEpWxdQ
BXDoUVOxnTL/UI6EW2CuXIUxaghiiYBkQfsj8j4wxWUdDC7FuO1q2ZIzUW/S5YDb
UEQV4HG7ByaxUOFRLrSKpV8bP3zPHMmx2x397/BNOY/wnCFSXiqDgORpcHdHGh1F
IhDb8tua7winWYToOs9Lu94gNJua9DwlTO1VSHTam0XRXuTDDVVfNv+MT8kiKQNk
Y60KqmRCnQeNkVI5wSU2lNtrg44QI4Q+vDcFnGextdHh53MlMDUUa6iGI5NOXN+J
XGT6aeGY+US5cHkL1ipy2sGtPiGE0PbxwyPl/LO7JiHgm4JiloY6wkjlWOB85RAY
X/93Mw8CwxhRTXsjSb/choMSkPRaN2iW8bT1rx+1oOd54YmlDtnde0PX7UBYYOGR
HB5tBNtqqLQYSd8lW4B2LKjNMSvFxLacgc0cbmevBBirmcd52nv13fhXf5K+wQh4
SQm2YMruI0Q/pjOfdV2yohmNPxUYYTSt44lN9l7uWT3iVtPYZNCYlsnRuBWQKTbY
FV0GS0XBz3eUBtQD8TDdH4pkHapL606bbMWbz+R2CMGGhQhlaUarpMW0Q/CMOZ5D
+dT0BdMBmgETQM1t7PsjmxXzel3q2WXdj0OPRkOmb0n5Zg2gNSvgY2jUekkgFHAt
FgETwW2WcV+BMRkR+LWzgEu2Fw8wn15FFIz2FKtPUScH8Z2kkJSNDJM3G9CkFQBw
bZl1+M2NN1h7VDfF/9Cp54CwZYClEn+qjn3cfiRDmixxWHf7ESEQj+t51C8Djh3D
yAquhJAntY4eaJD87FXxer9paopzIhijOqfWT0QJ0h7Bvlsh3cedDCVfHJevlk06
tNdc55o2uqjkTwklx3Wj9FPvV/L+3uyAgRGd8AlEuBI/Y14dCqSDKRo/fuQErDip
0UomxJUDBcFqPAj9Zofhd/CRWLTgOYr1vvAb7h/9PyjQiqOksXGQN+6q+0O2RHdU
AE+4gFmHtWNOISePs26sZL4VBi60j/xw51aWNV/BC4kfxZ0h8srUyN0Q1NI5bKPc
Twijwk9eIbrCNN8Q/ZylFqlkZqy1Iss8JFI1kb5hYK6g0i04jN86L3FNgV57m3Y9
ymOQOwcqtKS5QIJeTL0c3LyPQLJUZ6s4XOisTUoIGWgUuWGvbFfHY5z81HwKfVli
7nNLNXRRPowexEi/o+qfzZFt4L7x5woQloRk5FYIZ8wxrPGGfmRxBHIjqIUEnJ/w
1ynimZTAbZHlLNoas5KD58q6qKhHVESNCbBUC8CC0rrGEMUHpQxB8RNSH5n5N0/s
MEj+KN0wwHftaXPPcKxZ2qflRFmc98SKyGhA1nMKPqXOiWPffhMw4Ix5uYjMoYya
ec+C3RjJar0wYOjgO2kLQtUXu3rKs0ytmLblLPMlPhoj+5+KWe0vXKbqaM3CK1zJ
VxU+iN7JTkf/UacDYZCVm/GVb4vuaPy7sQrAGTQrBfEqVfg1JzcmC4+FQz8IGP4m
PG2Fhd5yBL3YoSu1Kip8aHhDJnlLQd2nF6Od4t7cYyz2KZ5KtxbPURaJhwWa2pXR
4V8rMWRCz38O8a2kzB/6+q/vddNf85FD50gY//bICIGIsiWJ+sXq24QjOYhkB3p3
e42nynJYVCafko/uRIgazssSrxE85T08GD6WrsJjrW/PHl3njzCkYPaxNbSAROfy
QvcaBdWqOx47iaOlAsiPvvcDDqm3a6tPfnP71y8/bZLxoC0esWlrjRa8cyVKL43w
yigHCkGXuKsiUEoB9GNpFAnMD91meqOPk4WyB7g32VwRKOgKy4TRz5DUwPBqn/Wy
0zWxZrttPIQP44jPX5+W2jYnNk48P2VY+FPOEmTIh7mOUQX16STKMwhOEVdg1YK2
irAbVyr4tZOeEAyzqwibwgq/lAhsP/pPdbz0ezdaKo5Wf4gk2jrw1Iiud4wH6zWa
iXJPP4Ke2lQqAke/1t5ROSBAdeOdyAbVPHFlMObm3rswxX9az64sWXQrbdhrT/T6
WLrO5lh9wvwhelSikycKzZ9l2XgUGk3LBauJEaUqauihL/KeXtNsc/MJ+/c8QlhC
Zy0MKhwlOSY2B4gTQdMbuYGXHPHLHM9qRj7ymLbfoe0WJseeE33dSlDCwjNMYvbd
x092qI0e9TNigANmdfD5yzih1fpSis+jvFb2BliCp+VpQZ/jeA0OhTA70BRohREd
YTlC0wV1d68TaFRbqHI13vIhxFUACpBP1RH5i2DAKjYlR7868brb/sTaeX9gC8gP
GoIl/sYn8MhCdM5mBn3NfGCZmoLKsYjSnuwFefP1Ne/QXRY/jij0uv9nvHznMlAj
h1Azg3Jzo1QfMzHVj7ghogKI0ASaNupz4PMJmy4dWv++42YYAuTpO6RMvKWQJZGh
nMA0HfQGGgln38NXsUMpsMaRe+SsJqOTL6LzN5tF07CMs6jfJPNu2+Lr/Mj8AXqH
Q1Lm1yEqpZI+tq2VeELqoFXLqLOH6o8lH46Yo4LNkueBqMm1zguT/SLiCBSCJ5fq
VzqJj/ulcRIMx6KpQYDcsyUkxzFRX2dBm2Ho4XYK13pVNdl2YJAckMTm6L7FCWqG
i6CCzvwD4AOLb94oQx3TvVHotTePQIgTAGQB51UP06Tc9q+7ybpWKDg/jt0+AwjP
Ey0EKQYhDXYPxUNO99xIa8b1nJ/z+yEq6w5q4lESUUl/OfVk69p9BoHaJ+fKJLTd
NIuz0ZGBUU+11AP80hSjMrCfoz6DRO0nqPYMaWBGnCD/mAnE/MNDfCvmIQJ7S/Rv
NuqpX97bI0bwijNjmABxN6IN/Nh7r3bN8bYuJGlw9dBtZPd3ToQsd6xUHTaNaECq
ntttgHi/KA+GDPYpfTh1wWO2C5W/S06QmvSqT46qN9Ha3o++NZqI9OBdAhAItIAe
+YzG0X0sTd+qUYktJJ2LIG95uR7dSfIIcRoE90aw+wuUlhGrcr7HFgGrWue27qXB
LqBeKVAQnTOI8+l+I4VRtMTYX+HBCoLtZEhiCp3qQnOTfglZeqy1k+r4J/4Kjdd6
cOY/1J4COdg9ItjlhxDc7Zkx1BCDlLHSEY/lgGjKXtQloKlo5G9YDzzoIJdYTiWq
GrfjsyBLai08KM3pi0Bwk4exbvZ/9H1vjSQhgc48U1mY9cABOaUAxdghtQ5UZrA0
G+lbTwy2erR29H3G7TJCe2lrulo6LtEyhkmBRfx37Rd5suz0AkTgr3j0sU6Qxv8z
UqMUmS8S/ePARn0x4kaD85KSa2sBK4W9NIMz8D5+tUrDGM5EUl7GUyyO+XGB4hg+
UIl1QGaH2B7BfxuHFoeGl5JxaIlXGQwBEhLfKZhP2nc2Cx4dx3rqpxC6QjfH4lIJ
BS6Mf2P0KaZpQaSz/xcY/l0JPcvqvbWuvhQkhzVTo5CssSVnlxd6iCRV9xbj1LH0
dytRToJ12wA3HrZ//fn/d6+DwwFGR67Rs0ROcclJQE95eJPY79lszjyJSnJk9sIU
qZJZFMo0viQ5SYFXZntIgQ7xOWJcTWMcVVROckCDwcJT9gYib0jdm1RGUoayAgA5
3YZrCpV3PtYSlb9eRHcOQYv2vTFnIyIMMCSRrJhN/IQcu/upfoxvo0c5I3lRCWgy
fvwMBvwaF+K+w20bujiNpolX2QKkUfuUDwkMtqpa+NpjnEFxydrgbRamzBFfshWv
wFdKZQMRgTM9NDRCJIuDdX9fQFj53/reXO2pJM86lRW4L3ZnpfTeBqu3W3wegSYE
VSm1dgwYy11LIDjLOcVuvGrFTqO5pzQ3fwXq0Sl1lXv83vmnC1ZxSYbTHcY+96P6
ew9P45GIS0MN1V6gVwdJ+pY78GyM+RKVsriRJKtBCPqva1KK9h6TdMgygjZfqyg8
4Dd0OXqC2ztyDI5TRfFPqSv8quzu/6eBfZuqoVfXilOSEm/j9Ym0/6sCtJcb/kT8
GcN9zf41BiJMlYniH+xdoXPYy/5+OKmcW4001le8AK8CNAwt5hiP/+GuEDhjigqk
dNXjXgZi47k99FuQeJCU84nDBONnPNrGqBW+mpLxXRQJN+8H8utHh4pTqVnJfYX9
33+QoGhm6HmEkszriOgsn2MTJTo5mHVxc481bKauMYhWnJlHMfIiVKfsJh7su+Pu
3jBOFaewn+/SpF1vXlazgSRIiS8w2i7HW6e5YukvAhWKBtlLR3bwvNZrwe7cYC9D
My2h9f8hJi7davqiRIBuQVo/L5padGubsBgMPbYS0mamVM/veUY+3NlzwJmAR6se
WxQHtB2XHbTIT4h51xlV+Hk+zUElI9iJcYK2olbLs+Nedb+51f49XYSEuUAA3KS2
KIa7sSdU8vOTyCNDkilIOBY+uJTbGgRG0kHWkc7wrEpu/Ojbaq4NALFIOjIH3lqH
l5FdmTud7gETP1KArSVYpmlnsQMk3bQCbmH+A780lyWj9P2r55g9P24SK0lrLb9i
Z/O4OohcQIaUbj6CEE1svGobAcOuaj9yzvHiygBvkPoaOKvh4TxTkri9PI2PGORn
e9lBS8jxX/sXR57zkRR9M6rGOhAodX39QthdNdHksUaHRJgdmXN58htb/HOL6h9D
PpoK8VTUvUNFSZOPQopt04gKcvYEMBceYYmS2QTfA6fn5IskuWdIxCNW5kOF0Je4
5plNyJqiuuLpEj6RsPJyzh9sIGu1bsnd6j6WUh1XFyjVVS1WH1lsr23gFZQ3EEoY
objkIv0VoOJ3KkvmtJNKksNdpotvjDZFbjarXUOpCHO34gVewTqMgDBnL3f+eKB/
oh8GtedB+VMb07NeRAYT7qemTdo17iXSI2OoQJYiM9C8SMztV9y970Slwr3tiB2t
aFjrCijhjyBVoT/zAx8jEuNSDS75U6cS/FS+vApG6ja5eyl3OjMWRW+2mOcrYgXc
0Kz5ai+t6EsdBJyj7JPPTv9k54imA5DsUK9Jgc4bNr64Als12t06O+gBHqKj4ped
+jN8Gvb5E33sfiamNJa4eAr0JmpfgGR2lwribKIBk5XLn6wlKTMus9p1XAy521k+
CH+cjdmAxrZHFbQHQ4I0xYuaRa7pevMHf7gmYP1goG4xkulOXDQK2HOWgow1ki1b
GFdN2MlDXcWQ3AZ9ENWMaDNr6jkHujO3rNJ1y0Ew7grjYeSrxnKpixhr6StAHQGZ
elGyfYO5nQrZKQGDU2i90+e6q+aNlGVDnQPmmJmm4rH/SAEYAp6rM4ih8/qPMeu4
9z9Vl8tvdywdd9g7gkWS4oHm3Fq0VJ2enYX3EwPh+aJWVfytJox4TEHpw5BCAtFx
o4pD2vT5dW8c9sSuVJ6Q/LUUk9jEr3smhnqiFfQUqAt09JRU9z+tH1HJHc/A/d1k
TkKuHVtIjDKKH1fJipTSz9I8t2aV27AW1JbAJwSj0hTsWCGGaclNQMyqmqVbTcc2
aZumKZdF4hkPYtl95Xw6R8GS+N2D6k6syLnY2fgd1q5nKfgkj/M6osQDCZZVEngN
0HOmf8Rzxxgj5AK4Ke53q16/Z6Mn8JixhSvJ7QT2SThBcR57CUT6z3CcQndNFdvO
4yXy/v5aY6S9wiV06ivPya0knhJhhDNGGHpIIW4juLITwnDReUDIHIlPb4hYGH0H
Tt1PKkqkRcHVfaORSwUEIP//HhJNwXe2h95srVmEv1MkSnReNiUun9yNdXp//zz3
JPuhjTMN/+n8Vp7WMT5UfX3v8uHtvYM8QeOomYYGIQY3/2Row94gjWcTi713NxsK
ivtz0VLUeaBuK5ybfW2hMYRtUqjscgts19FozoGRdqWv5Lh2Sy41+Sk51BsUhelN
Arqn6s/Rc26EKVSTAI6zPKskTosL09ECko13blmIbWiXZ+FlzxVbaiQPlBQfOHci
7uDc03tejx3brTfjtsFgHAH8AUIOIxBecDSuZ0kLwZSaTS8wHfYjGf3feXDmGvn0
07rNZVVOOd83CwAMZvedmVXMQod/CyeHnCBRHQ/ewKm6kUkEKt/4mAUrMbpsXWz3
33fFyx5bKkfPNDqrhaVThyE02dleM+ML5F2sFGiA8yfxALzTnBVrXnvQrRWViSSF
Pp/uSf491tcMcVAwLpadcnmDYATcCRNBBxFa211VxwCM3LtR3UL8s5DjxEoZBizS
rQFC2t0oT1OVcBpIj0II2HI0nKLc2lixfPlGERbyroNLLJSLNwfbXlkkFVU99sbW
6i4BLKLSjDKUaS3Jy8s3761LD8JiEQDgT4mYyRi+IFusdAPYaXbqlukxLj7/4IVG
ZLCZtI0K0cDWnF+aQyPFX+jfpuDXL5jszFaEKmxlyddlySYhiVrGtyBV2Yrubttq
ITgFXrVgycTPKjX75xzk7WwHXz7kmDDRqjEzhd/zn3OiMpKA7LseR4ayJatb3qBG
VbszMyHjS60Eh0vp75ftKchbCNUBSUily70B6AZzG0VrYgHS+VDWGf07btX0fRQ2
gNy2rHez65N+KbJPwZAsenv9F/XO/pFw0nDqrZsWME4Ml8nvBYxzvuQAbdfy7yE6
Vcfz/pOqHi07mFwml8uufZP2DO0v2/eQC++LkzzLKDjJpn3EZTxjcoxT1BGCHAx5
ePurg8xb5lD9D0kQItcgbaKTuLzOTF2jAfDKVcPBndv+Sg5CNte198y7jmu/3UQf
OSK46Co19gGFm+nhYOxHPjHm6ratbCs2+T7jSdVmpBWnAt1UI/gN1Ol+T+ZhK9fS
/Z7xZ15rk0z7YMU0CkXDCxebC7IhDhe9TnveMBji0UDLRylO9sBlAfHPYBzkBQZP
VmaTQUj2cC4jqanrJx2ayMu9K4b5yvgnMuOHBAPIWph/hZwXKuCaNo1TuTbQMnYC
JwM6Vw1krBpHjPqzYFxVj166Z7h2dPkGpA/bu5LLfsZP6l2b/X7hr1gLFJJROT2s
ktipsJ/lWTo16eZLgo+kmuuDzEkPml9y1CMf/QU8cR8K1AlE/V3ds+MfV1tVEcAe
BHQtF51fMMPXGwfy6vZ8JY4P8fnYsl7NIYTjSgxjgi1ObN+t2ci7561QzU1puDul
Tv1w4Horokol8YbbGfvZgXYrKhtJ9x2CbZ1Q2SCTEx6vu6XNmaDqBwhkrs2VYsJn
qzShjtUa98bgMEqf5vkkDncy6tyoLq+g8qnSbo+0PxhI6Snxbin/sxRIjo30yOqw
WqaEXty5YTUo0B9IrFvSFqMT11Yor9iG49qhVjQjI4xJZgaaXWtmI7MKoqvkLlRg
S5y05IuVo28Ift/WZuPQ89Ax4jG/qjV6Ccm0rWSijb59gYsZ1pDLiM3wB+ud4l2V
cblUpwWeZJ8UPPSAGHUVjjyVbQ0lQ1nykUor+iiufnxGuMMCVyfku6GAip1AfSLx
d2X0RDrmoKi+MgI53pBHRDkdXP2lkbo1TE9u8exGbVNEnQ//KPLX6zBnxuGVYbFy
VD4Wik8/18AxFQogsDDbFHP4JZM90gH2sy639/+f7eBwCOZhBD97IJEasAnGcWyR
PNaaLeGGRxV7jAuj5qDVfYNipPyNsNRWBrIOfOKdmMRM2Z2od4vcGkgkrY014kZ3
QPBscK+WUoJXzpfUYKvpVETolcPj/yUDI20+Tzjn2gaJyUBNCFlPlz5HZUTxMNND
PMKOucS5QuMvvkZoTVMVj5PLe4gxBZqhktz8ZQxeS3f7hwV6QfTXPKN/ydp1GbkI
42I2hGzGoEUgYaW2iLnjtS6L2DY2YNeGlLesOp0sFS46q6r0iZ84X8Vv9pStCCVI
szA+MEU3XjSvjEYxm2gy63wDetlxdKIDJNY9yXupeFIfGl6Z3TLqjW/3JIhKtPNA
GejSPFuYgRiz2tIngxnptkOLAeZVVobR+k0R4OscgZkDgYn8dPooNMuMpg7iKnEN
kgGO+2Hf2yqvndkwnGyGB/WH6GJMo1zLXe2yHvmz5x5YjgDgM59QOe6znIDY/V0D
gf2j0cgKGBBb6ng/eYu4bEjYOMRBm9+4q3aZFyg9qol3noUzUBUT7d3hIs1GxBmi
4p7wl8d+tlt33Mibpx5DHZzqvGKfShC5LUDOG6pTG/qt15sheJDoY26UNG3PFLvJ
J/rRH8P3d9rYOShJLORGBSaKD8P/U14Ovmr5pOAMKtmewAXUq1fkguWUpn9Hxzn7
jYCSMMAklKSVuG1CyUw0M61Aoz1U+IWGidA1tDiJN6KzDWld62GsyLY6/1aN4x87
+uAuO1uLOXYNQFP972D+x2dfp8BWG9CvZ1GcwZ36CWdxH5qwjrlFVeWcVjuz6u9G
7VuBBIdV3X0o55+F8FjurbxlplQqMmO6Wgw4ct57ZYPuskGLw06MwI50yq2kUf6Y
AIn0HDsr+fC05oLooaCzQ84D711EE3HKzdocZwdnKn58MxKmbqfp5uGcHdzXg3jF
NiBPT5n0tYHUSwCZgAXNqVOiREe3e2FJlOwfSYayEUYi8U1nPoCSmcB6mPXC5Ufz
uZjVWAzgxG/XD4DdWYmugfABuADOtk3u1M0Qty3iTCdv7O1SQt1owB2qrcLkRQlZ
S+ilfr1DEFBt8Mv4obqPLSV+qBG/u3ckVKhZLk8vkv6LOmszl2byWu5KwtNuEzxv
8/uVuFqqoAjigJLotg1MJzEBqAUGRevL/26IszNnoo61Its2/DsEymFYs/WTbWLD
5oo6q+kVr6ckDJ+xSQzvaaw4ryqUTVSYHvONvelGNq4ZbvXAwBrjp8dwfWczaUhW
NbN/OaxIaV+81aYRyOInHOVC6rNZdElSf41ZsHOS1/OSbE57tIb/zOQN2tsfKTR0
eGPraDIueEABOwwo8gH0nOHobjtocvF4B0SZgujfsxQNExZFQS5yfnHICk721+Ov
sW9bLlmifCvX2TqMIjhVpwyKd42SLHWTaAYcqX3QRjHej815q6J0HwetnrDKw9xv
zq4M4Xqvg5EYDcoBzSZotBDgrDS5Xb73bqDFYjSb1IVFET2WEFrQUQj/6zGGn/dZ
84gVQVTJQaIWkklUVi/cEfENlJaFPrvLpUESV5pOZvCx9pPUOcmQMR/fSwaVMyvA
dWF+bxPRrPQ1/r9CFwhscNiMk4zWWkTs1c2tO73BMi2Wd8mDonewzhBjYyJ80wAe
tIB22FmHKKbdzsYLGwFpuULdERSLGBQX22Y7OSIue7NxTn5XBoEjaT38512oOdwA
nFP55/Kx4oAiBIVRVXc5hj3VvmjO2spS9abhJPQqfXaBMXMB0BiZFvNsR5Rjg2rm
9bCC6EXelx0lZ8GhoinYKs5Ut+GKCTbRaV07FjBQEm/Vve74O3A9PFzXVWWuXYbG
1vLyAgtouHgZ+vX+mVYUku0XvpQhA5sCWXffmio+0a41ryKiCH1wFNaLvB/Qvpe2
LS2Zu5Q81M8uY4QpOzQJkBfV5EJoVhVGLxmFmy6VRwzlWSBESVMC46ujW3ihJs5t
K5GEy7GZESqAbARgj1jCeE04ZDezVUqd0+spy8sZqHvbJ6EDtex+VfibAfUBm+cg
ZuU9LPNEOVks5/D/OulknJFcP6jKkL9frwkb2s8cghyeAnQ8pHXCN3S06qzP6EbH
/+mT0Wcj2SWWRuJGdXRkNxmiYCIzs1skrGjivV3CS7CboXIyJH2/eX8yethTPQ0J
TpjVUOYVnN6UF2v9mcnZ2QZL0ygCTbHmVLwMvEcmoZ9xDecuMkBKa3XX2qVzA9RR
Xb69Bn2nibUMXISwZY+srD7gwCFaWuVN4aPp/py/B7qX69tbzq0fUCzO7CltuA+2
7+JAdiwM+OznB79yogrQF9ClMvXr6XL9HYopV4CNMQEIW4QriEST+wTMbotbQrVW
dmcZTN5q4gohmk3JpwHwPwZ0r56H18wyQVZtCTEpwG11VMdnUIrYpD/eJ49OExkr
2p4mtbObcoQUQyVEPtlmgeYREx8VnG7xsuTBkdixvBmfDiCEVZ9rT9IDC+bQpPR9
eP0vyRrDmHamznq2Tk4E9sOAg9b5SdCYUIwZ5tEFKJbnDeA3g9Cyd/hBSmjEma+f
ag0vN9UUnYyN46mxs4XAYKIIhk9ZiZfdgVPC8bFTvcIVielufbyZsRzOwk/m/pKC
4FJ3Cca9nHcXvimZ09ofeIQx8ME0TQ3Uv09XTR/6DoeRRY6SKuD5oUPHKTxQb73w
dg8X2aArcurhZZwb/GrXbqzm/jj7UB/rYYIqwUROJmKT91KkBBRNiVq0Dw2UfEX9
7jtVz7DNEDFpCXJyGhVPVVYtMPRd11l6ZO3x/GBZiKA3w4FPt1RlTmbXHE6RVC5a
3VNbMyzU86nUkad7Zalb3I4FIKXsWGgXX6G90vKPCpCiW1cpNq8HJ2EwK0Yk9l9f
sw/zWupaD9edMp/fkv1IV9ByL8lJm4e54baukmw2PSdbUg5g7c5PKCPwAl79VtgZ
7qzTN0DbOIWg0RMSWECS+z5u+Yz7lQw8RpvZywyk76m85ns3e58jKgw7cHucFMDp
mkbzqbqqr4G/nHBPPu3TXU+VVAW30nVofa/1GXOS5Fi6G33yfc/lPTZNfExlvhHg
sDtxqsBUqg5mqpNTpYLVT6JFZsHmovIN325HLiN7sihXpHa9M2Il4dj2FL0aYfx5
HPxQE51uM6xH61OYS3YKnoLpc7T5F18ncmDOfrPZGob16ngdEf/Io3NjvgL0Zgwr
TtikkX7aMkJRQRYXSdw3GMjedDq4oop93KSRVuaC3mC5pm5NxRaase+9+XTVt7eg
29gsZ0cXEh3np9wzMUMymFPfMuTmAiaG9vXZ4wUvUlH1M/mjCY4JiLcGBa6EZrxg
O24V87YuAmVkXlxiIK8Gt2ssF75L18nYHEibPWzCdZGqV+VsF8UqtJ4CwLswyt4/
p/KX+15rgqxdQg5WOr40bId4m+KkZJMxktOdtkrlBijVTfqN+n8pa86fVqiwFOlj
CjdSkOw3UrCWtpKkEqtV4ZbpbgWQiF/AIgsGfejT2Uuvb7CD751HpD5LZ51BSA1L
urNqh9SAm5kEJsSvAYof6nOa6lm1IKsJBlSJCOAVzEHmJWFlxeskO6E1hbPEVuMJ
dW4wUejih4B0BFaezhA2FfR8bMqvuIidA2NkUhmCJ5X4sjg1LmXcWbi9YhFfK9Fd
N5O6M7UGoYS/Mk6eJVIkQiIVM2dB5VfpseOkXA/j9d4vrLjNjcybh8vWhLC6KUtz
98vEOSklK131ndRwEDPVIATPrLzkb4iLkofro0/ufljtJ2Ac46XL7O9Kotn4WS1h
FXyY6FEp5paK+9+J1zxrg4FiTUvg3H6hnWwa0EWqUVIYcBCgQT60ouxy/R/vCxNW
nACW5YSbMYUUJO6p0x8gNQFXMEXYAUuBdXk9v0ZVgH6r5jrMsMcroD+IncMoPj6u
TYPC5M7RorcFB5QLDZgckoIoBisnjwVXpNfmQTwywzVgOAvtfC1olVbzQBa83ga6
VNXzCR/WFFB8+PytyhHcO8yNQw0UarYQ8x7g+hQBzF/kOQoB78wyetnQYaXsFNjT
8w6LnG+Z1WqRhx2dVus/YXXFxsC+CxfqaLnM92pJYAnZIIoC9zM9dCOq6Ef038YA
TkK+U9lTASOPBsmz3QtLGUlHEXZYSZCtMUwsJVerNw77lfl4bbh8XFpfhJbJSKZv
5dCaYi6OVwEV9R3dCRWAL1BdhU5URKFE35yB5pv93FQ9LapKUVg9FyGAm4DC26DF
k76EH1S/1Wmn9vWS1QVdPktTBBcXMKeZjDBw7o7ESqeMwYZ5yWFJxkEH747dsP6Z
yIVR3y8IR2j9iRKM5TQvdur9+ys5B2ZmruJfJ/PSF4YYiqmzeY1Yw3TJtvzZ1x6N
qNEaCTw4lKi21T8l/K3y+Qznp7zUUx9yMeETH8nTX+jxtjAESHU1SCPEhiaeCdec
UcLVyhqXXteRz+053AJKpBwohMgOj492YB9e5chaiZd1x3KvFKz65tobLgeUf4dy
LnhM/xjl27TcUFTFRL9c8x5LDGggnkcGHEeDos/7sT9YtUNu+IvhsYg1XWAHFk96
pQc3NrgSAoHLOSGSbbWqbBK81mO8QmwJ4iv7EvJhR/8FIA27vr++vqZWEj0nyERa
ePn3Dm2smz1GIpdfAjRyJSaY4m6cOOaqcKBrGx1w2BCDJc1HkMEb0v0BcQzb953A
J+oqB6rpa0CUZ+B7tVeSA8oS6MtzW3/AwU918UVZQm4e5rvK8s3ZatbmdF5DHjrg
0fpoMa5re7n3oSaHB2xPGURuYr916hSFUocddT74kxfqt1Thvg3yzEnuBicX/sfi
eYaj2/odameuxphe04W0BuXAbr+Zdvp4TZXSEMWJeNl8ci6NljqHCmEfGTy3WQea
sM9QYkMzJ1Cepg4lFhFX4wvvpqED+gutNfwsBm0HayGaERkypul99vsK5ZQV3HPv
jKg+d4yli+B9Ltmt5y2MKVzeBANRrd9Lubvu6dn6VFU58WBZiWQcM53UVzYIZwHL
Suy1ZoakUZXXbFjijHWL5d24NtGs6Zwr/MZVFTK8dnhFehf9Zqt/AUwR/bqaqCu2
dwNHMr3a6VQ/vQNe/sz8UYkDZ+X/O3EhCP2uiUnAKu96RPPOfM4oLK/VHDr2wIYb
vseQ6gQk3VGP4iPp6NJ67HOQAvOeCJkNuBT72VHUDCt3gdBHdO3dN9Kw5Feux2LA
+CicbCga97f3uxr7z8hbfWWgeAq21tFioOjM8p661mcaL7ZIdtdqoNnGR3z3zRnr
CU8mNjf0cSszi0v24/hfr8HNZZP+/4eB1AX3rrzLbx4yoj9nli2pMwsFwgLMvX/Q
IhsxIBS/MDlEINLKTUHMxMf2SeGvKMYJGoKDXV3GgY2exnzk827Pv3ZnLzSB0EbS
A3vEW+WZgddEEsAqk5euc3is0zGsaOm7pE6mIrUEgO3c/XPo4OI8ck1g5AacpGTI
yvJZj5SzhmVKDtdILmMIea6KkxMnqWeMF68D2CjK8EuCiIjkgans0NJW2+xOgD7K
JaKSyqeoKMVzDrhdl5IMDBLwSZU0CjcEbLB9rr/yHYnl723nVAXDEmKA6erVsXmO
Ja3EPBNrA0AkVZlVoSt3Jq8H+xbImoBtGDgIZLa9eP0cSZOjyuIZ2bPAoZiKOMBD
COch5a9goEsiWMxlINMVoIvmHd6eA9DJN1ZclKD+X4oT5RyPvIVEaP8PzWm5X+KD
DfMBKHiLvBBH120jP/JKpX6BWkbf3fVMZNwg6YiC7hbzdgx5CJ+yOZMx25Vt3hdD
8a979aReiMteYenoZeOAB9z+Xv0TAtQaYsEP/I5Mwm+DeL5pbdta+QGUn67MV0v9
K50T46Qn4OR+pAUDZqtWsXpmsB8YvHtMdG7e9v4tk3E2SclA7M7lc7ybQMZkrOOo
LIL6zHDUCwRgwEvP6UBmwOB3eP4ZSrNI7zp/K4TP9SoQ2XjWYck7vyQ7RTj1UD0k
mXcPJ1yo+MzYh4rjfL/7WxSPBTeil02T2TSFq8rC8KPE8geHCH1PC0gZpfRsFy4K
ZfIpTBjghJYMfZ4UxC2jbUhIuzFmMj7QcplmlzBH4J2ZYTjUFh+mwJHzz176a1NH
kj//jFlvCWCN4+Zfof087Kv5YGkAppygCD5dQQeHIHSmzXJvQf+afyVpde92Nfoc
pVlH1gpotwu6+9ERjiasmyFMbyhrOvhWcoNFZMjkJjDcpC6/1Ib3YmhWK/+z6orF
uPlgX5doCggknF7hC2tOJiOC2LrmsqwKkY6yKwDrejaAd00TxeagZDqqvndt+ekV
CMr06ETRwunD+2MGHQzTN69HQHJ05cumQWfHapT2aSoa28ujgKcjIcem3ReMiJ3G
5v3cOWGjMKCuyxN92LwlfSPCenR33d8rCzQTpWsTEO6h9rQcCczn+d6KuXRB/cs2
7xw0s1THWHFFvSsOlaPVJ1xrg2/aoTRRHpNiSP9SJ7IJW3+6R9pwC2zt2gRHY4Dl
r899g2UwmV7w/Xc5uk71EKw2pzJUz6GudT24rCjn7Aac3qZG/nCv84ebddOVLqWi
9UaWPlIrwBjQghMHcQdEmwwAzzsbUMZC6y++/X3o/FYdQncqGh1yrfzSxSNOiIhe
xTfQL2XFsKE5zZMYpFYwRtazUQc3UnOtgSXHQW+0utCcwF+8mOFXszOJsjUXnpn8
vepc9T4dX+4E5I+6WeFz3AluhhP5fRVbbH+ftEwD6roY5hSASG6AkCDRC0wjkHyw
WJ3DXfp8Pr5m21n6HO9V0XNxu3LtPD2m1ZYpHhkj1XzCrg4I3GAJJIpQAXhqIqcm
6nlgdJGnXx/pgJ7qgbpcKYCuVO217V6TdbDcp0YQgbB0TNq4LwhyYVLtkxyV+3yo
pzqOMy/qxRmqdwaRrzM8tc1hry1c/UTeIWjKCD+JMVH/9Rg8Cf7EXzJKqcQiWNmV
jufu+HOV9uyinVx5OXyO/25L0EUCB0hOfQQYe4+Frx7lmkIv1Foc6CDAJZQ1QePL
IM+XmXz5GFSzzr/wgfMIgzB/Y74acsLiLYYxkSU2Wvaa3o28B2FfxMsIErn91Zq5
07cbjDIyeHjuYZNhVTcWyCnyG+d0gSnlQAiVKKjj/bxBk/xaS/mH864TizR0I11Q
PoD1rbYlrJzy3+BOEvr5Q4czaeVy5hS9UlwEs8ah/XTAafl1BRMPcRNp3utOXF5I
aFrW5QY3Jls5jSlSqJ4r+1W9o5NLQ4bGDOCbAbijrHvf02a8MLjmMN1VylUfjukg
RBUH4kXnEV74D5olS3E2Zy07XELliL5krKXPGMg6bUnCaVEwdl0M+GfI3guI9jg/
2d+q4uvKG1BX1mQvxWYMuu50GiNKfUdEz6NAxdfbbk9MUcYEDGl5PyQBgzJa0mdE
dsUCZZFfy4sNN1K1um0b3RNW5z+MuJEy34O/JX5flWMoaVlIH8xiQ9M//tZRFRwT
SCt/TWEemAurTiTQCXqK98QRHTEYMZL4NvDop7aAIY/t1wyFNVyojkDnONd7eCgS
S+phJvPyToVZQO/5Ox+7mulCe5G8r0a42xdPgaXgziDqGzs3eeVOkoUUO+StTBti
1hlk9T+RelvcR12S81F4f+BHEEkPyzYPh6sbEBVVUDPDpdflLGxZiqfmpxFOIL0+
/OwVH5+SRXNUHwBdoJFzBwf2nBoyp+7fcblHEUeGaYHVxk0ly20b3er3ZiqGkC7s
vGz+B9JkYsBv+AABXbjkLfpaKnCmVM1ZpyyVTNM4ucIOLKeMKjHgh0phAOlpSy2L
tLHJ1Uc9EUvKhUU2WBKjv8iTukYD9RWJjMZwEPecXXkufQ9Y6ohlecIZdXTNACzT
nEfgbQaqJuMW9sDWCC7JU8dmXIjMRtutKgm3dSNVBVCGS/pN0oNzn4pE8QEVPg1u
3N9UzWtaDcREdAr0T7v+L6mGGcynNJ9Fi7HBx4eLZgP6KU79xXQZryLV5eg9lsFw
q0hRzF7a+y/El4KvzBxz5MGtj+AzXCFwx+zGCtthJqJkFwqDu7ywiSY0zBydyPH/
Qjup58d+R09OnXOaj0z0rNdtgMeDl6dZkrPCMBCxF/prq7m8EPbxEz/GPfEM2ebU
YfBkx/WQholz1MR76526cRve2d2zZDMUw7tI0OLeLIytzLiF09jlHF5YHfSs5CqL
xu6L23uWAYsTL7xZuatNw/IEyWFAY+Srx6kwEJobp/MRFHovWHoy332n543OEmw5
HKeEyVV2KaohDB3YHF/21ojwncIBelH2ENl8mUDo/+cgeLlNjEWQo+qmDQaWDIx7
4a+YYykKRYBURCfLKNlt4sQ80A5TTewj4vPqmyzH0gUoOQWPVwa0F5gxOMgb1kCk
oxC4KQmnDbZx4qPI/xL/FoZMeLkiLGye0mnzd8OExFb0+2RE18DpYU0ys12+eSht
Ap9VGzpZ/+QPXi3tPzplNK1BAksCWYe1ddSo+NR+m9VlplUycX/pf4lKlzUrnWZQ
cfqRUGsteMlSZy4niRrbspqlD+V+w6vU1CgXMIrRie2kPJZnpZEQioM8qSSusrBh
RDhuVRFqglctwt2MwL3BoNx864F/zDfYMYKwBqCRF/kqxAj731x7DUZ/siyo9Nqb
3gwaExAwY8QAYgRYu9WI4rCo9LO9xGzqKkvOKYa4OeoNTtsL06IbJSg6dsB25egH
ptIwPMHV6+df+QLxwafD1OwcvCd6bu0GJlGVI0dD+0DxYn1Kr3ELdNMUyypbB2t+
62zjH+oSVQmSQ3CKwpNAHQZNdJf/RyxU4kocLbXj0/O4wDaWTKaJcEFdLYDf2qAk
6Tg82PEnHPifpJfOOf9eGIxvb3NqD6DdHVmjn/RXEOoji6SJL0tuyIoA84UKfXpO
Sx3k7xyAfVgcD1/dT79uP2OCaRKjxM2a3iSWEZ32CTS9X3Fu8tiz3Fnyu7BJD3Dg
v+YREQbBSBc+HjpwberVy4V2CpALe1zdF26G6zB9acrDEDwg2Jx6YDR13SIpXqvw
dbuMMHaaNTDCCsyJftM6Gn23TQ91CLEX2vNGloGP3B9nAzdpuOkyNFdt4PKvNrb6
dwQEmW452Vs/FPt3fC7PmZnOuXpU3lSTP+9dJ0ToWHu9ylZJxzqp2BiWlj/7C16n
4AL7jYSTl2Bh+QpqMhzQHiQrCmw8MbPBpTD1zTAeaFLOAprtU9GwI9TinzUSL5f3
TTRXAbTwt1L4k+EdIptruhPM7AJpD6yEyDnAjllVYInegR3pE3WSpD7giN2d26/G
4QpNcTSnyeFJOaBUzYqmXQlchCcbZVCgSIpUX3ST9wCVxeC7mLeHf0YrZ249iK0R
FsXiuJXRX+QWFUNfSMkI+SJ9DcMx/xmRMo5PKp4RFbndU4RAsKaXTOwb4SQ7vHsk
Iaq9quCB1SmAI8kJ6RYCW6Lhm7/nd7HT7S0etZGxPS374A10C3npze9eIwoHz2fm
DoIafWcofqiYBTOjoIu2VQfkzIvqzW4Z+ryJRmntLmSkvzrtaIB1lkLKfUMzelBd
2NoDecxUWx8Lh4dFVL1OykaKw7+XoKgQ8R300gPK1NZ5ZL34Fj3MUsYIRyZ1PrHE
gIutaucY0nRw1OMxnmnBfiZCtAg55VIDsAmLJgcT18qenRPbiw3GkUbXgl5kLdRV
rMBEExLK7q/C1Yj9pr1mZbbGA77t4KHFYDqsSDZbPosAA4aKdZYHo4mXaiGrFFgs
xX0s8jlzKcS6O8aFktpl/8tGPCETyb1bxrvvuTtZMYlk89WFMeyjuxGPD2oPtzJD
tH+NWdIyw9L+XR4X4IXQG/R9gZDi1ct9MupnDay5vlDDuNkdN7B7CO6exRQXZl/S
OpGcITMQQeEVA12YTGMIyxcrx3ZLABCirrwPoGiUmFqjwfhkPx3V+6WTAH7FcTRQ
98HA6knxv2IU66bmsIgSgZA9UnezoIbZcc8YvId9qft/32hfWZE9GiVKNeIcp020
ycQpzYupVend+/cbnnTFLsbqsAYZg7IZjV5/joUjt9HOKkqrjG2cnC4LpDupLNoP
AjLJ9h1++ufGX0kAd6oJ3ds0jVNTV5k2Yb8V23FtwmvKn1X53m9kIkDnYNhpssYK
zZ0zLUTGkrXdfjXeAuqfdb0cMlePcoGlm2zaInEp0TumoJaJg09Ck1SsyZ1nwlt2
Kh4kbjkvcN4bL5h9Ew704JK6aqN8tc6v1naqfyrjmPcpqLW5utnt5Q5oLXWmz2TB
7Q8PHXARmBM+bskACntJTGK/flZpIj31vbYnJOueUEcKWUQug3Ij2u/gnloAcgld
n8hWVQJ2U5GHsJ/7/608me0ojiK1/xv5U7ItvNdYnsDYhSTmPbf2cwLOT1VK+bYm
zL1x+OJ1GCnKfpO0P19z08i5gRV0UDabMnlI9xr8VEPvaCzjR0KpJJkCHo8ftbPc
jf34waVhiBMhfUu5phG9gmt4/CXtaZzxjyliRnzJcZ6bJQMXjO15vXIQl3RtrBPq
+BnkPfs84DUGFi+l0WB/dDgfpE4a0ZLEGeApCY1Cu7aPw0J6+LLfFnOzLUEgohPX
+6mmVukciDFDty3ph8RNcNXDF5WdP6rXDnMHNjXQZYWAWbUdkvVqm82lgrEtsOiN
WU2F4n6XACVdkCsBRAqVMQbY+pkscfC/teoGZdT2e9fzs7xBloooNT3DKt1QOElZ
fwr2qDgoyZdiau86obgbbW+6YONgisSevm95d522wjJ0swswpkWUIoBfBP/ruQiP
cL8HaZ+S+TR4RBeAYLBkL4RxKElaUkiGwfX0JR9xaXr5CSqYsIFei1uSdUX+vUx8
wH4i/PAcObo8jywQVhRVX/cpp4GUqYVlFgCvfeUDh7eZhZy/KwEQ2tCV8qVhMlKu
6PYkub1H21drgCnKNkqPt9mJz3bauWdvi64z1UwvW68WXKM0en+M/Afp4faHlr1y
ZdrGoQdWx0nt5d3IfCmkeaTYYNCeaUCSblnuu7wra4dlQhHLQbaxUKtCZp6uTHIr
adIKhByxduQlguBnyosGlEXgX3OAy0rpudBa4/ByrpFs2HSlx3PzJ/ZSN+Eb4r59
FfVbMU/wHqImgDZFhm2Nn+2jL89TyPrHJAbEa+7eFOhPF281Rx4941obPut3Yhfa
vn4HwDNljyCvk9x+++Igx9GxJ/q03C+XbL4Y+Y7I/K1ZZvFh+WzBnC9rpwTW0ue7
aYpgv3BMY/cYwmmsBNo8bl8uoGyQmsUwNARk+Gi9hYDefFxO64EDNM07Uy053rdJ
T/gbl+vDkLeP/7BcN3ywiizgmI265m0Pd945SjK8ihFGHHBTxuFu7xgReIjmJoA6
VsZheLJD4PYfc/WKFsVfVfN03asxdRDJxbwNiRgxficJ6XQe2DHgOI19B59ysSti
nvP1WebIO0yvinAxWGi+OJBZFo7mwhjZhTlUbGIMJ22rnpqnbjYPObMHjMWNeAmp
SJWvCLWH3x5VEG4WlwiHyGehJ/OqmyJMvFcUxC1PiO5Vf1jl9H6ewGYFP+WOmcOv
VTnSnrydKk4H8+NlLIriRHwD3o2KbWpOodT17ShTRMs0+zhtErFy3Fho90p44+tY
iWr1E99zSl+ttOY645VgBBD81ppwh6CL/igqVPBy6Ygw89eH0d0/ukXoyd5++KI6
0aQRDJA1TmcgCI7OJCyVi7j9D+Pd/7qkrTDS4QxOcOUBMOlZZNIU9jkIyWnMHc03
x6okJR9pptP/NxZQ/AiVp9U+FrdcAcGDkvbP7brWU55pNNbgrphq+GiXzBBAs4h2
mvfdwxr9xq48YCKbteFyIkYeALW/r7tuRhAp/AswtAIQOD+ZcxzbIXiiHuD/KpKz
PXRwCy62llAihe3eeoYgsrSZYKOLmgG8FfkSklB37mUDiVD+0U5FA+mASl2Wr0UQ
fpyLfhCRS0ZlsBmOpUAQZfFmUw0cDxNze6CeAZMHJMGi9naImsNNVZOKmlx4Ve0m
MJUeT34bFJ12mSXddv2rBbWK9R2T8Vh2UUOYY2Iz9hV2LE9jc744913oIPsXao+c
2jWiuAJSBpUquaAd7N3rqDzglv+tKTU5JC/+wZ2lvvPCovBYuL4QQANz939MgH4k
WnT6Kmo2PSluGz9YrLsSZrmfp5O8rPN7p74ma0ztKUjxRDEhveRfcLs+RiNZkHo5
MMSuQM3gNAALvXxFELXEaHesw0Jh2dlGMGyjssnqIZ0xIqmoDuNCQfbp5a1NmusP
WJ+mQwfP2hXxjy12A8vCt/DUM+Ia3yL0MKTxMgdOGZkV9UzkMI87vdecU9OAJ12v
EmV3rTpbrFRxAHllExnpzMwfPlp2X3/wPZc1V4awWZjoQTQgUhEH0jtn51m+8nyB
lIRJkLN5+ZN7OcFtMpDQoZHsjltX0epQbWsI6lGTkCebUM+vmQfFTYCbelsBQNqR
n0MK15HDJCOSLX/8j0NhBfdVbGAEIkEswtXyafRG3jrtKzTD4AEl0CwK3jPyh+NC
j2e6koaJMgWS9x4aBmcd1yrE6Suz/f/e8NvOV0hVQJ9tcPN4kEWRkXYPZDCT4T58
PPUR6Hu/uAxA/M1Qi1is6bB4luNbwcRsB123jsTzlKu0ypQZsPojON9yTJwWAX5i
VUpHqcg2uWaQI2s7T/IkkOHnzGrnyNEIBOyi619FhTh5GJBt1WmhF9Z0qbkeP/eq
purQT6GQaS/cc51lX6bit067EEdAEMirX3t1+MDP29b2BFQXWWhgq+EklhrKcbor
8nicGj8sIFmt9iEuxaOeGoW29LAezdB22Ecx1D4FsZP0ADzFAvPnDMnKe+lkzqvo
ReyUoLHHdx32BN32DPTW7EDw/WKdzj1yeHb44La31zVZps5Pu0pJlQShPtsSEAEp
eTLjH0MHOOgBCpM+Ydt+bgBP1t2reCKtXiijGFXeeAKJhVdOBlL0k4E86ZccYLMz
2ETx/MWM77AAiw3qZKNFzidWfYewRNdT1zwR5MCVv/4AIUrpn4j/wqhwsRpj+EZO
7ewBeWFrmGWYSprLJHgwt0fMObpiDNV0Zc/w0s0RGZth2S2T9ppmgbr62NwUKC72
Bgw0JPDLA12M024RS4ci0i3jQR6MJTptEKbhQt20YpTkRXv8+W0BBNt6bzZtv71Z
6TqTIWqaANnSVvtG4fDl4QMguP7KjfzXyYA0BUABA5MaTWzNmkRBHd6xw/rWXbhb
9wi4MJFh+cVYM3jIFp3fCgKl0bttI3xe58CQUqw2pFFLcxWBwScifY6uKSCTmeAb
UbcLqYqjWlEVlmofhTkCBVCwIoHT7fwifoW/P4dCkvJSXmVxwzjEEo/h93L00QIT
3ki2q9cKw3p4WJXz8PYwd8enJr78jHKbMtBAudG+MAjdnYUwfSAy1zdhD+0xDnhd
2cevmUJB60TB9hhIaZAWdeeajcaIbNmIYsjwsIP9g6gIBJCem/DZL/k8X+2usg3u
E+KetSrbJntTkN8+MQVJSroH2e91eQwUIxDq/+aj0kNw60Gr1aDNuP1xnUU1J55n
Qp4gCyvydZyGk/HG3nHSrt9LFYNUhSlajWnY63LNcssqRATQiwFMcLFUnFxMEePT
NMN5lr1tsOuUdjjayxx059T8stSLWhjw0eraFzog7bwjLxTcgxf61ZUW8WIctoh9
jsRCm/iLjqk9WHRbEZUo2pO2XPu9iQ4C1BlOvhKKm/6HKWmYildSWm8ijFQ8R0Ef
iNGRO3ai9mlA93kXtDuSbkFDbs+9c/zt1xjygE5bAhhK1m+OwM5DoEbBRDR/BonX
HEPb72hazncM8e4vijZPgdDlSUBmbbhgYFYuh+A5tJrzCxiS7q7HFqjltxpJyGZD
YdOXs2pggUUhbRWAxRywm5TRPLjZDthL5U7zczkPINItVnCdXBc2Ejt5XaRXcBT9
gjWQynTCqtdkIN5J50EbeUlpSYCcvNVmTa4tvccmgfE50fCY/LCLTx+4VT13FXEv
erZh5+hqHPzfDhCh4BupC17ryf2UIIXUTPi9Sj8G8+LHoqhb11GRgAtpEJtMVfVQ
Xk9uNTr3JmJaqIwSwOlsZQCE+ejQf2M0h40F5FzKAAMv5Wehs/aNOaPMYu2iwnZ4
3UrfdenuEiwlH4phYR2qPfPE+cUtaNqmNY8NQiMiGrLLZPSi8UmHIMHgEd78pTnJ
dQU2f0bhYt1L5aM76qp0Z4QCNv+akX4LjRVcJB4FyRATBY5xnd1FVPr5KQhLmSkI
NWMY9PVVQpENfE3OGdp4ZhFF7rbM7c4tR279yfSncNtnGXnVKs208fXJ5JFkvCiX
DYmDz0+DSLcgqgU/E/cQgcmzPPLy3cAPAhISLyvBXbYlwwhztDlTcQc7Iwv61JSc
gd3mzeoO2ts1yBnfbeui8KejOTqRDFveni4Wq7eF8J9cR7Lhfg19GXckN/WK5IR6
dg2/mmgRiyewfRl+1+Pntv/KQRV6pKRtFXdk/KmiQVzf5gvfBVTObN27OnTAjHFp
bI+sp6txIiueyK4pYvMv12CaCwzp2q+VZbpTfTDktc4tXmXnG+Dq4jbjcG6E/l03
itzKZLbUUiSny3F4aV1OvCKo2hXdDVznqtzEfNgUn314behTBHVHzMWoaJxitnRC
gjF0nfo80Owuhhx5WQXggBZIXFztAHgBclRYwnnT7raws67ehUnI0f/5Kws5jXCG
odVq4dTn1AOtEgyY9FptpdpgbjYaKJeD4uWIqClx15G7yZRHz27lg4QR7BpQWmxv
qQblfn9JBl4N1Qj/DS6nQNU93SuopQFY7RB7CI1RwIjSfNU1gDteJFbQkNKN4mc5
U5iNLPm0envpJGVbHhrOJiuaVY97xOl/YO7PXDUKkC5LIxPevUbaJpL8qMJyMCwz
c0YvswFulADkkBbOb3uGOT9jCoRUhlY703YaGM0E6t8Zf1fQVQSkvF5jAQr6RIAy
hwLwAfl8wp7+1jtybXMDXLn5ig8y8HiPO9BpvmqOAH0oy4NxH/tXJXLcBdKA4t6m
dpD+dQrn8dxYzQjuhmOTdu9oJI5pHEN6nqtO2jpX7qvNioufzTFMsKPMB3jFjhjY
3BDTn5UizgrQCH4DpYKL+B1+KcQKx0W+y3LVIVEdIFDkgAXdd6q8wbXOh1Go7wu0
F5So/Rs7AXOmMypQuSz/D02vH1ZjaBAYhMWTzEBRk+Ic15znBYW3SaSZpReL0hxK
qdrN7uo7dIhFuGRVdjFb018WFMsaAExQLyq6126MQ0LPP1e8/sgmVghEVefzwHpF
2/jx+70hXyIwY61q2wjDGRnlEz4mDdRs8MFiOHJ+zceNwhDYbQcWPmV+BZMMnbOA
2fHlzlhu8oRAyFS8wOkLq92c1RxrU0vTu7XTaBsXMTT8aHOiK6KgvsaBeUbmHHJ3
5X27SJKEM7KI+NPft13Ti/LwdF90rF63c2EDbg7EGmiLTHApfa7/bBlN/joD81CY
aE6EY/B7mwxwox+hP39vzaCpQsAz6P0VbBn487vZcXE69sWs3iXga7blpJ7rQHwl
6NoQlEh6OHxe5PGOaK4h2nsMu8JHR6ju0SGsMGEA5oXY5nquM+0b5qsdIqqy5XGU
jJicJ3Ye/g6+PR0JvpCeuX1f5ivbSJQeZwPUXRvpGHr1JxO6+hFFDYnY9e6JVX/U
XEcqnWq8cNLjV3GBfrK/3qpB1mPkv6CAHNwwyG+FnVJeHp4P5hrdqVx+AoyXKvhQ
lH8AQKI2EI+MtDL1dCuGwXJcYjbh+L/W5OEYRm/QPcGY5KV6A4dHhgUFcW3uzewZ
Rv2cjjaDEmgIO6x2CrqP4GJd7wqsTb9Jscw1pi088l7XY6te0vGQRhxfpO3cdI/m
Vk8IEDss7d5q4sL72yLrchdlJpNRxkYF6KUfeLvHY2RG4Ddoz/CbvMd7NZnvSnTT
HTmeJviu0RN6Yp3y5shhuYqctghxQw0ucuNnWn9U+rT9085xKf9guZ5XMWWiA+b1
VbDFAq5P/n4i8TTgQaSlQiORTEREz0KbgAHxxqc42rW2XAhCmL+k8ncf47wVzdes
3WnO9stTQgDjTaF5h8kZHr04YSgRDkaiBhGaVpqS54gtsxKgaEqmF8WTIEkgnZJ2
jpczTBDVm59A25Nt2D6gLHchLR3DbzuofWpibFMiqV9rYjNSNyaQnzQHt95coOkZ
rRpNseUYvmPop+nmh0YivIWQGtI9KY85inCpthPjLd3zDEyjDRWWl/t+2C2o7nYh
IrfD7Ufq1moNxBPYgLVnTLF5lTIlqmLMNwLpqEYh3Ko+LvoUq76/BiaKkC8abfF5
qDlB+ra2Ns/v7NM/L+5fRRoReO6LYv3fGaA7AY6L8gk5+Qff+ja5kBT+pHOwDdBb
4soH7GLz7nfecsXB1PcmMt0drLQjQIIVYXiJzzZi+l+tbOoNDrcyoPnHF5vEWiZH
1UzO0lSSnCIcMpDyIls5vXX803Uz8wYIMTon2kgtLdVkmywxtVqOp2jAbHs8IwL0
KN6MpOQBm8GednEgfWzg61zQLOFQLVZmD8wlHPDDuRiK6QTIZN9IY+/Cs1wQTNwR
EEvDhmLkDFpyLjwupT1gQQ7AwuN2U+jlbDLhzp5JQS91MVENAhpLgElchC4cNLlN
eA7e4at/Ssbufu2z83VEB/v1yW2xtbtj10U9v2X70C168TNBrZdsTuln+i7dmine
NQ8rLzu7z8PpYbZiGAssLEyM3rfvvwkBHYyQ4cfoZ3hAhIyWmiz4UG5XpHI0QwM8
pdz9H8go1WSLbgZhywpI/B9HYIZn21A6UbGxUWYnaNCJvLte09LDymsyxrLRE5FN
diiEZ8o0I8ww6o4RbalQGf3uFvQE+G/y6Y6hC25SSHr+xl6eeExgc7WSILxgeKlq
pirWUbvaM2GgdA9nIQf5YYNweTR8DlGK3JfNVcLnNjNT3zcZuH4VHZPHUVtC9UnB
UDhTqtnv3Ni4IqXtkPuZOaCzLHML9kiUBeumvAq4UqjE1+ehCwaeh+3ZQOvObuI0
JtROAXERjkflxUOlPqUzT7H0rWAtTttmNj5J7RtJ2zms+dXId1ZPyD+LJqFSVcGk
kMsLXRo4ZLj8K/PH8qaWf8h6CD9cN44OU3XG+57d1L+YCx04jMPMnPFHFeXrCops
/xq35seeOiW1GC17+3V1XuSCliTUHmedpMy9uq57w4GHr6hiHDOhpEQmRNwmyLFR
ue7aDUlWA9mIQVdWtv+HU1kliJiDt/1r+9Is7suVSPdMwd9mgVAzxkkHJjjPYS+g
j+9E+/QF9vIj38NnLiJk8RO74d2xWnAZMFECVlwb8bBGI9FyyzjHlWMtCtZphMx7
6UrAwt5MdrtG2SY9LMAN/jHZcB7Md7V0ZKBMoVAjbhnHIDydjF8D+AZhTKOO268T
ziU+k/A54v4/yQS539ebogqE8/uQiVAcYJSZYdbQfdzXJWFoldcsm++qCvwcgLbb
QZxxqlcnjcQMWUjanUGI3NK+vxqhWWXq7CsGDkvKwPiVQx/K4WOQmsnQJ+c6iHyd
PWRrRC3uRYMD/FKRSF72+ZPWG413zCCPFCL8HYng+iD531QuKGp6fconEQuun1uv
f0ubPB1kTZJp2MKF6xlmjf84dX7bTivMbQHGaZ05+6BWNN0j6lwqQrRPLyxsoOcP
1/Ob6g7r/FTbU91WGmlwCbkwMtktKAtrKOMezvbYdCVCJScNvsgHUNheF3Fm1BWs
nvSlhRESAK8HkPbvHtXmqa9lPn1dA2j80xv11zFeyv/J/bLVH+Wsu73Au3oTh0q1
nPtd92hnkTU+RdkkGASRGi5YPunuVkWH+x+XfYC1NxJGO406h9G1l6CH5V4suHAa
C96hD/n7EgsZJP8o4f8gwHeueeOQKRhC9MUCdvCarMbS+Wrau8S8NJmyEg+BKCrq
kE0Ov4r0SqB57Ndg6WfVWLD4fELzJVrhHp3P3xw7GSzse26oTV4496zruYQ50i4R
IK/PCDQVVLG8uTTAKCaOnBcta5DDaXU3fl0p8R7EpOzvHdjFcdQFrebADNszGYCr
QMTulODDrBBGfzNgAkAcvLzKWFJitADHNVvhHgAKZLujY1V9NkK0MUKY4AonSW4Z
K6YO+GWaSSVVg+5ZbHfzcZaHJPIpufir4TbX0vBAx6mdmdFSQ6A8VnR6BDWV/DlP
jqcMGfzkTFPlGHEwd9jORccLJo0VpBA/hn8zpRcQV3SK0/3Q1dNXtpE+OKAv6j3d
kGYWwJ8B97bTYoY4M6StIPm9NHZU8g8nngcKor6Dwpj8EHhNC71g17sLPbs4S1Gc
Go2ywFur+wz907W0OirjX7axnH12n1b1zuorclVTAAgaiuxmvUQXTqjd6JgPLNlG
K7ZRw9HuDRcOLRNkVEbVeOD7DfEM7aQ7XVo4Z0vht+NEvg8bTJVtjxFAUgkNL3Z7
9W53OsDo2LJAiN/e484zQ2MJ0xjRTcvo36MX9KCjDC6vyHevUBKZH83H4ekuJcR/
YwkvlX4q+2ya/gE9+mDG3HxZr25HP9f0vo/gd/H/YMdqnXDdcV2cWKCvbi2Dt++m
MBcWYyOLaGMPqkFj58e9H+4tyqmzLCZ7wxZkRoc3Hcs3nyrfKxDhJQBxnsWZfnhj
3o+MhCoUR7sDI14+VPZwdWF6RB/S31WMRGvZSHYH/pwYSy/coWQeS+aHruQYAlQk
xgUte+iW+Q/CwL53xS394FcQlnWmw50b48AkTIT6T35CblRLBp0G7foM8LWpqYyo
J9/TjP5BWWVwcW8JJTqMWa8tzm0NYS/MA2AIjc1kR4kPHFiWvxmtU3ekoYH6VbsR
HyNleFjdhxh88zDwE91KWkqptVijPLFh2aCgX+jpmdZ+YRVrK0rTDfc3l6FgiAsM
FsFOOOZ1McySqyw3vFcyNrkSo5X85oiqizvMpntr6W1aYIJKNg6cba5YCaimw/WO
iEF2IN1ldb0ZAsDqnLwzl1sDMzi5Paf3eMhvGVkNekrpUnD0q9HJBtV/1RVtKN+s
nUj5xMvYnWm5h0bLhmC/Mbr7fWFIzHyxJetcKoVclFaa4sY2JJF7PTuKr6w3T3lv
XEqlVrgby4V/mMDMjdife/s30xxhVev46rWr6UAr/Z3GhAloiyq/z8S5RJrvyadn
2xxVP915VE5GFJqsicEZQMnnVmBb3BdEduqYIxMsx+rVy22PTpNEDMjuJLOVCYCi
yPTOEmSYSLHdR6gnbAgCDdyfGvCGLhcfSbdA8QtU5VIZgKsl0XDtRxuVmSjb2jEI
96zMbPtBBQX3rrT8OaytB2CIgaibspOcoIwmMxKf/n8P061i5tuu7VNRcpMr/Yh/
ogJlrSckO32bWfb9iiMyCTLSGaMMXyhoJ7i4gvW2zSYo+8DQN4PhWHNkWa4+kItw
k/F5AA+yJWqaFGbgyS2MoCYQQY1jqbEm4zNLK8degR3cQNchBAwvTYOnJgdRqwoE
mMUaielZJtf+99dof2ddJHLEFpnKe8jXwHhze+qtiU+GMsgFgywvwJkk9Ncu4mz2
WNL63XgO70Wi+AqnKb8Qamn/OwQOMdcR9F6mKCl1Anj+0JqqwfSNyLVdJG03CPGd
2v/ETB4CpqG4hry8NnCPBaSoryGtuNaeM2QyLtfUMmoSM8V3vUPPyPFPN3ak93Dp
Cwtr3QoYbQ+60z2guN9g+8XpFHF5bjEc8Ys69ScX6mCd3T3uZGu/Mn+/hUnPh+K1
p0Qao/OUIXAnsdBUYdhfai7ao1/5VwTiY5K9ZC7ZSPm/8DPz1HLcWnBuUKmhLTuR
fV9+YRzUZ3Rhlk3SyV3cT3dUrXXPn0/+hRH9H1y0PoLGJFC0+eLHkHinO/GZqLG7
xFmCa0IyBiKNZ+pozCuXcshRmPdNYC4OE7aIYes5DIoHNLnL0nJFfw7cYVScyXyx
1srL2YVdkX9fhNx1YXajhGpo8lYh0Jys6/kQ5F30EIqkemZWfewhH2Fl1fpMe8CD
Akuld3N2WpvI69f9wVx/DYzRVent/rytTCcx7mk9vhQZKRESe/1n7h5CdvoAqc6C
e9zN1Kg7dXHcu3fz8c2iuU8AbbU++RMXUNbCj9PG7liWdGa1j40Ta4/Sv75I4A5t
MyrhYaBvQ33yM+M0hwofSl1WNjCFMif26L0DZy3kpzKQEHY229fcJF/B+9a2Kv8p
FhJ3smVppwweVySBLK5wTcFt8XV3rwKGoNCU84ij9uleImCqw2G7Y11wn7NFk519
JPjZrM3f5o/yuczTHx39rTZTxeSSKZUFx9VZBLjfu20jXd9gDMMQrGgJOlVuq+b4
HnI25ObktKxseFZaB09EE9usUVqoTvY4cOzUgBZQ8V+fRTtUxsvHDjFG7P1iK4OX
jJO8xPeS7RSSTevfp5uqhzIyDWlIpGzuC7zP7KOS6OOX0OLR3b9+WhMn0jtNhAPb
12KfVGgn3JmcK5gPgKLOYBW5qcLXCwzIwgLZGGfj5rEbVQmyGLJ1mMVMh6nvFr33
SiZSjbMrRMhPej17nfHJlg3DkH1gXfdzIz8qYyzoMOPuLLMi1+w1n6IwlA5BiIeG
Do1hHxOmT9ZFzWFdvOwgP1xWPDscvVzO0Do/a2bVu+AaB9G1AxdumYnM4oeyrb/7
RBrd96aHRIFw4p7vdiWc8KdFBHt0tMC+8DpsewBBeZB4nube3c9EfSuKLpg/01N5
acnQKCKZbGfEHyRnAt7KJ7UJS2gi859foyLMxQd+GwEfFs7wbp2cwhCbbpmZomw0
oICH/QPkNZrqAGF8eDKIFK/xjyPG7Rhngi8alM8oRsledJOY+DOIT7iHtnR+sFXf
QehXHw0Ag13QAUOQIITfbrwyM9Olgwwb19KZdbNzq2uyL3MKMqTlo/AGT2MmK4CP
SuQxQiQznoZEJmGv10xwc3eJ1xwBug9tUDQ+GR0VF0usJlJb8MKWuvHynYZU7nHu
F5aZBjZGCxwkmR5bs/z/3vs22gv3ShwQwgUsL0zmz0D8ubRRrs2aZwKDjzkMNIq6
EVXHMfIC0/02Y7vAn+3WxQC6WN/8P8wNm+exMinPm7Xul4PWlHqcLlVv4ywLUTON
uJjksbDnopIcevc1kmFgzgB4F9V9rZhQQYavixK4f+OSRerXTA6KPf1wUIjCTzPv
3+lU2P2wO6sDDpuTlI+OeG5EEpDMxpITSpcQTFtaY+iY3h19ZRPY4/RpKY0ySesB
SDPFTb4SmzDV2LI+tsmGVQ7brJ5rfb7EIjpjaroT6bPw0eVnJDVNSC43lwdxeLE1
co8d2NFG2a5aQF9kJCZMJirpr1gk3xtQQEPUnIU2FfU7wWoeqqVDjfKFZmNOyGfO
a/3pDoLlozScTE6Kw7Pej7WveNvkybTm1yP61AlsqzQNFZGKz3w7sqjjbkeGPQUZ
Iv0KiwZRmU4EqXmNwIp3xE18dZc9zfOSiV8Lk8fCk6UquZkBFYWJRA0Em5rEkmRt
AsPfxgzwjeZCGrIvy6KAie27LM96ALqcer3Bk93xF9tr0cn+tjkSOE7+0eQwlzQi
IDBKEdptG5MKl/uFiQBkPixyvRC0xYI4ewpR11gKER5LddE2WNWDdPwL8Ak5TaKA
cizLUC6kiZbId3+TQroKgvoSblomB2wMGq288SRouqjwfCvKiuY4so6UaBvmX+FS
j73M89GAAY5x47uy8c5y+/N/wItMXBNcCj6blHJSDDY0jmJJ0ja1MBRepW4UruC8
Lk6PyA5PU8fuAFtH6bw2ZNflKapatSP95tpMoHgeLw6+CZ1s0PzrHQrXMdIx+DxH
oCI4cih6a3R+0OkFlH6nMs1h9e5SEXKeUGmbic/6A10cIOC7ZDAVCJmSOCsleNNd
Mo3O5pXbAY9tcfQPuEZIg5Ausk2ir5fF8uTMECAUzc/8Fymk72n+9MjeLQrWD1lD
zGh/Lk7ff4qnZOkUreCATSaI7T2GoKKduGPcsvoGGfo541qz2Rd17hoyya0y5X+G
KXEpNQBEV7LKLDytVSsy0Euyjmm+pynP790zHoK1qL3Skrz9XRyW0B6O7iQTBVzc
g2VHQD/yi8c5zWILz+8lOQapNsYNEXuzBzRau/tOhiHj71pCze+1KmN3gkVEbSIj
iO6iqngWFLsBPB2EIMGj27ryVRAK6BwIm1uXDenS2I0WTPzdZEgY6ymfOfuzS4Ne
qbVZXhtVFf7DBt0GEjEAHDRZd4+3cGcWU0eOrJ4xGIRBqpXDkloRegADCWQ+1lhk
pMfj1WfbL5semhpncXKyBKUXjXTq4h/wlUcfp44GDSVcK2DyzYzfuCAUpajsCHiu
/nyXWDH8LcjDb6u1ZeL1pP1LuvlyN5K7Bu2wXaGrQSDtrYb0GX/SWkJ/pz8wGFBL
qwN2Fa1J0QygsOa26OnByqNhdAlfH8+UaWxbFp2bETE+A63jFVwIUsNipoDBI1Go
OgoI5k4b+SC1ANnC1nvvtAG3boxHnZllhAzSeDxeUJ0U7PyOUQjvWHG/VuJv7uIA
vxR118J4/RixEg/eBtU0GQLCLTaNEe7IPZyqsgb8ngDCbUDvhr37hsFQ4r3vufNM
ZSdpmAdfebbLLhC1Q7Y6oumzavH0asBbz9ZXjd+tYZtmY19EQtDr2l1BsyEJKa2z
4M9P+cG6wtesmIE30huguLvUHW60apmQ8StZrhXFJl0qur+kubrwsiZu9qhSUCX8
iKyWHGRcqOmQPraHWJKzYRzM6oILgq0yeSsluwL0FRF5FAGZMeeMQKZIPua6Es2i
/t5+Lx6q+T0lLjp/vmw5hbKGSqvH7Vbgw5ML5s+75eVbWIb8RakbcHb5Dq4fLX3h
qygHZDEvZQf222USppdhUuJyu1pvIWuWBHULJm1c1S3BmmuelD/igtHy9/TgoDtv
nOmJYXgxAr6VNGL9I3Mqz3qBHwTvsEzdxqSd8A/bNh3tqPfv2w0hnLptWvJWq5WR
DEUhSmNwQMr2RoPJ/agCEeiDTgS+9BIXnpWfgcvKWnsHx+jNkEy07NkcoDUXy0J2
7IImDXVc3qjOQokkg1RtMS+ovnLQkHP3LG7kHchZt3hbQeYyygHnycDN4+Bsp5B/
/jC7WvG7S6ZUVBKh8sHuShOsvKX2MaUkXDoDiSwV6ybDFWzviLVQj9x6e/iZUBuQ
+k8Gt/+SqYEiHY63MTv0SlrrtmGg21hM1eiBUsCLdmWZzbdakdMOScneZBVs0M1S
ly9INxpbnHHfRJuScu0aw9KHhbovOiK6rgjfjhgVn4UaQUIghfIveLYgQTi4Yu1q
iWN65Ml7Qy4oJfROtAzBUv70YU6S9aiIjREMAf7K42A7ppbbnwlKlcnScto6ys9I
cJhcllpbVtLmz5ukg2V+L3MSmf1g+ReVJRKH7blwzUMDHuYFyIAc2xRHw68cV2pE
C8VXbv1T9+rKzq1XS1jcjNwME0cZGYW/vc+uo17T/XSqh+Ol5GYjADLaorC1W+EI
OqfOFnlI+ZgzDRPF33Wf3jNFjvZQkFZJ5LX4toTb01B2pM0qbOBPOSLFX5Pdz6DD
KoYaghrR3joWtd/6gZaWcNesJt4wPMXeCxGEwReGwWGf6w7oDN+fhkuhnu9E8NDd
mpWer37YMZekHpc2KAHNRUNwVBSe3+5h21qRFP0j7Bt0NxkuiC0qCWZHvlrqpn/D
Ncn4sRLccDOJf9JXFtlmDp0dRuTB18+EzkjNkbBj2By2rYIyXld8GRtSna24gtn9
3bQNOzw1l+uiTiPy5gaEsQe/276tlgvdm93/6qe1GOvqIKZiQ0EWxvil+/jz++eG
JFbkDjplQxKCkgEWdBQmJs0LDfoblrnXoxDVN/xdBDnFWylI0cGM42ghSDtmFuJ7
gRPzOEPiVjzVTyYFlRqTcKKHDeifiWBqlfTbrPQV61PC17wHH3rPbyZuKLJGxHEa
u227ofPrmIqW8z3FzyqZ+hjr+tCN0ysYvYFLkDu8lbxvfv5wgrcGuUc35FcD2Ztv
O9l5Nt67x+PRh03DiNVpzukL696ae3UpCnZyAbJw4Io7xFfnFCc8Z3V3dc9bCh+Y
spW2eQfMOgPkcZAeA72bzdkvuFQlBYj6a/5FUxUEEt+2CVI9om7sh2D/Qe/yc5i7
MPblYEIXXgwvT3UE6e2GAa9utEBe4QvpyfV00mKimxdW+R/s7cSmk4KSWUxXKxOW
W9YHCAcqs6hhyNSq5SaI9VFjmydobA1yhdUEowcaEYsUr/TDSRt3Ft4m8NvJahND
W7DgvACfQLVGyNaBnarklrkI3NR4VV6ImZGys4nSs9a5E4g+XqOOFh+5b15S8XYa
ESdEWZEZs66/CfymNbGGoDk41eQDT/JwxMyPKWkhJ8FjltOHyPlB2lHKVbT3BDis
ta1NJzv3xF545GVArse5tfE/M6MWga7jOskRZmvLnWODki3l+jR39WbZqTEwKLh+
e3MwDh0FILFwE3zqjIBJFpib++9pxMs5AY86+2Gdy+x/ELTQtMIRpQ1oWtCkOjpj
ivTLZWnp+pn48L9Icz6f50+9TnVXa4yqEFgHmxNcIJ5eTxHHKdGhujm3XiKeKmT2
UwN+AliAQxE7igJWmTbrYWmkbaH3t/hcgLVvrAepT3gaq5+9smbKzGmGwcXH4jIj
LtvWR/RbVd2D1wsCwfOGHXP7iGkTbrPlzPf2BsxM6dZ03QoGrE3B5TGeifhNx6mV
26MUQnU4IeLnmP/sn/b+hK8JAKwrUca3ShptZgsn2aLs0fe9GEEb7jGZuGvuWGZ+
Taq38FaZxqoOFKOvh5QB4mN/pYXvvGVAfg28tDmdtudxPGBSjTtbbPaEmGjLPmfH
w/rnx/yrpxxRJR3NzI+2KO7Jt6Hzgz+ot7RDv42gnv+pagWv10XIVp/I6P2KEGUi
AXhJ0V6PA0UiJTp74ywrUEmaHDPVerdqYPXv90o0ltbDFsHC+k4PmWQNggSkoaqi
G7Hmcknk+8C04dRGQYn7jnEgUU8TO/wRVc3BAZWdck0mshhkxXhQ9PYqCyBK9rnQ
m5SOGAPomU2yuypccv4Yb+qRhXkmGnJd5xfaVaX4eUIpIU+VMBVSZXJavTRXGjpn
W1S8tGeZH0MfX6lfwtTvuH086nHeGY+bAGXLUdyW2B/DoUpVl6uGcFtiEfNxTdkB
a9NOG2timcecsf8PMiop2v9tYPTSC2+6yU/tkYzOUjduVyaxqV8fpEjKAzBbUOxA
zFxs7a8BGIG8wPrF/mFj6Jf04ljrRq73pq+mJFRZ8cwFRs2yneYu8XhyI+ohmtbD
q/GrYJG0wGK91RxhDT+dBXKIlQjNiD3e0d4bEBnawJ68HOmIwmtZxQZ2EFWQ8WKX
oiNLkYPNauSAXyY9kJTpvhi4SgIzoJbQVmqYVfoeL/DJ6Ii8KKHSVHn8oaXkP4O6
wmbmExuzSNt/bTQJFNaWa4nI6XF14WQdBDD+FQ7CXW11DlBRS/liZpzjX3ZiXF7f
7EV7ZzDyHtdVe9ExKTg96TXA5mrguG+05ftNA7EvxgKofbcrTh5ZYuQdKAKg9/tc
pp51mN4iNIWJhnNZEg68M+a30wxaCifXyZ7yimpErhY7P4wCJAJEcFmJ+8vxGVyi
q00RaAetaSNBhyqT02h9yNZrcHB5zto/t27aQTGnTtgSAiBCwggUZ3nRdZvONQfM
ALemvSB+ai7pwGKf0gatWBvqmPQkIpGrCndGT81+8HXRgzQfXghHFIHMSRDnV3Fx
IcL80vihJ7ucVJZjiZ8cjfF+zJIiKOh7Q0in8SgpDQRmSnQ956KcHZjH/ONC4CoD
S828/9sGr5MrYkfygkMM/iUjH2Ij0tdq4aw7GQwPy1Xbsgw6CUW8Xa0avqVrg6u2
TDWAC7Z/L1iVpPk4mmy9plMpG4R0Mvx0D8z42fQhyihQCugt0riYzbHY2U5TuZe8
KGR9Sa8HwVri1SW/RrYt/ye28JQsL2pIAlaafybvk767n0BHggPFd6UmxGgmGqKY
tD26doWlI+MjFGgc6z/t17G6PYh/vwWRRAuHxGXfVMpNF9/tIQ20zPDvFJOcFzPq
PREJYk6Hf6No+OM5Fy/EIJ9mOGKFxsK1FyPvjcBWE6AI03VIqyhIMKfP2b8HyzG6
tt21egQxzsCGnxNzDd+OnFFTqfFfoEWMGjWEacm/aYve/Kw/yYWCTStAU1MVRz6o
TVl6NWksOCkRiurpxddkrFYAJLvyA4lLS7CNa+dL8B+2k9jizlNQNCoNE2mFI9TS
gGRMMnPUQ/8HakyG7Ro9SdHjcSm/6WxVGDwaBBTJ5uJdv8nnrA3/Ft0L5+t1rM+N
v4NgC07SAG5mv3vWmQLf9cXX0tj92ZARjxzzm7xtijFVhR/noLKOKaf6bVrBh19u
uFLw+qIX+JP422km3pQFBPt9GIVFJOfcAa+6Uj1uSdKxUrVYyqfkUFvr0ZSs7Ogm
ee+E8w5zFaIeAZdRaMIRvNSUDyFMOH/D+N+Cv6IyzwM59EgaXpBqbEVclwhck2yv
h6Jj1vc+srA0B2LW0FIXSo6fHzrN/lcifXm7OQCIb2IgTo4gwIOetUeFgOhcj6NR
1sDBgHbAgxbIx0ZHH985ZV76rmlLWpmgFyHqrw35sPjHppJJKmvOVLe9wtMaXmAo
novL7EqizXm9RNaQMNw1VzEx6r4w+W1HV78FYrnkltDE1u5uInjVk6NBHogcj8g9
qiB/yWG0njO2FxesloHCbhHTAPrBYfGDVX9bZ4m3EebLKFUdCrgrt4IRakgXOjCE
3P6yhird9m2Y7YH4VCiLcxPeAw7Y17CIj4xnk8UbG5CEWizeYHVg94AGFww+TBY1
if34f04UQwgWtTJy8f9hQaqh6isJM6ePEnhYoAUl1726fCL3aJ+lPXs6LwOViQzV
qy0AuyWa6WV6xjCWII7fWdlwsMXrBNK7BANO6aToT5ZSr+viLJh/s7vM1M4iJE54
uFz3Z1ZsQd/UWSUvzBkVEivIjemPBCGNijoRXF52t51EGuAabTpOYOVxYMO2UNwQ
HlRBGWzcKZa0HDN7fylTvxI8xacOLza/nTuH+6gbdWNOllSEmtto++ZYheSTjV/n
Rau4Y8I5So2K3H18xhgqGfLkx8saNgyZIxcV0rWcgyFgRgNfuvEx1ra26Abq7xGV
g5kIpMnMz/NUV5D2YRcHqUs/gWdHCXWmuaRcVskRNDBKJNBVL5NdsB2SjXHGSEWZ
j6JcloxM+K+QxfuHfM9FidrpGvt+ynmJDBjpSsgo/+R9g/w0iIqSRAG+xlSbjdig
Ohj7yLrB3AUUHfF6fpASUezdpM49cpRw/b1oFP65fhyAzrsrrrBLqXmPsh6bIk2m
taUK3hh+dIBtMGC5QBrvNGP7fX1QJJ27bFX7U41hFXEkcmrt3JNSbhoOHg0bWMUL
PDSqPjGYKokjr8H1jGlpKw+qNIZnsfMwm67C/WGGOfzJATPkRHATwz4D7k2m9Nhz
56bidr0Ms4X7Xlj/abPLiJqX9NZnJOSAlBBZ1PyFyC6Y944TBfhQ0rwTc8ZE/Kgq
uTh+2K9KbOraQNxD0EUlXp+kVL88h6RfKquh995C3daeIDwV9D+VL/k6v6s3EZgy
+/zFbkwBXByGLkMIeAtw5JxTAt3NCbd+67i2gcxoRc0nhYhKjmDo1ZCGIefgNAdp
W74wky550abmVaaq1ExQi+nj8CHSbfUkO6mJtngVulGwUzvB1Ic6WcBqGDBb5C9m
fsGU01Vc6LU55pyJQX/BsDTUNrHIoF8h3i8yL40wwNijVdzd0p5uyj10M4cr9gpa
RRj7HG3hqfBDaCtLUYeqil2HNN6HT7k0b9Bnq7dBzPIEWstcPKnEIc56nLOXvILo
4Umkg4/7GIOlv4QYjoqDGk0B9REm2jUmuo6iGMheBGaV4MORaBHkposc4YUpCoKC
CxER9jPW9StseXsTsKio1ij8wJV3OZTpNrzVH9gSaS4NtyV+ZtRs8Wsj3/cBqP1T
TXhA/V1ETXE/B4Yq1PPm0Q0pTY3PDTSnLQu77fwRfFz+F+pDn3nPgi32U7sWZadb
UDdfFfbu17NPDNAB1hDa8yDGMwrE7mUQ/0pXyyAUEOuWHAGMKqTzY8NkZLg5DMq8
mwExFAWU7mqHRmASMmegWmigejJwFhNpC1swdV6nSMOcdikK8H7cpBhe6t4Hz9T7
1ZEjZlEWnch1e310xtwx6fC2lwjegWA0oKR9+ONvAzkiRe2ogfdi/9jcd9I2B+mW
8mazOMdyrHmJo+cQEMewHxO6QWJ0ss3YhNJhHbwh+F3SOP7jZ7PaPVYMlwbVXW+c
mkgkTECR0vM0/6x0PQWAf1tkwcm06u29oy/EpFnFkrZQIHAbmp8372AVGJPo8r/d
fnXhT+DfHbeVUnDUmpenWn3PZ9v90S/N6xfHKEmKzDiXCYxl0Xa6pHkDwva3sPTT
Zkov99IQqZ+nsmfbOX1QmJUZ7BdWd3HwkAI8T5iAfKjVQVVWGNv7kfkF2yqOn1Za
VfJxxacu1YEgbmbqBFJuKwFWhIqgblsy0v95ayVXEViFbi4GUsrhX2hjEck4PIDZ
/p322QY74oJ2UNqsUEaWvAvFXxGPshU6c3Nm4Xee6n5FOky7A+yLkDerZd5SPG9Z
lUtIE1Rt746Guh18a3vHfStXA7Na+0nN2w4K47vVXehoqONT8Auy4vDSysL7XFwC
PC8dcKhk54i4ztW677D/vpolgGtgpJYZCoD3rNJgp+5fZ5bZcfY7cWCr/zl8Pf1R
7GLg2zuh9zDOKWKeBkqTiKQnSNokrKEMoCJzPzJqHYIxpBbU34qz7BGML3Q5oXL4
7i4SrEn8n5Q2JBtOE/TDAGfXe20KRWb3ucItrT5SxrvXSA5HGQYSDCl88r4+vwql
agAfmwCP532+G9/myELcXYdYFLOSEeCIZWM1/Qcno545e87mUwV9gQ2Rs504IhQN
9u3WIHt3DRJsD98oQeT5N/zepKbKhx9Jga8HNILe/TUKwPZhIor3bi2tgFNqprAK
4YVNDI49oRkiSTkJBoRf6POiMJ8PCwNPOkCVEL4Q8s4/p/KdU+uZWfpxoIB5gBI1
m+P2FAQO1Vdk+g2WzBm3k40mZjcX+j1/zr8QO0zVk7G2FYwvSW/uHzrTq29qUEG4
NwOTw3kKLdEDaqQTLFzpgvLZUpVdx+HAw6FMZCKwAuMqt0+0kWx5GLFIm31WbCFy
seXa+R699M5rA5bO15EZYO+b47Ni10AXwBaJPG5dGLBGSNBVIr/BGUUSFG7qPuyA
7qhHnB63xD0I9ZlE2tDzPzts0THaDX9L9aAhDdon9hwpb4sKMMhr9xVJgzg4XnxP
vCxiISZNDfuKXBG6CodKjNlTa56Hk4roaiNd/zpJjp1EySDozHulEdgbexjI+cNH
UBXu90dj6f0gs6XttRdCKybkFRd65vWM/mrKBCSQFycUbhrQRwamY705/riGAvR2
T4vXDg9yQPpMntBJslEIZmmp+j3iDxtYInypUZX82FpEsoemKz5BUYGCYQ1CfK9Y
AbGZ97ULFYYwPav9elMRZhXax+d+5c9pBPsQTCS60XlfQq7OA598cVN3UGt6+tmq
crPJwtgO0L7c4CpQApwBUIhk2kOTAWv4D0jHxpy5tmJQh6dQXaxr3WjUpyPlmle8
oGHTw69k0Q3h6TQ+3Ekt1lwBgMhDKzZ5tR0TuyhRxZIgQQxLMtRVoB+bw0rxBxYB
8kcnLsXdj9XCl3kOSECLJBvkqb9ig43XaN10icq5dFtQZY6g9fKh7CldQWgCLfBn
3WcT/FJazkodeuJp9Nswb9zKegQcAtCDZiNYCOWh1KNgAPvYTfnaaU5HGEEHUXXE
ftsFwZtzlEd30NTu8v1rEFVVVH5Mx1N1yo88X0PTICLOOAIg8MwK5ReOeo0/rM6i
OrmVJBwGwDqhL/ifOJuoOKyvSLFy/GSS0rwW4WVnFZSl6a4qw9YSWJRW0NJG4Rtn
vtgoEcR0YmuqEOojZCoXhImx+FokkwSAU2NM4ZueQ22G9ctCBqKFNfDI8mq8X7yZ
WCGO6+xeWfTPmMn+ZwSClwHYenMCwX9VdGgqnQ1uJ2X2zpEkMO3bdfubHqOWx/MX
NKvIdGOdLcUNLHdWEQhH3WBOpnpQpKbVTdW5hpIYe6tWVEvvXq+N9Afk2ESLXjfm
ZUv5nv83LDf8uD1ddvwG/iDlElTkl6rM7siVW23xgFQqfXS/dCpd/mrjSTLGmGbX
fOsyt37EkzEK17VZMYNyw+nPwcQWxXWaVVPHRWj8X4gbmr68vVX7q4zWrH1mjO5Y
V+RweJEGr//4c82kYRreR8kXK/5lJZQ4v+wGxZtFg52DLCSm9hmOoPfNvMj+0FmA
o1YJev3kB1LBAn44invjc8z+49E7BF9Wjnc8Sf0mbx7inm/1+6lEolWF3DFgYlt+
OTk0csjhnmVKub/CrkPsqegCHLK9y+jJL0iQsDqKfqOcvN+28FsuLhkb2UWwHRoh
Mzr8kVEJBwoYE8XV8J08hNkitEimXWe1hGD6veJRYsvOvlb/o8NxuhZxSB9ZIx5B
+g7pv/6JdeN8H6Z4jlmXJ7dKxlgq9vCskz4LlVy+wCbqoD/Ky37W2mFTR9CcaHaX
4820nttlFSWLbfGCV+ejI7wsN4FRnz3AA8c4R5G/F3fE+TRA4f3xm4GaElcGSk/8
cinCPP3xnY0CZRxZ50BGLGR1A3PLA4WlwB34t2FwdzZrTpISiiWkaipiCb4bchWy
a8IKSBt56OBjhDztyyqA16eOiKNoLbF0x526OOTeXMuaTvbEfaxzyoLwKUWcdS+R
zk77RX3xekMyO4lskyBwgksXRbaLLQ0JIpmAb9aOlusHBKYVBe8fjHTpDAf5toHA
QZlqkX9N4CmISPVeqwbFNkUbVkiUkiqUVjUgfzq0I7stjs8CjMcuLzwnS1P+eemr
AuC/ouWhEaCs8VDtItgLzMCtuFxz288uyXsW+YYM4KL1/Z3WzfU5ch6YAY8kdroP
mYtjThvoYcAre/o6OSVvOgOn5lIwXPF8+P3JuT4ssmSY1gyP9fyOvMNQAfmXM00z
VsVDGNaK6y6ymH5uCaxq+fiZqdXFQoxNvpp7OuR8Wye01g1YyGlhygFWuUtiqbjL
PEwvhfRj+m/XI1VIW21Gt8tJiVMEJ80ND3/IrZ4uOWHfO7nZCuUl9MGLHdsdW9TX
SsPVAosRYBudoleDS9RDSmB21ONZOPbNoSUA6RZCaSRfE9uZwdU6kulz9dQsHrUb
r6kyCrfM4/0dlwtYk/C+ii02YjSOtB4FqM9uXoIqWO8JdnZBPdFj0Skar++BRNAT
426p6WBiGKWij9rAoxZ4pUYVTbDI2nOvmfCQ7YbuRptCOOhaD6oslbO2/T+NfmgN
xcDbuvWfAX2EOEOxx9Qb7iHVc8Sb766yojd77X7NxHFragqU4EwUV2nXtRl9LdMr
1+hZTt8dC9nLclkl5Vcro6JTfZYmq1k9VVYpr+66WTpWKhsbDI0wAl+5HRZluNtT
MXoBfN8waKkKIjcBKsdLvU4q0d6d2u0RMWM/03e4wmdfmZFf5IzUL6U5HByxC82S
icbEa8l7IkhyH1alF2/xz/uhT+io+JWmlrjgwVrXGsQgi/2QXdow2dk7gECfUrzF
JCrauFYYqtR20hKPz7+l6nMVfOq8POwMlELD5gtfFWXCs/2PatlnYQotT+oO0bdt
Tm+D1LcAyH2pCbwIQxx8e4qRPb5bn2QgHz2y0tmNVbZZQ7jL4SR9jpOqasJ5AZgJ
O7Qe1gFpSjE5HQ44450XU1Vqaeyyh366sd/lvzHJLcZVkdogeINIUXHdWQfKlFm0
lE36UlhhtkUVJ3pOCQf1VE/d4/PsV7VVjpqLTR7XbZXu95UmGJs6bu0qd2m0REeg
tsl/l6Hv0EsSOWI67l8fuFD/bpGjqiF57aBfyLmEpRocdjLbbedEJGdzlOEKaJyc
XtXr4mNtQOxWr5Urz7nYdRobJV7bHpjtvIORcMM2L+1J/syFut6WfKs+9d1K8y1F
aOp6M7fqASl7r7OqoX+PKecvF3Tjyr/jga/FIJA1p9LynOxtroHjtc8g57pxnLqy
BQjxruR+Sr+tR0QGvj5DWGJcYhovBVIk8DpCEyiHuRJpUBlJuDqntUAEZCbjva8I
Uu4IjIrnhjUZIlFSevlAvfo17hGh3y52FVw2KtBGq+pdfc36lHVxRWN/A+MKEHy6
y/8Ixtqj9FRB/hTkKpUK1APnSeImS0nihZsiZZoBv8KTQOqVVTRzuaIA2GrQvgrQ
gPVgXBiP1cVhMfy3Z14MTvO2iuB/A/pgBgTbOnbOpz6PkbVPf/YXDwJLGv35/SAl
hf+I97O3teIizQ3bQKdwSfbUXWDqb7C/40zijK5OfK/2/oTPWtwk01b+k9crv8nf
0eJ/Eycrn3Cw3IPF3qZTaDyUBiXwXDmeiMknmgfiWNla3vRYcRc3XpK/lWWbcAUw
JwM62mcbf8pKfXqiqm9fkTR2S9Zbjwx19UKbpoWG189b5YRXpRVH2u6320I2K7eS
5JcTqOMid3NBw+jsFKhS/3rlLPi67zCLIszdXPV8uvrjlKfjVwxRNBVjWRFYy+z/
pkvqFjqpUhwUtdoFRkxa4xGbkv9uSDLsCcpdr+fLTcX2yBzlqX+IJFSrph5mu/5V
90dlBc5RfIuwDdYs6aS5e27v4kE0hzIHlHBFUlnNxoXkwbR5q0yOg7DGC5SKrTx8
fSGR3waREMnMpXVXxf7vRiP1vp70lAPmOCawoKmPxa8470qPWw4vVK+Qg18ggrN9
Y3VSPeeVOhRZIZ4lUbGPFQjLjH5oAFMIwrgJnlBEqnVKsVETzsUb34ZkTa6wFq5Z
AGtaahgGl2t4men9QClc+k8v4ghOHSsy3FVEEHRmmRBo0nct/C6UGdwPXpU/gJ0N
WQutKBRyjlDaTwYukM6VoUnbcOruqlzSnGeB3o69GmMs0QgwXVVYS7FzZXUjxNeA
IQFvEhNdlPl26oYzn60780AYIuH6nAbrqemfLpo3QFfPDnWnCoS5PViI1VUYsLk7
yLYyV42g4DSMXP1wVourHQmx9TGLYw5ceSLf+kc/cdzHrQGVXPKvgk5FT8IuVo4i
YmFU+ogbOOp3GnAyIcU0yRvnHfEcJhMPD8fEKyTdBtjlLl8ZIjuSeqRi/J8AHkIq
VNyw9ws/SW+gWERoTrwp/sGE2rlj5kBipCIARofE/QWsapgo4KoMYuuJpxbUnBUw
+if6ZtoleI8fsZeBRi9jUyh7I+GnwrRJxaIoH/n37DnAQOtnntPk3a7C68dstdwd
2F+ZUfb+TRvPGDFx7brT2Sfqye9knrChVgmThNkeAhA0yBF05tsqCgLan3XVK2bU
4xQkXRjxpu0ox3pdRivx64D7q6/5UTcwO9UA6DT9hzJZTXk63C+2hxCKtyALKTYa
a+WC6I/gTCcvnJzL112KcOifHCK/UJ7p1O1B5b1HXu5qRiXlzAeUY2mphTTe9jjC
vuUUkPWNWdtKvxv84QvsfVYLZgQrvGy+0xtJjP2BdtWPDUjuc5SDRrdR4H8wNvrw
4UvNWKBxoCLS78CwrYqxq2RHdWbzllyG7f2besUpHa6RLnxoIBigDKUt4H/OCZDO
PA/ABP6iObupqm87K71MUhmoZ/f1bLihNLtmZ/1nVlQAn1v2CFGVIh7dk+FTbceh
jvnoqV8t7YbJae9luzEgU9hqrno75NegXb+88T+IOHTMh9cHlT22M9xR9soDNJH4
l/VtIW7QpYwXZpiJyMRj/i00Ygbx152qjpCRMqWyUbRQmDXVMDfc/R/BM00cI6sR
6JR/l/0Vfjl8+h6H8efApLi1Er5lH7JlD8SY7vVcVLygmMGegKxw+WJsP58v6fZA
sOBVlO7LDwPwHzaDqtKHpdPvg5XsCL3i3ynlYEnPUtSbx0TQjE6Fozwsikndx0v6
NXmZfekOP4JfaQjmoyfEN/fkho4GrJEIyhAkkvTrdwsHnIK8cVcaz652lZ/GPLek
MTw/+BKzWSxiJ5R2/8PyLnhcrP98vf8H6S4GdMSwlNa/5KITan0mWz8KigrACPTV
cdhQW++LO4wKPz+e+dEvXrguA5QuponY/nq/1gVQ82n7/CKUzt4G86qfNrBFCTF/
MR9toga4xJWP5+TSbc2nmbW6PWWonCTmGh5A+NPFi+dxQ4HC4EmPNadMEcr1nzM5
ya9QwSBlxA8hSRx/XMCF0HGadWYCLxjt02QLzE8x/UNXl50WLc9uIUXL7btx2Fzc
r1LnJOKTPXQpLxw/QlGygKi42UtEwf3GJ3cYOOrInp+O5CXqJ/AGlb8WXXd42sdt
hPdYB1Rn20c7hWNgWTa9doklPDRvS8QfEWCZqO2+cG0GSOt32QH/MZtyK1bVHHRS
6h4uCE5eEyp2xB6dxUtNmpv4f8dkLWa6QK6ezLz2qsYAbjwkMUqj8LXk1tO7O8yR
+QWusvpDi37LS6Bm8hiV3Yo3SgZ8KwkQbOJNLWsa8U/10ZCqJz+GEOyeuto9w+MP
qv1pwg1ftgiYiJb9RJC7R/Z+KPqEytxNs2dQ180jU93+5480y0O841a1xqehy6kK
einNK7tX7DEJQ4BtSaXx8y6RPS1Zmrv/Hkp3HirjB7IE6YT52f9zuKG+JFeTf+E9
Z0xK/VtOYsf1YN64MKZWBasvB71vR6rV6KwEZTuQDc0Y5BhgSwkkQJ6J6NrG0f85
XMnui5dsHKDvlUeT6NNbPrIxxhafQ9CAbku8IG5aaEdAQg5c0M6ZKz4jbZfTKfyQ
TiqI3MDQUWkpN1CdnzEymsLaagFDuRPU2WMUAfkWTDlufIkJ5C0CHuO+MMkgZ2AR
XlKY3A8EituN+TLiwl1vXEbg0DWupDa8lPUm+j9UrSgBofUYtNZs10+FK/1HQXQI
CfTWbHiuds6Xc7efPR7bNn9g37XXbVAQUDj4iw7Bo28CPcpahG+4BdO+x46vT8id
jGpqkw94KqN/TpQjfs2BybJatDLWyPFXkN9KlvcJWOfp6F5WmrmoCwfqiiHtVx+m
qsY5UyJFqvzUYPMAG1uCRtJb5VwDfKHVynIoHp/S/+U69h2tMLTiCmpZ5OtqEHQ3
hmEKNPkn474bWNHYgw2O1FRaqB6jo/qW7qFsfjGR5WdBUJk/ZFp+CPtL5oil+dZS
165x9LgYFUhW2oknwc/xFd32Rf9+TaclhCAUbmMpDhhhLQoQJbMbDFEsf03Wn6kT
mGPkU5cI5VlqVwGV+ESBYWSMdoF8mFPgKinUtSD8ySmB3Uqz0pF5+8tr6R8kZ8uC
DOCbqG3UjtMvZuqKoEbD7BMkTkY8mVawLhEHP7GdUT/sjMxhd5H0yr8R3Mrdaplq
ukkg6cPGdZCEmkEWuVlZu6+T4hsxIrJbgdUhDZ2Dyat6Kb3I1R5og9tcTlw5obnm
ZRbeIVzvAMknme/JPwoURU6NUJu7y5d3Z4U6y51Dn7LJwurFwCXqgT72v5bCOI/g
/Dgy2M29evqrRZV5/jC4TK6tkUBpL1+au93Zs0v0b2/aJu5IvhMgIn2/uBgF/ttV
Y40IXwMkP42JixsRjRMqtFC0ikwZrqhIzx1QcS5PQJ6W88NBBkKYljOmC8BzGj3C
GQ5LuGnS6vg+iTrD78la2g7279j34M9d3etaXuMwAzfXG6Fi9QsQIY35ozO2HVz3
rWXIbSCgaWDhCN4a7pLzqbzKVZFBtuHCl4E/N5q3R4N+X9zhhlzy2DvxXIKJi8or
7G7Ko0QuIbKPmfQSoejgsudpCg4eOBxhihLFSxsmyzXduZswwype0IUcWqy+cayK
86fLlf7yBI0GZufiaM3dULhcpEEQNGnSdEsoufRFtdnJbycI7XTrNW1npZtiM5tt
ULjiwOeyRaoRhWbh9RjOK1BLyfwPa0J+EcfoM5BC0GFzhIi9DrfEJ2USv8QyZTT4
0FuGiTZLLNW9YFmO7scvIOVwlRV+5+1RnW+AzB3o3nl09Y13wXp2CA74niJrTcO0
jhIjEi1UPOgsyuCXyQVYU/y2VML5M2lt1vTxzr2kc16Sc7qLTpNVuVaiaS53V2rF
tGnT/P7PnTJv5PA7ecWdu6bKkeeJCTUv+nk6qaVPZQvZLSyxyGu/8jttnKLvP7oB
2fRthPlvHyFJU5CGIh6C5q3AkZY2atp8heGvh++FRZGnE21zJuz/09dYCfEsGq9G
r3an29IH3dZXXeCOFQN2Mi041BTWEE2ko7DotoDlpVqSVIl8BFL710lX3GTC11ux
Ln9/r915ud6oVdk5L3fBiL+DbxGxxr0Urhwtj3cpnpS3abr5EGt8XN8Dz3w26i6J
2bHoQgkJHvHfMLDBpVTF12JC3SftHN4pXcciEx9vtxrONuZn2iR9D8X+RDs9HzG3
YtxjBeN6mKxJT9TNAWEtePIFMXncWZ2QkoEywajtyDhdi5rqQSsCqzfUH0gwGdBc
WdDWPSINqkbjqho3aKfhi1CwfWJFufOLF8ebPDa6IJ/lFN4T5R/2gCpj+NN9LqJj
8El1fMdPqI5/qCOV28TCY13ABucDg1eWElk/RuKPYhleohc8lSIF/bCr3HX1fwtt
qr7xK1T9lTUJNxD9eAFK5QHJsYb7M5OA8/990DkhRX75R6ROH+ik565paGQnXIC0
lZFzZOMFp7hhxLexGEvulGdEXjBwOh5oQbBnejmJ1xxh9vZ2lEDPJO3rzwvn5E83
HnbSHEX+6jbRqnduJQldTO6SjTvZhnS9bUpTHpR13PtXga6gQNlj+Cr+lWt/o73Z
dI7QbYSm9+EGXqVzZLaUi0z5KP7ZFQNtj1NiwvV/rqGsv7KZ5nAuGb2qwXCDh5QC
1DNheAi+VIgfXK8c7QVnFH4aKNnePvviwFZuZlt1tEYZeEmifVWAl6ipCkIemk4N
ha/JuQUjgcggpnVULOP1cz10onPVFJWG3BtdqjCA9/Zszo/wXEYUylYet+CXx5Rk
q7DG65VocXJIkOahufuyZUSIv+wMkn0xRJwMdiY7xuZul2KlNWkBU5nkO66cSl7A
BDUaZISXT8SaeQf036teLJqprlFO6FGgdJPftOfuEhGERx1NXVB/LOiosQELOXdl
kIki9SFhp5F0nepzC+wAosySl5t8yHokiToexzFTXJGuEieFn8vhxJHDw+yKVEuC
ubcrkWgyxBxQygfkHXb9zh8xlN+hlUu0v0i/QptBeqDG5F895ydEzYdIcJsy/hVP
uN613Tcw4YWmNT1dlbfyihxcqNN2XqpgQtThgRiE3OMMtJC39vO3Qv5icMNahqdU
JHR1O/6onieAxBL5m0A4AqsiOVnVdGDoWe+MaU6CVzDPnJDtDHxsq5wY5Mzype44
1GVKmiMTD1yJMTSE9fe0xG6DEjj0W0fCV0N5L9zxh5lTE/mCE6KfylKJwcAjWZy5
o1xTlzGdo4QlnBR2BT3WkQ/HgpHfbhYwWBWXfxBU+6Z7atR7OAPgSeeemoEtISGK
ClJXgrXfDvZ5qzsjDnHWW8gmZfVhiSc5iDFHve5w1dv1pL3Gh82TbQiaU0ap9C6d
G2Ct77FKVFD8BI6dRTgAYIdspcbpmLp3isMWrWkrzi252gIfZ7Ioaalb0DWgT6DP
5eDnQNt+2D0Fza4dneYi83+4F6biYpzwBnWJ1b/pR4rJqSSS7TyxvGPo9opi2aaz
wTkPE7O66xch+eT57Z3BoALkYUvYpwKjxP6PANoccOEgyRSJQbA5eOxeXszc0tug
7oEmlSpQorJfi3C0GEORHmDU0qKp6N+8W8OYiEpBlp1aC3lzv5c0Ss+oaxSPGUi+
bXbyJI16Q+u5yrXtVjSZtm0pF3OvQKDLFiwSXsu9C85TXeuYur6cThxn6ZhoBuzm
JjxreqfsfmWIJ/zQK4jbu76DXQmhU9vHX79MyhVoQzr8uAQYtLhk/6O34XMZ04n5
JsUJ818uqAQErY2uG8/N4qIsoz9iqLPsV2x9ApoVVWZTYH/WTsHAodW19+54dDZb
jhY5sYeKFiHI9jtdo87xPHQpqGDmeSwMvWbJd2sqGDmUTD/17MIHlHxaZ0X+7Jxb
2E/dnb9dNjgoetZJ+quuWW6Q6z2gO+klmoLO21Kaawl3wUPskW0uOjOTWlERRJF3
FxUpXjn1kji5kMjubaeEz7pJsMXAkodsIvo9k42y5JudDNrsqdqaogirXcH2hWV0
KrSnZxVyM1dRQhHjAt5uey8GkestiXLV4khH9/1LOoqeX0Nk33bAr0t7kjD2MCpy
171AxSp8abIZQbx9EbKJGk7Iq4WnygpSc2S2vCxF75NJEJOxuIKQnkEsWrqcvE4x
G+h12ylymKZhuzIW2+7/CgqEe5axoZfChgTg3q4T26F1516BrSTaKPVwwruF7X0+
OZ8BpgbYLnNw6ZmsWY7SA0fzYWyyr13vsGBpyRZ2Q9lQV3cY2rkAacI+tU02Xk/5
3ynk73lSN8lxj+xZgv2k/s5djstB3ci3PYUGT3TxKy/bEX3es4KzDg3A2i/vG/s0
/a7pXSaM0dS+5zlAMiJ/f0PSnq9bSg9StuH4k1eK6uZGSzfiEcwZ2NaLmmnyrk+G
WipxNGP208oIaB0iSArRcW9LczWKT3QG0u3IC28W2BfKoUwbnd+TNQHVEZtnXQJp
TVtZGaMm+7S5hP8CjfdlGU6R8/QJUZd3O4E8w/UhAWiWDVI/OjHWW9FNjfBBYe3J
5WAE/WRVyq86ckkxPQEAaNWWVnJG2RMcuYrzxLfjcxwbZ3iA4zqk2FFw2lUe1F9i
Et3fnqd5RjReiu4C3hsU8KaXk8/7YNywpjLNGVeHTcCVTSC4Q0i2C6jjc7GXUY4z
ovxfQTTOcEyDtQcA+LVpWJ0RibBgbX5LjJOdtzv8vbw/HBYgZl7UJ2LkBKAZS3+m
FFazvUeFQJrnAoWF4HRakMHURBdUrH3HcJLglHDlVqEOyoByBxrUnGrf42+frsn4
kuiYfvZRMKY6aY8udi0wLqefuliDMSHuwEGEQkOCV7aKdgTnomzsm0dyQsSzW4/l
NWBZQVcPkbtU6WnWgYQqbssHADDb0j5aP4viyRjEjpuTixn9yPivZU9XU5lruj+y
Unx3bjg3Xe587pjLuBl1lvtxMGokIb3RGfA0CEHFb3nd4/5tAfpRXfdoZwKMzEzn
Y0MGUyb+5b5u76SC/ATDIylG2Dxc7hNR062JSy3/EErr2G1Wl/3gFRbrX7fJUeYK
BeK1ORT/yNEetIGHyQVnRb5dCXzXBcWbaOidY5veyIS0CtbJRLbbE45yLojYh2VG
hFIn9+uTV1PLMfpYi4tPqpN/65kwC2G9BfnaBjZEinX038kWtdsHhv1rXQGk+bji
lzbQtHLY3AsUl9hmi5rfMM0lvaIDXHqOXYt0ZkzKcOjFxui8T/V2NAJ7vsiWeQ71
J3F1I/todcHTTtySl2BZ/2Xw36TE1tG/hcmLtJ3IxygffDZRzmCLls84VItCViow
f8x/eoZbxBQnpSRe0AFlXmOnaMbquqxmKf+wt1iRNdWKL0hvRKZO9Lx2f8O5dDNL
nX1HEMg3S4f01VP29NPvCHC98Iv4RGRC79N7zk/08/84/4tmIT6VIQ2bczRSw50l
eaG9ZVmulk3oUYzsfNm3P2pGWU0wflGwD+WNnkflZkZRD0wlmGmzZ3FM7LCGBsHd
23L2uorQMc9G94xn4bLu9OsKMW19gKvgZiAGAUB3cTEPO43TmqERKuBxxNCPxSnE
2E3JAGNx1T8oqBYXToubripcQmgN7ZUD3ONoPWMglC3lTRXoqQUNowVDoxRTPbQ3
sUquF9Kwqg80yRvFTF5ZprYnqt3NavOZnyHqJC0V8tDpHu563Hpe7ZBwWCAUd8I7
KGuTr2XgiiFDqt+hLa+TOrid6XsT5QwBAE8gTw0PUH1Xp1jUjF/OfJaKDuOj3cjn
zIYqWr/Rj7bRQcKY7EjGp7xqFSZpL5LxeQsYi64+ZPFwIvlvJr40nWg9AKwhg+M/
Kyot2Ujinjp5znf/sfj8xSvyZ/rF75H2PpDD2smjNsOYTmuXa9zyiYmQLhDhU4Js
pr6aHVE8WN4ofaiL/IwNbdjJKkMGu6/U92KtMaXfIIOaduC/KYN4DwkGBT/urDK+
aGlga7k4b5jOraUQQWPaUFs+JH5tskH3oiagoGM8vYr/hU23solOcFBjsLeHtwZd
WibAlMkT+tzJu63H1Fvvktc8Psuiq+yyJt2kR/xmqF8TvvEM+67tNzbMaukLb7bO
dUlti/OzNNT8okaQQxbJydVIoRhqRNHRemWFPxJ8rIrcqRnGEYuf/ASFUkvm2Yd9
f8ZICJZWLQJMRSe+tA9cyJOV7HAmauhDhRtbH7xNKKWhucYV+1d2CPL/yPtQP7NK
YDxj4OtCVGMsUjNnnOzs3qJgiOlo8hwpeDeK6MF2rZ4EV0+onVpdwltM1FqOmxlg
hZsAbLB68OX7dH7+mtHtNc8qKX2CiNBWQQEMQoI7ytMxt23QMUrGkWtTrd9YLjRr
wrJjIsjTJSy7fkMqMOhEljG7RvmWXcvoAtdCkBWz+EHrK2YqPDIaOqevjJMhtQXB
nWjEKYoIoWsTyWIn78ayOn2vQZy0eK8BzuapSvi9g/e82D8QUQi32sXl6NblCyyK
5pQr0IWDryELUDiMODD3KmoxqNB+Jfa8YPteQb8tBkQBja3k48Q8di9HnRN1hmZH
UtKgb7XzQgiZnz9EBbhGIthqqSsZDHsAshINYEMHe/0LQWrBbO6/qkEn6Qef53YW
xcE1wVeW31fQMZwyHn86mVU2F7cFDDLb9EAec3AwStvQp4MEV33TlZ60m8ZVZPvC
fgbzgY9GQvYpJtgJ50/DM3VOgJJPWfMW3rrtB6TwMd/FV6rXVZmNX/ZjULVp9VvA
80svHVWJO/B5Y5kD0NeNrQW1NDf40/MISYOwrQLk1Gp3ZU6nmkufuQ7FbV0WaMti
SE7NG9+IRYe7jPw8OTSoQx8XRG4p3fUiOC/bei+qG3UMNF9RKCc0LHK62VB54bLA
kngtvn6rxrtFT3Zqn2WD5Daeirxj8Dpdh71J1zSSXltI38gFqx8IW1/uS/Bh1gVF
RI8rpFKtuIv2pYEIj5xL/U6bhiTRecKPGi2G7rRlhtbZagch0dudbkNYcQH15+xR
O2kFNbTwp1oBj9GKQSakDp5sN65rxVnLqXO34qeOcZGO+NPryo+L+ag/+teuRDk3
AFGVI02PkR9lEW0LssRyh3lnW/rYphQSQ5EalG3mOZzYcXiUEhrNZnbAd6sy6GE4
w1rjkHAzeZnKVktCb3XiFAIGo1TqfO2uaW4PMiU6WhSgfE7z4i9M6cBmdl/sLQln
HNK7eP2BxQfNBSlKPT2kHmZAwjrgYtOaR4qYTNzZLZqtU27oXgubtXllXmrspGfk
g38DEON6o3uosLGN6dgbHen7EuXWGygaQzJbm5sNnNmISPCUupwiDWkujkeR67u4
X1MqMruJALoiPQ7qRCqG2S5UdLfYWNxufoW9KTFQMyptQp5pSgRqwk1YqyiDF6oD
mh9o8eBKx+QPgYiFUOivipxoeyBv+VMrh/IffAJnHnDewigEW7dxqCBZRCFBnrm7
ycXMKlSqZ7PRbhxx8duUdwkeuk+syK4qTexx/CcywY9AH82ej6kBvKY4YEIZzwYT
hXf3UwQZGT1HGSKvM3OJ3r6nC8T83dRk+Qe6JNOS5/frrFX/G6nfs8bkKv5PZ2db
EjYYdvvHIex2j2UnOEri1ZAV1dk4l9AM5uo7CoF42nXjjadjCt/Z87NKDhGtvFyL
KUTCH7xq3MgBKVMXbfutUOzVQt79Y3jaUCZxk2klKzNpinoJ9koRtnhbYAFPspNB
2aHe7ZpJ+icsvKaijJ9DPNXINWYt0hRQwgsUNQFl9Q+VsXhMIPqqnue5DZ6xmFTV
lCDWZ1sX1nzGJZw7g1kw3FkMgAe+/53Ts2T6aqzd4sHRkbVrBmnkvHaM4SexmfjQ
fjgqTN+dQAyR/0l106SJcF9oWlUQIMjF/fj6VaNWk0WTtVG0GLPaGnXBbfC4lLgL
cHkfdB1oTYRJgzmCrZPoScUH4rV0irDVXFldg6i4vU+YCnlbtHbBAirjRLuG05JV
6yKSNx6WgwRQycPAEZt4yj5b5oG4HhhUOQLL0aBRPucoHSn0+Dgh+FSO4kbI4LNb
kyHm2TqjFV8XgxO9N6fcShxdBUaFHLR9CNcMSIEYktHm8idP4AgWslqNpLZS+G22
B120HieezkNgp4eXY7LALxQCHdBDE/vEjCj0tQ/b9lU0rEI4wsQRZGY5O3GsKpYq
ZODSim0+e/C43L104dmKIfqKb8YW+1IY0urDf3mn26vJTvkMkzIsVAt7QQ/LPCAy
J92jNzITMFNfQID/CWIRrGcFtC415hAWfMYp5vMsq+8J38buAObC9y81zLAEjfI8
1lVHwMW/a38DXZSY9rYe04xx3CZBCnhE+B3CkK6Tsm0xuNFAR4fzKoH2wvt3WSuj
t66RO1/L25TGx9rcDP6hhD+fP6+OWPox8U7MmkwNOvxh0QBHCsXAEiIdoNwIobV8
y7QKek8lRQ2U8DSa2+bL42s5Xg5NLOnwhVaH0kWyJLsIf+LymimDYzzG0p3kEIep
3sfyIoNbfLWDVTQZDz8E+wRqajYfmeo6g5NJDS+7T3IgqWPH6/8+UH/M0EHbzYnj
Mw/oq6QMyAOO4ZyQaPA9qmw13i/iMHOGhSyOzloBnhvq3PfQTuxGUWS3Bppl/0Lg
d1Lc5ikyyXWMeBIA12Yf3yA8swcNo7LicWTDGp82p0x/jAqpY+Xth+8xxFI2FHR0
MNcP9kctuLzNLoxWJ7GV89mvmJeWpBERkrRvvapOmKDZgbKE1M0bT8orIyfPr7a5
5PJrMew+MqnKgD1wAVOtIZJfvrkgXs/dKI9fGClLvX3AA59KoBf+hJ/WgH2bdK7M
m1h9yaUEeMdF8eMRT/h23FFRpLIjGSvTy5t+h1F2lbnfj7iGiEfZO95ZsGkgxrqW
PaziZEfsaLq1Ojq5s+PuwGo81n+VTNOqQu77YFNEXvLtzMCWx17KezlEO3M74trZ
DnYbRg1rLavKSBPhVM2Ji+MiU3fynYcLAp7DiP4UyU1D0WnBy7TstWlnq7S8I4fq
rOBXscfp5H56+QOlOB/ssbvYkjNFXN7FZJZZydUW7mDafWNdZ9ns3BBnFSUE7MTB
UNOHinTx17C2fHtZ4Qe1gbyLMU+DwluXx5vkDJBHGaEOT0aol+yxGLrmmM7FP1AV
WuBx89J4B6q/ZU1kweBxb+TRkl4z/4VHTm+Wt1OSAWURjAiBCy0g6nZ8Rgmc18Bf
Cks0c3fkXVaNdnObjoYHgeRNRVerpN0L4bEoO/WA+vkbXOe4GY6ASOQSwpUXuLCS
7Payn07wAWSvNM2DQrwD4bLrk6+3dqriaR5We3sKLiCk/7uyGHq2CqenCC+Ws019
DFTz/kr9BCtp7JCL+efqj/Q8yo7VgXUKfz1y9Cq9zDAiyvplMj6rzOzVvc2lDzuJ
lbUnALGRa1KKOsPy261FpjO2w/rEVfcfH2faVoqnN6JD7ThVsmifLVI3iYs8ZQGl
DLXRSSy3IAdMS0yN2wShWdRMXAfLfEOvWSy9z5mXmkHi1dTMieg/T2z/X7jAz8Ob
e3+sXEsBuhZWKmbbTSvXWczSX9xy8ks53fYIf6skum17RHZxocZ9AIocYINfci47
tIT8zU0lqHODh/syvW+VgKZtaOgii11Csh8dUDzD5zYl7KwQYr5RtW1tdp3fzzA6
cEH2oA8LcbCHcqrUgKo3sgCHy2woiR9ItT+9m5U+3GWqorJoglSEqz2P+C21zmHe
YtX/zzdE+Vv780qTHO8Rdst4rUWNelmoo8mEQFTN+bNjlCKswvN+Oo4igUczHb9J
7N+137ibf0omZXMuC21kpjwjDTZJoqxAK1QMamSbJ/mhXUy93G6nl1LKSMN/Jo8a
KTCKISfJdD8KBrZhOwj5CfMhp0kT7++82GPnc0RrrzDInseJ/9MbrgSamOb1RTZ+
qZ0I942ZAo9I1Y6MJInzm7En+l6D9T/KBIhKGSzOuwj31QsKKfhHqCi5KM6tBMKR
Auj2CBZYXafV3NXUVRae7KnQkagCd+Hjtwgl6ij44GRoAdM4d+zN5QXXp0/oPbB1
Ro9rLYZ9JPnEiGdFSm7NInzvucj8qpFZJfwUv9FqlsAZ7rkKc21Atuzwgphtanri
S78QTRv6Db7utd6rd0xN2R+FmieNdw5qEEtE4UFCT0REyJ/haBqfl3C0qGBA1QmH
iuUmCgNuvVq1QERgawy8FRgeF95hP3LpC6tf9STwnkuLwIRRAnWls0vnB4PXwMkm
piM5wuHJB6zf4LxONQQlDBA9mica832pmau7gTGSBrPlj+tTbaBWJyjUwic1kWbI
TWF9d6SiIkKCk90LsryQZ63g5bdP0QrpH2XZYK47ai49zWAQCToHxV/8gh6tnUYp
cdjZSTWroM4zg/DtRe7kFOYIambYUN8GtOu7f8zPk+v7iF2mbrC89lXCw6jDt7TQ
qtoaa32obNxcoWTN1HwAbIc6A4gN9kJSseI4SPE1E65Xyo9x6y6dXCMD1XNDZbvy
3kaVE8lJbZIvGxj2mVs5op77vQFj9L7m+J+hZnBT3IXXAQ/f3XTME+0LuBY9jWlK
8jXOYek3Fr7RVjzTJoNul1a9poKfd5m6wPjtA8YDZtAqxQPHdrDikrYJeoy1kImm
vQbeDNy6/T+Q0mZxO4Z3modkgAyRwcPKeh2MVb5xIram1vw7TQcRuFZ0v7LR3jCI
gv5W72qLugmEM4uVex9XIqOO2osaqmflyXYGCv1IHZSG1Voy6aBFZOfHGyeRrr0o
KtSdrBX+dDpMK1yrJ+LJrXvz+cH5zue3N5utJxH/o7vuadIuPbWf/2tNrBM3v3yW
57MppLaMIDUZrLtRgYJ8RMqZ2FX8SDwIteGXvzAicgmSxAX5N/t0CmJeCyvus9cV
JhmcG5FY6ixjXUu7O3M22vytrmMeAz60SALFBGuPwVR1AIBgx7F+BgBDvKBmSlNN
yu0APyGPOtGiBY/MyGZDDn83r1Tu447xbTzz0pVyR5RwIENqmq2JrLBnatnZpJ17
66sUt/sn541Ig6/qz/zaUPZ/8Y/vTq95lfI5FCpBuLXbNiSQJBqbnxAatgKXBnER
QTU0YQBrPW90cdxgGzQvRpoFvSkFB+DrsCsVJkp4GZXLafmWCqHlEH1fAl5gGpc4
UFAJmk+yYLikCEETq/0CQgJ2TFKuKRpVPNhqToPSwA/8lREAi7NZtU8UnJXB4iBn
S1bvYBqCKYyIQzYYJdIAz/MN5xGMXib2Qu/4Slkwq+oOUolHGSz7Ac5ROk66q55A
7gHoysLiCw3U2eG+lEbaOm9BeDls7+Rkdi+JB6x6nujAqohj2dK26M9c8Pz3gFPG
7FbxBPerojguj3jcrCSENITO8DZTf2N1abyWLaxvvWYKj/ZWq/HGzOstoPjwigKv
r3Jdff3MlBo7G1D0SE5+oh8CbjOlDwZrIP8ruVQJ7lY0y3jefK6mtWOAI1U0+6ut
yr1DUY3kevTG5f8pITFcROG08RecxGjX24zGVlhkjUP15QjWljFvCHW8NJSFKMlB
4wZSn9vi5UhqKG0c0LiO5AnUuaa7cP5q6+Ac/ZlPXO4MptRkhz6KfoGfexhHTsl+
Tb5wYjs4rfJ0CkIx48/Uleu2MOF/96mZ0FdHVraEJX3Ri2b5KYTrW5VSGiHnzrXU
wccyAuDzEay2uSxHPEP6/7wTGNU3ecFWLv8c46F2xpDdC+z0q2SLWwwKx7+UyUSr
dty3xXQrLweq8pv3roeJQEHvSienaDRyVoA+jv6tS7K377oKgGee72LfHfIX6faS
kvXEE4tpO4SLQQB7cE9SzIGtdjr4ypdTJoL7ePP3bY58EQHDiEn83hqRl7fKv3OC
Ay7OSJJNHJL18EDype2kfqpzAmXHC/wNx+kVUyoWJm/O0iJ9EraEKQDV2DkwSTQP
SinWSRkLOWgAD29odP9jL/9Z7IQZ9HfhgZR711lWlhuQ2awIEvVda1Cikh3qzwzh
lWBTWq7hHSfkqREJdD3VzwM9Wff5+TAtma5eFd38qxhSm79XQRNvNerRg/UdmWtU
VhlI6jOh/cjaQ0pH6pEnTqvL4aTVVvgKdrFY7MOncspmN7pn1bWAwghM3XV4apvk
iCqGPep1u5JZhFDph0smDVU0U7og4lxnD7odRBHB+/jCt6QPiDDdgOMQMh9I1Qbq
JeR7v8RDnLeFyhWXlEZuh+uk2qmDTrLeLxhX+iyEO8u+G7Rvu65cxuGiIDJq0oyY
Hcf5cyooh8/kVfWwivVsA0wmSUnBAv6aeEux8WTz/xlrbKKjH8hoCR8p5mYgcI8F
jcVdvlcdSPpd6DpgyntU9SnEGGipIZMxERqOyPSKt6xTS9z1IN54HxTShRW+H0zP
cKDwPawl+BYIWq4tZGuEBWO+BRxULzS5Ze0wVHbVNqrEa5jSHRtM9RO4Ohbciy9T
G6GaE/G+YZrE6IZ0p8LcLfr0jlhvrNNRuRcGkcRuP8CKzsJ7ZvK9JPWXSpF8PcSR
Fo5oNvscpZVQau5/1h7BSn8pZ13JC6tBq7FJLhObWFosfHEv/zMf8DEBHEIjZUQe
6wLw+vpV0N85mgVVNMBPPi79Z48KeQDaviGLd+Uknj1H14z0dIMBy0eZ8gKYFqas
iMGeamKBOidh2wNgzjVdWHy/ihmeQI+P+02HP7ZdQaDT3IdG/eTXNBQ/GbEa4CYN
y8b5uMMHDJNBqS0x6CchfZ/wI71VLWKGH8wDa3UI+HWlqN11/hG1KK+S2YEPDnsJ
t4Ew8FJ0Cw2+fwuuo4ojV2L2zMOUAf5L3yGgqRpu5oVv7STXtRgzyYJH6mjvdQk7
iTiQiWzWuO9C0DOxTCkzTgrI2D/ATWrsSasdl8a8sfPZOK5H0DN9+gw1Qiuxgy+4
UYQi7uoMn8KrrlFhENrhp2Iu/1O4ejgWpbpuwc3SXtsNawTS2vw/eZk/HwTzw/GE
WGx1o8xIp++t4crABqOG0AQDqB1i0Ay68mT4T6mehgF6JxIcmAUq4lbfdihzVowo
zhf2X6Co/YNHCHl5k+jjd4Qt/K9LxHdeBZ48n75gUosqjhj6Vb3CgaPMegGUgHZb
TbsmySUIs1Jngguz9XCYrG7g/vF+bd3wzZO9GwhmGAHYTzVd7MI4XhrhQzJzGV4t
CY5yNVku4lZUo4OLbJCacKf2TzGfcKkWTDpSBfUl7rEiDRsqf9mWfVXOeZnFniSE
LfoC3GIOZTJiwgIqq//LVws0CMWDcHvvqIH617P86M4LZDsWPSdthLG+tXDAZfMh
lmILlcNrsQ3HV3sXQ4WrCPS6+upBLV/8xBN6aP0eJoqP7AQDyQsyS/9U/Jsi/B5w
AmcMedhIQmHD22JRGA3LTEBdTnPtPa00bEm5GevYXpMnX06Y7+VxdAkyi0EFVZow
q1FcESHqEIE2yDvCWRiUpAHTlEchDZyAL0YTBfrKQw7a0eAJBbBiPZWZD6E/Hx/k
2MMZ6NiPNgaWKYssh6WVlMakbuGNibBvM6GHvs5lTQUrrHqyAd20++grvzTsyxC9
NADFuKUn0YADLsotULTxUaUWKbHCWqCdKpCa9+eilk3/1+kRAkJ049YO9IL7ijp6
G8kuc0JlDbCN2TD+qSXDDZQ3paC3DaogpB7v6Dv9cm9WBQojgDSXhinzBX4esM0c
9cnCsfd4WkM/mfXRdV/aA8vFm4VUQU2zML2qeH4PAkRfD9gjoN6JTelxzts7EYkA
kFsXydick1OyaqFpIW2Z80xYUC9By7rT6c8E+Mo2k5RvBMhJTz4atFYrbdMm/0s4
h3b6LgNtkq5eYKUGWU9bdjk3Uam5lNTVMuMU3d1LbFMgOMzHf6L+GK1plPaK7xJ9
awMRvWvFimSgQz336NCYVFtVtSD3V12+sDPVykxpsaZyn3bpzXKYZxepenk4NMyx
6xEKjt4dNlX/Cwb6RTpyvD+wvKUIkB0cGez8ZYHYP6nnOLvxGk9FN5bBRiN/MJI3
1434/7wL9JUHzUt6Z+zdA2337rxCkLBcXwnNCJmDZbarpco+XQsVMJORVRqU9Qll
9gitFfOv20QJSzkW3XrAEMsx9sJrFeWGAwz9ipqiSXA9nxu5gEILuHOK5gzYxDiB
8Z8vaX3CQAuOkx3Fga+TrqSHi8lAoom6DyIn4pO6O+3sOgynXgSverR907GwkGIJ
w/Z/fYbH/TafKlyIh9Bi7puGC45u/RztILh/bbselV/rgit/2MRPWPs1rTnJDW9x
ARBGfTf0BkjV+luBK59jbuR+C+3ltUQUXX6zTaEVqq3jl2VrmkoFsmjSFjvizAJX
NApOGbAPjOTVLarclOrmQBDoBdHfi2iJo3xkKZkkkI9Dfeqrh84HDgEaN9RBIcUW
U1UIfgeslCa848OQGDm2KR9Ah9cw2mkZkw6KMEsquzN/m0fdelJu1V3piEeh9i+9
4k6w8xq0naBHVdXGBFN7/oT7LfZNkkmH7FzOLUo4DDJj5TJfVDOzooVjnAAiwxZB
ONnOmOxQXP3CPoliidUEROKN2q/tDMt0lAKLSnDHn/ezrzuKilPmOH9WtvqTUkv4
mT0JufWIfKgngz4yo2BhYvQH1H1hbgoXyj8waGzFmS/bQXmtPyGLmsJB25xz/f7k
1pxFqLoUBoljoYK0ndlWEYGS6Zu0urlMAZf8hoEzLE69iTmq6+TWMYGgeKMKryR6
um+FXaxf6VOIauUCkz7nUq4OoBb6eVZuC5QcF7yFSnViCB3C6N9+AlqLWi+a3SuP
d6eH4jK6fu3DT2T7FGscY4EorFG4heaELXmoCmf5/YG+aglXP89vTcFFryVBIbFH
JA89JAvdrzwW6Rhvn+f40qEKGPU10VI0LzzNBXh2Yv4NMy3uM/dCBBRiWLPIsQPj
Y5kR7iEC9Ow/JdcI8dgTXb0CYNv03mlbOSBSnWeaEsFbwS9+4XEPi4pwVBas33Qm
EepiI1j+eGvMH4DQaBBznBPwfSGL5Vjwf0NzfPJLYKJwIi/A11SWpHM70Sc0HaKn
XxayoBgt21jCbmnMnt/kpz58OElTM3lS1QMFyOnzJJKwJCXJqSHLrc+hArCjK52e
3yiDzb/B9xLi1lg0mG/GMBUpcWj8ogAdc1ipg9ttQPUO5ZG33h6tvdK9DcaoTVH8
T8Z71azaJd7wUjN3Oyn4S2TtREIo+GccfGIioKxfOCOxgLQ0Hv6ga+GJeC+focNH
av8DsOw2o6M1/qFx9RPd088KDvhi3CEY033tmfuhF9O1AYq78nZCPL7KwM3JFhsj
kAy1lZCygvQXLiqhJlc+yE3c4+PWNN8hjlgUd9pERtseFVarwJZS+JlL2zA2B/zP
lCKSuICwGry5i5/Q/PpOG/UB7WesUApxaw9ZxHjv6DdHflkl81BgQ4BhP6OixTXs
FsjCpH/CQF4w1MYI0WKj7LVUCynr0OTHmoRcx2Pg5G0UMa5iyXKDBMpphQx1vlmR
gXsU7rdBgcHUdeMuY0R5n1xoTblcd0shjwOIGaKzvJ6G1CSwq/Yo9+p9c/Wg3UwB
Fxg5zRziUiqcIrcnaxlrqeJk2jldLSpgpo6og5jgtezBxuj33XIEXRJ3d/ZYAonO
7p8wPViBWZrZrFGU8Q5F4HHV9sQuvL5Qd1B/AyyG7Xm4I8ewdHVDxgN7UlcAm5GA
HL3VZV2rgT5d3+0C0Z+dpigbLbvshGLvI1R3qVaxkXu4eruk3jBdIkDNefXAjDO9
FTphInb1OxOLTwt10gtoYCYwFi7ZT7IzrjyXx5hvoE0Y+j8d8VM7TT/kPZoxjyh8
Jfgoh4++wVtXdueBhYa0h1iVHeA4afyp+qfbiopTkhzJvvSsRIq0q4Ry9rpGN/Bx
G4WHnRxqvc/lkXjws8tFwEVZfQig6DFLVnYk4ZttqfrUPwYNw6o9mxsoiLVhhZUW
gWsRuAo843Gd0ISYTzcyY20zHDuxybfz05aqAHtZeu08zWNJ/hcjKG3rLWzdfJFQ
/ZW3RIOpkXyhg1AsZOlO1YYUxQCQk40JhQ6VRerp4+0+2j/Z+tjvnDankLKen6yC
O9k45qceKJzq8zeDeZzT9QGxmvVopscpk5Y+NQMjOWRc+SAFrQC6g1S3ENACqpuW
1LxbPrm8q7hnsBfO4mtse56+K8jeThCjkYLSEtXciPVki8t8wW5H3BMKDDxz0h/V
4GcQSpU9x8wBsBxXjKPtYYrIRyFNys9nBjy+KddM85MuuqLuuHVoSLwB+4Fk7OKY
BP5oLnijgcc5qFOWissIyp9GpHYutEZwP/Rld78zrH0px/0k8VhegMZ0LODgkfuE
Fc5T14mpuBt8MyRSrYAkwesxrJRKsjIXw1uSs/2I5658KyYm3XtkbiQi8JNlg2Uk
478pYR8eeGmq25zkyH2hBdGtr/mW2LZ+3McJPIuzc7iQAssiSzs2CKkjoUgDQnos
ipothF0N2Ku1AdxdlVfPUeXifoiAK21vClL3ToqZddZ0GF9oDmrjHVCVyTBOHCBy
X0ObdWTxVL3vHs3+hEzszYxCCgZpk4cosoPrMlogm/ete/l3upePLrWIP3CYTUMa
06yp/Vmau5T7Y7+GG3Hqok07kAH9FwaLn8NAyI1qzqqZBwDgsDdRSi/t9PAmER0n
G44ZZOPjCOEIfD/E+gjVDnPDuJzDkjxSyhIFa+awAsPrIknFcSMgDJiUMdgEM+U4
og1Z8csRYeuICxwLt0U3HhYuoV09gb2se/rbqwKpyECrYOSHT3MaIGv4MVMaiQtD
UGLoHCeJIuw6hfYgppswTJZHOhsxi+EQt7p1g6I6Nb9UwRVLpxV79A8DThrNRJAs
5AsrsMcuFEyFFunG9WIcHKvJr//pvCVfUWP+MvRy6M4biEzoLDSGOv64R2FjkWXj
P+a6fmoyT66FIJOZe9Tn8jOpTST3Gq1/Y97nxXOFdY54C6mzFP/D1cq2QFKraru7
ilPKmpocY0WfqokzQBJfB1GL8rEuX6SbkTTZ9G0hRD/3NWWgx2maIi0WK1f1PXnJ
I7svm1zy1LtbJvNh2I3PBI8TLA1flgnW1nmph5ooKtjYxUjC9f6by0zyxxksqTA4
JP5eq32eqV1D/4i4EzdJpB7ZZ44tw8XwTkgRKuQeGwJPsDx6s5P+YxY4LYz3Ab1F
mEVmVIqDDDT556QLCHphl57PZfYlCoSXDkkHauNPGcO6Zc6F3KHFoQdVbxFldGkQ
m4jYa1tmYF5Gyi9SsIQse3qyG6SXrDk4JLGjTp+gD6PS+Gbg7ZyWd11kPlYkmFU0
0gp3XzN+G+K+1td741XymHCjHhNh6iWiVgySoccR/aAPCTjKT/2wyvhTMY4tLoYb
yVz+ELN97tntcVyMk8FoPgDFN6wFxPvoM/oTazuUKT2yrqk+eovhyQTwoMAUpiCu
UYVkmDXJQhthTrkgSWGAsh3l9AX3I7QMpFRkFTeRcMaIMvhTPVkTy33vqhZwkimz
qwmNhq8ziBqPnjxtdxedC7fn/vpMaDS7rqwp5rNKrUIK5c13NOPGh7+vs24H67Cx
gpR4dmTcrWgZSlXS54AA+/qz++sFonpz/y9KgMDrNx+JBAT8qeA0CM6CVcScD/Ix
V3OzbLSvf6uLI4TS7FLfdxespdjTlb4Oxix3b6e7dSU6f68ur0tuSrn1S6+GYP1X
8ADZ+16r7bopyotfvEpcA4m1xt1z/zHMQUd0pbaX/IFxkjDyIDjIdAc/DhK3pv6r
LDxaKlQ4sRtX2/vzU0I3vkBVWMB3Gh84KIgpOkopzsL+adTK70B/PTuIwZwdPpHy
j9KV7jgGbhCGEsCq9Oa7tNOMiv/KOmNlyLRa01Uab5y9U8BXfBwEp/YEWEShcNio
M+C9DrQyeXSHuw/+hX4f6mQXMVOi4+nWTTc4N5bYbeb+JyIXlGloH4MEZnNdkQLN
ro0hcC1PNu81AICJVYhtCFLDe+kyrM1TSefJnBWL40vyntry9pxVfgVqzQ691Bar
xxh/uDRbjulCd1nxEC5N5XP+co9wvbspFIfmovmYIoo4dz8MddLuzYy88KtMz1UN
+z91k1nJKqcEWIUDMEa+4+v5h602UOohLuC0FMVb034ylDrWlDGM1sI6ilNkLoAk
WNxYU8qudKTkiHGCY4vGG5PuvekpWQb7xe3NIlE1HlyiMUXWoEshKHi/ZT9CnJoK
GD4ctbyZeHAErA+o8dHq7urK0nyIUzWyo02vd0B3BfqJqmI2ymkHXPrdIt4ltvgX
E5t5EfRnTy4z2yxTSEN6VoGz6NemtQMo13Mz5dPjQvMj4EfqpO7i8kpg3gD8JCVp
Lt6Ixf9K6vS+0xNpU6+ohmcvuNIIP4WKbeg6yRfxwmOUF4OueAD+ac4L7Fmy0m3J
mVtBQQvzOyHsNn7xgIEyJO3mvrnVh0RIe3btu1z8tHm1h6X8wWd+lHXd5UlSlHUn
AcvBWD0GXKa1mGaKc1yAlByJ35NBf+OwZy2XZ3YOHKIWPTv+FXYqOjJY7WQRw1h6
6C30ryiqenlHmMo3d/QlHnv61BCcxVf8HyxGvD3q8O5XlMVjcCCHYFz1mhKMD/WK
zJFK6mY0FzbktSOreLbI9LmiKShsNjzU/ZfGCjDaczxRcedW60AyMwbtZua+vuFg
EjGH85zEKAyNcPibWMFLOS5o0nvjPvztRKvPTyF+3fI3PxLzYl7C13klKtjeF88Q
lo9ZE7g9kOsimvkVHGjcs8IkeJgVHLKrsSPG4bjhPxnA9xJZMoRt4vP9kpfw1VqZ
56WHRzLVnOlA5Puxe5rndpeb1j/hLKn68h9q9rwGcc5Txv4hiEzZVThns6nt6upd
xND1dTKI+dO3/Crzs+3jkHXjlRdmjox+zVuT1o+VDXuBQLbMokLOO8XjETH5vSxO
AUdQl9UMMNs1MyIQMqn9ddF7MzpdwVMzc9Tf1F0MCxbAdCHBLFqcOkh4iYZVvBXG
Hk5xSk4hh1LUUO18jgGCtfKH6lTr1gpEa0YNEuG8eKu4sY2XG0IWLZdsEXAtXD6X
OpUtR/3090bgAQGl40c/hQ4foKVxZvQ1p7wXmtlb2UveZa1yNRhIklgUuj1y/3/I
fAKjDhqP02RnGI0eDsWcJ7ekTwdVfhwmaEvPgtPOqDW/nOHYaKXW2ALEAIhnHbCl
qx47oxOPn9Ilw7kdr1guoxqPG1HVBdItRis7CieVPsrW+ZQyh+uQYtnThLFh06Cr
8IY1sNtZz2FHaCYGBd53tQ9sf4ur5LS0GC8iztLJbFNBXBiMEpsmNDfaEvqImv0P
QJy09n1alNUIyHRIW3Rx2/BOD2+MOc8QPL0oGb/oq+1uVZtPkOTKx6VPRaze9YA2
80t5/UbCym1jRjU2Wf0Q6HCDSjZnPA4CE9YicIFH/he+E9nP3TYOpNW/yisDsTDZ
h5NTmAt69YPn360N1gDAg8lZdpP/5B0DBIojZhML8JQYpIp5xhtop7hfn92Ud4zM
32Vr+oN/zPWgI8u3xDqMCskHzQVcTeKgJa6m5hXD2zaOnSHBIYQHf3T0uYnkY+Zx
68TVbKmFckqJwrrdkSxULIP3X2Olr0rADWnC+j9Aswpj/hEw5TeMiuUtfZHlH4rG
PP1vFHLjg4ntwhN0GhfRZQXS8deYjwLI/p7ygvQBfcIOcrfSJ/ScEWYe8Rk9SjiW
w7OLu9m7jm0rmKvPGp2yW2DojAdBe3A43ljdqd2cJSGt7iFN+FiS20/ItiJq9qVZ
Q1+0pnHTqcN9KOx36ztoQZVo+uf4vyW5VocjqejSO3OcSnPvNOmSzULTic9vAC0n
rQMZJNk2snmZTgOpgyw85Nw/VVAzB5Ou2UNQQcfTj/WAEMyg91RY+MDk1NVu7BpP
kl3PrRWETSaSHCDKxOb5gFev+O5oB2MH7exbuzKKPqhTUyyM0lcXmA6qS8mt9z9R
MGmLB5viHWhPcU8WOP3L815+m3QltF0H3R3Wk4rvfw0V/L8WkMqKE+6r99WJY4Op
25AfY4Ea9ZIH5OTs+PP/S/yTnLYheDY75K2ToubwHuUW+2h/e6Lt5MeCO4uGjxkE
K0prJBD8rNsV9dlIqFDAtVF/1eL1iJe1otRPP5yR+hUx8+8tLfhrD1XW1BB95rGj
KPQpYKrZCNvFrVs/iWVhYwcUN50b8o4YAF85UfJfN6235xj14cYGOhbQuhveVUcc
5me7KrNAke1XNFCmwh7CVGkw6bt5mLsmy+j9p4AQPLhA/U/LJitzVB9evhsk9vhO
soHvC+dqabKpQr/SYt7rGnjXOc0VdlIpQPeCkttj6q8MeAB5D4aXr4eCvdhS6MkC
BYEbWzAO1riHcNjEDjw2n33AtTjzb5J6/zMr/Y7SDtMwaN5mJLLl5OeIEDHXZXAH
fSaZr+JaCgr9mZqiVlH1FIFgxnna2m8AkIwFRuqd0vCw/5vkI9Jpxr9mdJMCE/pD
64ejKNKktiP3Nk4s3wFzwxCsN1NlGKyKaMIaFU1Vq6jKRBXyjMV0w3KWGr+5B9Vd
+aaoG1rtoog/4GP65tW50WXjHSO/f7OKxyunqvBKBimK/rP/o/NX7h+fH9gwotzQ
af2qGxYPTCaUAAzDIGw4HZ0ZuX3ezLaA4+lJ3CqwUUttwG9JqxqE1lghX5tU3vyS
CbNrvlKJQIhgaUxyJGUQzxkR1LAGYTYSidcIBsXwohkdq59nqDA6Sbg56/tn4rI/
carMarl+ICyHxMTjy/L06nvh05+5ki8dD2cZDmtf9e/Bh0hInqAF5rrJdMnDAmEe
II+Y4k1+FF/W5u9Ayonqf2bdUovdlOb0HSup4DmmGV4ctvyC3wqC54SFGtLcNX+6
4e6J/ndpMeJ9py4lMZTlQpf0jvRXGpZp+rTH/SkTJyvsaEYROduvgcv7lKvuP4o/
2rURoxyoUZhu9WWAauzFNEf3YuJJSGe6egXOD0XnlKdwlMqZQExOH/+Efbc+4cPH
7tNd1B5IZ4A2Qcqpi/tTI+LI/kTo6RZYSjSzoUQ2wH5UaOSZzob0lWnAcpI1+PqZ
w7pVt5Ev23TZaCKc37bMFgooKV17p3baIuxKsNWPjLTjbChbu7xL0St0LvfoLBMM
Fz4vUeSb9mkdcWNvrPmZkTl1uuDfORVnrWsXWkuVZAqwydFgvrhMHiTPiyROX3kt
kMVttRdOF9kLQckOwD2vpYUAVssUnth1d/HVG8Mzmgh5kfCS2I2sDgLKQ3QnfS5m
ZcCNSzS/znaeZcobiE316B+vbq+/UM333A5KZmV8L9/lF7NkxvwnnDFpjkwd5PU+
fgcAaAmjOSiKAAvv/VcGGWEhNxtz2TtySJ7+cmjCKPX4ozmqgpWAC0UHNwQgRlCi
VUgw6zKIunW9FsdqyUkKOK3FvHFYRMUk4WQk8xYmHEyJK84teYi68c2/0EkmJFuO
D3lLnKRhnyEXXW4ezGHT9A3WEainuw5TqBXrVW6qqxibjyVHn332qBxm9Fg85oj5
SBNgqjEoVHgSvYItS1NWKfckBbFUN6ZvQUaeVYcGtYZbVQ2ewHRLJi38dkBQ+Ztk
g0gkOJa6q/9NVk5omNKz1mLkuSPcvcxQkAFB4v23OCn/pldFqtUFOb2B904SOp/2
eXIiJP7xueJLykFle4OfHBdfJ+ZrDJRg041vsVQf6F8yNl2fMp3tArG8cbU5ykB4
Mve09CdfVAqnnvlMljocAHH3Jdsbk2qiYEU5diUbK0dTRK2hFu8nhH8VDBt9JFiV
6xMvTxEGxcXU5TdUmqkQc2NQACorIi0XLldcVEdeB2TQPdByZZtCR+cAFO2x9tiK
XYkF5FND1ksofg9Be4xygyaJW+mN+C57hx3A6BPPA3Z87vGK2Fas7DzF2Zf8DxVk
mmIZ47EBQyLcFJSwIKaBNYpaB6bdCCxIv7NP3RfskVLfAGG7S7zqR79XQzcmQgjs
gTLZFspFPVK0lUpfBbaFchgOyLgNlUP8KEpS7y0C2Brf3jijtTatUIj0dN9/J57P
rIODRlneXJPJ1Iqdw+JDJfz/0C7ueWwjWv6kv/IY5pGlnLmzklygCHq36TznSExz
O3pH7TuwvTuuoIvrd/QucQOXED5x118ANDscBDvMYe2MahiNmgsLaOORn+AuMOPf
CSI6QPhfAvBm82zK+lxRrdXHcJn/3AZthN/BzDQ0ZQopXeUNFhVnzslN7xvZKpR7
D3uQyIGu/waPZvlkLxlBDtIhm9j6s/jSsRBXrxxII26FXdkuVALICH+P7pwQuHto
N/ZPjaUHtnPTdPtvUGzhNawaULub1QSmzm32f9BIrqTNupnI6+dvkmwp5V/EMfKJ
m2sCInqkX4Z41yutZKg42+ELU1g5KWfopGmFn3fF7Pew7oxvWqPQcMVbxle+7r5m
c+Z9l+df0qruNthgwOBUPFn9e6fcno00fw9y4dOLAz2/IzxHvCzRg4SYpv3D95i5
I2HEIzCYes14E0k6sHoFFR42LeWai7n7qr1Bu3TuMzobadnLQjpdxqZ/R3JtFNiH
VNfPGiOix/4L940WoaFm0YZksK4bI95mWfbnLIUcyTJlE1xR6CVFsAF3MfsATaq/
zTs2u+3d7++WUjC9Y/o6Fc3j6PuKBD+j9TISONjmeK18ekMphWcIXCZgkgg9mxvg
DGUQsLscChWMRjD/lM6fON2VFPMYhW+2bgdzIeZW4MioOjqTkp/WnwGx675Bqu5M
qDhXOs5DbdScRZu96uAVSZ+y27iP6QCpIGbOh4/ph6Lzt+ZIyDdV4VLdvWEajsi+
9rc2Fd8ekc7+mW0J0u6PnszKdWft/HjbH/w1Od/piQg8+3OC61/hovV5t4Y9xX0V
JUo1meX/UX8h7HlpmW4FlmJTSyaeOGfcZNtIWYmmQ0u++fHS0duiH9LnmR0OdsuX
jPTsuJP2CMNZCfPAYhXl7NJZGTLz2baim8aaBPxoh7gYw1xHkERCx3zdY7W3xAGZ
hs+y9AORv0Ig3PHSrY5aJk9tNyMzFU92NifLdQyFRS83OYZeFWJSJGe4Y6+9Dl4b
fjEd9KYU42Pmcrvc98nZC2o4HFz9Eqlyt4YC8Yr/UzV7SEkH7kr2wp8kK3+Z+ZVu
NIgAYMbsg/qJqktE/7GXKN2ToHymE119Va+pia3yw/j5E2GcN/iZFhhlguQC2Cm9
rN0kfmEdGME2HZ2dZ3oP78RWGftKY8wljXW9JMZ1DfiHDr+Rscwg/LRltrcGpq5R
G1vqDLFIVwmnFGkCSasx7lSbgbLa5xFEM5O0F0SvF+Gzf8VIeXPdU/fCGufnVaws
DM/1u0J1fHwZKxapgjr9+JGNS+6QdFaD/pVS4f0OMugcN0N2mvmLhtMvRdQcVomM
DGpHni16mT79RcKhZEY0pSwXK6TxAA5/ySfZrQiqSOK/q9Z5ijC6zJyMER/xUtEB
Br/WUriAtNYIEHefCvBMRYHsV9eIQnkrJMJP89AYiMdvtalAP3ZMfLNirR4QQzbW
ZsB2sSHv1gF8fDVQUPGaof5R0jZdu9yq9XGEAAp0T21CFlluNxZWilu4zN3MGV6M
dBnCYkRktKvVgcgagZ4wrEI2rl7WX0C+lfd2R2ehzlOGCNoLxr+MLPZ3RlOTytBQ
qz4nkXejSfGAMQuKKI92AEkd0f4K2w9mdcRXNL/V7hnLNKontsap5uyKLcU7kwk2
taoWLBrRpfatTAkrW+YRRNTTN6hdCM97QtOoKBiLUMEqULiXZeW01AIJKqeZHvGd
fUGrwcC+C4q2OP4+zO0t4ZlMO64vHsXwc4sd1qIzVn+11bUwItQioHHW+vK50L8r
egSJuKaGKSf5Y7AnvDGhnyH9lLLxmVmtFc+/9WmsjooyZFmadpDvV+/chhaaGeme
UB8U46mZv9kXiNwfe4Z3T4IKUj8vgWHRvoVp6PNBHr0vlCpQNPMWlQZBb8eQ9T+p
reIB0d59HOjagyOb5e7ixYc3ORT0nv27eqht4PocbTETRNtLiI+v7vzymFUD2arQ
unEAVt5qHsnkxcuiCH6lkE1c3T6M7yRnEW2gbCsfESJL3DiuAg3bOA/dwYQAXJZi
f4zUTGJtQeGC2RTDwFMZ20AOWH6E+FVP7TI5KrzCCuPzNLWUH73EKLpV0c3blPOk
i0nW6QXmEOABwL0lgRx9qqDaTuGYlLXhj7FrZ5gRUsQR+PaC7zoDhzgKTY76SbTE
OTybql4cUGew8+FVz4syN/1Vi4G3od3vxXxj1pWFb6eCmBcalKYhejnv5N1A3/xR
lfOR3MIGP2p5P6Ff52xP1pPEVYmDPx1+SPIGgDUIv52n5PB+ZEUVX1aJ4DkyRK2z
3Y7E3btb/Ndk6Mf6TqYfhQ7KIhk9pShc5JeLk2e2V0jY9KE3eKmaVo6sCi26p4ov
FkagX6sqetYPPKik01iaTgO1vFFLmpmcQtQKgTXahLDmsHOQysuJRNls3GDp1qLo
sq5c6dIQmC0jb3gh6hiOFWEswZZwpF97ekQz1zR0TgD7rNsiWzF/D37D72f/abHv
W80MPeNTXjVNEhGoufcPiYG3kExoyGufVoRLFE8AFwFA7/K9HS8sWA+/Su11iezg
LXApd7HgrYLzCXAVS33pjDDrv1aGHBqZh8GeKr4U7V0b/ldo0rsra+Zdx/RWJ7ns
kfFPdridpFZ4y1etv73lAU5HS2crDswN3kQxqvcZm0GTBCUk5PGnkE6Q21TysKCe
Cgq2NG9AOccvqbiCOz2nw9JadbdYQWUDg6UftySdwCC22V4ACUUoeXg/r6oquLKy
9DAeqqx8Ekm0/7TOWGaXs2K/PxIRM5eFlSiYSrwq3uqCD0ZyRcnLr3TO2TrHxwKX
A17QuqM6KIp66DVpsCnsqyvZgNYV5+4frfLqEf9eYI8e/Euzb6+E3CsWbjp8P90g
J6OjZsC1XJqVakxVgJeSttscgSU9qvtSmAeuM+vsQSa2y2uJp+2vgn3pGn6n+b4A
rfy/RXi+/smsp7Nv7df9try/PSjWzr5Ql2SjogxE3NaqRSR0R8L77fmE7nGVDuJM
tifCUZpCKrBeXMs3yrqM2sJDfzxbuSQB84mxlDU3J2reIZKctiBFr10CC7Ejc0Uc
uW1SuV/Cw28gUQoZCZdIsqw7R4V66Qk2whISd5kXrvwF8JqN3pDO2oStjjRVe1o4
W8QI0Hp2Lrt6XAcpufej8UDZAXl0a6Wc6WxqlaDAfpBErKzdOQ2j2PWT9W6bknq4
o98djcWeTqmBfVcDeZffr2wvYwbxfEGEz5TnWNaxN9nu5uItM+2RqJMsgPMwthx1
RuCc2pqZB6i+dDzimk4wWv5DykK90GjEn38D8Gtuk3nNfdJlanT4CsbIWANtWxT3
zGhpZsbVE+uLb8uHrnXR5YGy87fzJ8y0reJiWNik04GEAwpX8/AI3CXK+QNLSS1A
gxt5Ka0ZqPfS7RphMol9ZJgsMV/bTquWc97tAQacKg6v7svkOnJWXeloPTurp7Tp
hxQl+H477e2CRiAxPmOTSnhwH+IZ70bFpCn3/i4Nf6OEnQha63M3IljFeDPZayd4
tqz99QmCMPxXHXLVQCyIC+2D+x4wXi+zSdjLcSrlEfW8NoZ3sB60Z+WHHUSX8R4o
qki+e+4pmcb7haUO2E/Ahr8y7Q12kt5q8c6lnuql0H+rdqAyHFHRahZlJdw7PT2C
cZ+U/JClh85PHQtuN1agIpQ8Uw3hMMOxOl8S8urPtE038IRm3EY47jxzdC6AT457
O3Um5rf8tgn+BTtKkDS7XNclIKzpT8naEBfBjxlq60YqxqvvuDmTViSNzVHsqPCk
9JJ4Og3djYfYBGKfBxDRUsF+UErSkruDhTXh21bR9+joE9yAddkNi0n3hxz0/2fO
NhFu2I+x07HeHU0HBG4oTAP33tUq2BNDk16hC98ahyHaB/VjddwIdftNolGuYAP+
LXWQdGpIuSieDAyOLAjRGdI6IcSPPVoGWcWvZY2ctS7yuZC33W5Me9dlAxYeLk5o
iRfc1yv4tikkIbkOCHiD2JZA0mx7NL928sSh/r82MUr7LuE7T/iupQ5J0HJXQh5p
3DztahEF+T96Dqdzn7XVGoVGsPn6d475Yuhiv0L9/FA6WuiPillnwCEUEtQr+nx4
B+cX0n63Nex3c2o8tbPRHLqZSJ/MUW7R1CxSUHLNp9w4RbAPeVZZbL/lL58wDnUP
wkRUIM/+vwjrAKqLnqzTUQt22ubNCAKksznU+yXoUvMiP7NGbesvOaVnVFY1jFHO
8Q1QdyDNWRrEnkpQVADXjjTE60yfRVmtNeSG3TpXAYT4cOWdJixA/B5TyL+Mzm31
t/1iHqt7u5mtpDat/zC07EjuZVs4tvV6AlsXPe++iynJh+RSEtiQssS7HAAUF1IA
FN5enYJ2opwL/ZIlvCI3X/nDKk2E0RWcsbvJr0X2M2JQUeIhAwCN44gYbsNIKvJp
DSJyWyt56l+lQVEZQ5r6ajPkQX3yKzszjXpfkEfHY+PpbKfBB82HGxShfac9zK0a
guOh5x7LvQYrCuWUAGSzMI3tTUM+Ily5jzeSk32ec42zGIM2mYQR1IfCm40CKqvM
9G/gdfHybYCUxXmlpWQ37ZllU5EIejMIXbyzFFLnbWY4O14l4Y1duF7yCdkJrqRU
H2iLzB66zmc1/RPFIvO7BJJAQS/nSkOukimqFFTMCdb99tnWCdbGjcaNUpEmJQUG
IK2CrsyyICMj9qbUX97oRpqJdg7nvW12BUhDQOyPwqe+rlpuRmmn6JpDRH0CBWFX
sHjXkqKoVSWez9KmcYZvqTA/+dg74IlW2h5yP2e2c1jwAXKVt77l3NLoIau2rmkE
MFKTth/DtjCBINUU2eCOTUFw4FrxraJbi4yUlVFDwVvBHj/F3ZJFFKO5zw2TkQB4
1uGEVT5ziX22Nb4XARt3Zip6q42ePO43+/HcTcXY5eKZ5SQOfevzdGeINBhyTFV8
4Dw+Il/+abM8JdwVUcqH20GW7pu2HtoPxslfjf91wDegfA1dbpm6eJkjbABbMA1x
asdsRiCSu7ov6bKO4UfwyhwdTDhEGJUblhhhdnImBuM=
`protect end_protected