`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
ddtXksX2+yylW5zu6QL2Lhnb2d1sD00763mmSITNX595NcHTEkwn0zB1Dry37fOW
FufOhVzEJp80NC5qZ/+F0Vk7Ik02dIR0elf3clrjeJRK85K4e3Hoo4xn7YbFUIms
l/8VZSb14+JVGURjfswrIyCUotIzlzVYZ6gzoZwDXIi5gQIBf/gI+KxNXPaKV+PQ
Ufys/12rjO6aI/pPlqSm0hCvftmBcnezN2hk1UeXgOIuKZnogjOsf0iJVX2aOOWE
6pD/psybjbnsNB6kH5uFTA5frkzIzkzl5d9+YDm9OyC+k84E83I/7/j+rk4L2dah
QJOvksSIzN867/4Qt8qYTQ==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="MvBXkzurAa5VTw+1JJ70nePUfoQXBvZOku/SMmg4TwQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
oRtzZL4VJ4iwysPsC8SXYCzXS8Fw2gtZTOskLcDV+1B9Nzn1zTyNtlo6lNICRmmK
ZRVu2BmCc2G+fmzynYlNTnSa7C0Cuel6FYpxCBlOuk3OF2tzAmLAuDyOH3Z1Yjzk
a0aHuoCdIRKv7BrZCdALt03JeUmXKPdOmIlkVGFl8yw=
`protect rights_digest_method = "sha256"
`protect end_toolblock="Jn9CQpRhJt4rnzZPRk+dOpzAubz7omckX1MrFd4p81o="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 25952 )
`protect data_block
gD6l00tciPUa6pDNTk/+t0OO0nC/UTtBwLB41d4inuAUA3i/ALrNyoJVcBnAmEQW
ptbcNp5fxEUJjnOxnedyZEuEBxWRieZFQnkRdF269oMnSNwXyWEtEi5CLK9qBIBB
i5upUAb+sW9DmG8z7yge3ZIxmicZ8qIlDNw1pAURuaEJgnn1x5xATEqBY4Nfy5sp
IJfG1X9ea3Xs4tPcovNVMkeCnMXAGirTBcBB0PRO0CqSr/qP+Bboag9WW+y2wuyA
Bvo0zaeh1fkeVNnfx7+ZI/zOrIu69SiK/gQmeI9GoJA6HdKEpFp7fGv3aqnGw3oH
36S26ZxjnrQ1GLgsvXjy6rMC4z+F/TSc6tZkFdRgYsAz7W0iCzr3iWCG9fGLo8un
wON3NxDvy+4fMBuE4g267RG0xWN1epDo94X5Gu7SP6EgTm5siOKNVKMbEEZvTOk1
AYlm5JcJdxEluspFwQeiXYL9qQe261eTEPZ0mhuXhysElxzRmYwzABoLCkiMXlBo
PvE6aGJnM/jsQvptrIZZ6h9irf/4MdKiqfjpokbsxWaIEIxUQBZpeEyeOwVP+RGg
jnwJGlmPK0pwwoGDFbBcffoNTOD3R1DwTXgrVxKK2WHTEraCa0YckMOWdFNDjp4h
WbsTXHfAs1TNfoKUQHHXbOX/fMnseCSSI76nTZWiexDH+Eng8njfpl+yooX8iBS5
dEwv8CybambTx8FGR7XR78vuE+CP0gy0+NYLUI58rgI8sD8EWQkdI1sEhOa0qzL0
VS4cTJPScfkGmFQJPjUQIeySeCMM7QzrZ1DDwMUNmF3RKu+3wh9KTfzZUE5vKrTO
G8MOQqSN+EaGHVC1Lhyd/rJQmn2dlkUthOi3RlormaFIYFnj7De18QMyXwzFklQ8
28sFiym/ihVKcgU87gTn9I2jhS1Jpt3NOI1ymYlPFKpkMLIJvSH40+7y/pWiCn69
G8qpTMtG9Fjrpk+KJRpkiaTcX5LllhTE0L7rSgdEfJWpcfpFIEpw3ssETkpiM40M
D9zgX6iSQ3o4iz/ffjykV9rJDxdOQjeezf89cadraSnKs/vKdKFhrz0CVBAGjZc3
kUzVafAajAa4En4jRk0Yty1ejQCvoXaLJslqwS0siSOwa0xt4WJtRkru+iR5n1hk
MQj+VDoCmIO8p3bm4j4bYGzk3w7HdPclRpCEDlVH+FNoldr/o/GXjXCyM7KZCd7j
UHyR6UnydnLLVkicBarr712S5AeQkRbYk0aNICXQSsDmXTy8vCt0YyqQSwRIQvBK
sub2XAzcmQUKNisCT4B8UxrzSTwZtCwZ2MOgpsHNfX74ehilNV1X3F2689fx1M/7
YwFMgK0eNXmuYF+8xFNtpx0ZH0eq3vXEetWdwjn/aV/ZRT19ZvYXbK4b1+xCNWP5
oc5t2cpaeTQOtpxNGdNJ9op97NP+qyH6bz0lAMXQbl4bLYnTyblDq49SjonNefHI
wn+8039OgB5FEA8D+X8bo2oH0Ecuhl/3FjNdxDWGjGxec2RbVdsROf22TJc1mFsA
zrCsdb25MuTy+0lg3OAeq9tekFqcAKdgw8IFf/qKfT6dXCPoX0/KU/k/wpgsipmX
dIB6Fn5aFfOAnKb379mAOEY7pUD6z6HgkBxoBjH0zP84gdI48sRRrtKzOVHUMEb+
Vvclhd2l/aPEb2HmBIKURnJZ517KKenlU8ObfKo54Fdsa9X90/B0d6N/mHvT1y9b
TCeAFR74p+5qE1wjaIn7/eUf0IbGq/ufIKjWV5mu1YVOM5Kf3KTD0IKMR2EBHQCa
z9G5+TKsTN+jIOWG/BACeX0/F5MXpJ1Lu28RJ/a+yNVLqnx3YaookNBx4mv+Xv2w
rC6jXxtbzcZ/I3Y4FlW/a8mJXAmEuR+SPBaryHw0ExAUJ3PmMmGNlyKbCxMsxV5w
WUQBKW3NMuZTGdVO8sByKcxTEPEPyt5FjRVfWNjw7FGLrPz/tOW8mH0bGPxgUaEx
xZm4IlqabsrjJ04qKG45Ba4MO3M2mQOCRMkVvJAj3fIKSRYK8XMynYpTDhT0oIxa
XK54DLW4vPygrUbmdVdLHs0fRMujH345pkIm7EK7cd5G7Q76meZFJP3Rz5WD0NTk
tnCQTqTWb+U2ItORr8GdttSeL22zY6hPTxYVvgdbm82hHbHEhHf/OJanqmGzRokz
BkULx9A7fHcaSQHg6pZL5iQr9p45YUXuVSuivOKwd2PcorGc8Y7eZstrLwQhnuzT
ZezRS1mOGu+yy/YiDgzRd65RO7q/2k1ZoC7FOvjbvjBYJsxZTvRQ0+EZBojikN7Y
+8M9xCiHA+cf3hkkXVw+LeR7FzGMJsPeX4o0OCtDZz0Kdohvd3NHI9UnUHGopNGu
tgBozF1fxcEDjBoHT6Yw2gIzevPqQzhjnFGo/6HMV6l8JG7QP/x6h5c1zRQmFqnS
it5mN93Q2/xxofVb5O6W2Rsum+yzaULsIDpGdUA/Vp8l9VLy7E/1QCzjVAJc3+pL
DT1ST5mPlGNwGc+RctT5nOsu8jksSb5ewOuwdBEwN+vLXV/JaefCEjUYxHH7Xaqf
O3zrFD05ViuySyFki7X+vLX7Dpxaedt9oSvSLuKis9VTTNUMaIhieVxggobwWtDG
Blyb7r6axNHs3rg/5QDfSVqF58HwE6DnYTPJ1I6T9kr+5OeJr5unX59oY8HaLVXK
aztIzitWXd4Xjg15j/9RVKlUdgC6ycKMtT+zAWsDQAxMkFbRsLNbURicE0jaQZ7i
m9oXeiM5dW6zdRAxandjPW4vfNAUTxRpraa7v6IytALizv9YuFLPcho32G/GWd55
ByTUyCXfCagXGUpFm0VVvq7363r+L7IsrKn4GYihULHl4JuOfa+JxN09TWEcFm1w
ogE4H4qCTqSoJXOKdpwxhMo8TataQVetSwsTDb2+uTha7u8BJS0DxBug3DyPczia
pBuV+cIUhhyfOYmG9joTZQ9P+pRasFJXCgfhPwZfS6GVoguZ+RP430Hq5HW6lg7q
vEFyBTgDe9mRgt2XtpFfuDCXHk8klBpaTruc6CP3oC79s22FdNzY7aS+Khwp5V/N
J5RPrvWDvX11XeF2ZvfgYOh/r1HCo3zeQUo1+a/AkzVyU4ipqAqnuvM4VH9itKwi
W/vRxClexuiXbSXDrd9u1X+rDQJiemALgE4BJBMMYDOgNwuPkK0LP2TflSOWG6Ku
YlmLItYuDyYLlH8AWWWaoALDSbjaPxz1kIxbKMotNcRGADWYTlQ4YOgkaXysA1EN
iine9gKT86bwKJXcy9bHgqhU5xaDt6fk3M525JEFARlstQArT+jKptLFRb8oqOhO
G+ycK9qsn6YitaAgAXs1c8/uCO++rqcMvOwhOtXq2CwkY8Hw40/DBR8zCCFLsAn4
rMQLkZw5Tp9RMIsrxyV9YPN7AOmzwvih96EfDYl7CX/DanGyIoB4YQ3h6pFZ1zL3
fZe/UhhCjojQ3a4vTtFxSghixeHtGLSu26ibCuFoP5Gx1U+KZ8+yFz8LSYF2/s05
O/9EZJn+oPvjfofGntxD7ZAV3sQ7USWlIamkx02TlkVJgpd57ZdII1IN8ATOs1p4
iTWUTkSznEzBwN2jDlnLy/1+IHhsdURcR+ySR9jj+guuK1GrtH7sChyIQwfK3Q3P
6DC6XSUvjTm6614jY+o66+RuhOCX+FGaoJm1XlM1ZKTSaduyhS0iiUbZzGhLuVSo
/63EdFHCn8e6VY7AqAEBYm6WbDc+1S4HdwhQtsjXZEskG5Mf7yfGdyeGR5dz1SOF
reCHuYxF+TtQgZPn8hUobXeFtqEhnCZI+wfjGbtL7AeCmOkgYWxEoVTlu/MKajWV
lfjIDixfuuN6KfineQONOyoq1z4bOX190Fd6dXGwg+W5rir2yPor/4SWH6eITGj2
RrdBfN5p7jTRItGwqulve6zgC5SQsv5GMJzFYyGzKsUB9SyBEMonHLDOB64fhmfB
YZPGulIt2D3A+QxJVaRq5sjQmqz53y2Nv6cofhy/G6HkIP2whfq2e17xDQD5YCmi
JBt6W1XPEqr3K3b+JNK+oU0Wtt/xEOlhhTQw9rcXDymAZpiVo25qbTd0eN0SHZbO
msk0vRMRhb909BfecYU8gJoq/UnoSIOzle6o6N0X0d6GW9WyPOU20AhfwMCcfvxF
BkR0g8KPgtHhrHyhIcpV7g0NdH9KRgBXByGco87SrQ8cxsCf6EkjJAH6pv6OKgfr
Jwi4VzhLXjvbKAXOXhAoDgHuBCtXWi+81s7oQ6Bf3c9fe/OK4e2p7bdhzZS1NhIi
DjACo6X2gehwiqUt1bmIySQkzFqgN+1X9X7FiFKmDSAptnXrIK48qzZ4UHUPJ5SR
tsHexn7Mr/6v9O0otX+7vcUqSbvWsmBT3COan/MQfgHPK0Czz0a+Tzl85xRPq9s/
yjOqknoG8c7Svm7kRY5N8jEPthV5qJZqUu9a69EPuBhvfEUkXRMoSumCfLIexKMo
g8FMJEYmK9ScBT8C94x05GlD+HEidz7osPOt0Ojjr/jc26/HVxURW/G2gC8yUIBc
VyweosYxhSO2sBpmVIVOcHF5uZ/eH4ffbJysEjVmeoTMPVpUDzXar9dA6dDyLuTo
TALKrgYt3gHqf8tfO6EZQI5v9r6q5RPrUzd0I3VrPFwNbaZrHoAFdvRYZsy0NCuk
T0HozNOqfmj9+Ymbgm8ndz89IuL56didcrgwFy8BO/yoHyliEz8eTEVz8/0SZJ/8
L/OrGYXDGFHdKevNsN5iooMP6F4gmV1Sg6e0txfdBevbFeKlj/OJruuqq4yf6gXD
So88RDBh/B1iBhg1luuCBq09KE7kMWZFRLaLzMEY6r6+8mpnCjp+V2UDkbPq0cCq
yHED44iZzkHMlLzFRef1xHSesMws8pRO/fzaE2CBp+wZxPLvaGxxUb+KY2PrNozg
8DME62UIdFHZiJjaHscQr8Ndq5iiTdJ9AYN+jQLTchKfTc4Gfo9Am+XxDJ2M+8ks
BgFwmXC520QY4XOZwWIHyToc5DBx87wGim+eMQ7fB0y3CvlxnleZrK+RoEhCIR12
UyGciMxUFyBxByPs0Y6X+h8R82l+QqBOKDxzzDo5xEBOTxJ/OjLwqwdBjdAj121C
g2Azw5RQ6uJfdVk8geerCDIG3MBE/kgVwfJA5o40gm2CsmikD9D2Nsa3zB7zqjnA
6ekzWsgwaT8HJ6HsTQslf4QU4ev9A5EWsb4MxfPoQg0rxIrk+hHMKDZ6OfjC+/JJ
B0M2HEBYB5e9v8dmHIzRqUjtnXeKwAtMWN/4BEmmccwNnF2v7xDAPlVLE01f8mzb
Jm97wO6cABaAqP3MIPugOi1QREphOiqXeZBoljfr90AckOdphkF8j0bOXL08edZk
lK9iLHdPKZV3VfNP7snJFT0n8P98pf1K1egFHKk6ZT477OEt6UhM9vAeDxEx0mvE
09Q5fvmTCjzCEsl2/vk+Gz4c/cBjoKcxYgmUl95l7a8HBIwzXC/oOWSsW5h+W0G1
rG/5rb6d1buPGOQDIza8SKLUSAnv/a5/eh+GRKYCt/Pkm7bWqUWo2tnRCjEZRF9W
KHYW9fZMSAqlQ9dWKMdJc2d5x0R5ZdX8PXIyAag899Q+XucUojaV9AsW1eSgDyps
tRncI3jmmiSlmNRM57EbDfvbHldyJr27/i4/iTdfLNmeXICUb4tYCDLfLSh/Dgzm
9aW3IF/FtD818dEe/zGVutK0+Y3FuvFdT/77nnK+rijZh7TVRdV7V9xk732afaEY
s7oSaDLqc6eLPTJE5Ff6z7lGyiIBCARXVSGCqzhb5iGpp3CDktbH2D1IvNtKIO8z
VqqRbBqPAIreRDdtqOIfklgekyA9zw2ajynwm+YeN8Sc6V4gkGa7G8bz+YU7wQCD
QQlWMwi2Z+J81srNYY3xo61G34xZIT52k/LCCOTQk0AaifYKRGnbAQHv6tpoYJQ+
xZkMy8xkQfzgu5Ibsh53fmaYKjUQm7/yaUKoqgxHoZMrQ3cQDxVkgxEQTjyL/qlp
RdXgQOIXrRhGtcgmn6GfeBmI/FUecJBmLqDbqm31ijhPBkZJXdzpXHO3+NUEnm+m
6SMWenhCRRIBhpHhDY/wFtOlWLm0YR4j+se8yEpEocybKCIU93r8QqMSCOOSYyLb
v8yzhk3z0jbzh+Ce93R8I+Rfnak8Um9B9u14VdYL9kgqv1LrKAE5ywOpBu61Yt+F
wNGCTKexnP5C7lX0iUeebmPzkGyhCbHcSyjxAJmlpAp3li4yUhqovMjPRjyf9tAG
7ue8z7mkCV7UznTE4swvnN5U9VKQNj/r6ikW1cnmNK5xFT+QW/EO5YqP/O2SKwrT
WKj7tTM3uuoY8wbyp2vThW+rDmm2DDglwb1RMtawgZj84WcPQ7pR7+IZflxuI2IE
oitxhdrQBNCo/UKKq36NmuSyYmH7OVu6H7ZRPuH4tccbvne4FYOUP6R/C1IHZ7FX
hCsD+WLxL6vRaVE8ZixUd36iY8CXdNUruhY32GW8qEXZXvVXA9eLFu2ZQbS4FU4d
XvUNPa+qqvL7AzI21Tw0CiSQq4kjGpavYiaVHk3IdY/y1iDjzX+MNlIuX/37CQbD
UW97hh3SDrHH+Z4faUAWl0qfy5QvxXfa04nJCh6txH2TvxtAWLrdmEOz8C2EGLy0
cI6QHfYIMmuTN6ON6HtY+ODK3NLE2050tzv7oRf8F6P60ldVwGr1O3jScyK3MqJ3
qzHvYGI2mtemKadHSW+aYsnmfnE0og2p0ipyGuKHvx4mk7DKXXIXAuYE00hqlRNU
RjBBiJi+nkxHJ06AeAM6vIbrvviIxqi424h1+lbI+YBIFTFjGToXVbuGmXRwTrNZ
2FUyueP4fveqJyl7Fdf2pmqLa8aRbDg4/6dfXvxdHHeMgwlLfVS1R6j5td7aiK/X
i5sb7OnKeHIjyIHo/uOMMaXHayTVcFxHnz8zZEKuheFWnVsVS6PY6iqGq2D0JB2K
km5nqOIOdfNqJgg9l0cCCTbhVAE2yVXxyrSTgYWs/nZyk7QMeG+XpryhUjSpI3Nt
zde9blTXS1g1UQ9hUB23ADRwbx5jjV9hXgOziLeJ10GtD4pS7nQ7tyjo64t8kros
MUFfSSMvf5ZSQELZFfEun2mTNVgsEcVEuvFVPfUgVLtr2RbMKcTyZnkTvEQ0wZRI
w1YMI3K0xylcWkECy0caOdKR3ubQDzOTtolaMCZC/QG7jVTQK0rorH1Pf2az8bib
HsO295SniOWjMKWlRlqqLi1nCgDT4NjlbB3n9Y5mGb6yOOlQiBM5cDxP3VkQbdEd
nGz/qySzrcbFxDUS3mCQiAil4aGe3H48OKZu//TOOa5pbe6wG21qzd7ZwmqBYOR4
YmWVbj32+w6QJneu9lg5hbn3AzafSHtqW1mx5bIyMrbIRPMRwkPHm6UH07U6f1R1
xlbtF010+aVQBOzss3m9fJm38SYKopbpInPKDtP+S5ye4s856ewFy2WyN94OTu1F
2c8y/OHSnbkznNG2R2yW7flRYcJqcYsbOFg9a/78ArrVcbx+KRD4kU/AeyfdmmD2
SmldfWzSQjVR7pWRMxycCd175sbafBVC+j1eey7ow9sZlqUeucQ6FpvrN6ZBsOMG
OXMA2WMR2fe9Q7GugpK5ri0rzpSUz7RgX77tUdjLh7KO9L6sSSo9ZxctP1DB4feV
NsN72OKbPO/Or0Fhw8Oti2dRjdSai23+DZgpkTMg1hYggexWDl4gd8qyRNwC2UG6
TW7YGy6AdwVSCiNop9qyA8aP6lJTWS4dTCX/jJfI03Hotw/bdPumLcbcEpw52sZ+
NIuzlNTPXK9uBBPBsFPsd0sIx2a972NOt4SAbmajo8VwWxAvVcGQkJTN0PeGZhrF
6SfWiNHtI59OO0gpNL2tZvq46LyoaUfAP8NpHQvcH6fMUXHU1PJWpO74zZH5ujGj
SToEo4YXxYKjirccjwoF8uQoW4zSsw+NlMX1ZFs1/6ny4oFR2Cw1AaZr7sCMg3qb
QMci2GCm6xbo2qxKCPzdLPcEPsOpZ5NHGDJwvQRJqWZE9SvxZbBaGLF4j+qy4f81
lnXJ1F+RoJ9UdOD3YevSqMKa8iryv3D9wf38MdPa38rYhBNW4gee+Amblb3MqDZr
J1S6g/3Dy1C3xJrjwr+NP/o6fd7igi0RRHTSYH3ZGF5au4lLSacUNdpBcfy3rjyg
a+II2Ixkf5ytbtUJgjkh8ZzKEyP5/I8BCb2iCeK19xGNe4H0n1UumtivqspcbfB5
YoKX4lH05gr5g8Wun1YBdkDE9fhjkrbRD4ywTn60rLn4TvldqSfYq+SWmJ9UY6tQ
uoFQ1pw500ptI9BnBAogCYIkrwoEN4DP2UyryJF1dwykYH8qx7F83aTw+tT1YjMK
omTk1tMg8zd/tPLKkYmI8gZF8WHBqdkBPrJmyQXQuJ5Dxq57UKEAnqvfftwPnnbS
zIfttf62+vlpS+bybzvr3LP2IDzMAWXC7Hq6GL3YQ468l9xcB6q+5QGpHpVo1wpT
odfWML6U8twQZ7/653hALvjnpsJdgms6OpbOqpnwpgOuP7c9rpdgmhO6pTUrJl5Q
pTJn8ahhr6KyV4YibvMOZp+maVXE72l+0IGAVzQ2CtD0EIlsLraWvqVJ166FsKha
I+gK/eeIeMYQLyg54qdudyeN2d4h+LrG2bDd9UPTpxiVqpTgy7CHoSSr4VG4bZI2
I5TuHH8OcsTRXJNE6R9Udeq1kHvFK/Ww1wToSf58aiiUYyNmOeVsfYZrK8tG5ZGj
tIr744bvSrkV14Hrr1I40ObgNTmRuPYLu4KvI+wU9e2DkHcAzkA4nYtGIg5MZhfJ
gb1PlT2rR/u3dCJ5jxzic27IDDbPZEdZf1sBOl1cgOYl2Vww/D+EG7DLrKkGQRKf
174DehHBxf+5Ez+MnobwCXBCzZMMZynoSo3nn+f85B+15rIkGdlO+qOV2OfGlcxZ
azdUqeQI8qjeec/ZR+3zV/dBq5sI3MgYSolHX86Rvd256Lb4rfz+STRaEQ5MvVRF
Jt5CYcjrNErUEUiqTLv2wVf+LuITiITUxCYL6KfmL6H2+9vXdqcHSTC2of7PqEH+
+r97t0/PXgkkX2qkBmQy2HXAscqIoHKek/9ysH4hW5hh2QKCD8QWJygjK8ybQSZu
JuuEwHlRTh2BaKPOp9RAlogf8/7fcmhU1065F/A5HBYYVjXPMxMMh/FbGqNKOfiY
za/sOAdyc3BT1aV4xin//VrLurugco6MAYpdCjRs7MPBEBcEAsa7qWenhDGoj42I
StEDQCqJXYwsp7zuZVZRM9xIwzL6cQbgeWKUn8hiVn1uO+OfBi/yhKIHpC+Z6ZWN
GCnVStMvqczsBhhc5wXI8QrvC8vmpNFwI5okor0UGCo3GOhga3OHWZYTC+wVu+f/
Z7AHy1G2aloX7kp2YRlTgzweOzhABxLQFCDLDnLAGqDKNSRcg8kplDBtxMcaIPET
iCS6kbj8hyTH4swpf0qn5IQs4HM1xna6EksPoEchd1tY9rMTYXvWFX3rbfPljFzs
x+VINTqOUljDrVqHtt4WwCXjXulB87mq8TaIcC3/Imic3OREez5E49w47Uz8z+BO
B1dfTnjrSMDN1QhSOd8avmiv4FpcRHUyezeo05dx8IPNWhA3gEGXll7UFAoVHMcG
GC3hxUjg9SdqtcHuXXtqkAmzy9PEHO/8O/EsnmaXcpxvE/MF3Pd7+gE1pAqbVztj
BemacIQSnK36wyCj8jznWPcZZvxNfFLz5VhFP6kORXR+aTLZVnKpcliebMzbYdCV
hhTYFGCbc+VT+wCuZkdEjqyLKNYXlPj6HqGo+Ky6uAWfh399ykmFhSSfg1QwIufP
UCJwMlsnxCCMNqS4l/xWnxZeHP3X4Y6n+StGxbCQ/PUyWWXsoGGESdMjweTBy+9Z
xSE4o/pMYF5ec9ettbujiHGhOFs0qxA3qyrlKbeozL3u7N7sZ0h4QHNXYVeHHlLT
ZqEVCW8LqEt/wIpGc46FyQLITQf4ofTm9dALq+wHQ47Ld/TGwSgxzZm0/SB6QNSj
c6iLfVHISey3R2K6iVuoae/7+M0UD1ah5WJTchZcLpg6ceZtve5/vnmka+OXzdeJ
785G+x0JRuaKy2x5AOv1QgILKT6b7/EPEucOxgGYaF/z2qe2w8jwCuTcPB7bv9zD
sX8ER3/oQWph1c9UzYkgqqrRaF0QP6573Jwl/Qr7az2Zdo5Fq/yFeiJAYhdTcF+4
ViiSXpA8SMFoWxJ4HcLnin1IMJcnwhO7s0k1LptkSKjhSaWv/GGaWNoiJHmQY0Qd
v3Azz3PWwvR/la2y5xjAYvz2IH1cVIbES5RqAUNXk9utXnQo0RK18PbISDNv6i8H
BLsvhZg/BxyxjXDWgkPvCG9908xKch0KCxneUEvXQqsqX7XJ5BlMLBOCwUhHRHOP
HBCxcYJnRnP+CGomU/RBW6WOIP6W8spnktGYy8M3PtiZ+e+DZ1cwhENvrzpf9Nm9
zdW9ZNzto4Ns36aI34vDpev/qhK6+Ajap+76pfblJiwy67JfMNteHjwZrDaGLafc
HAbZaa7/8LyuDf+5x0RFAtTVJYXWU/I5WL6O03jueuWQPw7gc1ZV6N8bx/8QtC9p
BXnVh5yPqowoO+9aMr5EIZjlXTgDXsxms47vMRwWbNT99r/jPYtpAsQENbpLakf2
Kp4raTVgzBOitAo6G7akGEHeuy/51Vx3Fvjv/MboSSMzQZTPUQqN41uEA+rmC7fR
LdxZv3S8DmN8YUafQ3ZXF31UOP5SqTRFIA6zFw90S50zga3F1QvgQTzeOmiZ9VOi
TKLbog6qBmRh72gK6RaNlsI+f03PawEwrn9bcuksOWMys0TZteKVX8nSJZuGiq9z
ifQUXatk9FTxvr4KpgDh+R8sq4jaQ69pVc/FCeAOxEPEuh10DrYOZo3wp9FeCMr0
Pj0w/OS1Iav7dZZAZ7bgwVa3Vh2EsKv5G9qzGkph8EB61R/urRmSIprChMVY1fxZ
IahokuOkZr8Ztjv+Eeh+3lam3na96CyPT5p5ngWGQlFmNZ2gqtuYehcyC24PiIki
prOqh0YzVlY4+/aWSNB3Cyf/MWLlcowdLmBcTpy8xeFLvZezfBVoKC2/81flG5MP
LcOyDAXEOL5ii0BWD6hUD6gJs5EKBjsBilLvBQSwtXxxNrLFDzcLqAXQeKR/vJdT
fEidb7+hzMmBBxVuq/kAnPwI13TE8NnjxUfiTREod2lTUSXGuRVMAA2kQMXr0HBb
Pw0LkZDZaLtGeasQm/qE/Cf6UMXwKNUzgjXvM/QaPRt2V4zYdh1kbLZ8RktDi/lu
nkdlxUHE2ZEyj7CQyjVPbj8TfGBZc1xjFUexy+QNo9+G7s4vjj87ZdHKSR4gnvJb
VFd6yNvKDw60cwsgqIjtP27wDOWJyrf8zCe6vPF4ZM1gay9upABtdvchm0KUEcHK
TzVyCRfTD1w/pgf/UvkeCP6SbHQZrc8k/9fwosgpiLxa1QStq/EQexK6/UCDzboc
V1JtgT9+Hyo1ETIAhlsK9cW6DRyGmUXULLz8oOGHfvJQv9m08aSyLW1dW7j7iByr
VBkuVTNa6POswgK2+3MCEnqHYCSR8WXz+jPNY3MU39JoQCWVQaapuecs1k/6nICz
jAwqq5eYAkhJOfXXjxxlRqOBHnInmwrdo8OCzv98j77LCQIzqHRTTD+m1LJhOr7s
uNduKiOb++18UAqN51WSCRGWea73LbafLAayUS3+lrdiWU2DyGnpLKMHEgORNH9/
BIqaxLTDE53EabyVvhqgH6arfVTBBWiMlSDTbhrKwyLX7QB40y/dKrWH/bzoI7qa
gFHwuthvNvcbXmbK5SmgHRrv5vW7LHbun4uiQwvNSVc0EhrIE+i+BEwFVjrRi8wd
DpXVzohV3xzaQsxKBCGjWpgHzVsg3TUh1heqvOHfu2Pi1bR60+v8AwuZKyKJVgsg
Cts6OTrlBv4n9eNqkCPVHDzEt3xlZdaeH/0AEUKhdy/7x1V64xJR0Z21D7R4t8wR
JZu5SgFMQyPl5QJwsDTzVWqcN7QyukDZhDBZPeYvk9xRlJauVszuClMKoMkGLG2q
s9ER16LZeFEzNe6j0E5ZVONANuiuweVHJlEGSOzfzM+9an/etDq/N3mXIY/+dWwC
C1ly0wwYCzBkupqw6Q6JPH2lrRZmM3Sko6UImJaOAfiKfX5+i5TeZA0wPlkoukkQ
k3KkGMjfS/09yYMrbAZDEqAzz+wd1d8rBrwvoxqTLLVr8CHPfEwhyleXrx1oug1C
dOBGLOAeTAshb2pSaLk2WhCqLSq/S4kNKaTtv43Luqt5fmjVpg8dmrmyRiSVwwxs
KjY1zWOHDsZfvyUEuHApkWI1I9d6yTByUzkU1heeh+inP7fsvgufC+NiYqiOqVOK
Or5t81UesHzBEp+wTkoJp9tGMkotE0o953dTJM7Hzgyu4vgojPT7kzA1ZxNvGdy7
3BYJ3nUZE9D5RuxhVlcHqAYskrL9fLo7NWXnh2X2OB45Y7L8J1STdoLTS2uunZuG
xUcQTT6iJKVJLxtPzEwSDK6pC30OKsaiJXzFg3yHu/IW6jj0KtIm72GXde0VFjRR
qYa41TUO2dKR1YnFD1bkqinNzBeM5QdtgD1evt6c4XuWluKZi2jCaTsqqfVdi0kW
Z+d+ve6xRxuKYafcmXQyvdQI2PUCjbsmcHLoaaKp2VHwIhl5YHbr/OKKGX5CEbSF
ml0NMvsOnqB/B11JQBM/mBBC4rqpPgRUlXlu3iQOqqSggKB2TrMP8/lk+MfFJY1r
tkcuRCaD+FdQZx90JY3c3MdMvTA9yKTotAXgSgWziBqn+OpldxH2iay/lU4Jo02I
Z8g8RS/bISFcUqznnrYzus2iLj50+oeR2O3+JcjdAeVErA7mopuX/np41V8Jylzy
TMbAY9pNOgOeRPMgKPbbkYLTT3ska/KsWgfdXSIVmLJxl7dZzY69tdwpizbiazSp
kEVQgJfpyiUD2eg45Ok9sH9na9yuaYrs+6SMzF+V4SlVzQOtD/EClx2KAFNdWq0R
eLaiIR2cteTRoMbFlV3hy3hl7TOdODJaX3fWpouNqZleA4cKJb59oFTVxb2NtnpQ
3vUg/iXgJrowchO4G/gMV32RoYDfNl2It/4+isP+UMEadOY82SKpKX+J4+GSMjWU
apgIJZESy8a0OIqMRpO4kmWyBM8S9+MWov/1P8h+JJmY2MhBAbxm3awLkhn4s2iM
uw4u25+dyU8PpwkLpww5LfZAsgRfxdnY0AKYlOHy2BI3CaQqdasBG9IwgaN8sWdV
Gg+544wo2i7ESavuqgH+33Z06V9GqpmwyHmQRtYk8eEd+hGG5CQax6LJGXK6e55k
AzF1/ws+6m2BjbsoCY1Y09IwjVPFov+H54AaDvMoRqzDWbugQCxO4h+pTfpuA8Zf
Br4aNTSBO316DbGY77MUJEzkHQXW+VKR/4QO+Eb76UOygn6TpMi1benw0M0ZlpKW
ddMdk81KxXTuChzoBlvpihrk0BWiPZs4GVStawywCitmL34BG4V9C77h92+cwOUO
56aXP1ojOzbpHppb7oWFSzT6umYIIPDYiEMI0PHqEHyLNsyjrbP7Uzkz9E2S0NEC
X3rMNn0eMhyDBx6TRKwIkSO/w51ZbKJz5+CkV6X/TMBuLwqQZKnT8WdiTjRgMpzb
eDhJ9Fo/yHNIhi9CbPluhypdeqDSGLefAD+OnwKqfaYNJQC2lWop3b0nvNIkSJk5
yeNI2jDPcX76Lhu39ctPoqd17AoQjqK3Y4ncFV/B3uCVNJY3VHap02IKRwqjP7WO
nZ4YbpJe6GOiSWBZAkfGstUnQ+37CX5eBfysbJx61oSto7LIl1acqaVWBImZMtRh
UIuXRY8nWxtZm6Kr8/PJrQ4W1LveeNiNyRnIi4tBFlmSUokocFwI/x0W7F0xGcYO
0R5BdmAoT1kF6U0eIDJHbkE4WG07Mnnf6xvDwbn13sUptids3GUYMR6cHu5efpW6
yKxva7tICH4quADbjhLyBdqvBCj63c5kkrVg+Kvu36LuvLmbXQ2ohjM14TpKDmQS
fEpAnLWChERgVnzypDaeAZYo6l/9W8KMX8i3R3uuE8dGBmQ60tKPTpkALjbHNH54
jbvZO9VmqLnKMTC08mwY/a0pMsPl6zSzNI0YSw9AR8tthWmHMMN0FyRTtl6tOM6e
+xgkVHCAnaZNX5qrAwTfvFpylin/wRMmlczDaZ02NDJ8K0LU70g7vpJsURiW3gfM
o9EPj4Q9AB2h/OkkqAmQvip7fZX9rqHBU9l1B63pwMhjB1r+mXcsTP10qdmUCC9s
Sei0RNCBpyoE7FsS4XQ9uWC7CbY+cZmlrUZarBUXvwu4XbYYBgv7OzojEJ6n1DvL
hRPtRQcgERNyDdckbvuMKEyu7MvG3+KCnyvcAjV86//NYTC+dfwc1mZf1Y1iUJHv
WSanTAnLtxhYU+idKIbXcc4fc9Lakh/QKnTA8VzyvC2P/WAUXDOQjK78IHW8brjP
cJhyK4W8l982xxxCIG57xDatQTyQ3QvEuMAqaaC8QcH4WB05r1U/r6mfhEpVszoF
TxX19mJpl5AJPzJazgu+7R7tNwZ9kCr4VQh96EDf/QGJ2jm72d87KQT/HrNNJI/x
7TOojXvSs2NgoUJahmQkoT2Fp3nygOkHamPgeMYehlKqmYdqRiFP74h1BdViBsBj
24vSFB7Te26iGFOezwbaOY7IY1sCu6uhI9AY3r2rnUwVSRdHVNpGV9do/tS1O1eF
j+6zZN5+a9AJO0jUqDbrJ56km2slrsekotMD5CYRwAZhBNEY9adg/hZxjeEcwieV
D5jNTGNMXsor9CWg8ofzKZOKu4GrzQpfTjoi7tg5kVYITRVEkRtt/XTi68mN0zV9
LfwTd8rac8wkb9aJ7P49YEijjq8Spjq9NRdP01YAM1yojmoL+Arzcsr6DQjMVaf/
kChm6R9XR7PyHjFbHzLxGshgahDKHdqvtq8WXxFbYSoj//fX5z4WM2qETEkVIsYv
cGKgbrAgDC1d9BxGKQnKt+2LkdJEScFOBFIX6J499jyPogEyOA3PAigYzxmWl+9+
XWSU/74BO8L/spYi6F0MgZF8Al+qMIXTRi+RhmeMl6u5+6qyRWOVUhqJy3OyhCG2
BAabU8mK/g/SNNqWZOlD+vynuN1C2Gh+WfhYkCYcW3hizuUe1xNqu6BSl9ir41NW
BUZcW1hdWJsHcbFnkW/guMk2Uv0S40hSm38xmKj3uB4Sn5ombFJd48dAfc/Tjy9S
WlQyCyd21tfqTSH90uaEybX/4+u2wOjtEwz9uKMZo5iq9Qqkzx7aYChE8b8PEnvY
VnWRDP2zUMpYU1kwhTqALNj01frBaJTzCVy/kxUPkPZZG6b5Z7wO/PaerAUblFAs
d2nTOjQrA2b7X02ByWkJxzZXQ75d6Z9IG6Bf47hdkhxZwdHcgQpYW4oH+HPl/h5P
qSxTV1oWgfy7ZwmXZFZINwf1w1aJpsV+H4eni1MKnD6zp4dMtcSmWjUcp9MhMPQ8
lAcabEoeb5i8MF7JVEJ3bEQ3xCGK09qdGEIC47apl8Ho8SJrY/pqXtf80LowMmgx
DJtrSDsRRhaSl5pOPt08QmQiGVeLyBhqAmIUViG1QwBB9DAzukryDUAYzh0F4cmi
FFoxzPi2B19nPPsvEFy+HaySArxRMvS/kla55IUMiusjeveKUGu3LccPRiv9QTP6
+NEuH4vnZNAJw44Iv3+Ddx8Y89Y9h6NMAONQNGG5zkyrEQLkwBV5h/x/vTA0RgCk
WBhKh8oWTk1v2ZtoZ9Ubv/Igh2vadGs2uZ/sWx1vDAwvaIWK/043X8aGQ7N0aU0/
C0rtmpGoPTTOgkhDEd1HU5aTQs6J+uar76+L6rLQKAQeLQD2gsXHn/juM5btzU+q
iZUPx89j2WxV/VTyH7vuPQRys0l3lxkdN8EBAyYC9WmchW7gKuN99X3KkJMobS3s
6ufhDrhZvGaYWTfyiBQty4vgT2HSkjxVH7kvd/s9KrSRHutrnImhLTxqSVPI+0h4
uX9pHUop3QCgHTm6Tb23JmvyxLqf78aX1tRSAVKN4syxR9UpWofTD8lW/qjmlcCv
4FVVRi6G/zKyE0ai+7WcIOcGGVPaXdtWHEVqT1YFyClFPYqzVLckXqELsrWbTU+Z
MAxOLSaF9Sdu/+HFWGyHQ6+wtChaRW1urrEKWwCJBhENLsXJi70P0t7KPvpu5bC9
FMSXAFox3dxwWh2XqcBGFoce0FDf/oIhqksvYrEpWx7ybetWyWeLubb6yrbQ1RBb
A1771xOZBHybeGLf6SchbntMEGOOrcLdVSdyGPYO9QAw7xqMSfpcqymhe7VQQmDX
EyzROuObAlnfACshCGN3lo5AbqerhWJwIzu+cFtqR+DDR2HnXvRPcQzr5/vS9pKk
Z3aMhLdMgJEEJXiw9SaZoBSejWZ/1VpnIKowMYouFuPLFDZjgWW2XCoa6yUOMfGd
ytW9KGfuH++tfbfZkhGe10wz/DeCTk8aJOuMwUjhgVBPhzJS2sEeqPYXLeFIDfJF
XiP037nNI6UyITzTH29HGKrsfy97VpnPyzxvHiXS//hbXR0g9CwgdkGosB411+D1
NLwU0en5T3wweJkD8lCLQr0zUUdV1lpKPNBaukn5LOw4bexL1lTgxtSFfWVN8Z+o
UglMSXnkj1BxcyHAWsxBkLR4cFhF6PfKEaDJZffqC9+w7LXsUMyjzA0B+t6NVQ/h
zeXdLimFFGchO2eRZvpD8wTO51C8Jr8WwLQ51qOxMgcu4WUjQ2u3GjY0nw3iy/tz
hZFsHVknBqTPf21pOJVwQ8EA/1ex9AdtysT91KQ3kBzrx5Nq7aiuvm3Hw4UyNfCX
P58IFTItyTae9Gxp98+LARgcUrUu9n3BLa2pRHZMDNMtSgFbd53LZgt895bLxA9W
kTGem+Cn94KDU7ljkaLFfNckDLavUR3YpCTRiDOyskLxzesCeb5sKGY1+Olw6qvW
rYEuxUSPDilmb4bCTpilf9e2bNC2igIEP2UqPqToZB6rkpm4C9SkGgJUS4CXGHvI
UykNt09ZTIqbEz0hMadfvdTREo0BnMpY4LBmi7sa+b6IvD0LpcBR/1JXHBE4YE8H
TkSU5xnQbcDB9Jy5ol8jVmbRVDXkU9vziQjdKTeU4T2UOpeVUsEHTFDV2VWjCZky
g69+rxq413O2S4LshlCsiFVctodIMZWGNaHv9+HJ1SmnpnrYJNYKJ4SFvCGdrgZ6
qnELt9U7avU4AXJ8f3TGeFcSyHcXMVC1O7Y1f/lDAMA0mcaxZHbX2YIa4FfD2UTM
zQreXp4er8YuAZhrvStXe7bb+LHJHg6aWC1ck5diX3Go9fEk2KLctuN7jcl8vvN6
APeuH7jshQQNQS3o8BEy2IgElL2dHM4V48TJYyGYdq4MJlirmvG14Kvu8CIrM9I8
nQMXlPdqkChLM/jwj0mXEsKoLe0PxzjJVKJM8wERXQxt3T3w4IYNCXICB5dd+aaJ
38lQMujjdmXDMy71WV7yuWor+3LwCS/l2KsuW99yFlwb84FL2dhWfZYjaBGSHml5
mqzWtpSO8D/yCJbk6xkKRk43LPGcKbMpo7D+pV8ifKsVV2Tbr+6T56cnBGFhT+yp
f0z1adls7dn1ih6fjyQQ5mhc+ykEyRHQEaCU8+jrcXwgVvwQ8KErpA3nIrFiu9VF
iYS4+BkUQiuUufkugN2z1+f0vd4PbCf6HmGTo8MF3poSOz64rs3vWhHFho+ZdBoV
TVY1oNBef5EN07sMzGwZqY6L/xaUY7U9JUxBRAhCoe7FMTVawgwqNxitc/kb4oUR
PuTUHMl2DJaLqa3mCpajWomQ/xfRAPRJyKBc6lnDpnrp0+Lw2iNe4f2Pot2l1Dfc
3D0KBlZkuRadq2wCsT9tEiWyfpRtkhRx4haEVm1EwtsKag6mqYlx/Jj050huZXD6
o8HtDVpISXWr+hZE0TBAwJToMoNC3/JyMEeQzaYw5lu6qofTl7hPgyasBmR84hjW
NXsJfs3144LsJduOr5NJ5Uzwckuf1YOVqv7Br8Ar3YFzGA7VA1JJmgHso04AHB0L
mSOe6aoQQo9BryGb2LgkvfvWg+kmUOpQYi+tKyiJQjOx9MW/T60rQgdgpMUdC1gD
7CrCP+TGBJzi8FFccIvBqQRMuJYdNzRCzi+oFWLI08zk2K8KJQ+EKeEzbFp+AxOc
r3yTjNGzQkYCX9m0PhyBmnt6dvvcWjG1uGSSzbI8V94y1psSZOo+cjPWdvDLC9Xw
LMxiZ/yPc6Zgfi3J+tL9J38OQFA5xWGTnWeQ7PDi4sTZ/3dt0tNTnvB6nC+sLuTr
XTScXbr+x03TBLvvrkG7xAKzyGXLexH69y2HJaO23u4h9Wc/5RSNGvhpz8Nj2tha
vkLQVY49dFfBTxVRyw37k0ptBQ6ey/uCeM9Esj7a46nS9qn4NRASBdqVVVG1btEi
zYG68TsPLbEBej5FCMu6Cm2fpLXOxhhRFKezKBKWboGoezI3SxaGLJWmkaqrTid7
sWnQMfQXDSdmdFj345cx1ilbaqn918VeyIrGDtH+actt1KTZK2myEUzjq01cKOfs
O7Ig1oSLg0yAK6zjCBgk8PPzPtGvFT0o7Pjb0W4itLbrNI7RfVhzWEfDWwBsnsix
CZldMKoFnb1DMVQWwKpezt/eUCizRPE/5Kp4MZbffM6UwQ7561BHW9ucRTiT0akU
oZYrfk/GHB3R1ZdFvRnVDVkTmhl1K5CWZlJ8Z6DWvtMTpbhiA/NIaGjGDgp58xaC
AwuH3mb3gnONeVc39pFe0sTLRZv4CfvAAi7fdOFdmm3Chi8LrS8prRWrKLaiTtnv
6WuGqllpUesg9QoWvl6Li4TLKafCrNMG4/RuuCG5tA/ODf6imhBceEFpibiHP1VR
GqqQjOEgzc9qGoV9vfhQ6bsZpc5xycmGfUGWLC9J6f5iUJqHF/8swZy64kCs8QYM
tSvT70wcU35QZRlJ1gm8BMYZNTDYzjhxuHYrGCunnmKNrFDj3gBFRpd38d1a7g8w
OtI/A3tIxOWgoIc/kdvJDU1uBCwx/tYTcnVeqJqQOQZqdWE8XDCrFHCQoxnjDCFc
ZaxqhXSbH0sqXiHnyHlSgixeZpjF0Jh8jbrS+4Ti77wgt+7Xqc8EaktAQ9LzmQws
QmSNEmIQQTI3GOejQgcHccLh+Tf61NTuBWQtTnfE7PjO7sHdAUBwOW/JQ1gOHVaT
+ncJDUlzyrEEyAJO9vmqLxUbDZk6FA5Jx/2fSV7Wttls1O2yRTFTiy5ggNxPiIUz
NIzBr6msYUPz+Ud4yOFK5uWrWdFFpVxw5VSvn9pzxJruZpSTkOQD2cAzDHaNghc8
lW4knJbEmUKxKl0J2kw3c+ORzBIyMXUF7H4QHTMtBq0e+Z80TXXqbm3w2kAsbQcv
ovnt6vUi3+zhs6paDEN4Z0pIzP0wcRd26y/gTd/rqGnvaA4iHRJ9cjmxA15VXi3p
2yeFGoXQ57zBkzuSk+7wHGNWV5akg+X1hPhEJ35byspsrna1yMP7AKhFIv8UO1Pj
+1I3kJ2nckN4yzMb4LYIMU2upACjbNf9zBZRri8mRgQnJj7NRBYOD/uPsIs4/eeD
iFp/Z9/uLj4Cf9hA066JK7t8JoPgibEGUl629Y4pVAMQ82z+SaG25UkZZMGgO7wX
8f8DVRck4ZC849hwGWkKmHzZri8pUDtMI1LeE9V3UX0mXPtc/qWfwSuVgAnGXgoc
gelNeWn+31u1EvHC3vSasvP9dHSZHbjspPrZmIU8czafuJFee/0COYzuBN7Jxjaf
k6xXHtaJumr+qX7BnOyTDvohZhmimFQYxG+K1bae/mzkNredmWfIsKByIHCxgy58
uxCW9c5RRNO51Pr7uEi35b7uG4Dhz0gdr8mjO1ksHRpJQCNOtYXZKpFr8Od4xX6M
NZizYI+PRAhcUiq/YwzoMScBRRYoIi4PWFv6erVh6ToVfq2y7mlu6pCm0Zg3Vv+k
+SkPKeeRFErnGiKNkFgYCLIj4H1oz9tYhGvLbFgRGHTUXkKJxKwUl0t4Z1cbtdui
W23eymovkw9UZMgc7fw2bVwR0K6+cAKI6apHIXVtTYOIJ82Gy4WT7BXhwh6QTxgo
B+Gg/AJyJFgzx07tArO+kNdJsODIqNAfzUfjZL8MVgzAqz52jXwqoTsapaN0cYin
Wy5S7WggRkkNF8jwlpsdLn99VrlwrPr2RFPc5DhmHdrzq/kBvPEdxZmDigYwNKYh
ndK6PCAxjkrJQ0E43Sr8ei7GArPBlzN+F2V2OevcCekbtmQsJ62Xgv/lQ2tyDVXQ
sBCNnRxUUQgd2NYtosjLtMP7W2Yd75wjBE46k7TkkqvaewnQ60KtkiSIsrZBL2Te
z+4fW0gf+wBwEeAp4B7R1l9YJUgtPnrQGCPyAN1M+TQq39tp0WZicMXRaR3V89qG
rfdzrWCbuiAPlQiKrV/N4jq53fUwBZY9MSaGt5OGuk/Ra44ggQCL6kQTKtceUmO2
kF5/wg+2krZDY+/5QKLC3AGzT4yQoaCbfUA/pI1VhGceQIfTp59ArdR2XhA6AVVa
H+1CsGXPS/bNmcBJxIbk8B5Emj1s0TySP6o2n6e0j5zqs9Y37NeLcYRHD3fTD75q
2++NH3eMckX6TArV67RkvgC38nB5EMwi5zNUTXhMSD6HWACu1cjGNiBlx09w0COR
lgAuT9aJEVuVrUH91oZDbpWGHPhRCOKTNB0dC2gwWTQdOcm1lXecvz74wTV8Hnj+
uwSPag+wspLQ1rin9Mwsgxqb0jBCvxPi4LacVMm6HCm3aydgZXXSdRUBB7/S6fEa
PgoGAqM7fR0rT8PBqXyGI01BT6HlQcaMle6o93F9uYkWsROZRde6UV2V50SKKZLF
L9rEKwF1Ei9Xv1sUb3XgTRJR4uGKV3awTstmrEpSRMZCJI5YFAtgQO1TYllWrJKm
FBaoxUvK9NpRsXadM2KSHR3DiZAeLHAngfZ2qOWhFZCVnnFdg4dVzMEORu3ejaFb
mfrD+QCERCCmFB0p/LpJ8Z4B+BQ4DgUPepMGuRP78D/MmUz6Q/NpRvqCh1KTBEys
HvI0hmk+ITV1W3goFp31dmaMR8pHH5uaIq9ewoSsa6/CVLUANN4IvNlFQW6CMH/r
P7ZKmG02uMxYgKMA2U0odNxVRpe24nK8+O844sGAYNKxy0cbxXTUgXWMPh9d4xQE
EiyW5huTWrIdR5ND5DLj5TqtgoTmR5Au8q/42gHeBDJPqUECIqe40XG59KPHmlOv
le7RTcQcmPlv6ogF0hqwNlYoB7bRUK6dSO1xAZpvoHn3/98hHuQSrV9QSsnfjShm
DvViZ1lRGcYTDOvlXJuZM/esdssOmbNmHdP4VRMImqc1OG2/Qxspubrv2naO05pj
IphweBgiVZrfz5qTDhVu7790pns/d3VGDocgHwS8QSZ1acmErb9E8BuhyxfSFxkb
yGov7Ci9g8aMcChiOflpaPANTNM2GyZvYhL78KfkaAEqfx+0PSDX5ZNS/AF7rjeG
VUvIb1gsYVU4hBpiM5TyZFM8R5z9i35BPqvQNLSYAiwvm/MFpFhToPu+2xFwgaI/
lGGWl5yhR1cGXbDFFrTPFNomwOGZhrZFnR20Dgzhca9W31QF+W0YPMTPgurPOG7+
8rbvcXRljlcIvvkegFkBPLTS/ObhKOJuZD4JwVi7kDtTCxr/i+TG3O+3/SZIdPXJ
eHCpJdO/HoNAEA/KQc9B6kTKU0zOAGRmMfmiaDao1c7+bvs77Ie65Oy91URBoEM3
PeuP/1BEejT8zMHer4ubY6Np1odNnwTqyver0UKysnbnxVFWic90X011PElJGcON
7lIB9bwk0Wjp/mraeoF+FG2Ir19ZrwhfrkrkoW5RSCmzyBiic/7GoXlFm6MOL/uC
vgSZWm+oYfVdqMrtT2ku34dFtYpdXQnrPoBfvPs24vIr00tIUfCMLzcz0QTokToS
aMUD4rxOW4Uvbtski3AzG6Ebw0oPKKFNd5tcR/e/RzeoeGdQYvsC5cgpQj+p6nBD
Z641SHqrQl8b3awSPKv/WRLNOUeuHobOlD5zgcCCdbDBzWaRLcGRlNKjSQna3qHP
gNL3kZSSbIpde5dBhaBS58ZkGplQQbqBtADvP/bmUeBUuW/wV/dsbWridBJ6X9KB
ybm0HWHEl7gZU2RLDPtRtbI6vND4NwaNFnoOWgEyRqPhIufd8AhHdXz4lC5e7wIo
IqWV+GLesAxussOvgrB5syaFXmEapFF6mIkZWJrAImQoAnYXgu9lqmGNZZZcdgQm
r+BhZYdmHH6Fhv6ib5NeYFrpAoYcKnvZ6e5fVvunl3XSLBglECkEK/05bL1QSJ5a
cRwbVHX3P0zaCFgRLLL2ZRQ8k3oUlMXbvBGJRPd8A9TEGnXab0NQ8wxHiH3qxo94
E1OdHIFo9RW0wKjVp2mc9wDWN5DduEFLixNbbj9O4VKSlFjVh8SeUGt6vht6BSKL
6ylrJBNHG4JkfJNnAGzrYxC3MYfILNTAdrsMaLcaqz7ORj1SBuBC5ynCf8ddE/+/
7se/pG2zUwCJfsIFTfL6RY+WrYRJIjfDAKXdISI8+uIw2/AeHZHwsd0YaBFIKhRQ
cZmrrK8efId7eh0l1OWJARXvjAv2F6BDTmnf85vg9c1Ko07JO6jTOT3ZxSjZ9HZ8
DMYOvePvEZtv5ZGfEW/fyOpxXF5XXku0pumk6EptmEKgaQeKwy1Kd9xzusWr6WUB
jqqDvDU9YxVfugF0yeURqUDViQNfWNhxfu/7BD0BEk4cnNhGfFGRkfbrhDYGu4D+
6jJuwmNeGfYPLNUrvLIJ1+xU09FzI8OHGzCGL0g48Dndu/34oJj8HBR1c9AeNAKz
evZVUl4smcsoLLAJnl99/JmVm20kTN3ufUCO7XPuuWbXKGkSsT5WLn57zS7fJ20F
+YJcTYFAovHTALNFg1/mw8dcfap01cXvYB5MAFRq65wh+6yHC+fMh53ST4xgo+3y
MXsOFqI3r3YfuCr8KRdm2IFZLwc0xT9voY2ihoUnG4skAZuXmftLlXBQNS0uffjV
oyIPte4JbhM5Isc51SEMUQfQ+Wto4HT140Kw+h2s6U2w4Fm1BeLFm0+T4uRVz9Fe
qDhxMA4tnp00FV3KNee823DHTv04ABgJJP1mCUYTNMZoC6bt0C5U1sPjDIIK9Ei4
84B/tKvaZW0rphkyy14raRbtWanVC+u0hYQ9FU72Rw5zGcCyNrwr2ybNQBCNUV7Q
k+oF7wSG4Q4xW1I07KeoJxiAL1hxmpOm21bIVRGiW+ruz60Ql87P/PC+DRmqXISR
ggDRhnPjqH6ywokbmyjYi4LDXp/0A14/2zHlCGKVirnCojhjmmrFhJDQkLjnCP0i
mjbdiZH8D+0hlaAOAz8pv6k5ZABrqTil4hqltB85kQzmFcSpB9GhOYfU1OX7EEdc
xLrYZJS8GN0GJX0Gh3/VoNGs0Y9YCGCDbMlMiWOyveo0R3WdmZANfttDSZ4ImSf2
hcWIkvuxdY0oq00sywaUulTsB26Ma6h38dMG3RrZeYqaFT4mMAncjPxtgVXXnvNZ
zTZbQ0UOWyHUh4YiS5mlKlt1l7E4So3exvaS2oEvuWIg60l9tyyZJZLuQ7vm1ANP
RiVEDdkuTfGOBwIkK5VSexpAv0uCXIeLpjugDhQLZzqNwr7mZwOnZaawS0qjGejE
hNhRANIO7+6N49ENThdP5Kx29dg99q2XG3RdjcFAD+nGX6wZ0seuycj2XOYfTWIj
a+R40K7baHb6IFHpGrXusPS3FpM9MbFDoIuDWYEkPCGz26/wTKvCbOLra/ramN8s
UKXqc+v6wPE8QLj47+9qBvULBJqKuP7JeMVptfqsPIBYEky6EuM/ugBvNm5LppD9
EKyXoJRWfpNwBJQ5+bptBNYK1+V7BQ13Xc9cfgRbWsqnUd/ZmBiDReSAF+O/sx8t
VGdf+OuA9gIQantxV4qiIVbCDPORRqN/pP7vYwc1trFdVN2T6SDSU/zPG0ZFaTHQ
evkaMpWDbnaH1yJD0bgZTSuRW9AR+egn7LIl5UzFQMFUxA2vqu5Ci7FXBmnCZHhv
+KzJzvM1ObUNDUCOnbVYAIN8kHiYcdy195CN8lh0TOvYzNN5LYJxatoBPkos61Se
BNF6JL+sp09TsN+NIu7RtCchNT4kwv1mYhczclNNGEO2JNunzLUQtz98LSJicfMp
MV8mCTe+P0jBi7dL+aY9+SK43/7ODmGqTkDfeA+wcUkNV+1qUaSMWlc9llT9Wlaa
UxiIL0tqi34L3OGCbr3Vbob/rCu6cgR92uZYExIhSjSdnt07ulZsXDGvMZ/ClUyT
UVwCrggNNOjC5ISkKtHB7lz3R3g4BgAkysGcx24XCfb7Wpw+aoCo/YzRPZ3J7a4e
Rlf16OYXgrfqnd8nI7w9oq+NieP636lrWvcL3ddricBgUkVklJrLHRSr/gHuLib8
xFHHP8XTyZQUHkxnobJgEg5s3107zp+syhVZQ/XYzkldjpIYk/5NhLif09Vz+SvL
XaOI05TAU30OgrSlcdu4LHliqp5KL9nmRxfJpnxvvNbM02eTKPxcLNyZ2jNX7dP8
ygXG0e9isOzCC/dfDlDFeuA/VhRidy5nuXUvMEW0ZfgHedoZtdgXCfdUKrv53UkI
ORLsvTGLpifiOSjxlxwDalE/nU6NN7v2cuRuBWFauqE/PhxHea+3A4XKGdVIAOD2
zL2jvx2drLa7RKAA3+YeXoW8f06Nvdq75UYGFc/i1Z3nRQSl/NSEO2mfn+SZPhn9
75pN3AylhS0jkt9d6U5nkNUbnjuSPiBOrIWAcY3eLEDQ/sQxvV1OrJMaMKBRQX9t
Mr+2gwTEHehh47+wXzl+4Yr3B+5chvXMmI+FB3GawxDIutgZKPrqUFJzo6LcKet9
74rFUMiqk2KG5swXEUwCvENbqhFej2JZcc4x8+9cmhLpmnt/hwjQ9MAGtTmobvo7
FKJWsLKhXLRm50VXVXeS+alUtwgil8ZBrErDycNA+KpXDWCHvt5gn3bPYCDFc62W
v+rlFGUmW83ZPgbwjdx0reRqygL92cDpKf5OjbzDQk24k1/XQfxWhQBsO/frLKRO
iL5485EHNGsHOud0qKHfTulZAt53Uqd55/E+PJfHwTZGw52mevoR+8SEBdzSb99n
TukoMDb4QUE30sPxoeBMdvLKHmtA1j3bXkoyytbzrQYUKEzMCXTxkJoSHMys33pl
mg6ZuJvL8X7BLJCxJod4LqrDgPnXkUdtyx/5gQZADw/HldYEb9zDEJemVx/4d77u
o/00MObS1cyB7XXq78gaPk9N2qpoYpGfe5JHHsZB9FKai7ATo0xlfppn5rmQA3+A
HQQHdc6bmD+Z3Xpvy2/kvHOPU7qKDaO1JTHyJlipwd9mtjFk5Yr/xsVFkdDaLkd3
Y1R+aSTaDiyJlKL7Kgi2SYWc5gciQJQyi4NGDNRNS8PMjCwrkHsTncHLUZK5yNZg
hmV0/Lx88rwhZFWr4Vh+HC/Cz5zpCuo6Jhda06VcSfO6B6Brmp845qCSI7Rk3u32
gFcljagywBYZdRMu/547r6QkaqCTxvbunVF9NweGjaga3b9kpqZF8cp5zjpRMeCc
r8syro+hBfssSeyAo/kyqrF3v4cb8IWIGO0MqqttYvD/duf4lak++UwgrMnkNIak
k1uouZRp5iMR0/PXowGnJfBUUmuxnQW4Q+3Ba1H4VQvsgTVqdpFgt+xDo0c/jjUA
BWZ/3VBQBYlh0Ndw0r7clRsZKBD95HOvSlP+A1/HdNgl6IWIUphxSRN35sI/Iwgl
/JV77huSAT9acraAipFcAXoeSRudGBSVkv5/DHYcTeCw5LsrV3b16K1E2cILPeP0
Or57nSjVvtkEOb0m2jJXZzAVi/7adtaL69AvV2OTsjvS+DzuNTHBuhmQoPnk1ZMt
ewO6XYfUpJff9amZg4vjm0MotuUAh+OzpDkI7z+3OoOuQyh9NpFdBR+5ynziYfD7
gXw7UQGCfFcU1RWvHeh9uZM13gaz53wCU9/v19yviI9ZT9QEf2RziSJsDpPlmybd
Pcb3PKQ2PWFc0+Lym6uK8p/8MJRZkj8TW8m4mV2qS1RxrkKFDFR+Xal0/TbgdVAr
sOwitsMZ0bWxJr4KBGiBye+5exXu6IUPsUKJ2see563WaLzv2Pm/85cIbjVg+UlQ
+oF2Hdo4FNm4ShAgudlA579saE5VxW6t0G6mHEi0ZqW6MBDbAU6bJoV9OKN6ZXdc
HeWi3pSj8DTeOdd4Bs++D/XUlJGPAxVFVsv11rc1kQ6h0DT63fsACdhgKpdA0QRn
rqy5oGM05O+X9DnyWTriEZFOa25c2u18Ok1Hsn7ytJWon/hT/n6tN2/dUIiabMyJ
RKW+yWyAZP6SALGS8y1m4TnbJQm5MJar9MH4dcWROHODVTvXTT4QUAGw0pdgTbv6
ljpkTwVI/awe1/RrRCN95RNIxwhMIezM/XXnibO4+lR1h6EhUl4/uTZNNum6WXnW
AL06Pb3BkldufiuFJlFg6Abv1iRNmhTvBHhMAszorc7O7YcnJhFdI2TH0IusUQdG
lD/8KBo+Oj/zWV//+SEw9BeYoHttBNvmvV3cCo3TuQ7Az3YtxR3DCQ/AkRNAgtC7
lPTHiKaKoM4kliTf6VrUWl0DjlbBn2pfxRMCT8ZHBzBX3OL4btPrU2atyZKLo6b3
TlkZ7Tf23ZYHPprlJiLJtHLi2qwLkcX8Rf1QHmP+wTvhDrVDw5IB/C1gVO/Mi4tB
j6yKFJUjz96WpFd3iy2wF8hwqJOfS2+1+lWJK/vGka2PkpTb5ReIOpbFQJsElj0D
Yfrqw6VeIAkLd4RkCSLg5NjnNfCjne8M7DMBQ5Hn8vQo/h+zz5Uh2Rz3BWEe0RTU
N9VpfC0SQ3xfgBvpvI1gtZ+3LPwiivv2FgAtz9DHVzTWyhJv19Ok2i+IOuhKd7t/
OqPZxifT8mF4gbq4LhTXfn9zo8N9KIkERWRZI5WknmCn/QoiOUcUfST6puI/S4G/
E1u2KZ6Ikm01zurLDfxZpPCwVPPyc0bD44jU7ZZztxGt9WwQvzZe2DJ9vC8EhnM8
v6VcYQNT+2YgzhzbCYFViy28DynmU85RaBMEGxHmmAPQrN/pWjgcCCuM7vapVczt
xGCACLXidAt+ORtjDNJ6xlA3GqlqwsxPZdNk2FtRyoTGAIeqPn+jSq+gSeB8S8W+
/Pe5IdIUVFNaAVWkfogB+aV8I7/NvdEqusGwcxsE60KowEnxsfvX1uvKS1HoRilP
/jxSbn5Puj+SywK1uO9jhnqwm9v9xLaC+e62wesXajAMgTJIkvrvw1LyKVokziQY
Gss1b2nW+bOHrLVI++GS3eVON4dSHvZhR16uvmvlE5+1vfiEBs1+JViYOZ645ccU
1YI3ls61HVeVPabwmE2Z4DAql6jqGB8yScV49eWaoZ7PIzXqwFuSjETOsDti4aJD
9+pqbVNdtApi0FIh3POmRXPogbxmhzzfx7yMBpYj1znCTPBEY0UnY8Tx5HptKnJZ
76hBy7SsRgwwmZzGeS2tycv/ovRmnXD3CgMWoX9vd8lT5Z2ZGjwjYqMTn40obNer
wra3272e0q9eZgJTENZni5Jj7DIGkm+KyjAx1UvZ4GX0MTV/6DpzanwKKNOHU28q
SDTySdRJeK1F0vB6/xieW585BHAeOdJ1/L4Ksj5iMcIR73vtSHc7/u/P96H7XgDA
v3GEkMPK/9ztyDbLdCcouIGJkx0varmoCq2VlZ1aucoO7hwhiezlAUNafJqw7uiE
NwZYilx+sXzBaZC8rK2CngubQgC4hrWTK4+GexUIW0Dzz6w4Uhnabxt+35KSZIVX
2ODwDrLP/5suP7ujq+4pnOzemtm9Aank+AU7AP0v+qRGeE5gglS5qS4WBac/TOMu
mDbX1paVVAYvNWYQcFyFdDMXOf47VXRuh1/EdiZzHmYc1mmFYv+ZUbOmcVmcJkBW
1Ju0MQFaxQqtkwSGM127hbx5H++nsCWV7pvf2hB3SRkWSDjcVwRXKHd5+ms76V9F
Z9QTaMQuyDXG87UdQ6gGwgjX+5dyVCJ/OVn9NJCwkv4zYsnAcfadJUSQJn92jxV5
GbjR8mDy/e2mpjNs728Xa/QtwUR2NhciWW4zamoxmyg8iR5CELB609L6ecEuJwm5
xWtaVxuAoAVHayesVNc3YQDD2VHvtDMRRPDFGwzAuYpW7DG84yPi+mZwijYBLzf+
qsrC+Tnpcwvyt2IyDlrVBsbJITDI1JrIcmaPyEu0keX/BPbCThTyTbnvSnoxj5m/
CurMhxKrJaPvjo88BLPFKXCiJVllq+1ENPbbgXrng81VzPZzr0sjiJpNd6oWmWNm
QS3/WR6xtDAv84EWWUONDYm1yLJ2JAfxF5pQkil+UsppBd2t9OCbo9Fs1nYV7nCY
UZohuRPtbOjsC1WJfjbL41NPPWrNlZQ4na1Q0iWoQt3a9FoPU3GNRINCtcLajRSx
1iGRuaeslTVkp6mm41kF0jE0XS1mSxHNlMVNyXLZXpqk5BAPibeev7Vi5L98m1mv
5jF5Bk59MT+v8/UX+gdXhK7Y4MCa+GqBaiM2NgrTcAYUIuLBxnocpc5KKLVY50j2
qzhH/jRUNHsqaPpv4wwmktL9ASkLd8tAXL/2SBX8wFzalP89ZwUoAePaoEk6WZIC
HP+0VY3WyD6xg3h+K3/BVw3UORuxqFbDfNa1XeCgDa0LFn6uRFYt7o6BnPVi/IqJ
8gpzSaAFW/OPUemULC4BJ1YQ7lev8fwrHJMv8kz1vzBaLHNU94OvD8ZXhrC2N2o3
qMYW3W/JfkeV7fQiA9uVphRX1uGBjNFp2L3BbrOeX18DNIgUthAX8jmBun1/B+NC
0O1N5i3a1ZxfQ6noy6YPRhC3ekFfFCs56O8O1spP+6ef8GOzQmvj6mJcRiFMHUc4
6J7ZMBl0TIiyjrcWB3jcAqvemdGxK0oPes/Cx7byofTMsC8NCMJdRzfnOhrv9A9R
EYjIsQjslQeQ6xVSQob/QqJ8tulouSoLD228sUievfRBlbbPFW33JBW0YC4uRy5p
vyDnccRMd3aY5lzNL22wRng3dx0Ps/TyFdFMVKlYYJdFp72+z8AIByMTszeYruok
BrKpw9SEJlWQx5NxdPwbMfO2KoE8OfHpc4yJEP+XnVPF2yypXPEcMiDgUAr6y3Gh
p/fnBfBYZcO7U0QzRf+RO7p9WhZ9l9EVgL3n6Lt2mF3XA/U1+yvRwcJKdQqmc3F9
eQGhqT5uqdClYx+q4OkX6aguj8sdYL2vCx0CfivsxQ81wS+IcVR0+l65xdvGI+/I
xfIrkH1FSxKqznpZC/IkLX9pdVIn77c62Xk4QAz6+2K4gxYAiy52OCPsLK3L12He
bhuF10mRhfNvoLoeZz/j+DAmaWLuypfJu5sUP8kaCkviF6/UeB9Vk2hT+/nWLD7w
LiFDDozuLWXFlFGuEu4XJTn6yNWUlXM42wXhe3LMYZ0TZAdNG9ycRxQL7Kck7yWF
pFPfrZSi2CjWQMP42MV7tlqguXKJG9Srywh0W7COPMv2oBK+2jrt9OPaBDweLQ4u
jPSqNGqbLTEvKTeqnf8CFjmJoBQMFeWPa3P6jfrAVID/K10nq+1CTV6H8B+W4gua
wNlCdTqcLEBk2mqIvh1TW7BYnWJcqZy6k8yOPiXeRWdNIB1Bpk52oF89FQQ5pedr
/CBenBAVnLN+YnQOrtnSkrcmYgK9naKN5DdtJxRc4gGJP54z4LEAu+2Cs433LhVg
4xSZUKRSn5fda8rtS19dSGOXhLTaDq06vC/KaY3PmPPKmnIHrHd8Oxuy7WeNB0dq
jY/kKrekbcNkuc27Nh7AEpnMr1o0e0zTF7m9IZM3jjD58uR1h3RM634aaLEhu/T5
o6QZ3366GQQuJv9A57FTGZcJ5b8ZsgrZr3bwfHTNNU1qQXOlwkzcC1VMEqgjoXSI
ndToQqQdHGK56Pe/EgHKGDs/hfcFQOsap34YF4C1AhhAK4lbVqDSCAuzFLotU6KR
0iKc8LCzwnSQqWhROO4x4LcSjTyCoM4A50vRrH55MaSlYSj6zy6M0B4iH9mVIU/I
tG0j7t4cB7z6c6gLOz93OEZRwWzUQIbEftpKmhGesjpv15ZusoiD31119TRIexP9
DkhR97EAuq1J6g0PmQ8bxbuE4jaaZHJrFTYXN2yVnmCDIYj5mFSU/EYQ7yc8qF8H
oXpAJMGNf4Yy4Z0mPMaKkkv1t+V7jzndtLb9StFcNKMSPZCs62gic1fK5Voy6xvR
8Odxe0RKBHPqRh+6EQOQA6txHwEvXcEVxsXFElwblNsuV/jZWLCWy/riPB44WAX8
f5BanK/ulHiiA5nQkzuwrmHizLAMLaNPYPwa36qrapxtJqrvnRAglQnUsPqx46KI
fXWK4RaGd5Qvpp1wLLEVmOzGknRlGbxpFf78uc9/TJBYm6CedolOgGWJLMdn6Omh
EHvnmMejV4ZzT8SH2I45NVinEyfuiZFobF0aItCdoU4DVheRbXDrdOGOSRe5+uSy
wOtIqXubzGyQehNfuIeE2lh+9wFEQ2wqd/wfAv8uzsccLjLJAveDiO65jr5SUHej
XuyPUuSy+ZHLAS5Xt293osOb068BF+UH/ZxQGo+I7u1kniVk5W2NZb+K++RMOHj7
658Fx16zH6WHVQgzlWWAzyiaZw8zEqF7W8stPZShYQcPTI6z+2en2IFDHQkVKAvE
vLCYE4MYuwIdQltLbY16r7m7I3YKJuH4pmV53rSiQAT86xFNKrXN9IGFVEWeIfI/
KKBym/4ZL17VaUqFZB56uTV1cBco/Q/gwG4HFRE481wVAz6tF+rb5qEm1P64m8e7
w3DtO8YgGmHp4xNQ3tI9JXIiHM5/pLzMYlAjEvWXivpgrB3VVz+leGMmqlhN7EP/
3mknl1Yw8onlYFT5FangRBei1BHjYFcD+pR3aGJTVH4AbaZoRrN8Gcj5W+XykBMV
P0poRLNwXYIA23opPLkevpZXKebSJk8cEnoOKekZjqRH/ZihDIF+RlTGXv4QftVE
i5IRRSwlZrvvOW0GcKv/m16ljYIlCxHDLHMT1D8iuInc0UWmwKKO8LPfeEcbHOvd
oXabdnCosLVrawFRT/AI/LlF7YPRoxyg7FQ5G7DgbMpB1bX+3fovwd4fUF2AFiJP
ZtoBxnnaip7gnDKz1yvOMud0iQyXQvFQubBsD65+9NzN9PGUoy9LHSyqf8Cm/gJr
LHPcU5PuLGMw12hifcdjH9uXLqkHLzkuWKk70dWxI/W1jqf5dqvQ8BSP+pGBoyIX
hlyLPRL1pK8HCSGRmu5m3MYBnRGDRJ+rlel+MXrsFi5PwV7E31uSVVt60M8EYXc2
Dvs1vXSyGRFE/BveDQFC47uQ/I1TR3XF5vTERq5OPoe4tJOMTGwtn7uNSnY22iEr
+xndX/rzxUTpJvM9p/1VbAuFmkFfkvyhzv5bMEBn9A+tKiUE5aAQhuR6B9XClsEP
AP0WTOkAW54j63616poKjFB3kLZ2SPYKbniUX418bfomrcSodLd5gBe3mqm98DYA
+SfA83C3Qf1FF0pSykjsRe5c7w6MYDGxQIUNblH+Bw++BnxzhRNfqeZm2UhLDMlY
jCwovrR2glO/qywLd+zhDSB3UKMaFy1bcNI8ChHt++eHA+fOxtuvYeBKQYRFEJpk
sodCiurXxwZCQgqUUpIlCX0NEiOQafD31hMZkC+k8KIZUATr+/tj0ysK+a4JFbLx
fUb3TgvMb+1ywL/phQ7Io3nut4hY8faL4bj4qD7xHy6pfz3Bi/E1P2PUY6/3bJXq
GOcJGn3EQDOor6gQID6jsM8BHzSdpjxq630N8LcMUJtH4zIjSh3RRvIpB39pHtpY
G2Dcf9DQYYsDq1l4VHKnQEa0Aodw4oNhK8Jx0gwS+hj9FNZJFDBfAP4jqLR1mofo
wNa8CAaLfNToJa6wbb1ZLPNy2D9Y6wpth3URPIMJMW3RpoSUvBrbZ42Qv9VcHCCH
0kzxSvg4PT0rSBbiJGYkv7E/zHKDVvkri66expE6KeJZJ4i5TpVtsoblMXFaHVY+
DtQib2C4An59orTWM/Ju0hhnA5uPHVRfcCGqF3/4JXnAAxOtCY1QaryWrViiqjae
H7vkqZORtA20ypE+ML8VzC1EO8YMsGBMSbRAiNfUkeGMPtmxogEBXg6TSWaaONpp
bP43QQSKRG5dvA3OfZzwGIM2bVhK8K3NkN3DQhvckHJImwi4c4M1bk9KeQdKW9Zh
ggYqu0Us5CJFuZg30GV/VKzNGccKif6qeEOGwQNVzpJ99yAu7rpmeVSI9t+u9Kft
QjjOnricZ7XNGzbJdf14QEVYMoXW/cGV7sQTJ7kj3hLAhxv9Ur6Klx27vRkhPNbI
Pf0o8w8cXBpe7SI79ZRFuBlmnNFDJpoIzz592DvOofjmFRgb83j7D5ebNZUEVx1g
Y/3PD1jw/1BjMtLMAJxUKjn5zvQyk+9bPkirim08+l1bpwTSE3JM7g+HJHX4b253
ZNEcSpdoMnp0sdCWPawO1kfYlMiNA8zEOtbVT2qHSX1pgh8teFmS5KBNbXzS7wWD
Ly8+bYzIw9epjqVbaUfuTIrWSNfoeDaHPGIA/s8PvTqEeqvWedEE/yoltYYHcY+E
4V6ATUAWMiUi4WsI9V1NjNPMUh2AzR/6Y+5pLKzpaKk+eK8fC+9mxNl3WE+505zN
3HtiIzeXRZEruucICx7KwgcLe3Zc5jUAQUmL1Hentl+37MMV1TkMzFlzwpInxQ7H
mGxBmU//7kDI45kDGwcg+MUDzNCaLB5dlsVOBSZ8vMa2/8II9ObtD/1OrIBTbubj
9qHXyjceWkCE4eYB6uhZP6W06HqALRxsAhc2skOvC21oh980SaeV59DnoVHwrlJB
Cz7d22GAqdFvLs4igtU+THEXxrNIs9bratGdPwDN8Ttj46o8F7Nk2bxhAp77hwx+
bKPxbrVNQcx3WtYEMhdEYzyG+33UBpB5Mh/DME0m/QoAZIpZAM8B/PwACDC4zz70
Hb6WC/lb+jXBLLpIFFJzI7Psdn1ign6xoYexorUCa+k8vTzMEDd2MvYEv6YbsHSF
+6XhIBTUpm1KiLaEdQ4so3sKZlesPnv2HkpMAMZiBCVzUmLafKL+nZk2/kAXhztq
T4gBqTb5tFgtm6S1ia1yklQC0+DePpYY5/S/ger9lgWD43nmm0k4IZrRR9MasO89
t8YRML/MKxNGEC4E7jZ1BZjWIAd90Ap2tw7Wbn9RvOx55pQSFp0JzredU3OxOaP6
6ZV4V7SrPQm8WiDrB2DCpzgXF09DCs7yxsw8Bo+n+6w5uWqQ0O22GEuXY2GBx2Av
XuT9Q/U6fAzQdhq8hAIghkuadeUG4nPbSHt+FlRAyI792j4EXBJHweWKl3nh2Ru0
9+oUUSW65bGgfZeVQ8Ml8H2Sa9f6bBtNQ9Dn6CWZvD+/2QRgdfpXv43wFPpR/mFv
6/vrGgjHbNtuTXqRYVSMXXyCorydR7+7Q1d0VsVIGJPl6T8HsJnIhg3ofCdMoB/E
krPV5JYnMTguZlH2EblFVYkExLsXq1viqDiCY/ydazCzsCDX2v7a6evlswTdF/GH
sq2EQDlWXz3MhyzQ5K4XLKTmtL7i0Mqr/8khfzrmUjMnNA97EUnGKvpeFIs+Xx81
FX46rqzzYjdRRkT5Pf3D3KmL1VwnhgAu7eEG77spUmbwvRrW9EpgKz5VUg4F0eED
CqE0CCUtxsRtpvLDliL+h5ZX0NmAwCzrqIN1lCrgcBJPiQMwwdNPVv9MszTc9l81
+iXaBXTcXvJjb5mlwRNbgb5GaSqS/2lPV4MNST4aNUHzAR0l9zPAlhpaJION7OzX
SkKCPAJ0RtuduS80zBWMtVK/R7VcNQ21OmqsXpwfdnWnUwlNz/UjpPrLqy9oQKcs
PLQOqPxYrAgdKnF8S5pPqMYoOI0Se2AUS1xGnEuKDTMPQZG/utVOCWEwwDWCdRWG
pOJYVVcOh427oMJdqDr8zjYJRhnuNPAuKdM7wahK3iKNseHii5hqfzD0l0hP5uAQ
EXpJ1Vj2dby5beBXv0NRUnMJHuwkQkEkXeMTxNZyRrRM9vPhV2YQ45uroli7zSUA
F1wXWVyh84h2/GLzFcHbkhN5oN9sm9ZOW09azPqYR02iGCkHj4olle6NKCgZ7R/P
FfK2jofO6/tMIcTiCX1fStiJLv/ueN2KZWSttHAhyb5Sf11GZBg1xJMiCkK0vDKH
5PWAgNEq/2ZzAu/3uXUj6hadOXwuJk9/5ZzL2UzXOnjOe3BhxsF3Lzk1Ks4kj0mO
Ax/wpj4fWsSxenZAwkqU+fJVvQqEhT6IKVp8BoS3sy1HQGDPCKZQBBDikyxj1/7w
VXvJfQhWUvwbqMeUUj9hmpw8o+ElcjEG9Jl2M9ehvbqPLRzHU58nvkiGmuuJCOI7
1XFM/3ATTG9jU5gRn+ucuo+uVAy8Ctiehg7FWTJTiz2RtIaLEbmkCLUpSGnYb48p
aeeNvR95MdfMOLU+LuMyso0kWH1i+Usaf8aZkTqxBj4=
`protect end_protected