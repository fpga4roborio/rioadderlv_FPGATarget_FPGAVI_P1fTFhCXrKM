`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
ddtXksX2+yylW5zu6QL2Lhnb2d1sD00763mmSITNX595NcHTEkwn0zB1Dry37fOW
FufOhVzEJp80NC5qZ/+F0Vk7Ik02dIR0elf3clrjeJRK85K4e3Hoo4xn7YbFUIms
l/8VZSb14+JVGURjfswrIyCUotIzlzVYZ6gzoZwDXIi5gQIBf/gI+KxNXPaKV+PQ
Ufys/12rjO6aI/pPlqSm0hCvftmBcnezN2hk1UeXgOIuKZnogjOsf0iJVX2aOOWE
6pD/psybjbnsNB6kH5uFTA5frkzIzkzl5d9+YDm9OyC+k84E83I/7/j+rk4L2dah
QJOvksSIzN867/4Qt8qYTQ==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="MvBXkzurAa5VTw+1JJ70nePUfoQXBvZOku/SMmg4TwQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
oRtzZL4VJ4iwysPsC8SXYCzXS8Fw2gtZTOskLcDV+1B9Nzn1zTyNtlo6lNICRmmK
ZRVu2BmCc2G+fmzynYlNTnSa7C0Cuel6FYpxCBlOuk3OF2tzAmLAuDyOH3Z1Yjzk
a0aHuoCdIRKv7BrZCdALt03JeUmXKPdOmIlkVGFl8yw=
`protect rights_digest_method = "sha256"
`protect end_toolblock="Jn9CQpRhJt4rnzZPRk+dOpzAubz7omckX1MrFd4p81o="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 5840 )
`protect data_block
gD6l00tciPUa6pDNTk/+tzLxvdHE2s3DQL3/JqqujQBC/Ei+vcAB8wM3doqg5vTg
mdfn9XB1bLOis2CVSfu295W2DNwHfMSTc/8BhCDRnTlLIX0UCJs9Za0+LoM0rMrV
T7EjVWppbP+Em6PkVKCwlmIQ7JKaifJ+Y+kjw9HCGboYo5074hY+K/CBbfsBQY86
Wmb41iJo9ZL6MITKm1koZBdlWzw1PKuHMSv+U/btQmDMTTPCyv6o7MLUHAcxOhcW
8nVqaB57uB0+mm0rOH6S38aAJm+M9ocjMZUCDPNLwsrmkjOj8nR9Bbd0lMLmadYV
rie8z/G7aDOAR/+r2glJ7391wekvgFIShMvxmoyVE1fFREvafVtZj9dnJAm3VLsQ
tWYKlBt4D/YDSL+FasJIzq6j/+N1fnoDMH3/MdNE0u3TMLADyJyO2l3rmvxl/rvB
O7cxen6q0O45ygMp2bsZizKbWhtCywcv/UGD4VPKdV9PxX12RlI31PEhgcjUWxtu
bCYYQgZZXY5Ucl/4rz0yv6gD9dUgs0mG288vkywliC85t3L75zIQkQMgKoxOqORJ
z/FlfAaMpEGEw1pD7ga0cPOSD0piFyOHq/tc3+p0nwCoKgfI+teMKCuDkCS5koTx
1byGqny+8r7iABbqHE5O87tDA4CA8TwlW6jvlxNKwtgCP2Myvjynd/2W0SICOgAR
X/eZKPQaUlzIEoXnG8mm4fCgX2lrBb0seKRBUD0kiYqE6jXGwGvHGEha4c8LD5jD
jXtpLhhZyGGQz0+9E2S2AWyNMRCpPasqoEZCSqmf/P/d3rdJru1yHz3IqVTEL4oJ
nFRnZuf8LOI6Wycet0iXL2jRWbP7fWy0QEUbUxs50/S6nnCUrpHWy432e/qc8Clk
iDvq13dgI8KLQt4fQH74n+S195luwtxT44GvGOladSWibE14uGiMqiTNokdMeNA5
f02W6gywzeYfr/wh4jzMeln4p3vsAih5COoi5edeFUArtrkdGQRpUxdDqyybALJ1
0+EMjX9oWbkLRMv3TiYOiBPoPjT8VmHZaLYOIYRV/zgLh4nwMUD6XXM6Hk3HulgS
RvNgGWq5MICdHb39nhHbyU1yytVMzPNVgmghZnsu2ME5z+iuT4j/E1uBvnb0jTc3
O3aJm9wz6wjIjfaSZnPBj//6iW/5a9iyvO1MGz2sxXhMdH20FBOgRGhERCwUcKdO
YfbgN/rW5md0xNcAlN0eh4vggNSVbM8OBf8OzVqocPH2G6Gf57CISFS8KpS2S2h/
T4DhgQYlmLL1XFXsvjkg+y5jmZTPiCbcj+bR9MFFxJtj8VxsKngOkdAtUiF1IW+i
gV0uC9eZ4/R4H0m2Y9hnGhEbkACnF195ej74wpQuq38+FtEraWkQP1XG7zVGEvA4
3eXxUbhb5CeJPVVzFt3TYlZTUVOu9xHps1K8y/ARWIIgr5u1L0jM5w9yLNEdoR0M
P6d1baeYOBT/viAo8ke56dHEJrQaGdPSZgz29HFVqymE+Ei7GvoYhN/KiCUI9Lg5
arsNmP/yVeednkQmG+kE9KlkNgJLl4PI9LT03T4gmuGI/zcJDJp+K0FKov07NyxQ
0d849GHbYgr7KSyxP9FiPZ9dx3GEf90tvD7K4ZplH8RVVsZU7XUujcRG5AENpEia
8vrHVSQICLnjhg7Giqp7YP9keOSJ2dtA1hatnT6lkLrjWrUwzdiGxGpF1z1pTRNi
37lOhJzFInSrMpRjbwBP/sog4ZGYEJE69o3mPWl5BLAJQNjiVt8vBpNp89ySyCIR
YgLge2y3pan9NHfme90LBV8ZSp9gU3FFNdts2k0BzIh0sMXfXtPl4tdicdr5k8T2
nETxpfg9n6APqLZNYOl6sQkxw3rtLscx2SiJ0sHD2mUHSYktLf2w3RRyf8XMOaXh
4lBeDmKQU5XMU0qnAikSNqmykQKqWAbKLPB735LKM4qtIwhzcu+/gPD/iIUiQVY0
oOkxbOR9T0EDOlWGyuCS1Mf41J/6jvjaYxZDPB3QB9B+RsXTBQ6tzTamFuwpeaY7
BqLCbW2BzQQa9OZNoFt+f5v3Rmu9COfSvfNmxPKBsTFWWpvIOcCKKg7uaPn5QqJD
/AfgphqGu5IEX4CG1BgtxE2xZgERo4v3+XFH1GkUfY7jlgiR9mS+nZRBW21d8/Ky
eGnLz04n1CC6M+6zZ9amvbFMXV80WMyBnsWQR8Qd3nYC5mllXHzzuVjfrAM8zxmB
mOEmxTwe80yHnW8ZmRAVXiRPHdmFoRAuRm16BvG4W47nw+leY45qWoQD/pjpa2am
gax4NkWxX+3EsM6/JwvS6MU0pOLurDn16aSnpAMdpy8b12s7W9dQgHEBKi0JDFFL
yBKadCvoouK/amvOvnxRiXtttyF0SOJJ0ty8Gajj/R+uxn3+fD80MkuNZMqWfS19
p2H64bDmaM7TVWqwWdeQxAr9Vn9SzO1PoOHfNzFR5uyQtslG39PzaTdFm2ZD2nyU
Ry4K3x/6ORiUeecYVxF5szUV5Gu64fz1rV0yOqVs6KkdpaGxq7oy0MRqzpD+RYMC
VNpb/tobooeITi2rGLZl8mweASbK13R7tnEUmko7nxp9aOqVclkbsyHUz06nLOGD
cGisuwc9E1KZxw4/4s5AHxO3CPKM2yUpfW3nqlkreA38imnt2VNCQpkn3getTaE0
EQvHt/RfUytU71zyd0FQHUMfRTAwXVQsZrAvMAMd4ZZqNEXsTflNby2oBr4quo+u
teNar1Fn/j3FX3qSBlcaqEdEcrl4YwbQVjY/2TwMBtq3JT7oSzfHdBezKAHiLBDS
bInvRWfJnGCY2MGYX7r6ARoncBHyd02qfAcM60IGAHwDg9UTmOgkMtDhBfQ7PlOO
lU6wyIZiR8gyJ5CWEqeuqBJTEFnyM4B5ljHkluC2i3dmGtFjaByRERHDP33jED/N
yevR83acRFjCslq7K5zX6QQUjXJZ/H9IYlAzwUHeByPjObqXrreqT91NICaCV2SX
CbMwuemJ2Zp+EIOy3mYTPKTzp4SdGAu2Klu29aSqAmvgFGhsM07MpAOPoY13t5WI
vvseEpNJ7PW07JbZ5Akc2Mc3IwqO7/qKmklYKjdSwBJFItN2O+TjX6/Jed9rdvlk
nIOPGPaBfetBUuO1XrDKYpPoUz+7uGr7fwol52ycTkT3wyfd7xg08vdLkn7kzWJz
nDuO5U8xiNZtFT2k5Maoh0DooVI3F8BJBh3DZZq2JhUxTofof0FXJSbUuCmak7WR
D7finYLneWBfN4OxAMkY3OE48s5eONHCvRwnzJKeGrr428SAfx65sQKcAARXRLWd
BlyJTGlh+Yg+/8RH6N0ZL+19HXE2hDYwUyz67sVdW5gqF9rA18MuuOSibDA1Jl5l
KSSoIpmnUoFT9WsEAd8PhPyPZ5RPaoaNnyurd6B8iGXrrtQPHKX75MBEqLYymDua
CwwBOzG4M0MdDkIY0VvK/FWcN0kYnCrJjla24kPi3BoSSWT8CFhk+XK0+aaGSp2N
pPQzmJruRSkvnmLP0uIxG/SPR9V7v5XVN5Pnb+/cdP029ISoON48QPadejO2CnsY
T0uwpnkxkxfeSHvTmpfPISNR1CzYmSqh/GYy7OE/34q5BE/tXeI0PK0xAwGGluzo
tzmmtpZRJtnc/Qx5d0odHWo8L27Jsl9IJkKm52zsQO67BwRex4Qc9icQk8zRjQvH
RuYWgVSDfGm2+EOseXCJRBFkQEMFJ7Bmh/BFLIfntvDn6Ey5WvgHHVgHiHxwzI2K
+sLKSef010sSSONY9zDzfUoIMwjq8QHV2HJX/qGGgrjfb4wsP9I7+8oi4jltw8t+
1uLVAbpy8zowkejwZvJQccjDH4ZpXu/+XCi7optrvtQSjVzsMawE6NZyre0/NCcz
jk9PZPNmBkCb22TXAJWVAH2pjMcR8tRiMFoLD6FUTD76mWO9oRgVNBu6ncET324N
2xjwdL0TDKTxh5Gznq98BPlXxkrJoO9AEagVMvLwrL5PnS+1gmbZdEq0j207zjHV
4l9sVwsTPD0gr18iR0xCqK9HzMmT0dYkIHcClJyf5paNH+nYkkKj3rVyqiDZOaGK
2biax3MzXDnptDnaoA6SE5/NkGP572dRDfWSGdZadI6Lf4vqLU1JFQ3jm7B4N0CH
zG6i8+Kr5La17YJGNKWNvVOt0hHlId3mP52/29Mx17A6upS59kR5a2qMnVyvoY0m
6/612A9skQXHV2vJO89GeRBdn1cWtJP6FWKscDoA2rzpksalbp2i++wVUI8k/wba
yRia1bd3qxU2Yb2tmnhlYruHc9a82cyNQrBt7cT8KC0XRYi50qHVwUvrh+5iX/qv
+uoddy2IwbWBSRI3FrbB3CF+o9ERPsmOprB8nZwav+3xTfi9JWvSVPbe6fXuQHzN
48A2BQDukeuiE/TlAHI+oBz07lbOrsyYnycZIlOQgPa1bOVtCJ3XX5oZQ3q16bBV
YFS5IzEXN3KbanX68vquijdF3bTm3ZtVF+UtRbfvG8S3llfMXcaM4tpK5krMM90i
xdX/TlEUTqjH9JQ4THW0tPI9RYpXmQ0vy2SHs0i9SIvUg4ycIQloezmQGfG1XUmf
8UjlMO0iGmpHPxtLBGQ+RUorM8Le8LDSH5TZWa8UM2pJjhJtgGMzs02bbLwt7m9n
cyvUc17R3PHo/EP51TcWqZqCAGP59cjfVG5nT1/FaX+D2mKqiejX8Svg6VXG/l0e
efuRi8CiZREifN0R4uqX9sOVxGJlmo7G1AzbpaELh6Ed60drob3SVtafrOc+6N1w
IBp1IRxtbEEsqFgmxwf7Ra9Vn8Le4BicFVKEjQlIHJnoyyHFGssGrdoVNejveAof
OP686ZKyl562PcUOAb6Xke9dhBU/G+MGFjXuUUx8oJfj9g8bN9nkL+EgLulFgtxh
APEwTNLJcYzr7ajJCJwWhY75UqCS/TdQCezwqUO1p3nQIWnpZzNwq/UwyMCf5lJA
T2y5nu12g7w332v9oqf+1NJf93qVk0g1He7zTl4GsBo6IrT4s/XNx+8aL3cW3sA6
WxcP29pSV320CegM2547ri7DUt3L14s11v5jxZPl9H21+k9MJMG8GOY+Knf1RVyK
2EX+PF8pW0HOTM9XojASXlg8BTgbOi5+yxwMv3PmtWj1FzctRK+2IetoTaXMkO8K
ZjNhJghSYI301B4TiZKct02w7plV9kwJLMlWSDSUvvEFwdJLyhvge1Jpqq6KSzew
1w5gkfeWW5j3YB3dbjivQyB7L9UjbjqZVaunGbLNWPA7ZxOSrL3D2seM+Zaoh+rO
Pz83b8h8teQj7q+JU4DDcjjNU/I0EvucE3s6/NXUUaMqNMPCr1KHRdmmml7Lf5Y6
rm+3rVkICU1YkVpO99NjNi1iI+CPi2U3rVNo4LdJp3PaThdmrfE6NUzMDiPHUYPZ
vMx48F1Rq+HkgOgpBcgfu1h/4dd39cTlKvQlxaYaUBMwpESuuLvOfhcFOq1Pc7AE
Hl69qgbGjIX10x7639YMMbUwLZFoZO+AStb7ECUby/tDnNlK8jwQ5tUQ5UTPyM7w
uhZHEwfndKn01Fq+TFV76fxKGgWBwEegl5qutVgbfoy/AsALdCcKTAe1SQS16577
M7aqQX9d/lgnHkY2P6b7AvQX45Fyr9YlSDz0r79sp1MhfbExeCwhIvwn8cxzV4m6
WfCeJVjrg9LvtldvB3Dzs8vnA1Z9STeGAQ+R8GMJAPvK2fTjCIvJb0pzbgDGdY8C
PHMtMk4jhN4az6Yl8hJ2wNKbWAFwpFYwLxQJjOIlhuQf3uDzahB6qkWqhpGRpULR
/gYHaqvkhT2rvoQaJVswb26arRwUhkpxAlYxh85Hq7O0C47hxwgtGkMMFgQnBFmF
p8eFs10kkKDYY5uFT++WhbobasqSCHymexXiNTDJXyVZduR0bsYGM6m5JnmGueXS
0UHmrZ+IWhLu76SqEv7rifhaAfWy4MBOrq34d+5rIpqL3E7ieVPA9JER3criTuAO
/03fWNin1oOzcdYZfXStffyjoBo5jhbksZbsJpfKkouOcP8syl5XjhH1oUg03TNR
cxd9+28lXQj17pxAgKBZXHnB5OI3t693RAnxH3A2Cy7IqDXh2ut3PBa8uIPg7eYM
JyNfTOYym8bGwTeqYF0YMYZ/RdlOpWQInVTrDtRc36RdtqbZAjew6Q2M+3LAMxRb
0tpmkK0mNuSGeLXotJhjdB1pliGMxxDq11TrSgXPojnIKN8y1PjK0SmU7jjAASkn
+1rMVjZrPCZgx13Yw6AL86SKh9NsOD7Gglm6OPkFfUIrCULiEn5K/142c1EGL4bm
KILdPIAmo45/+pmkFMweFbl0EjtarBmpFsckJB2EjP8OAKxSoJm9PcqzTuF+T8/Y
NTT12QXC0lRilU9zb99PszehiJ5vH18iMoAcg1Fy0QF0h/5QbIkgjZMFpSm8ePbg
0Em9mcUXFmq+PNb7fSdY3CNCO9uUWsYP6udsSdksNaUtqLyyZfU6E0/tvjnm4yGI
LzKXfV6eYbx8zNEYEREgCcnLa4kc5Hkw5ji6hZdyCFpschqbzqb79zu0RUNdxFuy
5QwBuYCUl535uEpnO8PZ2ue612AYoUUeJ2a5322qz6HcSQfp0xbwmijDstnNc6qh
LED3xFuTh3v3mp5zkM4Vkh6KySXn1cbxHoM52OqUi+U0h3jTMSLF5VQInsnley18
S389Ks5IR5XS4tUQpSiLs8Pj4iOpb3eZzs2QkTGKivRFbYvwD+jX2RYMT5kY6imo
VRiWbm2ujenQcuLTrZeQnp9DwNDM7jnk9wD5Gpxh291Agzouor5eQ/AdtZz7PWEC
1gVfIJCznb3YYnTE+W1vgtX9sZDu+RWXw66cCc+zbhCCsKnZAoA8xq0UVeac/14n
zQvKNX9rfw987jplg3L3jWlgk55qTDuj3pJoB7NBVfQF1fhX2BzNXXYsEpGLYvrg
kql+XWsSY0v9OXxCLIf8ts3kkV6FwZHsIJ+ds3j1Ml9v2o6qNCFj9fQR+Qaxgj3Z
XS3J9MfbsKPp/L+9irphrJsbICzAJhUoI9FfsJBe+sPqxRCLMn1Kst63QuJknz21
omdJ7SR5nXw+hJ4SXfuF9dyQ4dN9rY8Qy6uZzIXv6xaIdbBoE7L4VWpocp6SLzKO
8Ld2HGQOIzjbinCABuF3zZqWneW71sTs649iiThem4+qrfZj2jQ1CUJApgIVTB3L
x6TwYt83jQTvP/4U+VM5Dpjx+N3kABKZWG0gYYV4dXytNGAznHcVKZGycjIS8z+S
tMKPuwSlk4UlK032smRAIFDSc1feOPomyEGtGfwKUa4pSywC2d4OwPtX2xAgwKfu
oWCscm7v/sRnw9AF21uzIszJPmaVQxreAgZ3cAQ+jw/9Nu5gDP5hBs2plCJsxWaV
72Z+xSa4dHNehhnN9o8xZJGPqWMP+5Day3kPNsQrHj1iN3gWLGVrNDgr3NliY8/X
ZimeVz/8XZ6HeMyvYi508JVarfyOahjdGD8h3HlHmF1pcB7RYnB2B4uMQpE1DDYs
eZHZ40EDDDN+ZUTP0n13BmCElESHMUe2oeKtM/9TERuV335EHdjaBAfHlD3Vnl0u
vBaJOijswaiwZaVY0CpcXV75uC+mYBfryWTrC9LDQqfI8vDct6kozBmL46QDFFvQ
B6oZZYVF2gNYW6kkjo7rN+zRBeKDFsU64QkSnq4mPLeOu8Xfhmb6JWiAp5p5LkoQ
lLa2idD9RSkoR/ICIJfUslfzCebbJs4/r38d0NV/M1Q=
`protect end_protected