`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
ddtXksX2+yylW5zu6QL2Lhnb2d1sD00763mmSITNX595NcHTEkwn0zB1Dry37fOW
FufOhVzEJp80NC5qZ/+F0Vk7Ik02dIR0elf3clrjeJRK85K4e3Hoo4xn7YbFUIms
l/8VZSb14+JVGURjfswrIyCUotIzlzVYZ6gzoZwDXIi5gQIBf/gI+KxNXPaKV+PQ
Ufys/12rjO6aI/pPlqSm0hCvftmBcnezN2hk1UeXgOIuKZnogjOsf0iJVX2aOOWE
6pD/psybjbnsNB6kH5uFTA5frkzIzkzl5d9+YDm9OyC+k84E83I/7/j+rk4L2dah
QJOvksSIzN867/4Qt8qYTQ==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="MvBXkzurAa5VTw+1JJ70nePUfoQXBvZOku/SMmg4TwQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
oRtzZL4VJ4iwysPsC8SXYCzXS8Fw2gtZTOskLcDV+1B9Nzn1zTyNtlo6lNICRmmK
ZRVu2BmCc2G+fmzynYlNTnSa7C0Cuel6FYpxCBlOuk3OF2tzAmLAuDyOH3Z1Yjzk
a0aHuoCdIRKv7BrZCdALt03JeUmXKPdOmIlkVGFl8yw=
`protect rights_digest_method = "sha256"
`protect end_toolblock="Jn9CQpRhJt4rnzZPRk+dOpzAubz7omckX1MrFd4p81o="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 2896 )
`protect data_block
gD6l00tciPUa6pDNTk/+t0OO0nC/UTtBwLB41d4inuAUA3i/ALrNyoJVcBnAmEQW
ptbcNp5fxEUJjnOxnedyZEuEBxWRieZFQnkRdF269oOdA73JuXggf7O7Tl5NpItq
zIQZUgZPNnjcUXJXYQwzMUmE8uBf3IhZr3EsuHUlKISZpAvIiwUg/nODVNRJIQLG
wW9ifvVb1fXLR/7UwxajGZBP5u5i1MGzkXu5Jiu299LpMih2M42chGW5SVN0zDRV
RpY1fklxCbkl2GDIYH9TnUagj/1hwE33+v13VrK5oQnoBdF6T8cNiVUsFOJKCmfN
0RdwjAnErYZSiY7SxTEAey2QjmFh0AvDCbAeMP33zgqJpoRiVmefk5zSTOR0UnKz
38flxiYaqtAYwQAHEDfmwMq6+tKm6f91PJ6qv/tstcPRgLVULkRk0MJwjV4Ra0y1
/39HyMb/TI25yG9mWfrJHzl9lBsofopTozNqG1dwx8C9tZ87WTtc1tSq1JXg9zHa
XROMOuJg/ysGge3FCfw7V7QBkPj9EhX/UbpnzcjOQ1dWl5Ds95tNJzogP33ndMmE
M89Lpd5Uv6lxZ6+8SepQyAkQ4y1wh2tXYrtmT8D7+5V9C8Y/Ed9bd2uKQUnVVpbO
lpn0Ys6NJ5xhrHVEVx/J8ICytlx57NsEfjPy58eXx4y4aLZRstxkVCRCadRnEV+n
e7O/cDD9bWM1aBfBLAqwuSBQTmrQuvUrpIHW27f5Ea2eKrqDJWHQvE5z28+a22ne
R6M07eVS+h6voKi1wr1jC+9TJ/t88CpeXIbNp9/K1bWfu4AJ+11+GyqQsFKmjrgL
0iobZCfndqWJRuLQQKLrb/OMXAa5DUcloAwkSouKd4la5p3QQC41znQx0FdnjIvC
MuqhEyqRuzB0sbzBZ434a3k5/QC+/tRAa8SQistPdNLZW7vp9WFFA2l9QqM0cPlF
lQJoQHzyhR7Gq+Q6DRP0iygnRBBp+owWxVBNf7YFdzJw91ax6wybPyZrXDC37S3v
cjxoZZFDWD1twPj8UCmD1fIa/HNY21lK6E8XmQeGcODfXsjOTuLYuXz4nmMHuHBj
0piMF6HZaD+V2MDp15nr37K9AHsGk7sK4abBskiMz+fGe8RqTDks8PcIIaWZN6py
caUKm6eM3h6E6FJMxHyZtAqvecceoBqmXT/e1kK+shNMn70OsyLRaeTG96xUkvf3
3/1Qr5vCN+RlWoNduVE4keOZCILh2Q31Fmen5kZk24yndBM7vKkNO83fS6b5XBXl
vTQVuNwBMO+3Yc07jIJTDkymH6ZVzFbo/0he44c89u62W0rj9bVe7jBkYuU423dq
4w+DDqF9fwkmqOiPLN4i58Vzq2fQOK3hBNXhwwv2ulPQBLkKmQRHctuJikUSqr6c
KFtgqwZJg/YGCwCHztwUJGeCiU0FGqFXP7qP+IzcXWJbF04gRVYiyBFTOhHEsi0n
eiv3Ald8kIuL0KbMopn949DdKGeZdYNMqMpI+5vTf0FMyE/RdF+kzhG7dXoC2IkC
LmELYM7Itd42pBInVvAjpTXhKoov0cHuUW5IofmCPxjZw6YS9HboKqmIK/9arAJZ
0h6Wowyrm45W6PDJCEaAVJwPA9dJMWJ12JiNwVEHWT8eQH6TmmEWPvx3RqGvmvsd
gPIN3rtqF10so/cPQEDxZF+5kvfortcMzAs1ibG1ryUd5qUbxLPoiAAFQpoK9YlT
/JohkQoo3xgPsKMuYvJADgg1cPnkd0fBWNjjobbaA0MFSNd0Y651rSS1oJMrZpVo
eYH6W33geIflaOmwYNvKo0H1KGgX+HVxnWq/hgsrQiTSb7CaVTTGhyYHQSz7UHNF
bc0xUaaueal0ylu0eWLKcRXOETttX+BW4NbM5i528M8yFqH58mJXZhaKiLtaoRy/
qkEa3jC+PTYjyN1eXX5Q+pLXyilXVrXRAvrGetDcm3XTZ1MCNAqwKF68J1FbZEmP
VPNoXgGzltmghuwRyW0TsWo+JxhkPg4EZGhBtTwUPLKPVyDkADT71+7jmdmY6p5n
kuGZyYLVaxdjk4u/7KSfnydmnYMmNSMxJzLTJj0z+Hk8XTumYbFfC6v6w4N69le0
pV4LCsVJO4lZz3FCAhYVb7RVGNnL/1gdFm1rl3d95glF6JJ6IL+ZkwniOqCJrtSb
IPrSoZ+KFbMA6mJqWbG7hcysk664IRdEv1T71S/Kr1LHTb7cbHwh3R0lTiz1rRG0
6V33iAPpJJJQPvCBE9zNTQDU3zf0AfgV4Z+shI6pLdhkGhcw3cHoSKfm664inaj+
rfiJ3crNW7CubHYnCYwYi5fv8uy5VTCLQWnmPnL/xnuO7fxosUkDwhIdcskEDP0b
4Pqa5Ju6CyF+v6AOaAziMQ0PeRekHK++J/dL4BJwRvZoxWg+ziHAdY38UbxwuLPf
qJBY0dueHCTBgJR+mNoH2Nn6gHSAkdBWjWUecl1pA8VCMK1anEJ/gQ6wGE6/4OVH
TXHVAtBICJk1NK7XJfEsViqXMKoknNpKL8duqHeiqXIxl60S9AZ9qWEIjUzwrONc
b4BOnuE0RybgdeNM0vfmxxiCwvZ3Ooah3awVfV1y8OsCUSKmkvqR7CC9MZoIWKL/
8GJ27Ap4lNjNyPp4huPKLEpftBE3TD3wN0toMOccfJzO/oH3WtHfIArT1enuSLKy
dpYsnIEdg+9uzVPBVyE5vD+5Qj63fLvW/IQp21Y5Y3uPJosbFgV7Weo0GmEiEq7N
pjKTatzsIIf8BRyuHQD7oFaGX5u0QV1NGqN4BLwxdcTUBvy4DTuGNxVsAlSV9DxD
Kc+7E5NM3UJypaIcLHfl7OqCTK1yklUt6hrSdrHlFlPTB3u8KlyybtOFau/JLxG4
N0rEG8NW7ldfDYh78KnyYPiOcYR3EeKlJyWqy0eWUa2w1UqK1C4JYxD03fpczmWW
B5GGDt5ZLzH90McAuxnz1YNsodzjscQzTul0CU1Z6CapHENpo3KDomCsFI7RW+K2
eu3vxo1WNEaVEgDCw6Yo6o88IXQbUaUkL1qVWO8+vXD40+XXF8yLI35NgGhewsFV
chORO5fUiky7zt3j9UEf6ZI33bWinoSMIRoOgB8sI1EZCj9oKrEsiCKB5PZbyLa9
EErLrbqVWDGyhNYtBsdr5hgHQie6fAVD27KqpTua9wQFu9wnHbmdIJs2YTOFIRT3
tGxsWj9fNgnB49IMwxZplHWxqScbRB8sMskija2p4aEhyYiHsV66hq2Fhx8NM0h0
OjBWDrWP75O/CcPLluM1qy+ucXZZzRobD3wb6NVmvs1n74BN1mOL+8vMoAvRLaHo
6+hN34dp5KUn0K+GqcV9jl3GOUAj/QIEcn8ma0SQ/PWYwY2AvG6LHhHrxb+sH6xj
Qjui5HwmUpcWfOi07SDZ6kgtYSxE7ed12eWJAZfZaERzWSPwgmA3U8tqL3hoQoG+
ki2AC5Mwaen6TgCs23G1uOwIbbT+qtyfMcWFKDZjmqTEFuzh8khtL3WBA3dF1K5o
/Telnh+LbJVsynoLMpLgqxELARYOhDv9mctKyfKLsYQ8bDWPhtYtFB77eUR1UDya
GHmCPbqfhSP9WubL43ZMwPS3DiD32EQkmDV93scjFG1E50YqWINPmoimamIhia0c
/90Bsw6BRTh0xh2N33jmFUpjqMoFH0h4WUv1wCBHYsgDTBfQ9LV3ai+RSPw9Mywt
5Tt6CUoGnB6xQP5WSLDY55BajOwbnz1XO+6xwuoSAgCu7t8thkkj03IftBKjWnLM
kDWWMv3eIlpRfMSnF4DZLzru3T3LvgO1VeHaiEyzzXbiMlrUhsLJwNckeI9tQanT
PkGPejafaovoxAF4B47JwQ==
`protect end_protected