`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
ddtXksX2+yylW5zu6QL2Lhnb2d1sD00763mmSITNX595NcHTEkwn0zB1Dry37fOW
FufOhVzEJp80NC5qZ/+F0Vk7Ik02dIR0elf3clrjeJRK85K4e3Hoo4xn7YbFUIms
l/8VZSb14+JVGURjfswrIyCUotIzlzVYZ6gzoZwDXIi5gQIBf/gI+KxNXPaKV+PQ
Ufys/12rjO6aI/pPlqSm0hCvftmBcnezN2hk1UeXgOIuKZnogjOsf0iJVX2aOOWE
6pD/psybjbnsNB6kH5uFTA5frkzIzkzl5d9+YDm9OyC+k84E83I/7/j+rk4L2dah
QJOvksSIzN867/4Qt8qYTQ==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="MvBXkzurAa5VTw+1JJ70nePUfoQXBvZOku/SMmg4TwQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
oRtzZL4VJ4iwysPsC8SXYCzXS8Fw2gtZTOskLcDV+1B9Nzn1zTyNtlo6lNICRmmK
ZRVu2BmCc2G+fmzynYlNTnSa7C0Cuel6FYpxCBlOuk3OF2tzAmLAuDyOH3Z1Yjzk
a0aHuoCdIRKv7BrZCdALt03JeUmXKPdOmIlkVGFl8yw=
`protect rights_digest_method = "sha256"
`protect end_toolblock="Jn9CQpRhJt4rnzZPRk+dOpzAubz7omckX1MrFd4p81o="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 11056 )
`protect data_block
gD6l00tciPUa6pDNTk/+t0OO0nC/UTtBwLB41d4inuAUA3i/ALrNyoJVcBnAmEQW
ptbcNp5fxEUJjnOxnedyZEuEBxWRieZFQnkRdF269oN9xzEY1N5z8s4T+QEVp0rT
AnrimHid+BSnJ9ijmHjQPIc7HN4C9fMRmqB2k+NjtJhI1aAYdR9iKyyG99rswV7a
veaqWxFvFC5h1lTYefdkl7/ZmCielFP6TorxMAplyPgpShqY6GfrpLd0KzwANRfr
LGR4a4FUlmQ+6j6wtOIQmiBsoCVPk45vZ0M9Itx3Ski/WlF/uJqzr2XCRjJ+eXfz
FkuvbHWXlN8HYqEurPb71HOO2wGqhsMRSApZKi0Ufl29jB1l5JNbzO8KrURUC6x6
Wx0e7wcV6iB6x+QnkgCFGbu2QXiirE6j00C3YziCBFpeHJkQqBN0VqUfAeictWlp
87MCP7fgWlBfT2Scw053McIsMX+cHsA4LI8CqaETA51RNwS0xctnxCwrElqjos7L
OIdptgDSTilOGqhNqFAni0hON8IsDjwhMWEZx6JeFQ8lNo65hLKgZkg+SXPIkTOl
CCAs4Y9i3HpsX4L+2vIZUeOhDMcXpSo5qWk4QlCK9TMCf9OoKxZ5I+N2apirWRRP
vKkk2os+NaB8VJ7JzrhYZpwCqfZ/B3aXooqB2YRKjtwosA+tKbHoIdxzPTULLm4Z
/gf4RbCvg+/9y4dATjp8GQnDFc9N8elUOI+8iYJ+mCLAxrS6YRDjpHXsyYO26WJL
v9inaoyb2kN7FWWMk2Br1pkAOR2AitV03mfyAUv2/OihQpvjPt1+rrRR9cfYOsmk
G4tuL774/eifYvot+oGyIZULAoHoUKiAT/Lgd6+aocBW1Th9SHirD6Kzvk6vezHS
GQXtKGLi/IFX8wB/5rMscr8GbGIYl7T8/gmRGZzYM2Y37ab5EaFHABOswkfSEw0R
oSs/Y2uRSQmx1y+oxrFpRgDkOx5BpWQp+HeCkzgmpvN7rdhko1R/UlgHrHbRKNf8
c603Z72VnjPCR7Hl4CHIC0baxHkbglA7IiU4cuIPRkWS1D1UVt1Jr9Z0xNRfHCfB
9+KkTh2SKTNSLGcuotvtDsS72QZOXrYiFTvjSwO2O9+QkCRv4unOy1sO81y9Y7y7
DBGZwDafFSVRgB1S7j4xwHB1dGGIYXOGRseSTfP/4+r4VxzE6DWI/kuSWCT/FsJT
+f9yG/kdgkd7+K0srWKPO6jTaNPIf7l8Se0hgMEVYu4Ach+hxUDffSc4PGj49KLD
2BEy2XWV1u10A0vK6F2rbg6zHtInOWsyQtwQDYYNEpQI4d3kVxVUEZzcpe495Rwa
HcUrmcENrZMVDImM4okSH6oB4n/pw2YvZUc0n3TUdQ/En4BnzUTptvx6A44MdSDF
2ywEC7Zfs4EygBExdwgokanIngNhsZWLUwkbvs3KaCwbY6CGyPq2hWFOEOC9aeYT
obV0sq7hmhgGu272rpiJXFbSRGms6OuTp9v3WAk9aemvuvF8rmfK7Q7gTGHFeKnf
rh5p7Z1gGt3D5PAD1gohckMLARNQnIN9ukF9qX3jPyctsnbVOXEia2AaH4nDUkua
9xbuqjTL6ucAmtGgBmP4JqBunlBM/F2OKURHcxtFNA+HFRMO2tVWDLR3uj+dvmJB
Y44tKNJd/jql5MKF66Cb+uVk3ypd0f8VHM/akiTKFizYb1nSQGZD/zmmOe6I558Z
mXuwQSlraovOmgUiKpX5GjJ8uQh9x5je/8dgRAbuvD13lGzkj3JCaLhpzAUswynx
ikGV9WtMqIdivPids7dt3dKSax/3pMo1/pQq2e9PieOfzeZNu0DIwE3VVnrQwdw3
B3hRWZWoTyImOQ13rZUuQoh8+DhVBV35Zg6OqeeIzUi6e9Ma9oVf9tPUIUOeMhCi
gCx1eTgdrc/DZE7obUWFerTskaIEgeaK8UOqmCpUvr596BanY3JVVr5GbaVRldab
qgaWp9V4OUXtRUzcMdDlCwbquNeFOgWC+XEtqMJuYOpyA702+/JRYca10oectYff
CpT6RE2jzpxUHY8/R5w8pPYyrsqE2lYe1bEmp/UOaK+fgV6IQ1IRjprU9DBkhVIp
y6/azFQiGtfKLtPXVvKcgf25DCRNtN06Zpq5tJwTTPNpN1GX8bhcyaZM8pQt8B9i
T7EdIZmrnsdPHKkfiZdhBgkDQ4Ci7apfzJvxB6BL+BCk4+qXSQ9Gtz54M+JPXrfT
2ZcvnF3FXnrU99ADxYzbFZTfTge0EjhdEJhUHvqY69RJsvEh+pegNhZAKNNZyYQq
pClJ3+T36BCz+5MN14rPFcGFRZmphiMkoUYIVUixrjmjE5x6YrJPefixBiTtI2Lk
MsYcLYmYQ7BIhumAAsFoHO1HtqBO1RGrovX8r65R+PNnyMsfLcOKcMARJXdeIcu8
433IvutmALcNuqHQ7rqraP3vUaWdU1XVKZpVNyDhRJsO8VA6SRYhlolFpviu8/ie
EGRE33uArOKgXc9mrgBFuPqgXEbE7N2D6Vn0gMJ6MeGL/ch+L/+TY36pnVFo8B9e
MJ5ghYAaIe2UmJubLFaX/8SoHNuZTXR6pnJfNNMYR6/dk7tltI4rFCZd6Oi6ifNg
G46sXbIaa3Po6TA1a07DoJ0cNrWtBG2olucU26ihsHcMkmvUo8ga5V56fquvsp6O
xqVc6LIACMVQYe5kS9Q6kyV00TjHmj3wqNJRCRTe22amgOckXMzF2jwcEf62so/K
7jsT7uBhnBdHRr9bTSYEYpBxObKUKtR6030Gz+qVTDw6Kl4bPOMZm8ODdGpGt12b
GJzCc08IZmiwexSeLy5LOmg7BtIxvAdsvPxTx90mTH0gVYtjeZlOOaSpXeKyutyz
v9SIWQSjaI7ueTqcZ0MfTDhv5NAly2QPYxfQULsfY9OoXK/H9lfbdvR7OnUzYeiX
BLqo0xc8XVFWLei57B4ZThiFJn4YURZYY10Fk2QTqSilyVqDWntgfVVOYHx3ik+p
r4BA+MnKCHvoPUFJGyitzxC+aJsxt5GVfXuWPVii4f86Ju05N4yLm6jvVV4U00OA
OsGTXgNQq8lc49ep4VEA1hwOsa4kDynh+RoyI6R+zMLPV5GumLiJYlYknrdDqx0z
MbxmJrnt/ggUztPFgfvKeYRrVNtC+vBScl8VikoDtcOJB7imMudadUYM9HzuSQXu
Le7tj+q8OuhtYKhVYcegfgLAs6VKLB1dEw5HDzDt7bGAZH84eJUxJTWRmuE8qmUC
lEUdK4Z3DUSWBmJF1OtJZZt5hiI59iJeNIaxQ7na7Tsr5yDcIrJMcxfmKziM4PbH
lRfxO+Fxgo5jGUGNxXsWkT77yL4pJTFygSkS5yHNI6zs9n+JlaF2ge2vwJMQiJrL
AmKusVG99NboEImlALlPVjJcIA5aRdudo/vReDfskbUlA1vkwiCCmL/8stqsNdM+
3nq1eFr9rVIFdUE0sOKJYYqTL0Af13ReAdGVbQig9N1/nlgAcXxq9SxdzoPSwo3/
WH4OhZ9V/bz1P4pkP+fLo8K4ys9MVWZCZjzzqBlEIVt/JDzMzdRrhU2owxQdLueE
dTzDVus/IIeDvo0HHjCyn37hw0qs/iFBVx0gVGF6W9vcrzGiY2IzSG5D2rxWQacx
MZRE+yTv3P1OJqsMHekQONbGYBPkizygJpjlFyWQqZ/rVoSffb2/ZumcbKNzoD6M
j/N+t/Rm3WH/DBOgq/GBGhEsA0V3oV77BG5aXivBzztaRf/v9bvthaAAmgIaGTPE
IMhj8HIlNSHmDcj/weyKgl7zVHH51eHpUxZrizOY8m/H63whTEZ4h+FrPe6qnOS7
4wd0OD+XdaC+J0dEDsuBEVeKQjmaywWhG0yv5Q3cqK2PMPBD8iR/T+ujrZJSLMe/
kMwi8r77se9IG/CPip6N4+Tyj0mcBGCP66dI6X+I3+Aj8LOZGP5oTNSvhITJ07S2
bjDGh0uzK08VS0KxYEhfvWt6V55b+dVSg4B0tKLDQQrmaIl+gC0mkdOxMy4dsowp
cTHemF2wk0cwU3VBAq+8tdVU7Xv0E5uQgWTqBeE8d92wcOijqKbsu44m8BjrohsR
msDqZShf4RiGdGoTdTGGqRFDDQwCrrTqzjy5jHQLlHs0apP4gfdRUY9Q/oEyUEFP
uuz3SQX0l8e4lt1jktbrTQJrqwYMbKgTy0sHr3LVSrdAOGYrYCp8xmaJbtbt3COj
JcN0Z1cGyFyqXEvj6Ub4WgpSI2y2bmHFUlzwmc+dOI+8ZmYeozhmpDNhkRbwtUC/
S5dB1RxMKO/dFIto01XkJwtFeKNJzQHuP/c2XSL9Rr9s+mSqvai6ODqoUASwLb4Z
97UIHkgL/ZdaDewldoxAxCWEEB0ov/sdow4/N4SXHWrvUZeuDQcm8UjRE1buGGsU
qSR4r/olUWV0AxYHT/yRQanWfU9asAg2mewKH331/fHlzsUqjPPvDoYhl+wcHXeN
VJ48TO58OLkLikNjN9GIL6VpiJ/YxQQVFzTjAgVADIWbebuArTwehV+gi6XwV9Y8
ahjg3F7e6TMFlyZrleoQbfH5gJWQp54yNSSRqtwXgCWwrAQxbfJa/+w28e41/GNn
uNwRqaWknpSYaKE/bCBJORL3HR3NG4WmQaO9jVTA7e42Fy8cI+PUbluvflaV71Pi
1SY/DDp+ep91EGJP1JVifubh639GYSB8KbYA0MBe3gjtK+CIaQzp+i2I1RORJao9
yUIeQOouA+FA/pUwrC8u51XE5EFf6CiWC1I0uzhVsDTlMwKleTe71iOoO+MnJmgc
BhqDnPBA0JpTerRUOkjwYh997mC2L5RS44zhJb1WhQ6UJMc7iTYDCK6yXM14gnjn
JfaPTZAJdP8TUV0OUqgqyLKbZnL20NZt5ST0LH6yns22nY0Pf2Qzw+QH1rY2wd0y
0h3EWHAJOfDjeNlV4YeVCEKWBsdaLnCipOJTVWgT+8yXrf6G8QMkPv47YXGODcgN
7LDpCEhxTtCQk2hF9WM3s7rEeoKwjShZZIQHnE9MlQfPvQSj5DTAmtmiwzCo0YUW
p0NT86KuC8p1kCssEtrGBNw71u3h/Xt5EHCTcvkYUtEJjtOu2RdX6WcoKfPnQFTu
an+lhSiX2DUHxJni14GrZvAL85qMDm1JMMXXUHnvZ6HQLIZM3cCETcF+Vyaz+PpK
7Ya6jRD/dMZ1BwDvb54lIVISZC7QzUbBM6/iqACnSTSCEgZ/ojDpEwkTFj11nfgy
Qoj3u9xC8i4e8P8wuGM+vIvVWY5wDKoBOCaH12uHTmssPAfk3ZZhnMnRPu6LYzBb
qjN/ty/VwfHAdZytilqxOBNIUZRQPAatlTz3Whn0KJg5/uaX5qJH2uPy24Cdqji7
gz6CEm3RkBMKQMoR+BT8vcHYrK8x6Kw9E+t9tr7IC8frQI5PqI/43WzCOJpHAyJI
1zq6hTL+TYRRiHvaG0DD6+FS9U63voEW9eAZeFcUCRuUy1q9nZw1viKROJgny37y
1vNRaxkyY8DR6myB/hRrmr5dH0O1iNbdKAx66eCHyF4E6rHBygSnt2cZZK6jkT+m
+/Ym1Afq831ijkCibdvm+qbVGIpsnZ5G2zFTUU1krkECfHUlW57aGPbr4DUwET5w
kwpUO33bI9m8toBzjiKkDkMAOclEeYLQLPosANdWeUbVVRVRENb2cBcQIJu82PX0
xfrz+xQIfHrevdbZXXzJcF2kKQAN61+p8jyK3QnlchdcwCDlVnWF5/Gm4Nj8BHbH
n6JCnKF07atL8vJ0/XUq10WTI5tAKMNVCoCaXXL1VOTk1OGrQvCOnNB7CAObNOW2
WSP/gwrt8+zY9QGHKsHvdCB3Zm2vuwfb/uw8pE7wwpGxcwlI1mfW1kE+SMuE4IKv
4EG1JiM6nmRjMl7sphLA/myBD8jcKaVmuL6P+LJMBd0ydp2KX0P1iepgYlVbpv1J
sH8pOWTAUmljz9MJMZk16aZ8gH6/p5lKhyPQwNYVf5RjGB+QqB34jiuW+XLkIdfm
XCWc0wvIw73w6Ju5ZCLqbyL1zGXA8wJUkJprxu8fGS5wDBEgQe5T8u1LKiAF33Eh
Vgu5eaSJXJWOLXiaaS1VcfgbykIpHa2Nieo9HxNw4EznmRFp6KNahhzIkOypbQTj
U46grAmH0Se5ycSfbDuh96/CrmtHfiEh+IrF34hOMo8v5ZBQeuvDycsV62248kBa
WK1v8W5RW1WxljMpWaI3kPJ9w2Eb2QkCC/MP52u1SlCWu/OQQRLVFzU7NG5FSnYw
qnl7+4gZxKJdwZ3NT+vM7lJ49KUuvHB4W7W/gig4ZwJov03bCLG5UANCVseeVs0N
J1Hi9DvaYTYmM3+CBcVwRLz/bUv0LT9SLpeNaAOwB5Xtogk72tEHYX3+qG+yW+IL
w9bq/mexeiblipp4K7Zasg2zpMrTIhfL7f+29cKZDtteKfo/aAdxal2xrfsmD15u
/GJKh3BIkaeS2PY6OUSC5sxrv+JcX1KK8hQdUttR8sIxsJnT3/zVtmh3DSdL1PQc
ylkpl2F7vpzBd1GA5Rnm2306Ctlc3xpmT6MnJp1UVQ/cGw5Mm30AM6MgXE3JeLjM
Q4LWcNldWDtqunmbhKt+ivv7CKxvKgh/jhr3IakbeeLi02dcU+QSFoFF/tYur9wg
WQbUktJOEB5rSFQseYZj9C5eQ690HDvncG9o2HuRAwwmOi11i9WPSHnvxaz1hh2U
LZqfm3r0HEcq0MnTDbcqhwefNPWM4s9LwIytIkIyo4LGyxeVWesuGu4KKmXxO9jX
Y591mjP1/7cvp3RDw2vO4W57b6wvsyqv4s8wX6DSEBesWKk2+4x5ITUCA5/yenk7
K2CT3ewF0cwnc47IUGVD3UhOJzH1rtUD/qiP8jTGt1rbz9xNcqiJ8a9DQFXJRMCn
cZaVeKaf27ODQLoW0O2rIwKvEiStThXoCEI+lynP+5XlZBItmkhrKiHM8HLG3f3K
H1Q27XrNGLRS2VtUq2kmSDiNaXABdo+oRxMZ4htnwvHHcKtNjpn4Hyy8b8xRe8/B
vL8zwOl8ggdAaPzW4CDH6MK1wtEy6Hh0/JpsQi2e0MBJpvpziYgUMek8StwFAgTH
ey7NSqo+6DL0pGcQ5Kar+WyX10v7sIE2lD2R7v7zC+NXLYQMUKWKu6gAUYOhdBJ7
p6QFh44uUsLdniJ+jRLWELCDVVai0iaLFmgY6aFFOev0wJXIpgnu8Px8+dkZUpXv
qqPUjfDccNukCPbMoI6hFS1AXVIManano7gBj6hhwVbPjIgXgRiFNh+v//MZVzQF
Kj55kAHXih6d1fLsMCofgSdR9VPsPpANzOxkLj8TlAJHhqLHVHV6yqOyVq5cSXjh
YTeCzStji1fm7oCCt8WCi1a54jLKkzjhFnsGsCw1DLbFMB/ejB2D5GiKBVrsxp4F
P6gXqCvvTjTl1DodTkLt1nzTLRqwVqQ+zyGTNd9Yruli8wLQ2EK5CD0LVnjDlGrX
lwdiAQThCMnLFJy12ltHJ0EI68uNWatNX5DYUpZz1yx+JXIL6kEIVak47+xqFnJR
CBMB4FlNzCwPQdonHyd+6VN+FRdYN5NXyMh3n7WDG3+H5Qa/DwKcBVd1CmzQCMmG
RkNVvHEnD2N1xv9+7Y9EpPiiIIXbhBv+1D5FzG4Y27fiEus29dKgFQuwtc6Li8ka
BUtzKna22N4iucxJLj4LUhGzIdb8gM+74HMuUuZFKAMulUM1L6ZndLUl/lCYW1ge
OvPjpo8Acqa5JJrYsm9xlVMFdUHMhjc+Vh4Cd20jykFElg0cTnB6T2cCZ9Xzz5Fv
xEQDLYYMHQCKfwAhY3wuOgudNCFSyEzmbUjH7zyrwutaxABLvdvoEs/HgBSbtL8R
g/InIzXO63C2yJ5ezPQctJLOxqaqgk8/aIYzMM7A0JB2k4ZOEirXvJxOBnvJsYlO
LTSCjXuLtd06bnqq9o/LTcKFwYBE/N2/ZU+AqzQMvufKHggmPnC1lE0vZnx2ZPyR
D63gIDwKrnDCknPQze5jxGzLCpYiR0+4al2NdwFlBoOjMSSGhc28yuuLmZj6Ztwl
I5xXhnrufAdfWfnYfV8x0KOfaIhoAnNtzfeY4j0x+kzkthVUYD8Z7iQGg6gO4dp6
/5LPh4zXYlmAPzKZyV8kiKtnz3tRmM0fO7yEA1nydX8SL5+4HAdTu0S+MJIkrJSP
LLA7S0JssRixgE01Cmiru+tf3D6Ev60OHOIFHMbh8vQYiCsK2XiNLTwTz52mA4oH
tZVG6yVmKKWEXFc5wPyFciZP3D/Z9BKAD04tbp9GFrgJNmcrPwU3GGuwyZGoJ6zz
/DP4gI8mufVgq+pnMykZvoMTJQj+XH4n/+k3++d/Ijg5g4RpQ5u9MAW9FX29Jo8k
CcOjKj9SqmIrx3CdRI2PNU6yUtIf/Ywv5Pbc7z3iJiJ7QV+tEKHL5iyCZfrJsdTE
2L+2u0uzOBsqXqfBr9LFak4dTiT9nRWHow2lt9dSP0AtPZkPixbmEUmdkea+dLTY
1w/8n0FGYOMX/yluexVRPeJsxw61B7owLatS1ZQjcohwMBJu6KEUbAkWo6J049Ob
4oOmaqlB02IK5Yk8MZ/r2BQ+T+gpyZz2vOX4OjUqlG8sqUbp3/6F4guMtAXvox7K
2C5WTAfuMBDiZhuzSwEEyN8YimMApoKYqapQXShp3drF4XY73ZBAorU4Bn9m4fFk
j71he0dP8ljQ1G2GEtq1v/Ejo3xHbHDMB73qBCG+nkf7+mCU36YF+zk5S0SyAmQw
fn68BORJ+AkJCa6G25+/mqZr9kG/jtCRD0I26HZv2Aw8rAL2fzhw+3Tz9WSDn09e
c37+rnJljMd/m4rrHGIHt0YSh0Pyj3xtgDb2DdW0Mm5mIDWoFnTBpW5w7pK6+EjY
FaNYwl+aEfyT4/nhz1bII0K+dQNvQ7ZIh8ryyZCmfEWzgZOBLPk2EVgaD557/Pqb
yJhv5Mz9penE3pDIaxzvBjysDj1wWk8kbZIpYc7uC2oC5jChqThikMKYq1ksSLWY
mhiblczhgaUQAXstPjj6xFuCBCfH6OC+9UW2dpkwV104GuB8mC6DrFevRPPjvWRl
lOd4/wWDNcfLDOfO0bvujWQOXzv2QrhhPn7ERboUVvskrxx1zlowfs+u0mUzXbBe
2msP1a2kxP274EbqQPyBh9FhaOfnOa7fZZtJ/V1v+xGEG5fz9sE3E2p5CPKFRGv+
5mbI58/y4NnJV+ysdRHIErN2d+oy0OVyFvlU7VJ6zDr+I+nmvvpdsatnuLrD0sje
TBxfDNNhgga/SWqLfCQ3HkrYiWshApogSgCSm375n9Jxnc3qkstoBdURw1z5nn2h
eSsw+PN7cdtKXc3JZxSypH+rceFr3cprUuaL7+C/mMbYzfaMk0YV+mlZRp0eU6B5
g2wRseFofDvbPry9Dzt999+UpNWVfEW5O6dbtV9eGtzizlkp7lSOUgqbRdLaKqzq
s6pw0hhKzVjSJJUWfGkSXnba1gIVVKqg2h5uymPMD6mLbtFxswUUrqIrWHr+yGQo
TT6NqnyoLakYq6qUX+V6A5qcZn4Y+WYdCSBU4BWIIrAcZISUCqsNfnRHPrn3kHsi
mV1QZuRyNWsl6XUcsgJ8DFEbNpffRgbmwbYQOzIB+u3aZjy5UUKs5YBMgLXulcPD
HzSEZf0YTkZa8l4d8fUJVH+zCCxLlz0oPjNyKgDgx+m71VSsmqt9hw1o8i8ST3du
EUtj25/kEw8NSvkBrdofa7/Vdre4tIkE9LDSwibMbfLpZ9yIu/RLXsXXP39n1S2y
ipAso2WwCrb+yFaH0xxDQBZ+oRvzgr4/2a1bn3Wk3m9EexPBJEU3et6nVzTr9gNC
ysvb18LdiWBZbq8TXZfbsd86dQgjxz9RsKYI5kKGNqXdrO3Y1YI0FDQ4eb0Kf9GN
Kwz/Q3Bjs35sGOtUIiD6jUM2LkFMxybV6rC1svJJe1vUOJr7EiGkrZvRzYD9kq3z
epkTX7iOl7w7Ed3j5BCnZEwyGq0o66w6AOYolAAf4BH4UWz38p0sV66GENIfiVZz
qBK05RWLgScrT5qb1SRu2LbucBHmePEpngfWcTRWOEaTBcutVkBseA6eOmRc7BxW
beh7WsrX5H5ae4qxLKt2UsshTNGdPsiCZg041JeMG1p2pH4VLzJxxhg1vdqdxexQ
rQ0ZDp9QjFa7lIoqEqbUQJueXLD/IBwGtZLW0+U93c1nzUQY/AXzfUJm7t38bR7Y
mzRxo3OzH18Ws6UbpVc5JjRwBDDI4u2xei/pe6iCYS9jf2R8so3JeTEkL+VUiUho
9Gzm7P0GnDXDjBb6qyKsFgfOkncwn/6a2gS5iGrGOAlr00mWINF7YV0OEQEd0xeu
ODqt+kF/yimEIM4s9GBvOPZCFgZchTYM/FstXYdOQ2tuoTTWsLrZxzteluHBCvcH
vRHStxAccOItgStCBx+rZKSg6ohhImXU4vv5t/pYoqY5RoOb6ckMAvh2ah9z78DO
u6mMFzgz3tHPc1fBM8NJ4HvRK7TrmRUAP/FCL4hqhU28iAf7bkBGy23Rm9Z3tGRx
avo2gyA46Y50TtixhpuDkZ1PTVH/Fmpt1gKVo93DoJyUvAiysmuJIG0V2TrhiMQb
pHSIRNjSOm8KjlJnCBcDl47KJ1ZbAvzBbCn2M2so4fuWTGuw2B1c1FXP2tLcwg/A
RRgohZiFDPxPUa2xw7lSNlt6PIcmhZc44DG5CZ7ROF/KKQWHBSIAC+3t8DZ/1FNI
U2MsphQCAhfILyzXnZx868bDN4bAMsvTwdFXpNOAQf6h69hwT9nXX5BRBsxF2rfp
cCucDa7mjNSUc6taF3kps3a9kGc+U5t1cZw8PeLb9tbFj354viuO9a9JputOELhc
OnAMYcZ1cCayJ9mEh0bXDHFaODRE8SvSA/O2xhHzsQHI0jZsiykv7m4cBgbdnjqE
nztCL+mT0uTHvzAgg6mbwDHAM26oLb3qVwpOtSvVPSNBP5i0s6VmyjPpyPNVveoi
f77CuVGF7Hn7J6DWkz+vWwxU8AS4+ZYvJw6HYW9/bJvbYo52M4uSLVcdcjnLY3RJ
3hfY0u2mDli23QkHGs0odlJXc3AwOLUDDx4e3MNnkCXl2PSuaqHjy2m9e+cnv0VX
n4gnugOis+DWUPjZU9MODJ5RIRFPgYBlXRA3DpvQAunuT8vuJ1HmBmaGjkwxKgpm
zkPxrNA3d00EwICTfQ1ck8YDK4G66BhTJ7mfwedoh3agheTSklgdf4L5hSfk2clr
SyTYPQD0rW9/CvUCiUex0aCQF/uX6BWGh4ClTlHVrxA/XajfAfGoQFHfmpLoEGz0
yT+CfeLsBUq4Dxc28MZvy5WMOw/pgi8uCspNPjLEJnDs1K+yn5jkOdfPk4pr7BLL
C6abESOo7YPjMNK1bQAVtPcChrlO6huxmt3mPwtWI/mWsl83iNfXfv6XZePn3KuX
rcP+MHy/4m0zdqpCryxrAj7xGWWSIVdxWWQ+up53Q1Vp09igBhYCY8ql6HET7fcQ
TA07GbTxW5m0MJAoM39aFVkGS+Nsg1qgzX76HClmquKM/goBrceeImibelVcJtfO
ASBlcFfcLUTJ0vPLmuKnfTuYGveE8JiT1iR3HXKtkJhOrCilWKZQgyQKhlsy3UAT
pxsABQRHQOTCDGCQkmGTWAw9TurSRb9oIplZo4xNru5/S0cZigsXyv+GwiWcYHTr
kdm6dMRyQ56hzJP+FjpXICD330xzWb13cW7ZiSXd4EKNIzgTqvmhWPLkgkzC13XZ
8A09EidXVOAxOlPUk3wLfCsJ/0r5ztRBbMVB9Jd1Kx59ebTmSY/47OTDqgePTF5D
yqIekjHlDouwRUfKOInQj0x4UG47Ifuwuo3wmlfIBypuuEIoSDXtg6cUBs4EntFX
4Tf9ADZnRpzjc5jwET5Qz2Uzvx4aLNqYrrRP606I859EcMX9r9uYrePHS1e1cnhX
6A5FRLoHdSmiv+xIpLS6CXd4NWHv18zejEY4jK1ccM7vTeGdg09wUdk98axsWFwq
N+YokoVzqgIHn9M/T8XhdUN2vbdc7Bkf4PgbwcPBkecNxBnOYFoWblNyJY7TvJTX
x/lETXNXyKvY25Q6BRqgTH6l1KVouIjWha2N61Qrpz+b+mAC4Ob0M06bfWDyipnp
TbwLq8bGZl6Bd6DK9wqix69uR64c9frqpvypbiIrHv5dlyI3YigJ9PC9kyxPF0h9
WJseXMI/+9J2oPFuMj2z+4DcDs4u7gppvlHzM1qt+7Dw9+d/+ntjvkAJBWdWwiVu
HyANk0ZAXQZeKY2DnzD7N/Axiu1hukxO4Gopwpn5YWZZCvKn4Qkgp1Sf07Qm0Oek
mLKfOSh/sb/vf14mchcx0r13WZ36bCw+W+51aSfh1MJNSxvPlFaAMgp62oDMrbiR
zinh7yUoXOHot3Bov2j6ycTHl/BR8Z6rr4yh0VJDJ2AjJi+g0Ct5c7darquDjWXV
YAPH1WRbkmzx+zSU1iimljPBdDBMMGHzeI4GpOwHMWciUDLrPyWVFSup2MxMwQzF
BmZHy+B2bIf4tGSNQzcfSILrYOJ1CKxKy3wlLeG+AfEQ3NkANxw8drdhyH11FNAF
htNHiauwA3sHLiwLZBShwSceLJAhDpoEpoAGJ+v/Vb86HAL5D+tyS61hpvChsjf2
84kzAlLxqsZBddVwK1y9GXOLUGOXh840i0GGbO8zdvfP6ZsS+ZHvzrll2en5FJ7H
lsUhPEEB96WCEQ7YMRB6iubUlOwcSdD28QtWowfknWpD2P5GhVUchW/TUnVRk8jo
fTSqd5e0WAqOKDdv7zzis/1CfvJ3o/qPTseqvNoT8QTxkwgwDG3nE1AYFJ2wc0UF
yuZHoQGzpXcFRgYwizaB6g6d6Xt1mA4dQADMHSajsENLLMvGdRMr/6USA8Typcl8
b2E59ZOEQqM5QSGSVMpts0xVbkfDa9g83slZaApKX3PxueXXrtoW+I90SGF1nYyF
tjFs1GRyRp6ycp4qu6UXHT0ngL1LkAPH309zIWvKdsZgkaIk6Jpg4H1J3kZmd2U6
FQ5URNQl2nDjff8MTOk6rv1aN7at6+RNvc+og5Hl5q4255LVV0YYyRytoEz2Ddql
avpzT265lN7tcLwuqMi+c5rg7XJNcNqQVp/umnNpkiIHNV0KcM0PYJz2PPXsxcZ2
QpAcV7zFj2TxK/ZAJiIdLkvTFN2RZvIykY9v5/K2ITdRqxQkGej61zETDBU/cBq3
Kj1ZOelNA6rrRP0gChU5uhnOZEKhzSZ8J1lTBxhHzvIdSUVgfBkpbMhhfnYhKiAV
zcii9lvyXiIBsUIqZRKhYfoTqSZs7zKMt3Sn7aMz4HtY2YN8z0CJ17loTIkowVPt
pcCT/B71Yb6xpbD+lr78VWTWJeoKGBfsa+u09tuWdIST6xvn6RafRK8SvZyHn93b
2/bAn+uHumcgvf78iK1UXTJHF7bLH1EldFQlo45y6IGqc7SRkO7c8o1lX4yjLhoM
BjrOnAqANj0CuGm+s00ttPCgzddoxQXNAElYW96at3EHFyOiWFsP8v4ZnZJuyfiJ
aEOD8uk9oKitStWkdWlkkbk1HZPksa1SVtec0h1RIfuLQctgwuPVjtKtrmAHFEF8
coaM0VpT8+IIS5Lmek3lLKgZuDb3HCRncTBTqPS6A//YQxCDk51wWCsWQouT0kJG
4gmclFXJ9IBpi/9N/2ua4LM53IkuV4xafzSSWKiV5qCJskix+Nsm8p3l8EVg+lgz
W8wJIiB5yovmegLVQAhNs5JvJaztOfO/eeJttmAhDLiYZduqorogHm+Ij+gKbeN5
gyonembxS2baOsygwBR73AwMx8rZWRnw9ybrUo4jGYw0nNrNTePEySw8FUxIdyvi
KlDlLigJV+R3nJimPIziug2i3RuTpuAk+YH7HgMpBEh622G63xsTKiXiSUc0so+n
LQ0fFpyvEzjGrTMjrofdrXpbeHfTzD/b/QYeg/JEouwsDLEK5wkknIgBq6+WdkZA
1s4wDisxMPWpg3zyyY2sEIZU9mX5bc3TGfTd+d2npuBhMBYrkP5aTTisVX9PX9Wb
GSlocZWDcR7h2yFTfFT59WrIk2Y0jE9oOGgqJ1q/u3/kzMIeabUOQMkS6oDxKhNy
XVaALUDBbhkyLsUgb1PBHN9sQ9YAi3Fk+bcF6Thp3wxFnODOijhKl6LRrC/3H9x0
3PcNLqYLQtpdRrgnHroDMt23xrsCvA0FYAaufyLhuX4AB5AYSul8MjLWXLAwejSs
3VEvMPbFRudDM5n+hJrDYhbowYrDMT4CvCjOb53SJm3G5vBKd+DlZOP6I9kmdco2
nNSJuzaLF5VXtLXUtFFTI72DDtPklf80n+wGIqEzToE44Otjmo1t4g92kE5KzftR
/g2HqqAsU8KElpQoRDjxmQcz+KbtyWr8jLmvM1mHu2/faUQeK298E+tJtZXHuMjU
CDvpz0ktAzPTvBgaDe8eICnTKQp3TphbT4Ao+cMOxLDY+LvMycZj5WRQ1+RDl9ij
XN4e5pjahzFWm3Hp/iqHEgupHRF9YVQQM0XAkHfNXt0m2YYU9c9VHx5FVX7+MxJi
eDG2c6YKA9zX+ozsszqzn+3fpBJ8IfqYnwu7wMpJwviqxtwWIYlxdHQ77UzK20XV
5lE52pyGJr8GTuAhB7ovmSE6ddhiOR162yb3nnMDCpn5tDoEtELLzAQQ4T/1hWLF
2QucbKGE6SZzK5/eVMgK/g==
`protect end_protected