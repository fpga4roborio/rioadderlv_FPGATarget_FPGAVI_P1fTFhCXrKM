`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
ddtXksX2+yylW5zu6QL2Lhnb2d1sD00763mmSITNX595NcHTEkwn0zB1Dry37fOW
FufOhVzEJp80NC5qZ/+F0Vk7Ik02dIR0elf3clrjeJRK85K4e3Hoo4xn7YbFUIms
l/8VZSb14+JVGURjfswrIyCUotIzlzVYZ6gzoZwDXIi5gQIBf/gI+KxNXPaKV+PQ
Ufys/12rjO6aI/pPlqSm0hCvftmBcnezN2hk1UeXgOIuKZnogjOsf0iJVX2aOOWE
6pD/psybjbnsNB6kH5uFTA5frkzIzkzl5d9+YDm9OyC+k84E83I/7/j+rk4L2dah
QJOvksSIzN867/4Qt8qYTQ==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="MvBXkzurAa5VTw+1JJ70nePUfoQXBvZOku/SMmg4TwQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
oRtzZL4VJ4iwysPsC8SXYCzXS8Fw2gtZTOskLcDV+1B9Nzn1zTyNtlo6lNICRmmK
ZRVu2BmCc2G+fmzynYlNTnSa7C0Cuel6FYpxCBlOuk3OF2tzAmLAuDyOH3Z1Yjzk
a0aHuoCdIRKv7BrZCdALt03JeUmXKPdOmIlkVGFl8yw=
`protect rights_digest_method = "sha256"
`protect end_toolblock="Jn9CQpRhJt4rnzZPRk+dOpzAubz7omckX1MrFd4p81o="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 8208 )
`protect data_block
gD6l00tciPUa6pDNTk/+t0OO0nC/UTtBwLB41d4inuAUA3i/ALrNyoJVcBnAmEQW
ptbcNp5fxEUJjnOxnedyZEuEBxWRieZFQnkRdF269oNONyOsf1JidWjhANNn56il
xKZd5q0NI4VHelN3JW2m4A0qlAd9OVav74KKrkzFU7VPEvdWb+sX9em0/h0WpcEQ
Bg+jpEZasXTYFo/NHkpzntTIH4ZzDgvVuwEXRyoQSwmSiwcMsY5i6vmgAc1Ibj7v
ZzfJh+zqp19RH9VXDO3EHcxDPA2nR2C2zGzNdJgVvU/+hLceWqBdVnoSnxDgtYQE
QTH/NgiXFkDms8ZJ2t3LI1QUO8yPTBPSaSaQLRdSI7v6H+9l3M6OqKapYysOV46P
BXlSNAyUWJBwwGLbFLI8wAvZ0h/xWy+t2ZiqjeOdmMgNveEl/1PdPVWZiuQGsby4
CjIGaG1PTlxSs1oyyEUeYuQB6fOvsfRnwtygaHQoojW/JWxOtfCk9PWuSPNgoxtw
V0GXf3xPIf0jy5t01Dpf843vBrqpsAAuooHPVH6VnfsR+p6eKDAVKy16qHTg1hOl
B6UyR98Sao5lexV+GdQWwPJ1Yeh/PAtAWH5VduqqnNt4RLLsO31g9TvC4woVDq34
ctJO4SQwMhlMU6dKvXiA81n9WIO19n1NJ3RmcXM7ft38698AzAnk8T/EqaQKjYFC
YVwWB4KmjzzGHPwVxngDTGG6Nm9Eig0OEoqe+kLPR/kyqr8xzeI+tAAjlSwdxUvl
/KDGxljkAnUKblWCgLeasuX0hEgRD3yxU8/uFA5lZw0OSZRHXHzfe6d7gHRm3f/q
F0ptch8xkBCWK/FmQ9VOgw8koLEPY/ESaVEOdd91JTAdLqiOoQIc/PCyYmbfkOLn
VB17B4x5yqUShampjkh110zJn8P3wVq8Y+kF4fOTpfb36D3oF6MHDfK5RaVKHJj5
SANTwVrKj0Pt38M5uAXIetevaO/mywZz+sm6UZKMXovm9KTb1JyCpPKRJ146RxuZ
v5v8LvTQXsYGxb8KKF0FhI+stjOCJB69g6S6hxxF3NfSIpnN1aq9fGaN+49yp0Kz
HobYQDbbv81oDK2Zr+PlUcuINe4uU6OMqBw2CzvLd9WeAa0Anb6IS48+wGJvnWq+
4cUPgroe3fSCivQnqobkNGIkL2u8OI0e7fHQO11slZfA2ZYGVKjkC31mv54RPf8H
3F0YJTJNIl3oPuwBvhgoy+vRgjTkq0Pe2VW6EL5MpFTLjEFtj1C3bF66ceOv4f7l
ZWP7zn6qu3o/38xZzEZLKpsFmr+3iyog7RNKdliIyEVUALJWYUk4K/asI41LeGWu
yxmfc+S20qOuVIrzsBcjzRatV+nmLUkhqZMb2eLeg4r8kR3BIgtLZNWUBVawHZF9
eGMJxbzqAPtHtGY/8aVUdaURtlKccwOf9N5YcYLY82U4TfGuiP7zz5ysY+hBE8kC
faHb/f4KzLmZ5Qdeq3/8TUE3onoljnocg7RnuXO3g7Q/JtLzDHmVwUNFsU/KJt7/
jqBm7cjSuuAGGM//YKB3yNNGNXDY0XqJ9+eoFCVDoCgZKCgIqqTormO6x0/objmQ
dp/8yFHBi3Ehl8K9JKF/syTTlPjqo8Ii7pqW8inAor0YZqbvonfYljYINXNeBuEf
2P33nf1QoAThooiy78JOzi2FnaHb9fJrcgudGd+D3CcWv/jHE3zbzJSApf35oPsD
A5wGm78S3Z+o6BQO4kiLD4qNFPw0oJZQ1kjlznQN5fGiUgETB0HWq7QkU3OornZC
OCa7+CCp4Py/zHrth5uC/V/w2n2C+zR+FeccE0Ut5upMoPAcaky7KHjItwyE+TIO
pb1sR8TO6fYjmxcaFkHbNDb46LvIHoPAPVljS7UAmw3veYJgOg8yJhUi5WtJ2BIL
1Umk1kh6DSQwUE2zEUuesrTm/hdFlCm2JavYYQtIu1qLYOshJgu0ISzYF1yjsKNm
BhmM+BSHkMtRkUS+CAKM6H+Z2eefn9nHSTe9n/XRaJXVr+jdeEyFxlN4m6KXc1aP
ne7u6o6mBUShGBb1wZ6uChYvPKMx50Cf5mMslSUtjzmMKyMX9+j8PGgNVfENtR5t
rY1RKXStKqyh9lVunWG2TOS4J0IpnA6tvxl/em8Gt9Isl7iQBfYrzVN0JvKH4d9Z
pb2GJLwqYc20oL3k75tic82rYwvN949/2XsIlVo0slAlN6CCIoTk2wh0GTD6+LjK
3W4TaZUTIBky50duHt84fWkyJcsHIBw9q2F7qJyvsNm162p1TpGWZLNdCzii5mcx
7r948bQDuvV2QAFbLZtoI0AccADSWW13fxp/JlpbdQc7dXDxP1FRCOl2txXqvKWz
4xS2FnVGyN7q9z6L2iT+JNKqSzUjwK1Dv/2AFFnkidxsNoiVwB2JtsMRNddiLOXi
noUEJuNPMUhBmPgDS6mS5ublA8lmwmHy5jETHworYyiZtBuasuyVedAw767fHjnT
lqBuQ2LcQYaKjErozW/jhCVBUpoYkitEH3pk0kwtdhhn8XEdV0yOu6uFuOoiNach
b46Nq/3sAmpdooHE4PWhpb0G8M5ffdu+Of5bCwIuYGuN7B5iXx4ACsCHiQbD7GFw
i2Dsk68h89CqLIZKINIobxH9fOT0efhMCkBHMGh1Y1u0hpl/DLtbsTRL73snnEZZ
Gh60q7d8oSrS8a9OEtlwe7eOiJBTq4e0HHSPeQiOQvQsT/tkVeLiuWkQrPwJQyxN
UUnAwtwDgSX8wodYCHpEIVQYFzaqrw1rqefZdW9iqfHnJkAnPiZieO77Qs+3gBUM
mcnKW9RF05x5A+erYIsZDH6PHN3IfwSsqRbp9uFvcIxHXbVlQHqDWTknVpNxhZDd
d73OXL3TOkzQ9HKzzsKNky9qXeN/DdJtg+fLEBoHQZEjEpoYpG/72XRGaf/PMqqk
l6JBeEvdfGdjJWRTFJrTTjXTLHQdJU41f7NoStADbzyqCtXaCKal/a/ZQ3Ei1moH
y/M9LjtNrkRTT/zjb/0g3i5gQArq6wnlxHonduNHYjo52VpdejFGgLHBQKTwXYID
gVZ/JtFDxel1O2nc3UZZPELvajIMjjl9QdNVqA8HguFaz1ewd0YCBbg3WJrNZ4lc
Ol18fvpYNHHfXsiFDLZG5YUE2kQKF1wXenQAHULpEVQtWSUXqtX9Df73mR8vRqEP
aLzifBDCK3H+e15aGN4zDPz+BX8ZHGdiqKJFLGDOt0T2TThwA1XBryerc07b7CcX
KUI1Asyo7bjtBQKn1dzaonRxwe8gP/3HelvU5ocZ8aLBIAD6Q+VFPJ9yFTx0lhgi
mlL/h0TS1uTFSriigUAB1hUOu7yqCrGjs2ZZrA48YTwQMWNEP88XKQuC+9ZltaUB
6R1fzM9WAQibGGH7NFJlq8+qGQiQ/CJb7xOKVFD0WqstF5YOSkgEH6c0T8wGbium
LLQmlkFWykX3YgaU70hOXNKnDWlziy11AkrNRwnxVmdg4nxSKGtUxjlPTGgHzaS0
dUo8qAcN+Jf0zVe4gZq2qHgnLijdGVYVLloEd1ykNDvozdGsnjp5ZPK7xsU4cVq8
kRQLqbzcx9BtdlhlZGgOhA4eyG+W16Hq6N/1uaOwhyAF+tDjaiAmKvMr9mFbMxiK
S/CHO+6QYBKpxgy5sW87PNyslFeauAZhUEln8fN3Aaw5b2VR0gIpgp3cRKdnp6ly
DjLia/9yZ4iafytTBuR5+CkkHbxsHDIkazVKfWYG+DjrPXZCM3YE7r0TJl1/A1i7
wLB/PLba3nlM4s/2mLLg/Hm02qCrUpizx4TkwcH38FlVXujxa5hzwVpnNWmDDh0o
hPaX+/OZ7HwVLyYhuOSEA9LsmeFICwvA8g0PFbFa/sJueINjOJPFLAHX3+AzbXbU
91J0w4cpPTeTTcpyi11rjQnEieL22YFw9WPunAdxudRgNByyO+JjHDujQR883mM5
u3gF48tGA7RUqEuRZLzFF33g9JPviRIbffeVtHgnc17450iogTQPj17EG8WxOFWn
s/OEzIYiHouV/9zSTr4zrGLZM4UKVXOYRtMQQ6tSgqe+u1IJAFq6+6F8J1e8INDn
JXgRJ9JTkV+zMdRNPzsZ44Qile5J+7yr9a6o2D+NAMVWW5Z29qsyz8MQrIlhl5M4
NAjM+DQ4RShHbrNf554EQkz5LVTLC/xDavlShQyaU0roJyxRUStaSnmK7H4ccCY6
tHhlOjLpAGMklofBqFGmp10tvDBeWbZ8aQzHFMLtaoWoYl5kK9qL5YzzGIM+bddb
eaRrSQ+QPlmabyXI/V0pESxyIUyf5KYdmZsXDtYzU3cKkbn1Vluf4iOeCAaYST65
jpoz6xKGu8SrAJ2yd0NhhPtioauIOkxuvceKKHuRxvl9y/4Gfw4pyNJrsqty/h0X
CUujM+eu1UjQ3h2VOPorq48RMShk2QpEU+Bb3HHGcfFo9ooKvDcocsk+1ayjAXqP
NaSTmKHA7AinKhOWPXwnEvY9K+J/VnYeRd2bT4syPpced3Tb/Tl3CcdC8S0p0qq/
FSoSD32YRjcmA/bsz7+Xd2rpRuXT0aH2J70l9633lPnN3E0y0D/Oel4to9fqkrZg
YXoWAka6YqaxeIfWEy+4u1RlQu7tzeFVcjyHYmEEC7AUPt01Mpz3Fg+W1+awD+yb
fsjpIdmfkhN7TbzONmGdNHMImhqCa0Sm91RQlgXHPE4V+KCsvTSj0tvGRxgCXRAy
++sgAwKHEAiwAgrykJaM2losdDgvy0Tf2qj0JezKiNVNsXhHc9ONpWHYsevMI6mN
Fn9G69qHvPtNCUm5U/HlK59uDbwOt+U2caGN6ttBediHk9dLx+SOYWAnV2Rxxqbx
wMXmMnrP0kRqgsTaGPXC5TG0sOIU6M59UG1nsTMMd5lqcYAZnHy9ZYp1WJqgo8I5
zq4CBww3PSVEPU/d7X6KUx2Qbv4ClR7zy0sYDt0nrJrH2M71BnhY6IcOfpK9KDE9
38OELtiDI7aDH0swOIcRqvnJhPYpuaZ1F8CwJSEy9/YnC2OJjXbdz8+2RFKIpk5f
+8zCzHEATm+vQ33C9WeaZjltg3Gq/R3fzevjIzZMdceDoiVGDGqDmHDvXUSkopW5
WvxSe9r6U98v8J6gl6nYLSrGfS4o5YaKtL1zwwZijh9oKzDs9Q7Uvftm3tYqhqlA
fAlRf83UDl9EiUmO6LNbOvz+IIr8vXYfoZ2PMMXasadI7GdcwkgjNZYteFgzcBan
hInpZOncuhSEgktocoVXa4lpYX+WVevdvfCcp6FqSGP7Cpm60Am9OOA0BnpibsTP
q53mFeQuUsPEXXiTsdBKjI/UAMF/M/iQwUG3yUVBICw3seh0KAAlpfTeotx2t1q1
SZYOHqV/TIZcRwTc3FFebtmKTR3ZBmNkFcv6h9h0JgDpc9yL09iWBpNxJFSbTM9E
M320F1wtNkAOYdfrfwx2lr9F6SllI1j10H236TDClmdaEFZoBdGb4bVuBF6+oE4W
CBZXXY5P+YlOwpd1U52RHhmAzTrw4cj3LfUmp5hXgBgeFpGFNzcthbRxYVrlILl0
QB8Kogf7mOD2MmGn+oaGq6tJ9zeUYXviVsF/p7ZlIznNt8ogqGtes1UVSTmqEtzk
aWKBfrBLWmylLHOUi1TcJPKB7UTIsF6sK/ERnm1+LJueNIDGjdPDQacMSRlJinaW
FKNE43tbKKXAF8f0mmMmxBOXpEeupYQyuPHHBgPgq0o0vYYAGzgH3BKoBSvkaGI5
Mfa92IkmarmZxXZTf29p+0xZbfDeb3ckRhE3TcaQ0hXZMSFCgSRxkryRBx0uPFoO
FrvupvZjq9Rywq5YhC5k+gVgLgK9BglcxVVH3pWJD8eXe/0usOGc5aKuxPDua3r+
8361mIlxi13HdBzyROv4gj++xo1R/MgskfVDfLg8XAoproIfPAzifOyU1FCG2vVp
pts60IK/Vkbu5yFi/X1t/nNHv8AUspzOj+q9JSb1OQ9NrQZ7rIvLBtITUZHpuqRf
5JUSHM2hgUGlX1o/wb19jfj8gJkQotfJEyPEPaXdV8J8z+oWNVYY2QsuvAunMVvb
lZ1jg364qtRD/4xIoWJ60liDULbBQNkAcoHkelImGuUUe5y6pw3MNQKNRyzVIW5t
aS8rG4LKKUENwWzJV0mR9jdj68FRtwO+YR6n7y4nfx8o4Cj6PChRK210s7rJcFTs
QhjshVt6S+qGXQGFm5RlfH2CYV0WAHavrO14xRoLvftyZZAZuCKUgUD65sxOy00L
8mKXlN75BLaAxY+6yM8dyNQnXJQpnMNDjliShmWnCcmRbNn/f5aRsRVSiTcS+EZ0
FMH9Hq31jy354fFe4rzmfR5gGIR65mGEpN4G/7fcvcpAVXQzDEVOmP2yYnPrBDW6
2TOzETmT3KwUIiI4sQc88eV3IBCHdC1ukNOFiiIAuGAjQ6cNhSIsLE2nBSkOcSqb
4KIV+K6n8P6mEx4R0SyZ0n6eTtzDoi9Vo7vNymIO9CEBFkF47tATOZWjD/6CWSBD
rru/1rg/ubfE6OFCVLXFMxb3s2lSYZpYukZ4+BFeZdyaVSStFdgUGzJHJHmGjTk7
3PszE+uQyezuieth0G1LVu8H72FDIQe8m5IAIBLDDPMiVaRBw+fm8t2vCRXrSvKv
eUqJU7h9gYBz7phmbUcsOTq8okbB6kX47LxbDZZ6RFQFKCprZ0CxHZfNATUbDDR5
3At8P0l85yE284jq/r62ef1bDX1PG69DU8PvGlnxygGA9Y9mO5CdpDxfOasLCPW/
YBAYIcMUs1l8SupyY6Q+RWQVzm9Jak3VVNX1sFik1c10P9GBbBXEgu8bXW9ok/Qm
Iy8U6FeMmbNel4XlksAU5+0ybnnNOcRD4B9AiyaoWeaHyN3OG5YJTQliCwPx9IcI
Mo/53gW1a0pDSJYUzeKng5u+9d8YnHw7ep+PxUnMZmqtHrrlcfmMDxP97h0T2s6C
1RLWGXR2iezdQTamKrjhm92TVlWSPTDv0r6gu17IR9w55Ycv9M30+Gj4GAiuxTgw
PvD4/j1ungzLpl7deOj6C/tU5KcOKdXd01Mcc0zBRkc9n7FMJA2TDf32TYrmGOfz
bOzG5hWq4HkvGX2Ku2y2b7JwaxErNRhKEcG/3Mcjb2NUCkPZ25KB8/VE9JlZmKUF
7E1FOaP/C8NMfOd0FESzNThneMklFWSJi6PnjB+zX9K9YshYC01wsYjpK+9hmzR0
GGSBstsjKF2X7rcHhnzngXrkNalfwGCswprK+1EHh0pjnUg7Mvzn9bPNYcA6O8VP
JC7vJEaN7/cM7q575KtW1OLYxVYRFAF3/JzCDPL3h3gaqWuRTkH6TDOWhA9Wspru
n8jjSTOj5YOPSvgew/VmR8x+qmoalpUfG/OlmMK2vLoMfpbVnzB3nzm1RmfQ+I9B
tso6bdZDgno273gmDwPK60BTOf0ysuew7fA1qYxXsV+AWEmbQRE9oqBOQwB0hxcb
kLm9o/UXIGNqDh/1cv5H6m2DlswRX9kkliGVs2v3B7uMpTMN1Yuq/VcBxwZvsX9u
nVfupjxwKQUvVCCv1QbqOQC/l4FJ7T+loRlEnx71YcnxkvCxUljw99HJBjPpYo3e
iVXdkdz8iqi9D4XZg2bljPZWzyqv5XA/TJdzBPUVciKPn+Ejz5FfwK8aWfYay2iQ
D+JlBzsoTJeJZl1SA8RhnHBk6hj456qqQTRdqXlZCYqyLstMhUYV/OqLXlICdsiJ
SEU61hxezEljqp7V17KiAlqKYr5tg9brcbLH+Ql2c1NKIswaHNEOGor5gDwO9s7K
BCIcr8HzIFsDKED63i2XgtMRfTd78v3REnloe86ecPgSHFVf3ZuvIKUnAgi20QTo
JuuN3YXjy0rZOceQJSzh6MjrXXQjsOPdP1Qamfp3yahazBPqjnqal3od6Ocqx6eR
iIdCuk0I1S6bRndtznPHK9C4EMpcm63vX/+HIpZ6vXiYNet5cQdu8DThYrdvT2zB
CqzHn+5Y9nu4jKqzguLBbgCQ2evhWz3D+vIOnuLkTA9l5n2VKb9NC0QEmktmx6YW
HkcSXhsirUkaH6MTdcAJvhysOwDrlZ5AbYaiia3evmesqRYgzzRxwszkUI5W4weG
Mqe6G8E8AdMbazHSBfyKc8NRU716acA8U/RjLWunrJcsLWt0mzpHS1b/f1dJ1J2o
mVooOkv0ZAvSXjSy0Din/gBnDc3+BsyjmknQUaEBIQ7XTxY9wFYl1AJ0gnFOHK3F
Lgvgf+0uWbSqcOqPKWRJhkET6avypOb6ZPChA8kUzDd1BidyoFW1ozpKL6qN7HSN
PWPFIIp+jZdc9xV/KVTpA1y9uf9m/KBFFBTzkpKc+AqpN+ch9J9o0CEwngu47KQu
7MaHcZ6kLgm08/8qUVF/SS501Ax33U7YSKemUmk2HAJr3ONrKNgPvLyVq7Mm4qG5
TafZoodNRtadbyxl9b4kaX3bEruSYLtBJSGQ+k9mbI+L1RCzLaQb6ViTzMqJCque
KzmrFYlmTw7lmfnoCvig0HSq9QwjUtcbjydFaKQHR8x/Gc+VBt7QY0F0592q7S1Q
1htv1i7Xp1J5rkS/EBVWnvYBTcmuX8R/emaSVfEBwKF3tR6QhiNcuSCISVDtTsFy
Dlx9rhEKCoMIHMB9vSP+EWXRTui8jxrDYiq5tnOnhSgtnjEkEv1MV+jyB59rn1XO
+LklghfMDVSN7mwxchsK412YQTPIfeUvjFRsuGU8sI3nCkQO8F0HH28Q7cL1IKrA
gRSc010OrnKIb6FrxBnNyCoIIUxQpSz82bhXDCFRqg5AKcirs7X/qGzMmMqGL2su
inY2xVBOPphZSBrXZCBz/GR4TTPTFYiEX1onSjZmxIC7ZlI6ixzm7T3II/QOTX5u
Y9QuPp60Y+mExwaFwlDbr15MZEvw5xYHQe19653fLIUbXIvZF+3DtMNXFTFwXqIj
i9iZHcHMu9swrQcD6Yr1IntVUw6zSiiTOQxv/n2BqrpTWwYRFU22mkHhzWBib3oa
WiPiM+bXzw+MmCaoUO/VkP4zBbZdPr0etzvn5k2O+Zeczzv4YRCtJKogaEJFdbjl
sS7ZpFlYgxENRvXMM43hWed2DonSDZFV8noA0nU5BruNiA234EvC0ogwMb5SGmZm
mm8EWM/FvOBNNwcbLXEDcSVTHqAi5wKiNm5xXxmK/JLN3iR7ABw06oxOytIo5Glb
rpuqbzE62PyVyZdrnJ5rZrHcUf9W+2sXRTX/OQrIpLiDuhDgXwFX8L1gKObppMtp
xju6dfNUmiz14hCJ5pHwS67lA4PqKVRpJ44O6AKE6zn+pv51UAW536Yw1l/E3Uvr
iN4jtWzfA3svO2Stfk4s/Rv5TR3ZJbfDv+zVuy+h2MKj6O6dAptTCJw442RWc8KZ
2DILEgqxCpPf0wIccQi+l9y94CKqj02vbmftas7RKqJjzB4YmqNAVjBcIbgZPzrJ
UsPbIZYRYTpfR0NPaYDEEOIYOlRI0L2vnoIoS9uLsLfA+/5XHxf8MXtijuYc9Bay
DLB/z+3Y2m/0lHJ2j6BTVu/X4AGqOyaiqSppc1ozWMhpaAyT1ZLxaz4PY0QvNVjT
lZJwbbU+sxNNUFne3ekPdB5dHM36LdG7IXlmGw9YqGSfQUHRjb/Y/GPx4zG9UP/o
geuf+MCyi8y2yALzaSSya4dnz/o415ri0i4LMueXl0W/92CllmlMfEtQoxnm9FJ6
Ks53igvYwD8EwK3UQzta8Rpf7sCxsxY7hVQdRx+G2RZAyha9iKD3Zi0KlhF5McTz
EsF//VaA7mBW+SBtyMyXdoO+esHaJ0QzCwZWe7v7VGaXuB7yeGp8LeJvo5f7rQjL
asD/xnHShNjzMSmrchX70BldfrCp2HNNx9VeJqAwoKrKpbDp04f0Ro0RRf83T2W0
OkS3jI42KWKypWyxfqcGoiuq+lZV6ap6gRiOoQ1cuQk2by0ml+xAqNfwX7BLs1XH
8zX4oMK2HMdnl9ZPa09Y37cWPlbjTUPVThfOA/yhWCLlTpvzoop6opv8l33oOVGS
y3TBtShupnc0/KbD7BL+biEiY99cCI1XtuNNIcMj0jfsoMPmXqnG+bjSNnlZKPyH
lWcm7n1RRJyxkFHouQapJq3a3inf9GhVefOCvfm1KKKVRALsasajw7oDmIWjLcxU
KxKU9/dI2y7UQm3FxX88C8UsOuL0JaiD+ns3wHqZbPraJ6MvmoE9kHBjP9X/6N5M
CxxdDriNB/R9x3GzNqWa7RUjGWjSVI9+3X2n6Fgtya/YXPSCojUrtwOgriqfr6dH
ponP5aoiC+c0wnFwpYa0T62o7y3+aDwYeP7cf1GA9xHVClIDO8r43q4FT5F6ZnYK
zmrJwY1HdfSBcVb+xNDsEHWM1JjcBw7/IGESSb6j5PHtO5/1yvEZ3ceZxyiy5QnE
r1VkDyLm0apew+XhG0tAzTDyDJ5S+pRlO+J335bfXuaX05wDXuKb7xBNj5txZwNi
g16B20iTi4atOt9SZF7A4+MAdzR/z+oHrL30IG8Nqy1WJIEEQdc3SFZF6x+cggr/
iVstoCEIYoCnvnEM0bSi59kYr045l4EMijFzs82T5aV/RDQAyXiz2XaKX/LaWUZE
Gxk5xsbQc79A+FLl74ryvpLHXpEqA/xgnPX15F2oB7cf5b7c259HdsE4UmGB1SZl
0Ksrp6YovIa5rIk7C4vWm6bRlbX1MIpHHbfkaAoX0ajOoMegWvCiC4zCKXBJTxsL
0bCYYy58UYNDTEG3IAUwsG4qy8wHwYC8dTRBM9MkVkujSl4mA6iM1nWjIc0rPL5c
ZZDAWIvQ35KGxUwf2HveJlMzgeK02a6999KM197QG3vsN0OUvU5F87kXRaklVR3v
8vlAoqzyBUnSzf02NxLBA1R6feucJrAhX8ZKYEgnOM+1jwF7VVrttCeh3pMyznVS
`protect end_protected