`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
ddtXksX2+yylW5zu6QL2Lhnb2d1sD00763mmSITNX595NcHTEkwn0zB1Dry37fOW
FufOhVzEJp80NC5qZ/+F0Vk7Ik02dIR0elf3clrjeJRK85K4e3Hoo4xn7YbFUIms
l/8VZSb14+JVGURjfswrIyCUotIzlzVYZ6gzoZwDXIi5gQIBf/gI+KxNXPaKV+PQ
Ufys/12rjO6aI/pPlqSm0hCvftmBcnezN2hk1UeXgOIuKZnogjOsf0iJVX2aOOWE
6pD/psybjbnsNB6kH5uFTA5frkzIzkzl5d9+YDm9OyC+k84E83I/7/j+rk4L2dah
QJOvksSIzN867/4Qt8qYTQ==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="MvBXkzurAa5VTw+1JJ70nePUfoQXBvZOku/SMmg4TwQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
oRtzZL4VJ4iwysPsC8SXYCzXS8Fw2gtZTOskLcDV+1B9Nzn1zTyNtlo6lNICRmmK
ZRVu2BmCc2G+fmzynYlNTnSa7C0Cuel6FYpxCBlOuk3OF2tzAmLAuDyOH3Z1Yjzk
a0aHuoCdIRKv7BrZCdALt03JeUmXKPdOmIlkVGFl8yw=
`protect rights_digest_method = "sha256"
`protect end_toolblock="Jn9CQpRhJt4rnzZPRk+dOpzAubz7omckX1MrFd4p81o="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 15968 )
`protect data_block
gD6l00tciPUa6pDNTk/+t0OO0nC/UTtBwLB41d4inuAUA3i/ALrNyoJVcBnAmEQW
ptbcNp5fxEUJjnOxnedyZEuEBxWRieZFQnkRdF269oPUpLQJksk9fRXrEnuGVs+U
+OViOSdA+I95pLitSNnq6TMkexlf9Hhh3/iHZWcMjAzCaFwRUobOixTJC+YiSvn6
AOYjYC/sqZOkXwWqVsLsBXGtvmrpDEObnmm9pA5lPanSMiS4igffrodJ81+mgoYY
BrAYpDp7U8YDrXbI8DBoFjygMKVOueRGNge+/Zn/2l239ECu8eS9DuvAMYoP+XKQ
LDF9ToT5l+XLdrUEsUpfYM/vuKhkl32ex9c5P2+wpKAQdY/uv5mJcAWpuH08weiW
X/z7AborzavghIzKbQAquFfJVNlh7yL08NocRg6ji+sOr9fo+RVWI9jt8W+UqcGW
RUGJ+3xAyXS9Yll24gEsHPsxk0hRQOfzAKbPlsXbSbkcIZK/n5U+LneJ407/5Kf7
g1PNWElyI0Rc1Tn/tkM0SNT5+h5u3DCYHhHX7SzD5bvzp/pQk5hpjZ87ymzCMuM3
hImRSEEuwqdoNks/6JGkTJtCyNAe3E1XANVSTK+nT9weraJb2vXDG8q5CcG3k4ih
uXd29EYClUtNe1SDoUPZV2jptRwNV6ewtBTmcmoJ7MnZxRLjqQWNZUjrTarxd6qF
tXI1emrZNyORaRnAgrM20OdlNfggbcEq4+JN2IuEiJVXngCQfUyZ0j5XZEP6HhFa
5c0T0fWP9l3BfjUk1XhKsaEWezBpCcNyBFHm75fRG44+WBb4T9PgwfENa4vTsycM
rHJD+0ubkdzHxJKNg/rFIKXNSwySEjRa49gXfmcucAx2kSX1JsspC5wPZ7WJSsfN
SIQG2RvUCrxwaqjKs7qNlarO0uQZVRCWxWKqLAFSpzDpqf9YJbbbeU1hldwpUhf9
B5B54j+hSOEp7GsUALl6PGRCwUcQi7SjVydnNaZLe2J85WlufTB0Ckxw2hE8e+Sd
nlRfbCs1R8D8b7CBswe45lVTmiOPsxUb7cGncoQFxHZ6tXq874wp48PjUMfPkdaJ
OQtTLfD5BEnnUcFZUxh0Cn1G9ICYUvBAatxbOClW7sLoh1z/VpEHumjoCBoQvqsb
gWnKfIUaI/lQGCwapyjngEercypNg99Hh7x0ppu7CF2iohfwrv+BQwS1eOkiDnZ+
BL1m1QwmIDLL8+UO1Ydn7paZBpHX5OSg+9xNC0T153XirWJ5q4PKqv+blNaHFdBx
Wbqufv3MrnJ0/m7C2LkWZ8HiF8gCc5CTarQ3PxkrqQigc0grFIJx1DMWZwWoH42I
o5053nonB78TM6BlDVBoXqnOK1IiP6Xm0dpWLrVd6jURW+3G0+swn0qQu88foFJM
egg1OjQd0hWX3QMJBx1kBIodoSIDx+JWtUjsMP43W3fDSb/HLx2nlg03f7AnlRyz
fgqOqUiAC6ME59ahBv8uBKPYDqChg8NTSxehszeyFAOq5seHe5kevYSnVy4Pwane
ADQ1tD+ELyoFxrzO9RY3BPlklfk4fBVkPKIlYvdgU+ivstTPPX37AyYkopgUTVHV
wkEZLszULdjLaTfNQEZXplroD4l9ctkozhLxHDSprKDv2EpL/2JJMIxpQHvc0DKi
7e5Iec+bYRJ66G1pMNVHnx13UtlYx1yYxv7HrhAcK1zQJdqppFJQrkU2wE5oIEFs
ELHwrcaj3HtVi4TUfpJbMlj/+th0cmp1qdg2yE/1MK4sy0YMvL+PLDnleBg5oJVs
PvyGTdbuvkS1myFgUQ8Hc8w6YeUu9KGOnHRdP8tdz1sexpgZx8H4a4hiCOyzyBuU
BHU8OduAUNq3xCITm44LIabyZIoGilE+8+xQWVPnCMp/CJ4WevR0ck4sq1xtAYw9
4uWWVNi8Qk03TQk0KLuLbezUFpiM7XTpq9YRKWMalcgxuxFHVFrDfGvlX5DsKuPF
Zpcd4gNnMY0m5uHnxPpGvz9X/Wb7jOz1t6RHpMXFD6UgPurrF57YWdWCOScyDWqN
EkRfhWmIvpKf9zxo7w9OwdR4dfi1wa0+URbuFoupmKpX4bYT8kFeag47EC0r/pqG
zFDChpjwgKfNR5OanEqBfSrs7D4iOpTkB0zuaBlFK+Xxl8Xp4bwavl8N5BURVg4P
obSxzyHRKBv87g3930YO/3ASCkGwAUqX2NSYndF2WiMZ8QAAhRbYYwYrizv/mTpl
5RwEH8ot/8602S4gLleG5p3tcNYWNV7SmBTjboCtHpXB3AShgJPdry60rnvvAhZw
i08izBdLXs+YAzT6fMYmY1tIiPpm3NSaclIpzquhZvDMeGXViCJvD2jhWqICf1Kg
Urt/Axn9aOFLXMJLh6XuDcFzNH691bReI2ITtV3ot0BiMsFq8UaSDXYK3jeFDASg
OBupcKyAqSda9KYcYUpqWo1HzF8KqGJ02OZlr83G7GZA8E/Xcjh+yJMWDB753CC2
0CKqm4Nw2iQxTjk8a0qWM3edlDANQkeXuBRTup5mARAaK5CHs9MKCEXiEjXIq9Ym
yQTwRU2KsAbrgBbrntGNDs23xva8yq/GDmqNG7nSVmFnIMjjd3xOmvMhuwXkEZ+l
tr8BP6APuGE1kzFDTvn0lO2a576u8lCeW0igQsCTJWDK9uN7CUdHaM+6XRnuEyOu
Numk/6z9CQaz5sUZEfomwiibkwLo6SzDsyTn/bwLZC/q7voMvkUa0yxfpIfxvSDy
uIZcbjYoe+aAaEASh7wAOvYjYJOI4BUOIVOzX1yYoH7npB0CA6KOgs/lOuASD0cy
kL3eeL7K9aaWT4gsjt6nz5i6/0n0ukV2gWISGtbcq43IdNHfg04PRzfuBEMmjR1N
87rsKoUcSbcYW9pJEz/D2hi26IW0MundiQq1PIXXnDCpuLV820lXEPKDxyoze7JC
a6g0ShephmHexdww1SU4aFErR5dSmyWYWsMuI8wDa9hgtmL2N1DCjdep7d+03cqM
6pBQ06soUlOzN6eKubfL5bqo6VwFvk+3lZXp+FDRVsAWKPkhcdOK+e1RGE9L86B5
/ATCmrAOlTCwsv8tvGNj3qbgDkwOEV90S/mVE0cJCREwqmzM1H4MkgR9OKq3W5gX
EKbj9YVxuHdUuUFhVULPCdgnWZHFqA9JBwwHAi+GDkHQ17i8d6ZeYuAu+qiBCMFr
u7yLSa09cFSQWCJQ6HlMO4mTm0RlMs2d1ZtvAq5Q9l0z3TDaAEGbKS15fb/cu7YU
uLs/31QFzz0CAwxYo0G9dE3g/X++E9s7rCg0X03I1to0l2HbbSbOlpfQmNSn5x4o
jDSVRQ51UL50rg8wJFA/JKBzpro4ACFaL6vfa7EL8VygfigUBrcJhAAUQ6pxwlWV
Ky/vw0C56OKFwP2QnDY0pHlqBJgNvm+MP5WI3l06nmso9NwWbZ+u6M+cKLLZDbgG
iYNhvi7HCAZp59o5SnMG2E6AFT8YCOo/+yUFbPJzI3br7GFwF1sg7N6O8GztthyJ
0iZiOLOqY3a2Hox/BNeVgQcYRtw1WSTO1DAvSRfylPOwWgsqYQXeoPpGsYdrLKEt
9wkRNjL9U+TKL6xpz46FqihTWIfkkwbibzBAPdeuXZGVa2/57EEw5ZMuKTY5UVXG
UBGns3boELnL9wy6SL8J6RYWIUmG4SUR2SwoOIqXryRZNkTSphrSI8Uci9rGjlH5
rCTUp44XmZMNQMy4HoyH5EGxExFSE80UHqKigw3Rrmy1BQ+xSMmsz6fJ3wHPWmbl
pW1WR1NT6TAYg+IXHKLqV3L8P0iLKeG1pwLRUtxzxlvR3b0wHnKZLICPqFwALQIv
2pqni9W5KRMsX2ageRwdg3BWPza8qyaCTCE7VOCxrnHybJRM29fYEjmPXUE6pXKr
V+FCqTTqxEJcUtCcsg3iGEyFbGuJYHrinEDw+sSakc63y3P70wevXINFbGL/TRf7
k7o9RSdHOriSQ413UYwAs2eSUN5Hb/S1wtr3OesdRovh/JIJ3D2y7mBvY6Y740YW
pZ2j4DJdqOSdBzOzORbGMBIx0/KyYGf/YHVJh55hIntidX0RiNfvUJYdW0tWz1V3
qvU3MFF0uBJVykGUs8YETyeXR0Xo/jHrYIQ7ZZTMn1OpEdHjjl0U29vVHxEkiJcX
sr1LOFejFuhBT3+pED5tIhbT5wJnDmq446r58EWf6dwB7KQKHWpa1a0eEODoyhdC
XJ3x7qAbakZACerxtd29+znq1qa/+4X9iBgI3XxSYzIL8IdNPXVYr5HUXmN+3i+l
bz0iHIPAIEtQQ4n/32PD4ATFsjrZyQLDq8M/nzx1CQgMo7QviwDS0Efi+PzX6kI6
PonRVMKmC2yOc1EbZu/R3Rl9Pd5LyWqozPg3/MfUKogiKC9sk1PZP1Sym6WhsRGd
SC/7z+pqizx3lkpGBGuVYRqhCiyRYCQCQHFFxshoF7pqypSPpvW2usVQP0s4OcQy
/etHLX6qz/ihii3Zcbb1IEsfwHZ8K91un2kgxxhxd0V6Q1P3F9yP3sJ22LA5Thz0
szdWv7z9JwUCNbs0WUTXRzfpeBNABVwAWRQUMQKFxNWDQdnUMGNc+LS+uM/dxCCn
admlcXdZqtoIg2MkCpiblL3MscxoRNUEavd04yxfnp0NO4ZuT+ofD73xnQpk2Vb8
lZqWJuptJSMclcoL66mfn0r5QpZuQi9MSyEmnTHw4vAPDr1hEN8aM4RxRP7vhuYl
7wG36aKda+op1tw1Z5hYObJ6q+SDQzDiikpUneG78/XW7z8tAsrvd0TcVdOBCDJk
k8hggL4L9kT/RZdNNbxLP45FdSkETapaFrOcuWqrTPSBmPVcxcPaeOX8VsCXcIfO
i+/69Y5xYma92HsJxn5US+kcB83K/zXFSViUU6orPm525atgk2FhaPqArnkYodZZ
BcSEQZsgjnP8VE0/IpN6yurefXcCf2VsXlTe139wLBRTGQa6OMDilbAJ35YVyWRb
ko5owYiATEk/+vUtxfGtlhn6cJI+Yszp+r/a3H7zVszwwQDHB/SY2+2/U7jeTxoA
SPaEDWzVFySIolxFmv7E4LDnoqr35HtmVI31pbGM4P4ypO80pgEbeoOnBgjBlq/2
CqWP5xN5PRXkITq4rwk/7a3ricIhB5xxH2qOleiI+A4UyecYqBtQApMy9eOYviq3
5j29OiZVoRlN8ztGiGgqv0x9GsMeHLGKAO8GNwkZ0tZPaKmtqNWS07NUE8NZIn5a
jhGXZl1/udU2RHViVoegBnHQ35GXSpbpNn6hx89MzL+fuYLsQDFGd88fgsxx1rnT
b1WSiRiD0+OHHuigsauMnjccD/JvGBHGv2aD7ZoUjWE17oWjPXPorSVtVvbevJ5N
GzNrFnEArHiWU6bEcfDm5t/3q+HBB+IvzHK6aI+hvYuLi+ErQ41z6cYHEVWcqCQi
4QBNOclSeUj+p6vsa8T+d0u7Uv3RXQz+LhKakALd17DPJ2RGvYr5kbd/y9D3KfJY
6zQ16OdWP7R/GhcMMQXHRJ35hETpP5hllkY/pD+tjczdf0fBddjZAa6jiD/DDC8r
jFiOyv9xebQ10fs6epZmzvDM/PeQ66VMOvYGv2ymmRmbyT+g729xsbNM6md+uNYp
Vc2E39ceodkrtO5BBdjFfN8UxkQbTjQx7citM+OhSf5C8pbgKWcqKMd+taPiGzo1
OkL1hv3C+N3IwswAA67Y1odDj/+FbihRG4T4Aov2KHSh+/lmKSz52Q2ifqeBIvKs
YxAV6+m8wg7WNiy/EmseB6I7EeHbqL4rW5xrrtDAlG2X5ctY996kXurseKF9Nbn/
D2nqc2cmx6YPc0WVE0lQu2KJrJ7iuusj6zr4a0r9OyAtnz8LIXe+iIN2J4qqHpls
BrhQwEMO/tWhbwhvE9rR7EQyO5Oc7m6U1aNDGOUn4rWRCTxXHXrO7KiaFId0kECc
8zv3WrpDYY0jIIKZTw21tfiZINgfwhyqzqKjt9cA4YkMjAE42HRikIGXIx3C5thm
B9pIp/yX6qkmxu3VijGd0lCFTvDl4bvgCHhvVH/w81I+vJ7UKptokaslAyevalnU
ztf50MdrcdG1elwDdXiq7ookQt25HYJWC/5XOFk7llWI/+cxgnMLXd1b4ACRhQuo
Q6yzOTrBCwYDUUaI3GSG0BC5Hc09ffNKlcaFlK4VakvnDoXqO8FE8FH8ZRGoaok/
jpF8SAP1A9tQ5J4k2MdMNNpt346Vub+9Ma7dRE4iWg4dLrT4tVq35ug7c7M//9VW
b8fKAE2Or8Or9lA9PBKtPp/abMY4v7rJlvvQ2msOT35CPLpGGSQo0BfGYyINCYRN
FSXQz1FpZFO8BVLlibi0KALa/jaJ1ox1nX+lml3lykGM8hN+ZFlwMK/+vi/YSFl/
HFbewP/p8udteUMoJJxf7SFREdUpJjGndD0vEFCnURrDYC5BInOGemVjkguUi3BJ
b14RuTr/7aexC1aggt57RG8yIoRIMakypoRPS0Vp59WXSS/V+5W84N708hUN+yp0
tb0Jm/gxLasXsF4UO2jXQ+29+In0jTdcfLHDVl8jDmuI0XHBgsbzvcoRoG4izSk0
YREZ3/NvPCesHIAv3jM8ShcWu46wxpa0BMBKPDa5HXeS8+TMdLoBzxt+bGKjBax0
5mah9UdAttU0XezyFESC7nOk+D18gZCXYCodZguTlvT0d6FdYFx7q8uGg8fiEQd3
VU8FAZJrASxAVSLBh3kI11JvnSClLVBF3j/Yx3xV5XWkrGokT16pjI2diR9oqHQE
9H9IQbpDDGJbfXlNyzxN+cehAGNNN6uZo5gyRxFqoXR+sc28B3tK/do8QF8BKEo3
BLxzMKlzC2XzzSgatDJhIk/YY5jAPUMrrT7oTElwAmmBo4lSkEr+LA5vVmx/bDOp
st7Mi8qc9DVrt+tZS0ri17hHjOWRfz9pxHEzRDbP3TYpzfL9kNheC+xcQA9UtbQ8
QYCdGi68i0Lb0F84yj0AcDaEeGP4TOJbhGcmLFdJmtj33WULln8fiHgLw4nSeCko
lrOSmC43tziJI+fhaHolV19OEXsn2YgXfug2ZM/yj5OXJD7Nwk2tKCfUBLTMQ4Um
60EujnfBNvzpshejUJipMG0BKxof1saw6OnolGCUXoqmLBWrLFGEN432v9GqMHaN
KaAgd+L1/jgx4nJMpbTQDZ9/WNAyGZjnz/vvVihrwnC1L5KWpEuBsRu1pCwzDsMc
qMXKP5F7Z6EI2zYJ65pUsW/dJz3/RoJ51MH6pt+il0/n5Ett3SJGwaFl1KamciWw
iacXfB92hu0479UlXuU8OTQ7LdT0bHmdnfNjN63iS0C8kK7obfyqiVxH6VqTU5c1
RrBxzcNGw8DUvYlJCBOy6DrZ5cDgQXb7FbPlbA+QLA8cyYHsO8lYW/ptyB2reMEB
FlYjuDc9Pcf5ssPHmVu9Mh5KpmmGXVXuVs3lbrzl3jTqbogoVhdYosRXCTDuq7R/
1Y3zvKFFETUyYCMCr0LDfsQFhgZmfbuyAl80LmXRVnmpVcDsZU3f8oadhpgRZTa+
coEMcuYCow6K/ZhRE8fdHGkQh5kC2hVOS4lFH2xjY7xaWk0s5m5IrKr4jvFpsLEA
9XOWUqsZ0cjcNBdIK7VDdvIZLVSsZ7dqkBmQClh5K8Oo+wca2Yprt2R/jd6gT8fj
Hta6S2VDaFwHPW7ODP3PUTNY9ms73ExXjVfqN9z0aHCy4fRfj3hD6Cwf2gMo1/Yb
2dtpgv8domWGye2gq7MbXkt2glDptNwhdOhvnqBBLcdNsv2F9WZt/XMIXOuyL/7b
5UHMKYCjKvmDmhHtc+5Ue6bYPRccq8CNJugw3z6ETw5OObeO3lcxI0cVIXxV5561
Ei+kg+eFhIbuFteqZFP6Yksbn/dpBrG1O/BGr4U/QVvLuAFbmYe7ICZ6IL/HJDvc
soXpw348KAz+JMqxPJWT8AiGRgA7To3g5kb+Y6gbDmSk5OZ0ioKjTttdKBlx2zFc
hjRahlipox0WVlyHBnOwtEbrTH8Hhf1Ou7dOEheBA3gRWYg2rpuiSE9BfYtILVQc
6W3ihC5QqDMivFTxsT5ZcYDy3cy7+DdU3A6suOpuyqgeQCXgPd0sSAqtFPQk70ib
WHsWv51M/b75DWJkPzkAbsrsw7oI4D43aLhhevm8Y5eGs37d61jnxmVjgIvLH1nN
I5nU+Ua2BnbSXGbHD3YCeFUNXrJEyBhc3RepK1chov3pEhX82KcHbuRhoxkhmqzT
vY0zT8enWk74fGcY1wDruhJGLCs/6zk7vr3wPiEsDW6NP6+GqMgTrQs76tiVS5pw
UNdcXgZSycKEWpt2b+zHKvaPX2wdYTSOp300IfynYezyE5EdvX5Jw3Nd2A64atsI
KckrXRIh/EU819AZo6lPv6UetlSirfANQaTlbMv2g12qHBqcaBi1LA7L8q7PpcrD
EKHLBb1KQYUfNCirVIWlTCFJUk/1hXrASCtvxiZ8vl71GNgcp9zTfKI7B+ybobTn
UHldtPPf6cBNJZUx0mscrYfTxbLANukGOrhBC/5j7ML1pyEfjRcyz7PygoH1q1om
pbvoB0TR5Nmgfvc9MtnsoCVSkKi3wzOi0T+7gX8zT/6wli6KZjWPpjD7rAdYo4oQ
dg2bbAm4255NQKNqozEngEfTCMczqBFnQvFfwSPcbp3GRIJkRkHldVoXISlMK8DX
TdZwy5wdLXKRu+pPn6LJl9GiS2KVMUp5NfBD//JphxwLgQFNAwJFfm3WQuxzKOs0
af8SeiKBgUtuL2rVAVdb0y/vn0nF7xsmXrwJ09Zb884SecSsinA6uLOEAraiUpAP
gOqTc0I1D7A3GDM7dEWJ2vpK5MAIeJWWvRD+1zgDIdNkeI+ZipEh993NWFDJgzBw
9oe6d+gwXzyb9exoM1q4grM9NUqKS8OR9bUoYmPcEn2KWoaERDznX9u4A2JAByx0
jRi7YxmULzWBzLWDUbWEeGCRiErICe4dbzYnHBORidkfElkYHDwMobvBD1AV6cok
cgXFGsZJ+9yAa5jUnRL4AScb1W2/6+3Qp7z3lSR78BJM+vmZw+vdO8yBuzK1rUIR
weMlQsE/d3HSEpJR5iJbnjVzE3dFhzfsfWtMOJIxORPlx4Ja/ofZyeAh7O6rw0I1
HP3lR/mAQS76Un1vC4Ac+ynipRzV7Zr4WsRyANrZbcGrwb4XjpVpdLOOHt+RjG1f
ObMBP8HifgoEEhot9dER5n+R/zr1KnOX78oaSonbOXW+OgWcpel/CCuOhfUGDiX5
ZTyEzOiY3KwbZUgqmickPs++IttUTd8MTO0neTa9OUqs8x+q2whOUWdEDiGVsbf4
GbURJLaGlugA0+uiUSj0ura00huxOZtt5RyLX+lR7WV9sWGnm3sTjqf3CPnEpjfI
/tZRf09DmNKOmaudSBI1/yFroWlV8whxX6WTsHdemT2sHaHNzMTzcyIO66oq0ZUS
Oi6CX8+e55TVDQ98plgaDPjVyOYeFxZCC0B93O0Io3EkJLNyavr3wj+dtHIZAMFd
0omn85tspGL1cAd6Qrj3cgSx+atUPXQiPfub8Q7+IlOL2BH2wrcak/MpfmpoLrZQ
kip/usEn01hA+sSly5t3035uLu0rP8+EByaieA+H1yrOw3ZwOOXVgDMTB9DfVJim
0dGWPem0X0OuJBD6sjAPtvW/hQE3nZsU1vroxpBwmQUNtw4089TWjgdQIk7lxgwL
j2q6c5D0ImQQALHu0kqcF2/DrKViyeaR5SGn45QEucu35FeWXiylII8dpbjJf33V
M7MbdmL4XLp/IDMSDSXpC6NgH291qHnxQUpRlokTZJewNT4A3jC/4ZnRxQ6QY6un
5sNPVe7Sqx+pPr5D7uZWoveRs7iumV47eHU4m/szxjvknpyYMLOTMO7jWpxhNn1R
zNF3LO/BF6dLeEOONDdI19MBRZivkDjrZFrU3G5EyUAM3ipzdn8j6uUKviHFqu7Z
OX9nlN69xWjclOiQWPImlp8hGyv3Y6tOhEE36tXmwaYdP7nzvMfO3KTAUdDFQLkc
I1x63o18E7bhDxmu9SMviqwR5EMQk+ga6DKa2ut+kWt4dO9MtsdeElIqtuc6SZak
iCirZTNLpl3hPocm8cWdApZmql7R/ACSTbcF0C0wkTKBKnB6lebX3BahbfoyFyGk
QXn/g4SCOwBCZNHKGzt6She1FNs1e6hWTvwkq8nWJcCAN0VEeV3ptyH85em4Evk/
LFKK5e9TeBhi3IbaontWj3i0tTIkKS0vmKo85xAAV0FtMTjC0EfFR3tiz4w49fb8
o4RCV4SjUKeRmWZE4s+k7QvmTbB5FpvJhzRYHtUVxvpXTo4aldGP8Bn48NOUztiB
wkc7LnBoWFvwc+/AgZr6Oy3I54Vt+KNC/OZ1322nzLrGA9jZVNYLnWcME0yYVeFk
AUKc1zNp+XbSgfw+0aiJOlNkJZmMMR7E0Q5Q5w3yI8ABiqYzMlyUmPRC+DeLsGo8
5M6szFdM4ToUvHRNr+2/yaLmUVzg3eQa4Wf39JTXoawdCnXWUww4vwskq313m8Bb
Zr9pCq1NBKAcHMSuvTEqQTjCgPbh4nHhFgPh5gOsk/0xZITvf/19xCguId6fye28
TycVT1L/ScY9YU/sTI5oK/odK/wSlrS/Vm0r1TKc1NS4dcey1GS7af84JuxYjZW3
pU63C1lMczOGff3NCm4IrgLBOdL7gb0RWUOezg6n6iDVvIyYPxFfibDufTp0k0dA
8qo6slRPPpMSdc/KYOGK4l6mkqkVQ+dAEOkeg2TZKK7Doom4fnSKlXvzSKhKUqYy
YzSlVnYttRaDQ70C7ijtYrjTG3qShF5gJU5t6Dvic2vEZmfwW5MY/bs7uZWEdbZS
5Vhb1f5K2rUHhkg35rX8XZzbXPz0xG2Hue5xvKBDyC0AxHWS7oALVMLochaffHSY
xUn6HwFVZO14gxoyUA3RzFW1xF/keKJYgdyyQNfBxso2MCVIbkZZh6ddtp/qW/32
Z/9FRfw50MnFqjAXPMSB15U+igOXY0rCo0r+b2uWXDMsVSZxmeMr8aXofO5b18uc
bu3/hEb1u1EXjmhFEWcSM9aL5QmcBIpvWi5NRMzY11KEn9XS/9/nTJtOqEotGvPj
FkDMj+9DuXitoUWcKKc6GoNxSyYC69vU1mSRiu3Fs0VZWzrvS1KowX5CK+DgVTRS
fmrKSEQAdnpH5JBHxCapH+iMSuuHxm15Mm8bDxwOrSAN231e54A9X7Y1M7xtZftZ
N9EM8mgOq6Mz29tK2RgpX9tV78Lb6xlHk1KfYrSOZr/kTb+z+gjJfNggNFbn/LmW
smkWNbKhmWtK5OEaoxzZH8OVGsoHeDi5DA4iRSxqBt/1Atpu9fnVYjrUIf8fbZ22
pbq+x9SzmFv7uHFFZ6gdStEmdpsMHn7PZBorgh67Hgy1GjS8EvgWeRRbaTQrMOsb
wn9FSr3bfk9XL0QIYEKie0uccxi55AzAmT+GRlaxu1/srTjtLejCvhkLeB84A+uh
ROdWpXphVOfmAomuklgZvJcQzJ5IRIwjKuhUXKYfyNuFg5yGpaRA+nXT+pzSzI2I
zRy5lAgctCw2LnPbfxEni5Qa9IdiOkq4BdQaj/7d8es/STeJncUMAexiFh6LoYzo
glE4nmlcWi/e5Bxl/8w4GexYc0Plna+dmQ2g5Rd74K/HP994Pa5swJ33ZHQCYn3W
c+NS88b66+0yHRl9OsRVnfGp1tx0JHW9FcoO4aex0w/3nHh8KpMDrcAJZkMkJU3j
byZD+CRqAbgSwjgDPBqQlYeipy2SohoxBp1AbmDXVnQPtARN958PBE2S/+6bnhDf
SSXDPkOU6FtmF3upZdHzv2JJ4E6ijMUHSMOYZqqEOSzYl5fbExDsG6sgPDJ7R+x2
lZ+PuUPB1kl3pmP9fyB49XZCIRg4Ny1wqvdUk0SItt/Zj02YMvRsbV/bBe6U25eA
rjYkChFp44J03GVXbZ8xoafK7c8wT7OUH9iiQNckXcXJCV3Vn3fELzu/Xy+GZHzF
PKPI7T/7z+668f0s1W9smsSOoQ1kp4ZXN+dcQYOu+ZwkaqDYmp3rNuEL1pI+OePX
rNXD65GWkjAs0QpLlmy7xBW0nCdOLNzYc2I7HpTQNBvxMaT4JrTU+trUJLa5eekV
GSQf2UwceH51sP0+9/l4xegFrbsvxsgT1XUMuvmbya63u7T36NOVifKk5cabvGBW
J8DYozdu9L3INKQMgOXm96nF6h4Xt79gNHYVYwhcCDfQ1LZCKMq+DVdifOqqwdb8
KJaTg3dr6nwVB0c7utMcvfr8P6tSUrRbl7AXMig0NUjjC9E2M80y5FsgRELSdQ3D
QnMHhi+X2C3Xpsk/ihVbA44lmpyQyYL87NRLLniL/lqvg4pM8cwR7Bk3gxz4JqJI
9E4PPNo6S7kcyS9b+22ef+Ay0HIVA+KY16j9itpVgdl/haQ1izhpRE6YPCjfvin9
cSUtOKmvPj/cQsXtfQVxWp85u174hUB2edo89TQJTmxiZwKMkhCEpdZRUBcSI+1H
nBEptfKiF/tvGKS2Ef075ziLR2jI3jQ3ILgQ2cFzJ7tpmEPn6tphz71TXtxqPsSl
MOynMvv6UakGN/HpuAJCiY4tPCq0uSijeGfiyv2S2DuI2n1FfnP8Yaeaoc1ZPXpM
KPghLuDQxWDEX2UErluMe5tz+z0wXsjonirIjxgY9bK+9PekTs2i2EB67kh2MvHI
kr3iVvbeG0FlfonTBJzO+I9Us7ro83NBFEt3oax1GQ7sDEdRAXBBzWyI4fgkarop
YbEh5uYLacJNHEeHHVt4fsdksQf3PxfnauFllC8LE8H3Zw7+JzXa5i6c14WlgDtP
16eWG3WUEG0E6F08G/1LUMVKKqOQ9bnhbzINCJDHjTj+dCWClu9Fvd4DOVoFV/Z9
opS9qXEa2+qTyfU/+TiLkRUG1aUkWV9a2+dplQT1b6OsPFU/RVQ1Ales2pp3PO3d
tbWdd7tX8DKmAxYsiVj+n5bEYO2PBAlmeAxGbP1/QsbaOK82od+KQBdzY2PELZ6h
13fiA/gXBbHlGVDWQoR1TW0CQeiz/6v18OoxGvPOBit2BGD1qo6JOC0nAfwEhcGe
tYx/eye/7NvG9HVDYZcrct1YR6Rr47TpS6Or1UMz5v/X0kH2s4e9dP0Gcon9VVaG
A/aY//dewxFDM/4UONGUafUWupwS01QMR+0QLMACE7QzmKUrKbtBnSuhKM5yY/az
XnGweZFG9hWBxpOnp98HrEz7dU8D8OOg4SCLCmyEWmYnRh4SdBJBNwOMNR5GJQo3
KAcXF1zIVWd/QmdyWStu9/3fljOwh5CTS5Kl9/tcq6hNrh2VRiaChdBnV+nyI5S5
2lfMX79jMJenPO7OQ5WqIL9mpp9d5F7GMEYl2eQfp5VCQe1TC7gLXBHLg7FXzozh
FS4f90zhVkh9Kkk0TYYFsE0ktg0XJ9EujGcxtaYpGwyHbJpG5mTL9+ly+3tsec0u
714/7FDLV5Z/XB3TGIge60U0RTu/M0uuaCOBd7ej5Se7Y6vVdKzk1ljLJLygq3lV
OZtqMovs+TVrYvBbpu+RqeSHQ6gTwXj3DeAar/UY1USeAr2BjtnDHD8fi9t+DMjr
dq1+xaKd3ImrrgJSyJFjs/dBlr428fffKV7m/KG65VfsNk/S/bXEjIFzDG2U5yQa
1sqbE9nEQrPG3hSjFQmRuZuKmJt20s5VKjClbXQrBm0uKnPvg5Nc/1CqnXp9Jebs
NKaQkoPhwELEjEVdcBoga5MQwod4tdx8NgfUc/ds0u0STnP6Z1+YG7bQNhNBuSNd
aMUgo53Txc4LcoPK7d7Kvt6lbDUgQWziso4T52IR/NMaXDho7XQ6qsWuMAloC9vM
hIC3IDphzsL0i6Q8WSPyyJHqUIvPOS94Q/vHNJknsBiu7l24VZmjAsKaasX7VHrQ
gz0D67E9zXsDjoHDi4WQvnZgLh/R/is92GpiJT6d1MJnWQ824SuwibFZoYtMJkbj
gC/9yl0ak/cQQ5yL6/x4hWUR7OwgjT13HdBeF3iC9HPx2u8q+dXQ0minkKCfxTnW
Y51ufxtiiH3IUBEE46Cnbt8KGFLwHL3vxC84C9EUi1uQfOBrcnq+cUE84z3qHl2d
1EvVBWvVznXjZb9RVerrlvP9lbI1GX6o/FxbpB6+XpNM8LY5NDil6reQZ3Kn/fO6
HKwHJcHGi1XMctxu1dG8Im/2Mz56nkyj4jj4GoFQr27dCtkv3VR7ah/BQ8fzfzmu
IUdWoxdqEZ01Pc9DO8A2M9AsP/bGC9PxeatVu7Pf9jtZkmJ0qev4cJMS+WOO9z/k
XFqzhSZ3LRa/s4ViyVgwzWTBA5+36cxRWTvhfCE2pMwc5KBj8rSfBkwEPUsezS5T
oEdWH8j+DjbWLASaXdwPmkRjdIrBa7HctEuNm/6AcoTq5X7kkKyajcPu8FuE1WsB
lcrEwa28D7pCV1s9jIZDX4bTU/6phoTyMBbblMOrBS6518tRq/KzPoBGbyrGmlCH
zuPE+6GLap/c1kh/u2GMI+MlmTUmpyYYJy8kzMZXJbltQ1PuJTo6SzlDQz2yyLuM
cU976GvbpLjLE/IjVeNjKD7ULRh48Dbj0upaKHu6xENuOnJ8wKYTxtHImoKGT1AF
hWiXrCvg68SzDCPU4lIwrErmgL1rwHdxAfckbheSIZrpA0pIOVoFXBHuxaPB+AgS
jfG4BBKE8rYNKTU1/Izw3yau20boevDrDHeuqPAOuFuCztIfvV4DJCpG9BIFVDI2
dniybzCrLr9saGXy/38UdNTHjQ027KAgrZFUx3gtG5gM532siweQ3ipAtXiA0lSo
K79M9oe6Hqow5skHwSDxZ5gaw2zke2uq1GMHydk52zptJiNpxnCGoKFLn6G/yv7h
7jHvxY5JFcVK/I9a2p+7uzg89uWGO9uWdBvA9GXWd4L45GemrmG3TJK6Z/4I4Hm4
T9aKjcaEVn2CyAC3nDogKgfS32ofCfW8XB9TiFK62LGRUDG8uJxYag5UYUwVVpBD
Bo6KaelQHW6+MybQsJTgAAPnqCvLpskxPBPBDZQhjG/q5LjFQzcR9RJIOZMNCfgS
ntsW6GeKu6HcbFXm1EupG5y+hXVzCqnr7ZN9PP8d541M72xqhIaFG1KTt+Rc8eaW
SCAVfX8WGFfRd4CrcpP9vpn5lBHw/X5xA2Nr7Rf8E6qFuVIZNGAr4ZlYTnYkI1+p
cib44WQ+NSrtdaGM82cHMHY8/KuVEFcSFFj63NOBPxkGqB7YDflMmJz1W190mBe7
mbkqMW+pEFgCHsl5Z9j5XnGmSS56gOAlZaBzDH1FG9tGinpY1u2wPUkTT3Pdr9V5
nBGcFIdBC8/CmWB4deRZLFflCi3SbtqtOHbC44gVwNf2O89I6yjybOdevP02hyZG
s9eNuy05H1vnUCBD0sjLax5dZdgK26W9JXMy5pq9LKVID9t9pa8WCu1DTz6HncAY
LJwCQ0ASi4c5CyI/Mf+QF6SIgoo4ReHiNEHH+kl+xL3JgiKzsHufnC9X1UIBC7Sp
36fmAqDp5iavEQa9by4zKBl6OHICyI0W1NV/S2FGE8asMOfEvaqEFJaNxcD0WuBP
VghKgB7rq57tzGppu9CmpTJpe/ZWu0cNabQhOyjGaKvJ3XkOdtn3OMXbniUxtJLA
0bEwrmfrXVqRVUB29rpy3NHyRU8spU/FhoPjiTNF41R0y9lDI2QseqWWwBApo0Jd
MPr3RFslS8y49X/x5b4iBFD16RimZZW93rqdsTk/VugKizJHGyRSH4fHhSuAL6DD
pCOEjlpFyn9MB8T3BFWH+FZzqu8mna9xgklziYM6jT7ajn+Svy4YcFgBc3F19v3f
Xu0EpB+1mZ7cWABi+6Z0nwx7ZuYZCsxYdJWjh4oAaDG3kTbmc4Mny+Wg67/nHkvA
GJqT8xXaU/q82yf8nyWS7rmlA5cBVmD15+CMeg5Y3STKfMRtl4mBPWE/jdu5P+ia
vgP4xoYI0rbHqaGmAQr9r/x3D7MBn1w1Hxmakt3lTeaKwyU77HRB1e9tbEogi9Fb
jlB9ufsZ/NEzGnDKks3PZBst0Z29Fom65y6Ea5nofe05zrrmZMCntlSfD6FC3TD2
mN29eUnauKjWJ/BePvaBS9HyPkkQL6YzCyqMrMXjgnmsFpZ6zOPgg/Qk8ZtHPJEH
GXgyk3D9XpsBj7J+w9yVnxWw+zw1JNVM1wQN/m9btqxJm0fc96C1BiZGfdZI4xeT
v17UPIJi6omGWXBmch7o0Ovlq7S1ZUSSgd/DpzvgOqxi7WhYqbdbqvzpv7mOtIcG
+/qEOHUz97pjeeMsyZPvMSRClanDRpifKOetBBXMsuKAJH3ei0L+T4CCU6oJXK17
2MWvJ+UlMI6J3mmJz9/sNWy3eHAHABy13znifVYZe/J1iby41Kt6lr9yyTn8whtV
CwNoaDRD8l6zCZs8YtRH3kUyU9bgFjdJFpMozZQ4KeVWoO3Ja7wmp9ZjSKLqXVvg
85DvRRgqGzhIkdT/4l3OSZ7d8gGaU1Ydr/1h2j5hzZgG9dLdP2qj9Qts5jwYDUZ9
N32BfN+/lE6m1nvXEOknRpqYV69mtRDZNYHCQSWL/+RxGTmF9z7ErwtDprkKFAoW
faM9/BbvUAZyiI0+l9QsAb83E/qRiCLm/AuwjnVbXL7A5bVZG43oYb9H+fBbWcK2
NPGOdp0ffwzrOkyT8B2DYTVOyglIM6JAcAG32fhXL+LDF8ucqjwgLdYVNzp7Sass
TOiVlesspTTOlCbNPouYKBk1glyHYhM+jXPlFIN1KEodmgKzN4ZGyKEejUn/cr0Y
YbsNh2a8PJGMRiWIAc2f89N64UsQS88QTclY0zk5LfzF2lc8YJOMyzR0mQssQkMP
k6CCIeE2cZJtUyAAQvt1Z+HRi6neVg3DIa4h+T7adNGvQEvENu5WItjak6cb3yQD
JuXWmc9dej4ndogtD3wGe2MhM5txqNRArBpZduSRIoB3EWT/p9yXFUwg4z3PyLR8
1AScDGo+4cRGBYPCCtOSi72bQM3KVc94Q1CjcZeAY+eoZuCDMnftxRltBww/6fPU
kP7Wo4+pKU1qGrklRtFJo5+bZ/BcCHcz5dXcEOQEkc8WfaE2cKDlx9BA9X5RoAVE
CjPm+zgu1nv8jWjyhh5Jl5LT0z2KcTIgL41pVPWP3JS31qFrr/yhOBxgFXSXuooh
MP/AitKrjImrW0oZSJOiEpK/sBOdL3pnAXgTG4dnssK2z0mOSoLiXGIRpy3it5R1
OdQi0XoDsiTXAJu9O4YoXY6IdWQYdby5PgOi8mjA01wyW2PUwndRprdb9F7CNQNH
tPcL4ZMcAgLWGwuzOeXiO3CNqmqSRZnwWE3MIzfWFUYreGnYkbbfgMC7Ciw0+SCS
6yqR3ZCVSa1yxVsDobD9sSP8icMkRyrkvTzg0+WMinOLLTdoQCmAhjCkFfxevYpQ
vOdMB/etI0SP9ZcwuYtAZhvrBwhJ6FxOZ1pxqge3r4HMh52e8Ty+7HwooTwj0Ri/
t5dBToL+qO2q/eQwJplXSxNYnTxtAmiX563Xo66xLzJtjo0e6blhrtu+WClJaLUP
TU9tQ3ejD+f7cRsxiMk5EW6ozsyXbngE/mJcsxZG8rb3PmQsoJrT+fTI5nhCoahW
DFkeisxUyVdOB8VYPiTRaCb6yFXkG/dQW5yZA4Pci97/YDyRJkwf6kWUMcbcsmXS
2KSJZ/iCcXq01PrHRDlgIdN//kSPP3+bWbW3WPzcx0fFHJnmJqzAq8RUehqA0B4j
ttU5lI/gAt+EchhN2rdMwuEorYd3Lh8QrFuga8AqiBRKbSiBOB3XqGfw+23AVao9
9gmuLt1WmUA/9nM3T5zjEYrqk9eqmIxUJ77C3H8tvt5GM/WZyuZdRHh4cyHhvoYm
5B81Ut/QXhOOEkAb5kBahRVCeQ81ymONHjNgznlBEsTyNcgCKqUqyziH8Y5p2hTT
K8n4Vxj/7C4WMM/GlGaG4FDmtazPUHwtEzo0Tg8B4umzpRkN96x298HsNkX/qUHe
8Ul+4kxbXAIDQN+XmI47lz7fn7geIoOIjFvdEtEY+gwruM3Y7bPajjyZi6cDAkgb
/bzC/o/q8S6La08idVkzB9Hahx5ymdgpteZyWlvAANYAj7snHpaIYJXgecEGAaU8
JoMr4mtl1gSHOz3kQKAw65YoQCE96yByPPwHldomeZe+QJkE5VSbEWW2gS9fu7Y+
q8cbKG3PKFhtefzVHLKbKknBPNo8Ju0GXJMSlaEftHOMzVjObD/LLgO2m560Ro9E
yMYYljeIe2N1NQJwcB1u/IXV4qdjH/iGshFIhD+aLmnrkD0UL9TDPnBlQWCe5CcX
xciQ5PP/NpbD54LDRu8hGUUShFRbev3V7xScnNnPwVZOS8Za3vlR/KGmq8y9BZuZ
OV8yTNGxuhXpCW8T2O6l+DPEwM9mv3iuPtKCHAHd/VZ9dausPbKY3qxh595hlbz1
Yn9rcsmK6NihdkUFrPKkbIWWii6oFIJLG6Q4LU2VYVzko/1SMlkfDewhLlMLUf7m
bcyzf8/JuNDLoKTtkS0RfazKsUeBwfUAsQojolLtAi8gnAV3dOdY5Z5Ps/t9DXWL
+qc23bWOH31OlIQR6k6aeST6gR/wI+OYNsr1qga/80BhTDpEqsHD47jmzEpZKjH7
Dhy+s1z6zri0DF2fWhOpu13dqrdBPMYQR7/hfIY5y95uzCaOaZP78AvNFUhGHI0Y
LeP21rkJMq9rtlNPBCczCITffWHk6f+1ev/Uo6fdZ+O+uMTgDkTgCP8EI+FEGiR2
Yom5t/1m+eTtoMm43dgvMLkKc+tqZszCqQUkG0JSSeqTBY+wrCLmKhTmYIZCISvC
354IQ7lgTEOe0kZGQZferSjuZ56J7YSlqi+RAK1xjvP33JQfRRh616lcTQ5T8yQA
rFLsbIuQRNDtpptZv0MGmAKceznaWQMD+ww9fDY3vlbsercOnSCMdA194z2wyQSL
eRfLuUGtrsH6VLpKFQwiJE99yc3m7d3wbLU8BEn+zIiq2E4dMzbrFh1UsMFTGhNY
QXvHZQfVQ4VmP+Z+g5Z+mgqCO4sYwztaHJf5iw7uni2hUovZINoAz8BzyrVNuMx5
5b+W0J8moV/5BPKJcFCKzKA0d7fnWwWWUeVQDaIpNbmBegDoPc6DQOfg+oPM4isL
19yNbXBOHf9Q3cW+MBcGEQivljxd2vsHAsh9abNDdaI7kO1JtIAMYmh/rhzmfdiK
FTGbBrnECJ2ffFCXMB280Qy60OPYE98iR6DwVrr3eJCZzRKGR0ctKaO3yth/AbDL
xY+vsAWXTA0E3jJfc7yg4+f3bRZpehHYNtxqbDUQmCMAe8xJsCxCshv+LDmSGKcB
tUdWTgdaSzF1U0FxM1k9y7N4JBqRPbTN3+qBYYK3V2fTZ/88nrFqpJrcjQE7RVDj
M1Jt5SVVqdjILO1w7QlLNjrzsXqBXct7JtK5CgER+m+83InubDPXbAx0bKaX1hS5
ZU8g/g5Vo4aSDN6G+a99GVGshrXnocO5B2yP7P0noy8O2+epDvpFHgS+u2Ne8KBu
HKwz/g/sUE7kQHqNrwri9KLD+m1cJdVW5h/FRedIJGnL/t4/uI5svnTs6u9CP217
jdlSrWQ41FtSBasPUvaSYzBmiwEEcJD+VcKptmlvDLcrVW1t0xWGe3/a13HWjx05
/Ms6Cy4ERTCZDOGvHea6ptGuoc/wgb4ZKPf79jmO2Zw//ZLZFR4jZpDjB1pGU+Ea
jxX0NeoAE8A/NkiRXoPsu2KSNsHSBLGCoaisfhMn9R6jt/Ba72rihvWkHBzGUhvK
PaS1nZmrPOX26Y3GnONpl7oY1wzpA5CmiD/7Dldzke5yEiEvBtJfNbkrsmHfyJDh
5PB1VZCYqKE2vnVGkw00RmU3bqPBlSYKc8787iT9zP80ShZxSqx87C8DLDHMsetk
OLKh3sHmUomVZtbfIq9E/GX+G3sKRt1Md32meCERF6Iv3obMsdEyVEUI8uslXRzD
zKyZyDiwmOStUaDoLxbqseU0Z1DWpHspE7YrKpY+2N4O0ZlDfWF22RDUrbl/UTlC
pJBnjgjvqeQFRM3jQl3Gp6NT2331ofm6ozjkvk+f3vOvBJDyEZYWiexskXngvTXM
fJph8orb0KbYs9FWVF4yHRBONKQJpRMGh+aTIM2/QhiM0A3/YyQHoA2d9Vi3cHNM
bhVv96JHkOlgSTrw63naRRFVuFYdqeMIIrzIlVUkzlJeucszNJFoGF14a3eN1o4c
W8BG/JaxLBZBT01PWO+ZE4piWplg6isyxtJ3rfOEpobci3o6J7tFJUvzZuC0xtNS
OS7hYriAw+/GmjIs+zp00Uy38lNLdnz1wO4FB2A41ZT0HRCM2IVJo0WkrXLhKvCl
CpXP1iRkloqKGb4N9FNwIA/afH33f9SHKnLZWlixo2/rXvXQ8m+erT0xeBHXWNVv
Myq7yzRXJIqLks0agVrPbTVj3PL2CWVr8pXymXaY5shM5GwBXGMtUum5rkFIvkRu
ZtYrukjd2EEy1OIKIZHLgkd4h1YMMixvNIoy7VHuL4zqlAwTRmcbckSfSAx56jHN
Of+Hh9wCsmzEjPKtuXe4qSm4FU6okpLT5O8M17mmF7qXUGx21xuZg2ngPBSF6D/y
/m3fNt2ZHw+jr/kacdmriMjCGKXFHbhEqtcTvDvfFAwXMDTmRw00+/rRKfSybq/s
OYunp1UghbQpMZKpU0ayJxCgMGtq3iL8JMiWvddLPjcrNZTIxjZ4A9LUJuvFga7b
eaak0coxryoH1R6NtwYv7a9LqpGghY4lPNgmgxbeGB983NHiduAZJGTzjq028OKl
xupOqV0PNHCUeKmGM9sJ4kdnHDI8qhiABDSAWrKpN1jxiyyl+SYhMGTlCJIO70Ah
sXNqxMsF3Y+WBUdWftHPnLcQD4uWQts1vMkQ71ld3hNcMxQbT6V/ahLbScN/mP2V
29537guxqoFGnwLK69KhJVtvaGEceJCdhCJp3c6X1XCEYDH2aYq04XpUpPRlHIpG
q+nHw4RH98B9rxZprIF/GEfoSSBoPu3qLD7ZE7BGPEZeyKGO0pTmVQYgZFE/99nk
za7tsGGXe8p2j4LKkUc9WrVAbUpLkkyEkA+T3xaV/jik6TWN2zU4TUWrs35tCOsZ
aYpBtVSig9zTQi+Cq8nqJvQ3V3fecSQ70WmPOtlvOo5BpC5UZ+ygjBQGpWViaeHF
QuvkCDYNAM3PRUGbxO9xCxDzwRtETLlCp3wZpg8swTY=
`protect end_protected