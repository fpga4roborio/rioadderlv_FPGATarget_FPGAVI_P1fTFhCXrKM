`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
ddtXksX2+yylW5zu6QL2Lhnb2d1sD00763mmSITNX595NcHTEkwn0zB1Dry37fOW
FufOhVzEJp80NC5qZ/+F0Vk7Ik02dIR0elf3clrjeJRK85K4e3Hoo4xn7YbFUIms
l/8VZSb14+JVGURjfswrIyCUotIzlzVYZ6gzoZwDXIi5gQIBf/gI+KxNXPaKV+PQ
Ufys/12rjO6aI/pPlqSm0hCvftmBcnezN2hk1UeXgOIuKZnogjOsf0iJVX2aOOWE
6pD/psybjbnsNB6kH5uFTA5frkzIzkzl5d9+YDm9OyC+k84E83I/7/j+rk4L2dah
QJOvksSIzN867/4Qt8qYTQ==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="MvBXkzurAa5VTw+1JJ70nePUfoQXBvZOku/SMmg4TwQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
oRtzZL4VJ4iwysPsC8SXYCzXS8Fw2gtZTOskLcDV+1B9Nzn1zTyNtlo6lNICRmmK
ZRVu2BmCc2G+fmzynYlNTnSa7C0Cuel6FYpxCBlOuk3OF2tzAmLAuDyOH3Z1Yjzk
a0aHuoCdIRKv7BrZCdALt03JeUmXKPdOmIlkVGFl8yw=
`protect rights_digest_method = "sha256"
`protect end_toolblock="Jn9CQpRhJt4rnzZPRk+dOpzAubz7omckX1MrFd4p81o="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 25616 )
`protect data_block
gD6l00tciPUa6pDNTk/+t0OO0nC/UTtBwLB41d4inuAUA3i/ALrNyoJVcBnAmEQW
ptbcNp5fxEUJjnOxnedyZEuEBxWRieZFQnkRdF269oN5R7TgpawG28ENRN9A8e1Q
YUShbExxEEKiPMrwzxBnh5WSbGYSKQuEiD53ZHcXo0D7NjoIZkVb8E4Ip+INy9Sm
0Pu8l7yz1MkcW0DAYQ6uh+HlqoEhIQUg0jiHq2LCMh0Rcbky65YFE17MsIaEKrsy
kfP26ibHtGlbFfGTRFIeDMrkiRl/1hxJgeNSidSmNznC1Bczzyo6vpH7CVZrVkVi
4lSQVwOT6Uxypdnyvc1REPQ+6PlQLr1d9RNuRkAQUkbP7NVKdhSa2Gn0mU7Kwszs
7sceQ6rU9R0aX6rXGZXMVagp9c7+0yeO/QJdQUgs2DXrtt5C/3IdkXQuGT8TNkrZ
ebByLxaxpEoQOGaMtZLjQ3hZPjuyE98YqX5Ol70Yt6DutNuMDQ0cKMxeG/UcWtWy
fPjKrWNILwIpuMRanbFrrmTL0uUtdY+lDLSv75gvmIYNvtfkr8oxJ64s5+c+nIxt
8hXbumGvL6wb+9jooKRP+dLqLxIRtKQ0qyIYQvu2ziAs4I0GOSuutTfqV7pzVwWP
uT+tLq5P2COtV3WurreZZ2lLAcWmgRGiJGMGGU1nH/GgB5wGkIFGd8cbubo/mCSF
euCZV75IKvhwSGSoBYiI2iitNI8cs/JvjNi6JQXhCm4zbIFly/529NGnESpYjWls
mGfi63bQOC21kGG3bwjkrQhhIjo+ekdu/cVDANdR39ElyQqZcxgkii73Bfv5c/UA
Qe8t8ZEfBsdI2ukieRaTnL+t9q/SGS81u+FGka2f7S2XAfTTN5YWuWryHRfRATLR
BfOjropYEzFanaREmgesgEH4AKa7aR9up1QJSny6f2EQ6VMiw2eCkJOOTbZA3fHC
17yS1IYwXyd5H+qoMhWTOQVUF2v+zeu+oDx+NNf+tXMNwiX22Ch/LIie/M1YcmMm
bAQdKmOEBEbKh1RBws7MVYKehEqkggJQioqDRvvK6zwuVfAsYjJXmbq/aGHUAako
d4uWchKdqeFf0CvpAODeiTBcOtDzOXVAWOYkDZjwKH/BNf10OE1+3C789s4t+Unh
sL35j1c8xPQsODKa0hjU241LiSVN3lHBz8P3xoqv4enbDkij1qYyoVKYLDTuMeGP
0UOf+TDwqfIO82R9ETAP9XOOAqkQcjmr0nTYS3gk//2ormIqRA1D3ysSg3mFsvcg
wCdYnybFNkMW3vW+8fcKB20Q2gty9GT/GYe3Pd+XPYirLc6/fi9RJxCwQLRYh9K3
7m2xo8lLv7Kptisf1aRumfdIOaVIALPKw8Hwe71tIDEhTm3k/k3ilyAoi88CDjmU
yslz/x7Y/vZvz+2STfeof10ZeP4PZJ3xGRiRaTP2k4337D3jz0rjJI3gmiIwKsNp
ygYQ/YjpNOd4DCX/cJK72YdgV8TUeOpDwCHIKDAgzctF3b7w0ngLJCpudLxpjI/d
cyb5FIDIVqS/fCKKznX7mQQVIVAfIGV2LlpRinRQx7vYmilMpdQ5mtwt8Esz+ueC
XlSTDyvFUNbZVNz59LF7HUraajKbpj3WTFKt7lQ8wuxegXWWX3rpFD+YbhKuS63O
Ee/YG0lI9SgT/KiVxzf2IN1buVB2tIgBbyxhICtEHtQUpCI4X9dkhRG9WUKlPGOf
GUPaA2fyNzo1da+qtzmmkZLuYvfZRK4LtZvPvtODCAwyJELArjktinp1QPYrdYcL
jNlwPjc8uY2OqCMefu2+/G/qu2/NU8A5EJRbM0iyiyZ2TKLI7sNRoH05ZzFZ0Q0t
fpLE2le/sNklsdzJ/IQAz5b7t3Bipw8ZYfrSDLrn6JcfmNJ+DRQQcAJwXWLUi2KE
7gyDWKfEhyYRhv+XmS9d81huUjsMvjDxADH9DkluXbTIm2o+wWiAv+3VwRrWnC9U
4qxmxvb6OkhUgUe6hGXBXdrOOJ8f4g4RRbCWxRp7QSi5U+qZnBr5KkgI926lWJK9
HMEZSkF/tcoGZZyK+3lZcRrwxs/aO4osgp3IJtuacdvWwjX1n/AxWd3Nd+vfRpYa
6VUatdfu2js6ofQ1O67gEhrXYzvwS83QnzjDPGZJ4NZP7RWQQ9KrwIaThIFYbu02
QqpsCvtwTgJ1Wd5pls8T3bZDwikH9v33nXCxf7SarOEUhLBufs7PacRZjgDIrAhl
cw9d2Xwmxji3GzvpmEcLdAWM3rCKf/f5f6ARuNHZ7kLZazkCMdzrNXEbT0NWDb/b
2IKwiAStypgdXbEVN8ADjDBDLuON/4RFuo/GskXJP4DA+D5WIBPaXxT7OmLlLhZp
lCoigCRks2BG1hlnxpDzoHveA6+FsQBngNCsdVaxT+Qtb/ZjZQHHjHIYUBBnPaUm
sOzbnQ9mPqcV8nw+ZJgeyxz0spb5obVteec63lAJnebBh8i6W8Rg0tWCx72C3AmI
QGi7lBz09mwuSgjj/1q7mXVQQYCWhCXp/RhOD9kQ6Brglc+0UvvuynqF29Z9MMTr
k/rZXmRl57Y2CwQ05W2R2fQGcJdyh2Qes0M3mVbFCec+4M1pzcfCR/jdTyPhE5eZ
ozYHx3SViOSuxRNi3OSvlHNg9aS9cxVX10PnxMH2jeserCoKUOEf0XDrRzDRUoxW
+x+KtTvcN8rf2u47rDvS92Rk4IU2ZlmEKkS2K7CShDrH7H+wom81FsNL3QLcLWr/
ml3G/udHSdw9O3UbKUHHdN6QvGoIwXGIcHZLX0lpfUt1soMxmBWLnGHP06sLrbR+
5NYBOwdB41gDenRWGzkCZQzo6IbCVIEURFgEEZC7RsoPfm6mJYvGF3BpNNztpWao
iOQXPnPjMshOOcJpm1SAfOREkzJkhIXMEU6i8H+khAaa/mSy9Sp9GICpaqAMw7mP
eALDvYkmY9Z134dqjJxo3I/T4d57kH78tLjnSYDNdtQzH++IZTS7ZVH6chLpCpUX
XlqXCPddcSeDGVnGy6ejeDynIebJlpF7pjBvckAumlgK9wGGY1iQdeUm9Q1bwEO+
k7eouh0HeMw+bEhUIRCody97zRffNuoLZJi94hRTPxbbhjepYWqcCasEXAzaapQM
w8amwuhmrYQAUfKNNYr9KH44XgsHhuJzpFtBUQU/iF/WMsE5nZKTXA0Xoq/5gwWZ
qNkiSsOIOL8bTYH861sMr+RqL6UPzo5m7/PtCYlFytvm1eWpp+UhpV6RkZwgUhE+
gOp36tfiHSOmWs/fUpbDNjOp58z0Unr7fvqpZKxol+uy3SfcHrzanGpuuZ/whbnZ
8ARHAaR0AYk4hQgvzEGLswn+J+pB87ltyDWAqM/DyvFT+a7kFECcefR5lsqHSBpD
vn0mLTwLUxQ0tgLCZXCWl39GPR+ikqc9/agP967K1G63IFajRfm+QIiDD2ZSj5nR
2W+2BmjoJdA2G7BDf2kh/6KZknMyl6QzwwAEXimuNjUNLbeoHY6BdmTzGaLrWT/H
owRLlIab+F5/8iI4VCebEcIAexuhbFZ37Czi+7RkUQchP+yDHRdfXFaYJspSR5do
q0Bh+5V4BLSd1XXZOTsNv9oafxa8E+8AuVaE6NhRDVyS4sVo3ZSJQk/PkHTxNnmj
uQRSHTslb3QINdgofbB5+TwrU3thuN04/4ti+LBgj82c1GLFTArbPrKmBzPjbb31
vlo54Ra0C6ytIUuew/kr9H2yidK0nS9Y68SXPijQ6avbUJzVENAjzUaW5Gioexyq
feKH4D2Xq8E2pqCSNMeHtHJRFDmrvrh1m27pzczavOvfNUy2JNFWJ6NJBFESiT/9
xXh7VeiqTgxX4cup2aFrE6lUgnWI+n9LuGxpQdVgKdaSVi493OEwjvdgapyc20ra
DI3cIkW0af0IUzkVZgb8wCr0JSVx2Z05LkM5+6GHgAF4Djy4ps/BsxVI8g8doMGb
nSz8xUNrAmm+wLTtf2EtKux32JMivfoyB8vrvmuGAdgFa6uJkNtE9Cw5frLWIrq8
MQWgOm8clTYCFp+DRQxDyJFV7zKFSsedIG7qF2M7q/vWUtR9/ywYHjsJ0Y5gufdN
nA4m2MMR8L6vUojgenJAjhYugkuszsgaUBb1ICs9qta/q84stM98StdZ737nUhpZ
LKc8ESxTB9hlXe12PZ76w3+08/hCxsVyfrtSYpU82qS02lO+ZKRCVETdHPbMUZvq
ux4bwTdiyrnCSA5vEPSkRaU98yLiNR0jDdf53kXoq67bfAnFqGUYMK2s37qjVPQk
Cm2v1BLkJiCu7O1u2NSntCsdXwlw7dOCRa1NXHk2lx7CWtYuAWOyMwvu7bvL5dgp
GXUJCWgHKZ39b5cNngNgfIooi0Kt05BxUrIzoEZelF4KQhECZm9+mISuXz1zQKMl
ite1U04EpnoBoaAulSgBpD/086hDU3RKl2scPugiPTWYKIEkzO4Nn6VeLMwcAuZ6
1dkSWnf0i89XWWxVxc8+97wVjwecLsX/FAf3jTGseSgSNq5u0jbIwbVwXpLGNdZG
tl9608aY8kV9lJEmRtXCyK/9WtWrd07s07YhhsQufFUe50XvbW7zcTnsfH7r4cvG
OTMtCxh0xMBBImCFU2Dngu7PDDZXIil56IWF59wtuIPaRE5VUDM5+k9N37DAUMqb
StH5M5S7Ypy2ZnE60PCmm6dTl4Jvp4hqCGq2KDfJYcmMJT37OPY19BqBy9Bcbw0L
v2aZ6Zp7h4cU6eQR5q8Yt8cYtpcz9ixjdvlHg0WOQSfQRiRRmu5FaZOhn7KYsZeK
St5tWT1egjq1BgHEAVS1FV2Z+snCJKOrVIfsmK2NQ1ZiVsz6nDgOav3UOFLYLbrh
u4eEoaHgTGOtgFgzUEPaR5a0NYpiCmpsLSoYegMV5LluN3c55zrHRdFun3qv9FgP
aCyiSNeZ5H/cq0ChzS+wM3h43YfJc9ktESLtSk5GOFjoeZ+Av+zR9a61jBG33Qqs
HILjCs/5VoD0p6Ro653Gacx5isTUi6FbrwbtPrNqao3kE6WhRYezYOEqsV2F5wM/
0RozpRiQ+AzqLGr54C0oBgFXpdcCC+xRmtIgtX8KB4lm0Zr4zvtki/HHLJ0wl7M1
UOfishCXgIu5ehzti8e9r8a5/lU3Flu1aFc6fur+yO2VMzEpQs2UfqIDMhI1H37o
3OghpBGyvraS2mep53JD9CqHSgMWzlAq+GgIdWV8IHzMHkFqdlvrCBzdEIb/3/MU
DJF/6jV8OhnLSN5rRwoF4Juhi6nfXVW57/KiS26Jhvd/KNk00Ptiz6dTwAQUMQdw
YHvC70eGtl1WF2pOf4M+ZDmvljjF2246Vpca9engsqnuGbaIB5QOrMxvksJcFAYD
Co8x5Abj/F1XIvY8Fvia1cIQ/QrN4Gk7FyyrXEe2s4FlkpB6HwUrKLcCbgxaR395
jLkjGPXnuwgBLZ6A6pO5625rCtiuBizFhI1AnHh1UZod725wyaBKiWehQW1cfH4g
VUfdwf7+HDJER7N4Hv+ykNfi0VaPd/Ipz5MWGB9EriwpSiBEstjFNLwjtI0N8sQG
nwZuCP9yoZtMOcCietTN2vMBzkQNQNDGfnFSE4r4wrQ/kyAFQ6a2QbXEfkxgNN/G
nSWC9OekyN6SCjr9r3WjjNheOpFoaZGRBCIRm2e7iq6BeLnhQWwJLNlggS418tJ4
plGBWpCTsdbgXCcTeocbSCLDNJqU8NYJasXsXNQCVTMElF/E6JMddPjYcLGDYUKf
H8iTE79RixuuV9vrLXwr3eUq5apQi6QznW8bVg2zPO50KOE7oq/6IobnveB+T554
UaoUwKpRG7zOnwWe/yuYIzeKFvqko8+fMER4HHl1gcAIL+yuj4jNMGeiFJmdp3er
N5jDpfd+47KMI98IQ1VGXDQqgJxKS7CosOu0Ws6SCuAlHlIpZ894DYdqwP6JtMKh
WxawzI9RXMIgsKq4KouVWHkFYLX2MSDb3E5XdIlu45wkY5Ac8yu3LrpldYBVGJgn
tvEPHUBtskr2v8GWL84guyQjmLbogSnjCFKTAVb1N3vtIeAjVPQHbE3EGxdMOszJ
hRRB94FbQFwCr47F8wD02hbpCdolQeR29IRIL7hIw8DvtkN0zwV7uZxrYDC0W8/v
5UuMadFQDADyA76Kg4L2eC+RhHnTUkj61XkmOqZjLde1hAr/x95/Th8voN/vJ+y4
nmmReza9/hmr4BZQ/6CrXUdhqRf6Jcmrlsgav41A1tV7W4LHGgmh1qIQn3Zkzhig
faoJx9YconOxYe4kTP6Beqg2NZhG1R1UZtV59WpGrXAMPDAkVBm7tU1lijmieEWt
vgvbysqXj6qbJAEAkYz1yISe6b3rX17kI24VAit5Hlq0fUNYmk0+BiKbbclbnyrO
DpDhmFhjHrQyRH8R82WSNBRtBtJLQg/LxU0aHV0vXOTIZPT5AoC6tRLfbQSj4oV3
cgWVlrR08VHZ0dCdrfrZShwezkzrr3XjWTam849VrIcektP1lligLeWY3ueEayCS
KlsaPQoZ1oKGrqOv9WfTtA4ZzhTNqY6Ov4NV4Y4kH0MR0rs8rX4Cn4HZQPMep08b
KbhRSdV1JCq6A7XDLSWAkP5nxYlGrB5lWb4VFQWWnbGLSklg45N7lCv+ZmPMVc83
B9cRujIXOpf145zku5BLHeHHZsrGwIrRbLhfLiiHfEMU8yxeYnIpMlPSAwzMjWZT
uKAzNixBD1kR2WFMZrIBTHEOxePoPqsJoFriELRLtAAbyg/KBjhdu2MTbPs4nYca
y0BgwTJLYpLhCCJwUTZUoGOh62M/m1Pszgs6QnRQND76qtEPLamQJdFO/RccAXxf
WFXJcnJ+mmyP7W8hOstXC0cWZo4wbagoTAxew5gE7oRwl5HEsAmDgJ9oMTWkhgsF
IRmLrBo5KQAQA1qUQIrROvAgFk/p/qvPZoPezXUhugVgw9prmCYOC7RHxMnapZaO
o1mkblcsEb+uAi0yHzf7Ewi3fk/K47kqFgc3NSed2h9j/+wHf8sEQ/6kcyvTN/DO
OTm0p4rfQjonCD+sdsFmGcwnWGdocC7hY37vWxnhmCbSAPUFw3i+nlhoCLO/Y6ez
kHQZ2IIRwm4CBknxKAwE1Uv85sfuf75bK0+j2nI2jNev863jX9FjkPp5ZCltRo6+
9YcTO76KdbPQ8u3CVV/37b9sO6h54IymvT3NSSqCXeHFATSpn7x1E+RDgeqIIUtX
Sdm3OjJsQjtidsUkj/pb/312LuhOT+hzW8+UI1+JdO1o822l+g1ZiWUoThFsDfjB
imgTgZXkjbpzse5Nxvpd1Lqzb8H2KAuYEMlZFAUsFcbxrkH2eKLbks867fW1pnW2
DvhCNJAyW/D0EWBozKM/R9uUDU9CrXu/w3plgqpNbCgrvxPcXuhhHSjmcrTsBBq6
9v8hqWgrEzMSwzg0qsnFSk6DPOf9gSE/Lf2S3XsDJd9JSUh7jPMYvJLUOkqQ1Qxh
29H/KCGCNLOIvGGWK5/bJylGpwzpKW8pBYjxO6xVtLKOX73GpiBLxqVVlqtFS8+Q
eG99emvkMh7SQcFD+Xjgwla/TPYNpXnczrqbjiVG5Fnb3E/QKL+PgvmUF36KJTV0
GKoXjZXqjeq1m1jpLiXtoKINe+r1VEkirx4XhD04MgZzhxTvcT13vmB7dW8iJc7n
hqVrvdvc1aTHPTP1l2H3gNEgBHapD7eJZcaBo02GxuNBLbEwR+dyrr6N/zSDTG/2
nTE9y7zdtR3FhuAZ6kFNn8O5WU5qu5bqLz7yhFEaQTTYZueTho1FYAgb5G5Igv/x
OWkZFyunYg335k3cj0UbqTVfEKUi1NOfmdaPzowGqxOU+sknnFL8TI72sXTwEs0i
Mmx87JJNpW7ej7zPnJnvFw2DJFvScjg/J4alQqdUei1R34uBPgxiNDxSZN1oPsrp
jhJl7/rpddzxwHpzdzeUMFeNhSPrtbHy8TQgejigyDg9rcv4xkwhQL/YvBq4QkB5
L4NqIyuj2zvZBkXDaRRwvW5lDfUKVyTQ2Ra16pkLF3NTTkVv9NFvJaZS67LJTfXU
zwVQogxWHAvsFwm5/DMNjcnkCsEMgGN1wyOG+dXVomFsKA1JxmLYGaH5cEpgwtpY
Rjbiu05h61aSYYdADiF9I5woykJ0gxuKD26HvklDpWLtgiDgvKHbeN1plounXI4z
3jXpS+mLiUFpO0ZbXZPt13+CgB6m6plvUbt//KnaMZaTxJugkPtX/xUO+W11msR+
oBRZcePnIxcjS3Qcwt6hfes7jj2CwBnsZGM+0/HKai9/Ac7+m+PE40G1wox0pMmp
jMNec3crc8yQJchfJekZk9pNApip6tDttyQ5HidH0moyn8AatOH+aq1KdCZN+Nz2
aKNAQXf6EwiJQP+sx+XJgp6bpQsg/yXulZTvnOg+6Xm05KLXZbC/lZFTPfAz+uuq
bBRyMzoGDeBAqC4VotHxXxDO+YusflbYkjniZLmJ1B5Q1MkCuJCeyPd2alirYzyR
TvxeqSmMIL1pgzaTcvR7TZXbw6AdAdLjCCXuCz29wfhgkOoN9pylHejZcQrgVp3s
NXth+q85fZ9JSuy6FzUut4Pt//lV2PYSoJt640cNu4/s78foqMDmq9BU7Gz0Ho8h
gDZFLjgpuZBuawjbZ0d0olHiYTGI+xmEw/TFkdQqcGRUeIrYA8d4lhJviZ8OqJyF
P2thn4QI4E8o3m+rCPo1jt24Z71UIkKq9B84NQ8a9wgnL4Vizim4gOusmLoSFGiw
HTfQL+4UXf13gNxOmqxHkHrSPZqrFQrntFOev1pTzlzcH5r+TyACBpNyEka/FVeS
ImJ9k2Vx3Oo+XfdBhCefUN2Cv8J8EGHRtyIzv8pVP8X/1aT642A06uXKQfC6Agd/
YUFtAP7fv1ljE/7UyhxMX6ujBRx9kft9fr+MNZ2o8nIHTb9KiD/rcIa2MvxYuaCH
yHOvJC5oCBKtmJBXa66gpJy749HOB5JZg8+WrnBcWCZ6k1zF0xrmQlxBWWkzgrue
qR4KtC0FW8YMNOV+5qpjwcrbcjbIrpWzbPbxeHKKHzHTT1PdAua4DiOCFsuv6FqV
OvPfR7wOpllmGQ25ynosZSf/ps94/RBajbrdY8Hp55wPQZPAzvYFYtd3KHl+7o9G
M28ABX3u2QhzV0Az33Ps6iJWgC1sNFwWxI2lZYs5Dhth2XDRp0olQukyv7CxkFtU
VVQm9F4CZm7t2QbK3YflmBxJKwnPHFDLGzy6LGZoTBufTTbiHLOP2OA3I0bywfE1
HhuDp3Hfy8efKaFBSF7lEFcCW/HL+lrlq2ZP4FKj5xEC/g7iY2OESGt7131DUuJ6
JuhzM03osWUyqn+SR2WEYOG8kL05dP3yPGZeAHxs5RES9NeKreut8k/fWGZMQTCZ
mSFNMkWoHjkVqsVNvErKx2nfnfQoZaKhoxjWJoQa3L6MA3dbi68DMLujpswsR0iF
GR8/eeLkC1BBOg06XOmHHVpihVfsGTIYF6Nq+PWcyAZjNnfalPzKaq8y1/36KKdg
HObVCbG6/kBrxS4Ek6nIObI6LggzFqzV3c9IDktjCz86VOB5lFK03LmUEdAx9clc
8UUYjWaIDRmntSMPg83n6CpuOOiwrE5WWqWBnpX5mJUDI8pVmL9id+FdieJDG5Io
eX8hjVv4fxgWf7MrLzG43evSKIuVN6FbpQHJTz82kQ+1VvdK0fwiGCTplMFYbAAh
s+i9EEIVl49JmLjJkM/FMUc3Ef3xHAFSPEFJFIE9EyHXlBgcRufYFTQ5VXEFc9Ok
5o9yUc3O6vWh4SI8PyqF1Kb1Wx8/EFjUZfJO+ftI3BxztAan/APKED4FR2Zb4PpK
FtSVIFtmpB7lMGUpMReJkOih8CLR4qSLOycMfu3p00PBE5g75x7p2UQxt+NyWvI6
idnZCGGVjH3T9HjSYgXPXqs1uFZkZ6xOtvFCGk5AVOr0hGO0xkz5V5nVKDIDTTeK
vCvAQxDvAHNP0MA/ik4QMKfQj3rsBFcxlQpXLZ7CsLE4RF8Dk/pG+JyUB5S07pAh
1eF56gexFjhk6cHy5Nrcl6fmVUEOi/Otiq0o7j/RGa1HFuiPVKKCafeM2nZ64UY+
um/XJD6R9eqxTvx7FGmddCzK5YBzV3QJ0qF+IVK/udN5sEfrcAXaLMGXwl1k1ody
ZWAiQgYYZPIVKG2Qziv+Q/m173VMRTwUGd0exuFFcEDv62cq7iTHU7bBfYXasHHw
A63FLCHKGHl9vMdQBKV9qp0cCXhip/cU1eEuJFLF9mlPxlmLDRUdG3woQLPi8SUG
AhArB07BlNbIz5TBh8EMvWTC2K3hHwLrI7VNEc+98u+bFZUlgpgbW60m90sxXuUd
pGSeWROiGcglJ2OPkczAq6oCK+32rjnU3crgro7nlWSR3/dzN91TvOwBbCkoTzNR
mVbQrmbeb4CDNw0mycMI6/oo0jnzXKLu8twfKoPQcpP9dnt2qHMZxwcHp9D5LuEx
Ui80Py9mQNLGlaThmBoUXS3+ZLgtNKkeFhJpTbnVJ/fmxz/FVthogUPaFnLNvd6G
22teeZ/q83VYv0RJJ2z5eDTsMJ6GlefK/KOUyAEhWXxO++wjylIpRd501ssmBUHT
sk4o7N5dpOikkoCCXLCvjmDj1iV5aeOXFU+GUhnrEjOI86OHiZ01SBv0yMemAs4w
WTcg65dJ+odB5ebh2pIyOrU2pjyDnVjHe6+AI3BgpeGvDjiV6VrfAXp63PN7GmlN
9/CRfxVNLgDp1kJjOleHy1nVdSXTXf4dCtN5fsq0dwji9v9D2sEbHwliOsMNe72g
YoH5/Xz6sGkPMAqZjuHcyNVGdFeczlRYWNeVrVF0P3P3vMwiPUbi3bPoBTM98XcY
ZiuoC6TLRNtALvX/HgHK/bISCyw0JAAQmfei+3ocl4PyG8x/gJyaWnr5MoFyHlHj
M4TIHXYIxU1CFx0LoWQ4vpassoAqTPoaAl2PTSk67hH8Q4DkWT5MRSLzUb+gS5q6
2hMZ4FHOMFStc0Y/MsG47unR2QBCmbNUYGXtmRtkLP7J0JL4Lq+CH3E2Z9a10LIX
JaYHzX6xiUHRnTG0Yj+BDW0dTCITp0GB6ZtuvoagPki7qYM4P+eux0cRjGq53J/O
CBNybjaLepFGoNOHByEkDFxLBMIKK4npkA+Kxv3ZdN4/JAizTYC2oG2myzgMBOFt
haHW7GD5OyTqLuPUyZX5yRJ5lKwdVZFp1OzVNHzKhSrWtDIg64RUMeM6xuIQBHag
23StGU1DxNWJI+LlH++OnbUYLV8TJFdY7AoEELLfar5QYWHc6d3rb4KMzudOv9yK
r+m5hWYRiYAAlRajL+VzGIc8PiWYxG+MKVlD0h1X1t2SSDX9ewUTNAwiCkoDHq2h
0bxRs377giViTiKxBzs5ZfTadHvZCt8KhgL0s/fi7WOyD6Sf/BbNFBufK5gULqSr
ExBXxpag7CvqHVYtPLMdmWcNZMGDX0dESgeot+ipa0waFfh+EpsP3OvVpL0hmhu8
Qc5NsjeXTcO/C9PAzkLQUjme0YJh5Vq5lty0goQYLZ2jcOlXxcsBAhfHolIaKzPh
VeqCr8VHOFx4bGOfLcneCJEReaLX3xCApJrFZj44JUMRmQt/4pnVw+tl9xYlg3Np
1CnesOW7lLEDeApKbIUuXYDn3kKzQtyB37xM6tAE04X2zFL/KetgUmbDD6SrEGHT
Nx/AMCrnaHqYAjitFp7RZ8tP1At4IdwFARfU46w4SMZ4t8HZeeglARoBODQj31m+
aSQ0kDoZCa1Q5WJ7ZfuN/1Xy4EKO+iUub5HNwhQ4WrkqA8wTDos+yvOQQsYB3WRn
bJ0aZ4RbdMVSdKaO+Kkfw4DcrdC72EQ63/eaaml4eVRzLflpQHzp4i6AKAfokwKw
8SPzZzi3cKhlYm4NVg+0yFs2Butp0W8P1LtFekQMXAKhbpIn3tUe4Yc2DeRjOCkQ
BTiowWO7ujTPi22Z8uUXX/V3j8S/h2/C6Ur52AzfMlWmT7u1Nk+Mr+YHbd6pl3YL
RM8C35CZi+Z1T/GXiVrzkDxNYDyBP/Rml8oVagZICYRYsKP5oc0O9gqwTY/iG3vY
kn8ZsxkE7A6mcQVjdmaKInTI/YFBRfj90SVgRQ5xR/CmZuuBrEQmt5/inmNSg/sm
q5XRcYorgcLwZcWoEfhB1ddRd8SRVk6UJxLBuye8hyAOqfY2IgbfOyFeW32mT9Ht
tWOAm/lS+tJzxpuztVkdoyvLMG7CZ7pyhkW0IdGJzjGbmSL0dYhsH7GMX6Vvp25r
/PkgOqOmrvKoIaH/1cJQIiEpieDfls6qrBnEqGxrYEGeEC3l8HXsguWV8CdVTnVO
X1ETnnUMC4N1VsrBI6xJTpG4pvGB9rbLBHTBA/aGFKoQFxUy6X3Hqhq/2FoT/y9G
H2QFw/w2CaZn34Lg4d0GhNQb9PeD7CiEFECA+jHKIe/cofPc6wX2Ux1sEm3PxEfw
dIOtaj+zdbgzjEO+Dn4L15a6sHmHRsProLRYo4+k7pGDVhjamP7iXk1ylKctK4jB
1s709Q14OGiBks5d9pOebx1xeM4IgwZySsciVWnypZnm51Aj1Jbtky70IT7KxjyM
qj45JEzesmzBYvr1E51WLIcyMNfZNKh46TJZMoqCnuibpO3PpTRhiQBhgEM199Re
jf6i92zgbgXJyjKx2qgpFG0GflCTh24jek7bJX16gBKkJcQVN+MsAKUkxPFhHkzF
7VoMPBW2PV9voFvRso1cPStdq+dsVtHAJn9vpM+3ye1NpoY7ULdGHpmd0OGXO8MW
bAtaAn4WxhWmVyz8wfPiuMfU+YBnyy27DVBtoGSFgzQIL2mRR8pSz0K+MbaJRmPb
rHZmYViqnuPj3mNjJsQMVpP9CAVOxLNdxErWdNJJmMsmRDyX2Ty4jvQYUAkZWnHt
enZOk8/qMZWL/F7NdqCOffzplO/OOhlQ01fjTmh9Ir26F8JLrCJs/yngdH1znstc
JJReFjqfPE/Y0+M9/mg7LEo+XJ+FN8gGh+JorwUj7fVY7NSEjNct6XPXJyHu0jG4
OZRx+AqkLFF/jyRTNzyj+8OHdUau8ogGsUABhNb65xuQ/tN4S9UtDLGn9pEgmmjO
PpQBLk42gRFr/AS/Lns+C5yDY3I6e4txOWbuQYM6YEQnPbbD3j1mh39oEdxoPnjC
67+B/md1MtV4WX22BYYFcMtD4qDzfeeGr/dWe0GrSsoC57HZd0D7Ky602G1M/oiu
XtbhnjYQMX7gNSAumDG2qNv8kqPudN0sE5KyOO6xk8iQSK3MeZRalegQA24DcEgn
68M0jeCo+G4AjfJ9axP7gkCxie1s5aYplnSTat3yrORV+ThuZSIsghDm+QJgJ44M
BIJLgdhVls/InBnl3R7sno66Jh6L7sRLSFIKa8bzyJ19BJa/0YPpX58WeXHcl9Jk
811ffyNIr71SJSWowy2LJA3VYWjdqCmkjjvuQG3wYdkGcDs3UpChuJoP/Q2EpHJq
Buwr8tKmQHXmUERYb+8ja23eVHVMzTSSm8uPUk3b7RwqNMWt+Zii05gH9LzFKc0G
FJw2dnQ3dBtVZ5joF1mkSZV6Qqwh5iQ2VP9dfxgtY1sitslHCs+JGw+GSM3X5XrS
+P7w2oMhNJ1uV4+13+WS4ZEqEUhhvL85VHB7tnfn6LOplDtjrLZ/h22L+P08KnJS
DnezULKQxl/K6ioAWbJl2HfyKQEyfOS40RrfsGCQflC7RMhBrflcP6otPu9+3KsU
/X8s63dflEw2GUy/7aiHwkP4d5q/uOAY0agFI3kKbhz0nb5RR+/Q8OFhkmwk8snG
K8Fv0fkhZ+H0yUPDoVCyKTSrZQeee9a8OxGZyobUfXWPlRe9UP4SkhnSbC/y7P7r
awRZi7NwkkLyt+RYh0IJtCHWZUmEwNQlcVyM0WatkmjuhdSofj2iyTTMNnKHAlXM
mvOJhye2bA7KWYmRAq2LumolnxPqcDWQFlirzRTFj+fAtAPwS6uIPHhsaK9K3PAQ
wURTbSzE2etem/9iKraQgziy1tt99zXCzpOBDQjkzFm5hs0qbb4wnsgPPci4VIqS
ZPLI1irl8DP3gnweXnD4GHVPc+Q9/Fxx5KKIZF6YAskicN1twVReDZLJE5v8Dn/Y
FotD0qqcc5pK2JeZ1TrllNzSvZlB0dy4GwNEJEIlVJfgxLKxq0PYSv/uZG9+Vcuy
WyF27+sUGotkAjz1JpvJhOZ8lC+L6WYygbcJd7K/QYQ7rUuxBEdZ4v8lHfyxJWtZ
nuuuQDm26BIgaHIHAoBzKZzchqX4ROSGXVqJEwFH0X/J4PDOXoxrMKGSKB3Fu0FS
gvmsYKNwDSps7Hmqxtb7NUOdcaSTG296eNdU/u6MEaod1I3KcwOXgPB2XmdTvgoV
Zk9c6EvhJYgBDaYkcyuN07SliiPo9Flq9DMozGrB6a45zlMdswfxYIZtUiceC+hx
i46wDtIsrCUDqB+k2HM06C+5UiO8M53A3qjvzMx9Xf452sAw6DFHu2Ot4Ge/dv5M
+f319RVSp5NdHLq1PTuwR2EvFBMT+I4umdLWg28wyPdKf11uU9cOdet1CNtltXAn
/jfmXmWM7DjQ1cg57N4D4kGps6UL7D7n/1YNRj6Dq5XUM/HhrJe+wXDX+/SGQsMh
BpfsB9r8vF2nvCJm312H292J3t+K59WahIL+0qhXcuFRd78OmSrSAvPFygiPmtEJ
lccv1fcnkAovK8duVvpNkeVPEHD8By/Dyk6fuqh/zhRyuxOqndg1uhEWnncj5KFO
4BzvlJW7q9SJ2XscWWyBPjrPijWJH5S4ZTd4YRNkHE2MVW9+6GP7+I0qToJ9ESkR
lZrd2YyXS5hU7GmMQ1RMXJF1ZqNTBFIlcf5ZuuKiKUIRMbXzmUMIeGyUn8gl159W
Yu6S7pnBj3SCH+0JMBMWu4nO8BzWNov2zDwETWme6JzBTaSHmW6tH1qmKFTqZhW4
prc/nut/FbgNjYognMSPBJqOAqwEINldcSIV4hJU6jlRTl7eT09O0ipp2akR8ryy
ACL6yvKrjpRWMASqGszsaAens6Xq86z1y7zDAEWW1dkQdXaindH7dGXOhuam7hMW
tHBzvGyv2NFT0+QvVL1Nf46DC29fk91OHDmlNgKvKOlZ2v+BAO8daNbNmy7tHaIV
crUTJv/mJok013nyoiOZolT6i0KY+36ZDkJ+KxbVuYcujYNHU/07095xHWh7XOT6
/lGWFvh53Ic4rt0Ur1sk/VTnStLLbqjtn8bNILY843jfwLAWRjuZht746LqwAGjC
sbycI28OJYCoePXNdThB5UugC9Yv2318DMr/a37CQeJQQT0C5HwBsLyMvYvtht33
A6mcHO+AR/hUoPrtxyghLwIVe5RTnuA3cAyIf5pssZozc8puMlgR0pqvZZSutSN2
vylXnVrVFYZaHDWL6qfyyUqKf4Xj3hzy28eg039jKp7HDgY7ICTgM8w/8PA9juwN
SGiPH7ZL/KfP7JVzpWi9wjLxxjaCc0Onh10fzoxZgeMW3N/baLAiveKZChx1Vdpj
BlPBtfWunrxGOYPWcT4rQEs6dLGfDAMWW6XS7+fVSF32fY16Wi2Rba+WTaGqDqHE
iV4IGPjFTEXn/DMbdFdwRvqgVq3u5QpxyHPJ2wnpa1WFjq+euqHTVdRlf3Za0dGg
3vL1RFxfRU1SX9nosOI9S01WZGxMjoLmqbrb1Tvz+ZUGZ/uwzSbEiB2kSCB9iiKv
2rADGcEmSCOzoigpFFIQ+d9SPai7NkVebGhkuxMtrNLhMRW9zskyYq99/0aD+wOr
9GEVzuDeaYzNK72uMBsWrtKMSaMhvKsLExPRNecqZMylqjh/mYT3PdURop/8mP3e
F9exfqvSEqMrRojWmYCNQonIE2yCYuzJSskTcMB5xIlRA54ossErfRw8Mc8DIBB5
gx6/j/ou18rxrf7jqs7X9+ifhPWeeC1NnXcQKfPYy8XINch5wPRC7ZRnDWKYg8Wk
+F2qZC1X/waoiqi6erVadUe2prssv7ew1dzsedNBaZ1p0g/Vgxwhohvn4iG0bkgM
YWH34iPNNRKJW61av8FJ1apHBMQVZKm9UBiks+IfYRqfs4BaCUylUpYqj0yz8SLp
oec3kWhgh0iN5HndU5puZfZnS8me5d98rRflu3VnUmcMDdJMrSO6JmeyomzpsaS4
dO6KMRFc1EWRqr9iHa6AkmiZ8hE492F8AsaHAAOxdNIw6MSB/q9DNsTFwULWrt/P
+UNy7Xt49ZG7LnEncY4BurWKef1Aes+Ge2BjvtY4bmEXY+ocROUYORgRX/Clu1BR
zzgo4qdq8sokr9wOJmeKaExcB0F7ZHczslVST1hMdsFiE6YjzeZ+Xuhx+DGO56R/
45UOBkoaS76EVgbSGJtHTp1qpEFASElII+4aMUAFcGzRwcJG4naAmM9zcfn7ngDI
LE4swvT2M45b/QJriSdCwpd9fVV1DfteCX1WpfZ9E3iHJa7x0CSWmFVu2xcKq5Jm
Vufh0hwqhAPN3lRMmjdlrslBoNS44Tkul2hCLjuhmJVAcE8zJRPAp5VaSYX98fla
/EmWcWywcALz0bB0rvdpsUB8dFwTbN2RVq45eyPJfW1wf954t2TCPZFnI4frwDqg
UAj4gr0PVYk/x95aK+HXA15TInx+feS7A1qMV3hmHlN/0vbp5JarEYg9pdZfEA8/
26t4L/eG9e69NsEIliMu0tgMkm8bX0C0gYuxraeN7iOTRONq6t9NVPI7uiHwDZBN
kbcKiYxLLBZwttGDWQQr88n/0SE2DeyCN6fq5YxWjlKbUp/YHohvauordE1H4xEh
f9rJa/oi4TxsSEVko5D7t9XUlW9lb7rUpj6QdXgXyw6F79C10pwAWZ2jSGmUrKXz
KtAZvQrtRZ5t8yIK8hUHmW/7ROUEE7HEqnLEPlUFE7iZjXCqvSOVbfYTYvbJN/uN
G4Y0tAM2UtxxdSDGgs0R/QZhNHkfImZD1MvsQ7IbtkIdG4RdDSpAJ1bXJYKfa8+n
lCNk3EsoAQY94fn3mo4tQ8VFzwjAiUFszBspdWM4wE1S+Ha241GbwKa2I3EsXbG1
vLCa+FfBTngqgH0s7ZkXgVgepn4LpPZevkYJz5D9IX9W/xf+D4hUif3VbsfJLkws
ySVL1MzbK2qVGKeGJssfxYFbmaC0N/g02qRAJ7cf1brHq0u6udU5qTkk05PPZTcQ
soLMF8jo/9UinXrsU7PsGCsAm+pp+Ic1GTbi9jGdjDGfErf1N4knVxIWLkVKWb4N
1UyoGBcMOnVy7Pkh7h9e5pYLM3qOBjOl6e8wfhyMxjpTry+YR41LvoubLQR+Jage
i1nMOrDn4rSAR2Ty24jBtH97jLLdtIVPagZP3hO5T1IcwAkELqrP+7ddul3R0vVW
nsFKTP89o0FaBl2hZU3LTVZLXJ4GWqpaJjw3mkabOONpVMcdphJY42eFFSIojLHf
pQsMIgHScaBraSkGKttodN2hGY4LsC4GXOulB440lTOvYQyOzrgWd8Dp3iL1ZNa1
tMfZnQiuOLj0Z375IkE0M+OLAF1z+unAGIP3L3HeGCz46Xoc7gLaD8X03YdSClM1
Zkk5nrrn21qfSc5DCXrWoyuMEIOHrDqXVSoPIHDhyUYyCNpjlD0V1PHMC139Dh70
n5Gw8V1+BgIfrVZUEJSvzIC58b06wUnK6C0QSA3y5yEkTSmgBeNLFnb4hgr6aCvr
jqMDhj8g3Bm8ipSR9mMcMguyazL80ViMjz5JeJPc18MkeugCATZZ8WmcyH1L6aeO
ygZkArgwUsKLVOIUJERU1E8E+l51QFGHQCyq22QQXAP6VM2eH7ZrPiGdJY8iARnK
h25Qhi3edpJ/zYHGwvG1nZgfRNBFdIT7KBdsLk25my2aJt+gp+f3EWmrEYblyNnl
29G8t9MNn+GlEbYA4OxubLFwDibg/hY/5K63cFYrEsVVxWmpC60bJ/ZtIvwZd+Iu
evaI6u/Z895kpS9t8MnRb0fl7lZ29B8MEiuhBnO5ufMrLERAFG5Ppsi7kT+tkBuY
MXYQeWKCcoyCy5CbHjtie9UcBVoKWNwu3KXwwzUdHMLmWId2NQC0uiDBuu1Exdll
+DUqIC76u1HTJMyV9ayP9FTnuTnMhRDfmYV9cf3udJ5uBzcDjHvZENHZ+xSdDQIW
wnYt0JzKOepzj/N8h6z4UDCBj4lHlwKAJ9to3mS3jKAlZeef75Niahnr0924NSAI
27+rQooNzsK1jRiHxDEywPnN1HgJoSrsjm75lG//dP9f4hZeJ2VW22OJl/ZQMb5p
8ElqOPGAT36UOZktYRLy3PEIp9BL79m6yygpvltFcy4oLYM8MU3jZt6W/XdqAEKr
hFOPx7reaU73CboTIUd7CjO9Yqqmt41HKpGBn3TXKBrNkG22bJ8IRyC3cdXjAs9D
YEYdsYJ4zEqrWSJA+CEdfZdMfh/NmJQcCuXVP6oq6SVLi718K/8UTSk0EeegH9Iy
GJ5qVUlGB9RdCumV2cGWxDGalq7epGi6sBCEsHxlJnxMv8QKiBoSDa1OgHs5C3WX
dH21al4fhdIeSUbPYUvhVBw/oofYEZY0rtfojxkE5DcXLv3Y7kJ/A2/2qfcFpkgP
E4M3Ionghu87ScII/sR2svqZv63TfvkAQEWyhlF58Uobx3I9ydpSs88Te1jFejcu
s40JibQ84x4ClopRYRC8zkwEyVqo9AOSCngR65fpMsed7W/ee85Kg3+vM+/zKSZy
HaFLdRKqNohJQSp4OsVpNomXzdjOuR8VDWLKbUk26Bx8taRmex79oEhUgbOfg5QW
vtWjedGzBFyZv5LvxL+cS55s091fjNoaw+OWQfnTe7VyacQ8GuHuJtbC1UrEyfzQ
AJoFw6SrQuEUJuk52xTBa/5sLCsb9Fphnlopun9ckZLk0KWgVNFF9tksY9d0N+CF
ketj+S8uGaO4V34aOTMXLAb57GHc6KOrr8yT+KLnuujCkapciKeIpdLL0ilAAtCn
9Xgob6dgYvDDF/Qh8GIcZFXPVW4lu6jxbI2Y96LBxumFJd/rw7CJltO+lJZop/8Q
h6C42Nrp7yWUOCeE4x3J7BTDD6bkN+++KecHFX5FdoD9JYSkhAw7ZsUMyDM5IJa9
TlDn/KQQMHYjmk7R1Cg0pZh87LLkl3nLE+4tT6yrwCTen3uBQ/MfGriFBfjZmVr1
/gwfJIJb359XQZBhVZ/rIPBuoi2gXPxtrf/3Oh916bPJ7PhYdmydyKZ/PS8CMPca
SPCq9yqPAEVeGR3YdvRwkXNt6FdyooKmVOq0GEGzX2zBG42OAqc4S3kfLMwIlwJH
wBCc1FOdOlmlntYrHcvlWqUBEL+qnI/cGJ2qi/vTuTBBxZ+Cyvj2uZdPfZWSkHwO
/t1C3JLpHQL+RZswr/uSJKITq76T8pQ3cnxIzORkv1ieMaok1GwDJrPCb9Qnd1Pt
N4PEFgLnHk9mxwXSE1LEkrwztIwrPwbsg42lsdYmVfBys2Qa1Z5BD6v7a2QftEsP
denTIsVE49qxS/2/RG3HrcKEdpywzkib7FgINX4QcYxRzV8m/c7BOQ3jEstVfcJV
HoW6dDVgMvj/g5breNfUuKFxqrbfXjDY/MThXzj+vE0un6Z3aSF8U84MBANixSsz
+qH56T7J0TsFj0qojBE7k+NLLBhgOAqFfP2APpfVV84+dsSWHMqy3kIGLsusPdxy
iTzHsw5CPuOdf3/nifRdfOWr2T1PBvUnhVGLK9SEPbKXpakP3/Pi+mvcaTouF0nn
6S5zYZFhUOD5kJt+wnmbB0Y4gWPD41yF+p7tJF/DptmUzx4WzScJuZ5eBxpVospe
UdqW6HfP6vNmKi0cfylghezF1AVKyjH5THZ3kgluqEux1VtWzDqcew4rEYvPnlyP
PWGbJUC5XQUMVALnkmsKwfpsyyAK3EMTQDZfm0QiSbpyWR+11/nQLTTTfibDN6Sg
OHKGBvuqPdXlta5NcwhrUkLW556oJaLNoErrezSFLhUzqdeZbxiZHbS4QlLE3rDp
WLhl+jIzDtZtt7SEyKpNVD3ZasELrA73Jw52QFk9X+wupb4xSJmvRB6XgFpNyLGl
McJp+WPUWkqSzm8kPwcsiQ9ZqpcqMAlQXacGlVROgiH4K4f282cnEN7Ep3FEHwWY
As2f4RADeyXULs5EtpeogY8/5cZN+Gq2s+1VQOpBspokIej4gTLvWe2XSuiZpUYA
KgTykwwqkn9b+t82hn3meEPieiiTDnHotjjnIrhMbydHCoaTK0vSc5+BoAM53fup
B8JtoLDHjK+aGojvnx2TFZNzm87/kOna02bP73MDnMXmLX4W1XmFHZydgBVnEFkS
/P85gZL3jDT5H0mElVzbXnNHTPLZhxHNRnoXBRCBZgo70/GB4+9GUm3M/hqU8jVQ
SVfbh997sGTEYyXWD+tPTZ5r//Sarz3YJbVs0s54Bb/O1cBQKVHOWHp0Z+8JCkEa
1SJnf9U4BB4qS0hyibLK+0QQViPhPnZ6LqC1c+cXJ7mgNFk2WnqnbbPWI+8l+t2b
N8WIseBYZNX/EMrGFqruNPbT6ARyrp+XgAElTJVjC/biZwQZcrdSnv/LeYl7E4nw
P9NZc0+nyTrdkdSEMLk0ZY1H+vbK8J6dLXdpbO3eIojUP9g/2nXERVvOi17FXYgh
wl3kuMh2gxywLbgIIuKSDbSICiKxoAuFDPU52BLNmjka+ZOu4rJEK1ikC9DMUoTE
8F9ciM0x8y2uDMG3FuBdXXpXCGpZn7LN0oa4vMhJ1leJ6onyViJ30pwbBpKVUCfy
8XvCZt2whwBNgIRXtM7wptHlLOw1TQmRPOCs6W8o0dm8jldzUIJNZH5W7WDnFDw5
83kd2pKKsy1SFr2gu7tThE+B8SFHFGhxlJosKikhdzKuBijA9YFD+PsqBZ3LXoR/
d6NU7WURm96UFAg4Fc4/gELY4VcbUE24ITIca6jO8hXSu4Euj/oMuOI6d4ROxdZ2
x3iOI/QvV0NjcrIZCPo2QbsahXMQ8QNDijh6EsefYJh1gjLChXLNIefRIyROrKEa
B4B7QcKx2t3AFz5/sOCWaaavm1gg4c2dvU9HadxocAQEdWPf6wtgOAHUOgjlvgTY
A2CqxN7x1ZjfZJMGoGtsbPzSb4NByCh/6SjEffCDIhZxXcfC2IvRTW8pHpSwH3d9
aDtb4ue8ba1p04vG2+ii7wc7fGv79sDqIMfCKQBeSrFsGCf4EgM/iAyPKD1LmYB6
esTQi7nYUH2oKtpCS2ZnEu1qpHH2q41qGjAWyNPY+X+e4d03RLjOY/+ssvRFtaso
pudlGwB87AlIqS0iElY2NBsx3EYrha5xLpuoEnev+GFcPfjdeA3EEDsvJcxOJYtH
haPQV9PIodF/3LuxB3UFtQcd2X5ygrQcrJubihGfmcIoVwtR9HW6k5FH9fz4dtu6
TsHjYB/qU7//j1DpZ8d0M/B1x7DI+cIZ86ktklnXwq5Y1iKnU5Ny9JoJSDtBsPn3
vLQwiHADGZR+sM9tzSmu5gVY6c/FpnmLjgAMdejumINLpFYB/WzemLs6KSIRhXhD
FnNaTwMmnmWyejs9A4b7oDA27K7y8dmtFY9wU4cdHugExHjgPcCOUbGGsIp8kl5g
AHHFV9yaI6QIvSKsIiGl9m4dGn8Ws2xUG48rmtk/LiOI5Njr/eRRNljAgIFSt1GU
iV596bK+fxGQLSiHjODEcrGDAgloMlCe8mdy/KsZwEUruPhlT3KuuATK96/AI3AW
+DLthZp4nE0kCPX7judNzW4l7UtGow0aSfIVKboKviiZuo+96vpznhJj3rTcvbyb
YIIp42bnkLRZ1bjxDb5Gdi19XhRruXApY/hhDnPa5lSEDI0YIAjh+cLpbv6F+pMh
DcOpQyfEIHHPNijRJcUej3cZPcbavDZL5ogyEMBFl/2DgE+m67euv2DvgVbWJe4g
BP9LcCfqrQll+G748FWiTRB/jTr7X2n6O+LPFA8B+lVY1I/yHcEZe1FqNMH3a0ao
D9c862j+Jhrz4/ol90jEhlBg9CS1Ou+ZFQd6mrJIKITk984tC+kU+GRu9m1cuu7F
MhLE2cE92zXCzoZwWypH1qGd4nEZQGC5BPsJvnoBkzlGH75ufChrlFz24MNvxCSL
1ZguW81+ugkE8LYnKfBKzlp+e+RR+QayEHP+nwXBTgvoA54FrycWQaBHzHWGM3Nh
9WiNEewXxqCEJvv35CSuoQDwnThAZ/Earlx10JHsM0YTNEcgMRGeth1eCwSo+SaS
RFjTUCyD1d/hTVN6q2Zbi+U1/kVdbScEfzbxihKSenQgoU90MyRqSgmvE7wIq5pk
FCn45RMKXN8bgvQhgHY6WK8WILEDW07ZcbvxQwG5pLqsTB/GL8Mk14PC+ga+9+5M
NNIFdp553iCjrB0uThVqrGC6VDW6xnxChEK/pmOsJ4+L5ogpN7mEVYv4Ii9pW7qE
Q1onP4osfTnlMjWxSVDFsHtB+igH98kQb65AEKUcbGUMg1i/ZfBbrFSuGIPwjWKZ
5iMesXXCnis97IkC7odSzW7KAEHJF3eiW5Vds+LRWMqR2Qz8NvOAiTE8ywVSqWSr
sBJBidxWXnDg0vblYnyHGmRWp6+AGlz8BnukM+f8/noLeOYgd4vjHaDQXPUqfB+l
xpNvN6nYo7f0V5GPo4/Fk00NKrK5NZNqRjBplK4joFP2fgqNv3LgpjinJnt9NlKM
prB9rfJMXfV+bGJvOVJthQiQDCLcupUO9tiDQWQp/KKUh9u4iwMTPH0nZO7TvOjn
RyXa9nEt86Nzsg8asg0D22PfVh/MnQdvcRG40dw+O0SwPfNUoNgUNvR4XHK6iG5H
Ek6h3qWJ8rEiYHAVpVIUza1jPs136enFUGN7R2muqI2PbFP3BctOSF8/rIOoA99G
3IFk7rj/w91qzhYue9IP32xh2Db3qf+oUehO5HQIg/5P829EtItvJvsS64FnNUZv
NZAYlml4uaXgQ1XoH3AHQDaHkUKKw/Kxl0U6qrjpXgGozCN/4U+vWYV0w9EgmGad
iXkT1uASn9GFIzNn9xN13jqPjbQWIlzkGr8imeRk+REOKix+oFdOMBau4boKK/Km
9MM3R0e39SWv/06aydrGSPpl3WxXBP5KSNzhpU6JEOaNAhayEI4YW7tbGavrIrB7
K0qXwn9vylkuBphlavsZTg3gyLsSSjQJtGRrpYDh2A6Zn97seHxdivbFUbKbWamy
bJVIeTdgiCk1MqD9/2xH+UA3INZG4CXNRBu3CroYuVACfBRsXT9sjNCl9ann1EC6
K/0AgnzwfVWGOinY8NjccxmPrlmCkj5sUORQNMwoUG8SdZozrdmhIVwAguc2a5MB
GZbJYpe4Dmrf1bvTC+A6tPX6YSDEKCchtH4N1dIrR0VarAmDFTlNmcxRMrnmjgXo
OFQJBqFmmtpZ+KFTNaRCKHgMzULpgVttiDCO1d4HxTrk8THLnBZCJaYzkHOP18a7
N4kk7SllwNzJeWwUwLV4kfa68QR5cokaN1Wr+nKvbAUnflxKYgFwYLOyEMQxhJm2
77Ez6ZDzSOx+XuWIS2VsmRqjDLip0O99HBa1W6n3VLpO9/+n5vVA4n6NREz4ryF9
MzDAL0v0KvDHMCECXB9TtBOV6GPoDeiaf1WfzOf2sgGHeEMy+cZmRGIFfBf5EXSx
+IG+AZ6vKKOvPNDx4lLB+63S6VaD98ComFQMjfPMDmBpIvzh6vQrutYRkBqOyxT5
G6Vfh7H/O4xz/dFB/1soyHOc8f7J4fTVv1U3MMvSkUsRIMiDphRxd83FGeJMTlVE
jG6LTVjG79lGoyfyC7dbvTVoVZEzfMsQWbCrBpZDzQRHSyY3uWdJFQ+zXK4rgYw8
MD8upvH1YYBwEe0Txrnt1I25rXqBr4buYadBFtg7HvlaMnFeGtQtXwPrzYmTBCzj
XgUp9gruKWiNvGGfLm8kcD3eni0ln+IVmtnqMBDyUCATWhVs9GnrTcQvX4tulQ7O
EBZqVVYGsNHFGXISssX+zzfHf+BAmlnSeG0ydY0S5WOv/EPND8cWAjOc6EbS559D
QEJ5DpPYqX0aoDKydqTQSPDI6Y3Xi4KCRlhLHPNJozgzvXcYGvvJUkjyWN2wTLl/
LLLfJf0hSjCPfOtBsd5AHnSXjRWzEC2oKxIlsqXyi8GkN6bgYfKHr6rRj5EhJQvR
KY56HeH6qH1a+T9UnGUp+VHhzPMXPAWdGrpCLqsMBsTTye5Pdn758/kBUTRpQO1R
3NsNnJFvFg2yayFJ9+iQ5hinMnzlPwoxMkb6bHNKsQn4kT6iEpGgW5wLYT/OLNNp
/pOCXEVnaVBdt90V9hWQN1fsk0eIKAZkr1wDf4XwveGoRoeXoVKH2v8Rp6dcEYv9
xBwHMg3JuKwgza7lgSbIAGcVc3Wo2K3I6oaZ7UVZqnIM72oXfc/wHR6yfv3Mr0F3
ORGr0l2Mjstdadsdv+l4ecp63lX1IjaMjP/VgOL+IH71jNdlH/jheZBH/rex1ViE
q22V6YqDGHbxFiqgwWdoFrF3ll+Q/AXC5zkG9tiJRTKY1WtkBcoTwPA47c32hDUy
ymnOfCTqk9Nc2LRra6bMJFEK6gadlAnoqgoeJjQwNENjVCPWLGrZg0PKMUtJb1kt
p5IWfxzdzYilVX3rxsahVsTIKAb4efSZuBewGdbmsGG/WPfR97+v5Z4xGODuj8/a
W6etiZP/BCTFpYr/zYEbQkYVK8Dww/UEW5FtLr5sSBh1m9/83ysiXwd7HU0TD10C
ktTDL0mYtEwUK9aHFr846DgPm49WrUoKMh6F/5StIwE38GxYDoUeQguInqt5JvXn
HY1JuwyFbdIumT+/RI2ozuvqaB6Rz+ar60XNejBb4aIRWyYT4q5MwTIjPTaj2wJB
BgGe7L6R7vVGzQ9qkSWH5TrSzRt2IViS/D4JMfw2BdkiSIFpWGWT4mV88w7qOOo8
1wUz46p5a/Y9ojQ6kWetO1/GxhHBfs0opoaUH+VX119KqGWUlJpytaE/BfA6ycz7
PeMnYIdG8wemvkRO6PQ6p/cbbvI/2IlxJYe0Uk8rjmit5O3gz99ikT4z2FmgXxSx
Hw475erUxWifF65b1djLc5j1Ga7FSRsHm5SRpfsWa03QpAGI3+Y8P6f//GMe1l3h
4dnMJ8/aBw6XQG4Ee5n83YTlVRQGsQLJkj+nO2ZbEba5yVYW+I2M9PR/OwQHZDPJ
AHEaniCByVFk3wrvXdZq5ToL4rzsxpifXTd1JZgfe3qVYDryUcwrf4K7Umn1XsZi
kgL9oDpy8cTKg0H9ROMw1fkrJ0VS7snKdDyQ91uznkD7NSWewhM/SyabC1yJkzno
3uBDnmZbSzVd6pPoXR75UHKeeJAXWT6VXrmPymmjz2h76OpUWi2kB0+qqMQ/off9
vzkpQ8EgGi7S8A1S28TLbK9UZ1rPq4PLq8muGWLCKZDba84bGILMSYVsqZ64vjaB
pVFPHtuUFg8osP8Y4E1uIhWa4Jnz6FJFM1z7R5zulcEzZs1trYAudyERYoRStnIP
O6HTuZUz5ljnn9QzK0rVsHhcCBat+/TyNJLp8grYJzbCOesZivxVROrq9+OfHMqu
Qit0ateQb1SASgNl8gHVcOGDYCVwZGRjRHjm4fR8taCOM3qwRvaEhqIqIkQJ6iUD
gmYDMXej8p8j+83Y415C9ik/u2ez5joigKQUcaxmlo+U15Mw2anE1jrvNKeO4qa1
ndOZUHrwr64EqG8JxxT1ct4DkCj/lNCSnstckx833fXF/OL1yxT9sc9AVSVpvT5c
XexEmhbIctZRWkBWW5Qbsd7y8uEzM3HCsSovO5tkzx/JhH6YpYTLCVmRNxJx7Pys
ge48g1/H2FjYr16fE6mteIhT9BjxI/nHl5mZ5ShwG8o/W/YU968T8kc/0tTwlTgw
bn4aPm5/B5jDLVEp4J7gThq80Feut1mnwSCdUnDjj8GguuC3fuGA+P8WE0ihUPyY
E8Y2ITb2xd4jNqbqggZ6C9Ewjb1Bb2tJfMSO6Acd1v5RWV4BEePC1T1ek2dNHCw+
wumVrKKAfVDmAySLLElHDX/pdxijbyjJGF5Z3B1StK1Ce+7TleYpXUR7eez1MB5z
Ij9+YF4SkOUlaltlo+nqgJ5yZrW8xN4njGrD/ifWnd42CkfA0UKQLGlgGv1XzTkA
+1gNETNLI83owD01y1aqCp9Tseixhn+rszb6hOkBPAgsYUhQWS66yAvrqVcwKDXj
Xa7+pysvJiOcvQthqVeoedgclD7wUjuh0nGwXDRCaX1QWmSFOx3D6NXGZq/bKvmU
uUvT27RQheQJQpudIf6JIrE9owMThYrw0CcShv/w5noNG8pTpsJPVyi179H+Ppqq
85K7gJChi0eIPjkiz4Ts3GwU1dys5hUATQdnu4Hp++ddyF3Vd++cYyr5gUfAHMYI
3RbdRRGlvRPIzyjl7fQRWsqqgSo0Lr4ZzjL6gUd/yVhUwAuEBpJ7qzl1sJviFKSd
JQdJM/bxWQriNa96JY/H/NSfUcnz8Q8ZTjOLdwwOokoFkVvSC/qGJ1zjNkfRLSnI
2Q/azb8EPaCioHIRCg6UH/Ja9dGQnIKKDUMwvBamtrLD2B7u3J+pMSrtDVVI/nh0
PLGozuObzjJ76ASXR/EO4TPLHMP2nf913bHt5rlkuc695+oKmftyEkuoreb6Cx1V
JIzi77DdrUquZj0mVSAt9uNeGhXJ9WNtVeGtVGuxqwImLSzihW7ojGBobFjg+43b
Ks4CbctVORcHrjfCDnfVvp8fGyHetXTifI76uUEbwczj3oIR4BymHf5YoUxmpBSy
XNkNlSsBRjREGKtMh4DnJsMgoPlD6WBLVLYmI1LM5PA/n0f61KTqfk6ysJAhMXMl
nHY3cjNNaFKHG4GDK24XeGGfdPt5gXq41iqSIWuaNkVwjRcAk0UBBBeWi9dozmcR
5bvO26wxL0JrGzuNodsdhZ3vAQe3yzNqOhyuuUYEWwJaRAbK63Jh7AYVz5ThGsQO
cN8OX28DrZ/mNGoeAovKNKmd6kon6kmXF/NYwzG4Kk7R57g6ZRaBgKe4EmUue6km
610cJVTUVg8edLqIbvgk1bqKI9+3Gi0mOY/+M4cus+Z84I+72p5BSuK8cx0mDe3q
Oa2B3VIO3DGfTPrZLCCKen8W8kaX9OrcfHIEf/j5LTQYfRmb5V0jv+QRdCOQfQ1t
83HdJx4SXTHyaT7s7GNytFYAm6q0qYW/8NPbK8XKEO4ePfPiljOVVh+3mA8spyIH
UXRQCQ5Syptb4yUu8uGAiEF+FkuvuDnn3srqxzYXyirf5eyHFTFmhhDj+5ixbdFz
0H+MEkmJqboNsdWN3CYTGvDRatKVmIgA5qqEtMkzPWSTCybWbWA0LgL+kgogu6cv
ngSPUWlmi/dBL3zSLByGuqXjx+VwIW3roI77wAcjIuaG2nexkGU9smCq4hbwTHn6
9y+H7KkNUfT70gLQPSXdkV/2DyTJBJ7BQ0RSoeGnm5crTOYaSbssRvRWuJVH3tEA
mMxzxRIhGB7NOXCacoUpYHnPss3asyHXGNyEhsuf07gEOR9wNZ7WkshDIlNeZkXP
wCU/mk0HovLScAuh0mPlpFL/L+Lsf2mC8m00KNMKRcNpQwzxZNyTI4bHwanXEYuE
f0tFgk8d7iIhzyJw55WxczUg/37g9H1rlebQoRXJsTyLz9S5Svb8PkfywZyG2/OJ
BN73InJcCtdn5jzKld3+rMm0vgYeRrKKjxNvz3nd81rbNoEOKz1DfS7HSbEMg2so
rzFfX+OAc4M+5Kelt/QG2JzeNDLafDvjHBN8L8dExBgFDgRrSp6GaH32TYm/TDLu
OfUnl4aV3wML6noWsAFoeF0e0bE1glCDfZx5E/uA7e1Okp62w4z5qzWTzlluDLhF
jsw6si5Y+wCdothmyGYoVRLYxjxQgWmysJVL2xWK/G/cxqwX5WIZ26cW/4tODLes
o/Op5LVvCzCUtcvwm419ZlaPlrn0vLy40/MUQlaTCsm8wUoWA9nlYDwx47qNF98/
NwGkwGScFiqhlfTgS855KCuQKHT4/BO42Hklg9VLwimORpe6letPhhtKu+2CNtH1
L62arn+nnbUL5KVgtUO28HybB8ge/n8Wss/vGennUTldkXyo9/ArvGvsFvc4Ov/v
usYMu4Y2sR1g8LgiMzS/Qm88EB5Sa1mYrVjRm2/kTOzXj/hq3gaufAbk9oHfVmWa
jrDei1WREPs172thNYkInDRlkU5mK6tHw2O7mrOlW1vrQ5WaWnuvJpseevqqvoj0
PxwzmVKpM7qcFDLVb3hFrBfFFFmQOMZZZ2nnQy08oyYU2glEdUVkryMYD3L2PIJT
p35vLNaA0LtjyQmQUCx6Orw93b9f0mGxnhdjdan4tHzXss0PeeWVA2n9UJiYkEmZ
V5JOGOXaAdNOFNj55X6ecFJ+ZwY/eFNeX4hnDTP48rrQF2rA3B0bX5mT3ouYh9nl
LP8ugwzwqgddK6d8jKpXfAT3DzTolvICC+LFruxWVvHXZRKIU3UFo2CQ+FbjN4Yv
y/Fr/aqZGYq1VtibktdiUbjeLoFN3FxpUqvIS65/n5veNbyHX7YPavcDj6LAvoQZ
Yv/DvbeMFLQojLhbsBgBETqjjAfzxj/+5/4g0HAJvkGx/cIkVjg7gHp5+D3YLDTd
revVH4cAAPNtd6lCbSu2W+Wv9ulOQCLNMkXEFsdCaT2RBsc9YD9OYpfJd46V3tjM
k2tsy3Oe3lCkaOvXuLKZHozvDhlwMQq8Z8VdwYLT7YReDF++wtox/0w9ODOwhpy3
Enl5yjmwF9K8Z2nVbMH/rUnEKlwrhNxP3z4GVHLa7eclpEighifYh+PzMlBESPf+
c7tviR0MxvVW/68k3DayaK9Bq0ghWTFV5tIGat2Cxpj845au9ViS9D6NXbIj6q5D
5tzF9MSjycOweDaD3RNi9o15zPxC6/l6D399aE6sAafE+QHEERnFtBb4gMF5XTrh
5FDIgeIdWmJjOn1FskEMK2p4KxYcQuK3NC5M8G+V/Xr3F7EPFvoXji8GksTrdhiW
M7PcHbi3g6vgXgQP/PQp7uVecIQSBrTYLjK3uIxW4Hl4hljV10CO53lytoENnsic
xeK6FnPqGeb1t/M4+ET/EB9Mkwev7L2/72QRmSHhjI+A0avI1pIBeBF98gc8ODn3
w3TlrBKXL9LFJJIpFKZWd6qoy1R9k7gp0X8mAetKlxHyK53LnY3hlykTD3bO6WZG
LZQhlJKv9VdyTJjFi8yq1Qy/twojkSRAjpk7mLtN2oOXUxtN8jBtwL/t06dYSjs/
5/XZi5NgBbsezPkSgqOBkv3srF6Pa7+28bESofC77iEjQv5WJCO+N5LZhNx9SQU9
DYY8XB/ZsmFcOvYfBB8t4w+ErR+UiRQFBG+SG2/Hdv4IPDIpA63R5xfaR7IKe1/p
41r6TDFojHdNiWI66FfQg+p1OlV6oZQRgsC3BXK+s8j4YPM6pHlh8v4YuwWhDRHD
i1kEQvU7dmf8TZ0HiLvC/vwQcGoPKJfuUkL25iiHg0mT14+O4poMQrr6oS8AnIBn
x8Dxvn6dbZ+EqxV7kPVlLOT1R011iuMLB+ek9Gek5kovLvQdwuXbcahbU+E0GwLk
fe6RDCS0s7sfvFPaJK+3T0EeiRQVMzWGz1T5YYTqnq1a9jMX0vsLenBLoHx6hOgs
Dr3t/ctoqqBH/xPYpNICvNrmuYLt3PshGdtwCr5iUYi0GkHlZVZZYhNQqK4SIeXW
pc3XnCfJ71GN6eXkyl8HT1Kn0SpqZ86fkjyeteVmUuFeG3Nby7hbizDlFuXNVGqG
RD4Ybm1sNl32DyLygypW2WXaHvCLlia6MsLqv3Fxy92245mqbJp71mrV5RblpcTo
MY2f7MS9WsKyH6kf26X+oNnOewXEzJWVkbX5GuybjMGEiC0veXSF1dwIMamk+tRb
gGq+efYpa/2oXVTHrZOKHx3Bd5LS44/WeEwI0owDHGoZ8LXi2uv/uG7LnvilYiX0
I1oMbroO/yZBTDRcAV0L7zjscnzsVS1+A9rAD6bJb9aFakzUdChWodYeCZ/p/6//
26n/LS2AUPB6eBx1YecGQR5RiNenscJJXIsHbD7tPgngluDMHw6lN2XahS5cwSx4
Z3Ic+fCU94Sg7lglV4mec+4fHRZFMzYxRW3LsgdYmEMkm4jldYlsClGpHzeUQu+f
bOh2O9FWP1qHjIjWmXZUIosczsgaMAIL79Mr/EH7Y0gR0lYpjvlCs22SzExnMEEM
IC2eN2pN+AWCeCJHj3dgZ2CwairoDRC0upomcOe/8N7OR99S+J1ehq0Mg7a/kMdM
BrktIyY8fqr48oyER5JG4l+Prhh9t9iaNfcUDo92UBr+TryvJlluAOM44nTJcaZZ
TdRzsBOAN7ihZB65NPXjhQHl5qEbGm8WQJixOepWe0QQwOUDDnJ9eSYgXq52vyqn
2RS2kd5gETVK3rwLppU6NbMvU68MxEXBNuU5rx+hpECzp4J5FAd/bQ7xWezTm8Ps
DAXCNS/yJ6NuSFi+xYMgss65d0APGVEca+OYkXV4qedRw+1fGwrTl7RixBf9YY//
J1p5eP7ihG+ZmKZnQDjQPxnQ4SghfxyEeeTl+p0Dx5jOEuHelWLh3SWaYcJzhiqI
1u5/5Q+FJ3nZohqIJTtFYsjtWqKD80zUyBw+NZcLQwc4uQoETJcqMn8M6kAB4yqF
zGxwn44n9eUfljLSsEFW6Kvdjgu8lKN2N35Imla0LPrjhcHjqLlyLFQiRR0eYHCl
HFOCb0IJ59A8TRjetE4QtPINioJw4j+X9SXlzFutxp7Tu53iBEUyjjjb1p6VkydL
7dlkymdRSsESf39JJXdfuZUHsn0zBtyEHxtQotd//d3EZ57jzacpa38rDD3Qne8x
Bw2bt/iN+mMKanCKMd2LNwwRMs+gefA+vX+vOjxbr1jOMBoMivjGt3JpQsDzBGQU
+lEKpkm/sQtkUA/GuzwH4Qrr9n5tlFUg2c1B966ybC39MW/6luEe0epxSbrU4aJu
WAn0Mt79oCSA2ZpQPOAJzugBEwWHIMsko3J0ocSvI0OmWXCIwfbhoQGzUk5kR0rh
kyce8RQ0bJWXoxn9RXbsjiHKdGev3IDL3JjtrrU0cdd6bzl37/VQH1TQJlOwMMrv
4fkysLwTp6BDkpghk9mYvN+ILfGjMVNdF+7iAF+vwaURWOSYyBRI9sIIV+0y8T+R
wULttWZZMv971nULVmtly+FFIjAcYv9X4uVffU6i9LMOnCRpcqkU+Y59uGqrpxgB
udK2lC/3AR1E1UEP284vqQwz7s1YKF98My6gG+Cd3WaMYXafVvJQzpB3rC85BCA6
G1aDfQ0Q8JU2SNzhpq/rgHKx+h0DBVinjzYw49wTFdwv11S32TO6976+9NVc0ZmJ
OXx9isYmLMtFBRONLsqp9bpw6LtdNid8YV/bHvX6ET3h/eTf9zgvCSPRV9vvaQtH
qW7VvKde9uuGUrrTLLOZZCPBqKuJ2XFSl/sfffjorgKVuS5GpRX0Saj8njKmsEp0
FPcsbpvKpotQ3L0peevDbDvRG3DA9YA+cih5AGXkqMDtMT574zed/hiyBlZcaKLr
xqwkGc0B4H9/uJbXcsJf5DbRMTEE54YMk/2Cvn0thRmkwYtVqHSzHcdvYoYVrhwn
2nEBwQ4gvK2rMhyR3ISLfJJJTHk4jA+PkCIUVrw/uQ/IOvJxgNoegyz1qRCfAauI
dHx4sQD0OrWdQ1h1nikIUHaG/eWKv3Wys7POOTZxmpf1Sluzi7000fJKrUD0WEec
qommhXY5sIjKTUrcRVkkZB/XJyWRUDHASr05JW570pxWx0B/1b0z7UQoXi0vsGGV
1JhxMiY+PXJdBYZYCY56D6y3s7l3qAKXDfDkuIk2YWzGgfH/2TWqELMJTQ6uI+OC
r7rr3IogJkwe2x/aCveFCc2QhpYeT/exuyCENUX2TOG+6dSCxg/0d5oxXH+bhErJ
s9RxpXk6WTz7QEhVsswUFt/qaO5uVvraYbMBgbAM+OM8TFFKv7puFD8b2ZP1JcdJ
7q31w118uNtkRI6gvYXfHWKliTilc0GAupWtNJfGin63iEEU7bgHSQVsfE+A8GED
go6hh1wPe2g+bn2Sr3bYfbAiVCT2GxmdtYBwVw2U8Oi7EGPXHk3hX907p5FEVeXO
qhd5f2QaITUvjvL73jMNAEmiF/OR4pEyycvEy9Ns5lyu0cxqQMlZYvKSL0/YOqkA
SqadnEzEOukZqd9wKeWYOic79dCLmgPlEp4F3astVyMrysDNNeN3VUA40bvCflse
Tk4Wx3M3i7fQmy4H0WsL0i2+PvkqbqJbUKuV5WrDns7rEp6SssHAuSsuINy0Nbis
iX241yES+fYU+1Xual9+YT2JwAeaBf7C25BZUnrAKfpoWpbefN0bWP0/L+vMSWlT
4XOY3ePjHac1c8nlhHrUaZPXrgsao1eFQI6ccEW7G+iijGyoNCk4u4Y9Y2/sYKMt
lDOHIkpeusEuug6B/6UEUAiU6wgo6tRS+sdv6XIuopjmjkU6fRg+BqNHyrSMIYE/
UHIPVhRgJCj1c5gtx3TrZTNg9r62oceRpFD4q4zMscDL8c+XP7Fcdxx2ypW2Xyrz
bKPt0s/YeU4GZ7YHS2xJG3i/z3hPoLHIImEuFtIhhPpMipNklekQhavSmPTPPN4f
3tnAvoZvUq5Q3QbSmTIFYpxJs2F47J39+fI9YJQMIiVk9QmchTRZ8VLnQt82NtMI
9m1108P+t6SZ9LWNRPHPl3CQvQTC4G1Yu0bnahPQ9UgCrern+gpdAgmPNj6kAYmF
DR5UeOwG3WaWAYPPNCqdD5t4fMMJUe33sEJzlzIChPpps1IUndS+5KzDH0OBJLUV
OF20TZv/Mp/kam6Tp/uQ8Dm/3giYz0LAtvXfveHwId5e80Z4dZ6H/Ud7FDPO3C4/
TI5hdVpD2CWhdWDxA5tpGcWbwob3d3ylEEWLTgfAPQkqMwMRMqakS68wNj3ayAvT
tPPSokBIB/mZzpAOf7wkhyVi/Lguq1BvFw2pTYhM1Mnq6bmBaJic2yY6J+jIQG59
AwiX5icyPeVCcuKEVl9/JwPdIADqeCU6SzVKCeMLOxs/uH/h3C/Kk1wFrF91sqPH
ird/w4VYVKHUbNlvtL5eMgGqeWTvpVQx3ee9zY3D6+SLUXqkK+ZQgCbeLiv5y0dU
y7MPozY0ANhI90D+ZZ3B7x7XvcwhgHoeK+r3QFP1TdOZ+HdygoOdGzgTWGxI5xZL
DELpE8Zzp/TvtPNciRzSnzXmAHYuSIbk37BDrD7fIPkMFiebMWV30OZtlSZopz2H
O6N1WCziAynu5/J2FyHcAmGpyVHJkcuX/dV69uZD3DDRYs5JRQO5Ar+lbemyoam8
HEUjojBCy3qHRehE4O8TuNLQBDoFZo4iEPUJGz46zDqY/T/TgYONxUWvqNC4R7+2
V1tW3Y7E1bBXfgnPwDJiD42dhR07eBo3Sc0SwsqRPKYlsGaUNqmL+JX7a3ticape
7FdKEnCusxWd0OmGmppEMvLVMbeg7NjK46mHP7ae47Cw9jOm/PKRQkiAJtLeSr/o
ic6sR87Csv+FEMLjX18ZTsXwbUG82+Jk3dS4nlx8rQVGlqMQtDlwioZEukGHBr15
I8en9OUniyZxYjgLenzBRj8rtp2UigW3LPIo1g59mEjz/nwJHB8Vp5UscItowfMk
We72R6zEn0oGweMSuo0dMk76f2EkyEHjAuLGgK4P9W1F4LsklwakO6vKYlcWiwrP
iVE71tKAh0oLib/8lCNnvWlFELV3xuPIERwUXRRhV9WYudQwxzQztglMUhyjRarC
5GJFAC37kjf0F6OEly145SLrh3xKTARkHeS7fgQy2/zVRbcBmAYanKMR0ea6O76j
tns7yIhM7GZlb6fIfns7qLfRAcjjJojnAU5kejwBMgbej5sr1hkOUJdjVlc0yhE+
I1kVOFfQehoAHnRd+fLm8iv48BSBBLlPnHuFMvoIlR4K71hMPocUOYC7SrpSX6eM
u2KJsu+5aaCyxL+G2/HlPZUWezbSalFsKBiyIWlRkE1OM16aC8y3oRWtAaVOA/+N
1h4zENat79cFrDrw271lp7gfw55WKyBblgaNtOwSXfQ=
`protect end_protected