`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
ddtXksX2+yylW5zu6QL2Lhnb2d1sD00763mmSITNX595NcHTEkwn0zB1Dry37fOW
FufOhVzEJp80NC5qZ/+F0Vk7Ik02dIR0elf3clrjeJRK85K4e3Hoo4xn7YbFUIms
l/8VZSb14+JVGURjfswrIyCUotIzlzVYZ6gzoZwDXIi5gQIBf/gI+KxNXPaKV+PQ
Ufys/12rjO6aI/pPlqSm0hCvftmBcnezN2hk1UeXgOIuKZnogjOsf0iJVX2aOOWE
6pD/psybjbnsNB6kH5uFTA5frkzIzkzl5d9+YDm9OyC+k84E83I/7/j+rk4L2dah
QJOvksSIzN867/4Qt8qYTQ==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="MvBXkzurAa5VTw+1JJ70nePUfoQXBvZOku/SMmg4TwQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
oRtzZL4VJ4iwysPsC8SXYCzXS8Fw2gtZTOskLcDV+1B9Nzn1zTyNtlo6lNICRmmK
ZRVu2BmCc2G+fmzynYlNTnSa7C0Cuel6FYpxCBlOuk3OF2tzAmLAuDyOH3Z1Yjzk
a0aHuoCdIRKv7BrZCdALt03JeUmXKPdOmIlkVGFl8yw=
`protect rights_digest_method = "sha256"
`protect end_toolblock="Jn9CQpRhJt4rnzZPRk+dOpzAubz7omckX1MrFd4p81o="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 19600 )
`protect data_block
gD6l00tciPUa6pDNTk/+t0OO0nC/UTtBwLB41d4inuAUA3i/ALrNyoJVcBnAmEQW
ptbcNp5fxEUJjnOxnedyZEuEBxWRieZFQnkRdF269oMiAhD3m34gROZjw1MVMPxQ
1FvHM4crbgZ/Sn1EROlYaiSFmpCwe3d3aGN8fiVLOGOqXpx0Dr5jHhbDcEKy2eTP
3VTY5GBZ26fi3uEytT6/PHBnha9PazRidtlTy8mF3IVBMxjnhmY8iuJnF8zuqvRF
IMvDnFL0QCqss+C5wlpNTb3ywsT/cN5djY/eAZcxo0KJETyQBHpP7wcu64gsYrOa
ODwpTxnbNEMQCK+SgJOZtRDb+4NQjrEik3SpHpW4hJfgVXGhuaeKWTPmdyMoKNyI
WLlBnhiP6ptZxKOFWABN4x5Pz1TUXXDbSOK0YkDQ9U5c/SiCkCYJjUCd9yGXlRUJ
rQ8Y8rdgxel49bkcO5Qm/sytDv2hF/2UUN+5jHJLica/S7u39LpW4tzioKOSeJoN
ysnywNAfmFnecAVylLaZ5eoQhqvoreIFa0yBlGhdPZiC+YdFC4Rn66obbJ03zY4U
R7rQAOeN2zEubcDEUSTHADELp2NILU41RLqLv4POWOHRfU2fhzG8n20c5qj+RRLH
I+R1JRvnq3jKKweVe5xCvRqkZy3rG/Eb4kyy6H6UTo64y8YvUcb0HJRfGWzvuVcp
gTxzSbYU2Xq94xD48+Kl0zihFZ6E6qAxW4oG2aNCNOV3+lL5Qy0NwVWVbSsGVOsE
9IW8nBFbJbhAI61EzwPw6We0kxozl+SY/VE7255ViObx8AjNjinP7j9MbD7FXogY
yKRTMw9ydtjRdda4c+XSjfYy3KdvU3UK3xcm3nyYxf9xMp3r3BCAjDNZgyr/j8bH
1Rr4iSl4x8kyXkaUU5nqpQSEGFrRDyWDYSLihKOxETElaFbC3yIPpX0kxBB8gz4S
Z6NOAfDTadh95ynj7pl+0/f6MeUhAfO7C6POHdRXiabrYENhyhxTcjkjDRtRX+Yf
qvOPEO/iaLWoCSH+Yhd9VWpFwePB8pqxg15PEBjCaK3fYJY0cHU+l6bkhdgIfkWp
99JC+7rKfZUPS8AKV9vXDDWqPbxH1a5TQzC+7kFw3JBoiR4KIFaiZCAMTwO/8M84
645nJP+CjkZ4SwA0nle+3Q/yGk6VCPYLr7t0eLsxKjnm4Oas5yhb4a/M8NHetc9n
PmSg3zOfVpLBb/KFO8sSLnCB/Du3Eg7lANUoQ58otj6DKUUt6HUCaXfwNd+FoYtb
Er5kBS4/o/TNw1+yAye/pUfESfSYCiDjXWqi73pkaOH1gA6XMvG46/UVLJGJkHcP
2kRlOqaVM59uZIeLAAyGuMn8H5ZWtZM7Re3vAyBCoot+BY/BAljSJlssjUS3bUiz
0yBMFhgCiAvtbKrEqk0x48uwupPErXN3lHJcTmGR7+PgikidMpzKw9gGtRYf7EUI
Avj32WUzW4qopK9SHtzWpJy5EmNwBca8RPMTrJ/hcC36UAEZ/ZamnPkCQySaTFhx
jv3faMU1CZ+3SMP8TInCsMDwiPzX//++W+nzihmCSDFwA+NS+W5hAWxQZou2ndyW
3Eg5U/dL/P9Y1pFu2bHzCuwSKfqOaOs7nGuZaiv8FV2qtxGZ0jMRp99p1YNqsbTW
1eJ02sEyYUk9Kn0lr9R7aFT8spvcjA0bwNyqJFpOsgJicga2sD77Iu8Vl1d/XuZN
Qx6NsEPC58ZYrJi6Ht/z28sLkHJYU0LY6fIvBI7IyoICXAes/29qU1rB8YefNgrr
n8+PyJFXTi63GE/z5RAhBfBlIOb5i36CfZBOrB1lgBvud0FQcgJHKGY9UVg0nvfz
MwbKCwJLc2alb4LYEpVomNs3O/wL1lIQqqp/GvjBm3fEP1PWTrPPXH3fp76JTNyB
VJUkg1HF+hIt8lk3jUJz7f+LZ1v7kwAnoWwJB12uEom3T3i5FdGDr1MgGxcG7I67
sxDc2NnefcNaGrm5N8ZxbWW7ergHr3q7uANhGdyNv0ECYld4SX+xDYWVEZh3xgiH
ocCrvbvtE4Q+65eRJqHM7qR+XLfUizcOChwg0VL6VXEAcnxGX4e82hdDwb/juAkJ
KVWRK7Rs4XzWaaQ6eZ/l0I3UICZVeC61+/ZxfqZCVI8TkCDnp9Dp5ENBHrEC7IRz
bv1W8R1DVZOS2+mQZKzDmRs9rzuGFPalYx5t5BDDMBP7uku/JdGjXrT84ttLGWpR
ON0dfjnufdr5hhvv3ljz4tRPleqYk46R4eE4BUsCrREmGcFSHe2a4JKp1/353N1B
8LiK+dDveT95YVdDOQ6WzVQBQtKlkFeg7lnDj6IbDC96oNEgL5zlhi3hI9MxcNrv
XiUfog4ufwCHQOq43QDokixlLwKr4HXTbPcNOhW16pUe+vou3oCRX8hOqMfLS6QZ
eNZeypAjkBTgsGNin+/FfaYrk66bbNRMWsxTu7D0wr1G/y424mBvOYYF72jQduBm
7N7I/CDmJqQd6l2997Nk4TZkkzWmFPaYJ5/TkOmlgMGIDrYumO8e3xIP3Q4FusBn
nVdzBxz6N91j5uF5PE409RiHISjqA/M9vC7/OT8IXTVVvVk9KZgGfIOtYNdeDf6f
1WSoIEsNCKc+UIjph+/imN32E9n6R77Z01MLcP1Y1mIHVBLAGfWcwjLsbJdC358t
MPGSwq6KYZdJnr3Uclwg+qhsD2Hwk0AP3jm5H/5zSkIHZCF6x97fGzhVWK6rhSsR
m2oAa+RuhVVhY5TtytZtsGwKAb5pg7CaIwwCr0hxi8PpAl4bPAEFqiWi26g7yHIs
mBhlX26ckgcV69Zss+u7cKDCalHtK6dsevGU1marUlc9anUgddOgkWi6dRRb32Pl
BZ/iz8VG9hkdPhV6IRObQQk5KFfeyF6hthEiHAmmdOHqwAKa3AnvE244lTEsHN7A
2c0P1z1qpFXIK7Nls9/gTPFcNukoGI4FOGjQOUkbJqlINa6h6HuiXOiZUmi/xJuV
QSUiDNYgqSRACX0N1jXQFPZCogYp/t4qyNLFLH5HFp8CMXkEOa4CIqP7rOq9gmS8
3GE+hUsOX/nHsogpeBELPr8iqDlqseaOMsXzR1KD7VxVW0rEl64ScPvgH7GHdzZd
KleZu/jNxxp1WKO7wvVHoZNJNWFk0jONUBXaEq7F1mLoE+N1AO6tnbWVF/SFfT6S
28pr9FMI1daXlo/Nnh/whuIWM4rpff03rYK2R4kFbWBGUYSAT0TfQGmpeyGgiLRP
itdkJxGicPW7fYcTlDMPb95Wro4T4CBfaklBbFuqikzknyBf4cp/ciJz5KZi11D/
hMO4QVFt8oqioLdXj9ApyZih1YUUQT6NcfLGuJuym4xp0Ok6S5TD2VElc0tyIp4r
l8EZX29SNRrvYlBxux+1NhLUfOZ132n1bDtUlRbHda6cAkp+8e41/cVxEAdxwwW7
1+UOKvKoJJDZLia/l8AliF9NMk+0sbygEiglWW3EuFs2O4KxB0Trc4rrLrMNI7aO
h6gBOAPrn/BFaKJeaGdAdEAjNLO45LaZPSa7wsvtSSq/H0V5/1z9N/ZGcnORSB5b
TEPYSoZFYfUBaoNqh+ZhauAbMG7LO9MbJiifv3pFjs8R55fEKkCHSeJUyLsOoJcn
OXtqgYBR6bVyuPTFz+OtbooqBWPN/NsVyO9ycS3re6R6rntdGGbgOX/RRY27nahd
Y6oK52zFQZfZ3HH4oMHRD8yi1lsYRKabyVWbG2RNmIylo+5C9P9lhraHdzET7I7H
1nRKekefhTHN5SELYQfGeNE0GZ5h18A/f8ZdJ6kJa63GX4qv70ox87978g53ZWOF
pQOyD6Rk8dFfneCXpSA9etlOcKVTH1F1OeBC7zPjOo6rCFbUz3IYIBPQG5qB74RA
aTSn1h0m8xy5ece7q5xfuzhz4SkCx9eNZA0lbgXExzLvgV2U68efpTjOx1gAy8lL
pcV0gXQZxBypNKppLyabNMNWbOQNiaFxRTPgxlKq1XN8a8Wow6YCm3RGxgYHEoZB
AlBBzQKM3YXB4ZbYBBUNYDoxLfoUtfLB16VYACOJTMmLT0PMeKhoh4wgIQijsN7/
yfYWJCd5N9WP4ehavL/mGpPhS7F84wcYTGswFlL3DRgcCg6DH9cSv7cX3yOfUDze
WODxHp7Uww+/qFPiAyYy8ugoiNvylzQ6ULUeBLcZTuDa3nvzQs5QT1SNSjOyuCqO
zUUYud4ZKDnWUUXtouNzLb1xLQZhZXdnm9gdl3JQRHqbze9IQRyv2XTNF1kUfQfo
OpEcgPblLEo7YjHumbGsLVfLas3uiIsjBTo096bxz2L2xzDmGbSu880PSIlRuUno
KHIEiINxBqDQ1F1XwL/iok5tVd5N1sbz0t8SsEGnfnhGnfjxBTynxk63VtKn3+bW
jCjuZlBx+0uSJ+BDCbkRmY0gEqvbJx5tHDAf2QEIjFls8gKGbahftfkqzv1T/RJd
GkTuYiSagm/cVTSVjsmkNqWrzbBccZct+mVVu++wNIZM7vbEGJe3pB2Xj/8+uwKX
qW6w5kSuRh7E9dpeJ4VMPi3pf/4TQ6e4eQhIxIvLtThBI3okgp66EpiSlHLzWTPG
kOWMXHe92jFEBNW7a5lGYxHv7b6eXCMKRELAONQ7MitifHtoPZ/CZA94u8lo95Ao
09oIysO0rz0PVooHl+RLXYWCFfLamThIpGFqRNgW0SiXyPp7lAgR7EHqP598xKjo
rpBTz5EDcUxyWIg2D1FPuGxRGBesIDpl6S8JQkRLpi9MNfo6ZG0LXL/FEkD9heVz
uir8C46/vdA36HosNCD9SSSaI3d4Kb8HPxVhI2DNZW69la16xf5UrvsbQCKSwDzG
tCsx1Nfhl6/ZL0RW1HELlMpzSV8GR+wmVZkDUfN9QH7+ksPMkjiEGsdVqI0TSn6l
L60nwK/NGT+pJQ9FhFaKiZM0qgRC4QBFyJ8NhyiQVWGautNJNuvR2J9d/AK9zXtY
CHYI2jRz+gn4OhbRufmTUDhhVbzc48FnwzfchInb9jH6IFa/MDRSqw190dvJU1Yz
vRtoU/hJvWyLXVaKEKn0RMF3Wf/Abq8Urt1YO94iwIHlVwKlfbIQvry97HbIlY+F
nNGTBJ/3SOY3qxFZEONnUV2LA/cL8Of2pUCU0xtKU7C59sy/HBDpG6MqGwIlpn+v
vdbuXUSIUTrE7Fm/JVOfMlBM+z5KFSYkbdaMHXvZPnGbJRAWqNq6OYs7WYzN0RNt
/ywjjwiTny7RGEP8KekWVaSoN79taxq+YjLuIPCNV0Wqvn18f2KENCVx4RkkhuTX
qCTuhDhMGxLJt55MQBT6TgCpM4c0Fp3WCW7bzJoYT3iudYcLzNbvBihqGEhrD1zr
KMopDLSMgWK7KZM4Mxro9bX3v+Pj0Lqmvtn0dUQGVjHbJBdPxJa+jnRSptmrjS+a
pOzaDToqTRoneeVzlRxU/eS8NBl+4QfC1QNQc3jsROV266dfgW+LXACaFL+9b8Kh
AGreJbA/KJBhs4FNn/ZaD6VD7zvWz0ZXDIMGk9V2PMe6FQLZh4TthlBg1d+JoVXB
jlWXblZ6gEB/QVGUpUsZoXaksOSllkW5jdVM8wgPBI50z+ZZcp2llLGQJffBcBEj
lOwgmTLN4a8XvwCYnoXEr9+Qiyo/A5WZlBW9qYUZtGftiG31ACQnUmwbQnBQ6bF9
mgLIIsPP+6kCde29RVwvKRzI+F9vUCLGpBSBz8OgBSQQOUiusep2Be9efh9gcHFl
7xrfTJQ9aZjqS+thGC0O8hlDuDmzB4VUIfVbO+2RziuXMJbsh5PIkEa9KUPf4zZe
btedzzS7QJOPy6iVtwYxP5ag+DoFNzasRa+SbwtlrYanzjpE70DTqVmABkR1Zccy
o4DOlhOYF+4Y5lN/bNV2CrcIvHU5wNLbEmyAKxkoGv/YGP2RdTR0+aamCrIWJB6U
a2811C2LNCdN3grG7X3oHPtrpwiU9Qa2TYzqNn/ss4HP35gT5RjeNlwzaiGhzkCP
PwAfFP/tEySI4OmGu1EdXayn8NaCJVEiDGt8hCEA4Jof0tfcznRmHcw0NY/IHOKp
SNoSRORORlzuHR2I0wSFAcEvmauyrH2WwArG7+RjubNmnmOF5OeJ7l9YrULzerGP
ZvuoIq8qapIh0mRjwLWWDxY4nNvroO+Ryu7OdAg80bYDqPDi4CbvPjWFBqrzxYmV
xl79ouh9CwaAguu6SVDR/nEshyLqMV7RpmPPQW+Wc6dvmZaa5tpvcTH9drSyW8ah
5ZxffNbgeMI5b63grcXBt6y93/MO1OJIxNJSkZuyOAcn+WBae5Ig3+S1PyO6rlrC
hwR0DO4qUR31R9sxeqQrmMtr+WY/lCV4MTkjBvQDu334dHR/L/byUQY3GtG0qQ4r
Ifm1Ymz17qqNqo14sfr9rwRDBkqp8sm+zDlbXgYv8D156SbDQhVpKAYb+VhRjQxR
8Ff5VVutwhekEJcoA6iXrFV8rfwO30l8jKHxpc46Fhk1F9LNomC+xYl2aK9RGHVN
Uf7OZKm//hQKnjMZAyj236nEGaoxukRloVHwwkeQVbwk9KbTkLgLkFgoOZk7zNll
eMVJLmgQA43c/NKhz8NDthYWG8OWZdMm0iCrCk6zmzispr6yCx7CxEWMf2OMO0n6
/3q2+Dt5i+nF6AbnotMef/QxmLZTp8FN0+wfng0wbIbmCK7ib3HB2jTbXAlFmv5s
9riwxDt0+I/iNnKrtYyp7svgx6ngJQdwl+o+HFQzBE/Zf6reJMYpVmxiC2PDKKa4
dtUUbRyzTMx5uWZrb9nL8IeWqhgPfBLfnFC8dKMjQo3Tp4ZfTvuvtiRLNDIUNUFn
298VGDJ/k5s9vNGHkn4Pz4ikfAEU1662Sl76UYM7PHYepiN4/U3oebVEwg64cWar
eKR8wCPqQ+vgVeNP6TBef6BVBWX2UTsX16hrA7hkPL6mflP8NeXL+44hvGJYh9NB
UjNZzyCjIaPUKU+Qox8cR6V3Mh7gc6PiXvYvBTN+C1HfNRUWIa1dQjFmEayl0mwo
lAFks0y7scU4JOIzrMAtoi/3UrWCDQLkzdmZv/VPt86/e4S/jbTKZgDUItT1lgqQ
VNNsWmwSn3QUGE2QXCOjms84hEo7jWtKQ/mSfIO7gVos3T2sIm3pf4E7VvYihQRo
v2XvjLiY//sH9zHzGhBaCWQUB1UiqtcqewBH+tPB1bId2ArbSu6LcWkqlsd9Ek4J
pG9AaVx32EjNgled7dk/V1sQUEV8+7YrNsNhE/E/JUFCOxHB7+OnZ1QYnaIC3DEm
MwvmtRP3wtW6U3HmoU0GC1poO7/Dd8+6n4UWR0OuUcS53KSMnQvs2Ngd7fcdM6Pp
aRo+Dgm6nsFDuFf3Sm5bvqwwHLc4EOSyBKRL/tNfp16CujJsRflWVmvHdQQNuBLA
QiZGnxew9c+3XYZoPGIpgR04KgK5a7nh+SJnqd44RnvVwHEW74mvVbVWMWZHFLHP
hLQ1PF1JvmVIn8RxqFk1IHY3dlgw62e1F8ei3QrEs4yzsDaomGHuTWUSzwcpX1zK
Qw+O7DUoeN7/2R8hMsQngsjRpcjJ/Wty4JWXvJkPHrl/eQihwEeZjcZccqAabMo+
qgUhC0WWpkzjlqtChxzZIaih2dZxLOtAN/EohPz+iYpwWvTBwNhLHTsVOSvnMD7b
U1ZYOThFVHvpY8ni5wwX6MQk+ih7mR3ieT1vMDI89sCnCjHpZlS5VBiIMJ9grXTh
BxpqG8iNTHm/xlP2PIe2x25Cc3HwbvRP4EACCvGchD1mXsL2QY/l476yooG8VJY7
SmFhxGJhJmJkEqH+uUcHVb8l5rWk7kGxlH03IiE+FziddYdiua4uGwTtfuaFSnH3
73lwmnNmHA9TGz2ADsBRPfxv/iEB3lzjTvjn4yuDckZoTGieHJMqxQ6drmORPqdS
Al4wcezIiyrhDpUF7RCDMvXVcnzygQuLWvMSSUfmSu6hFlth3UR0uWj55Hrkio4I
07gWCbXMlytxsx835k+vXyMj7Tz7g0hokyGPzagVDMCnhABqiFXCkoGOJZ85HLuD
UXUmUtV9nNZVW8Hu24UF5nq8mKwnxpQY4Uo7MTqIWVq5dcXDBQlEKgUhfTr2ppJg
1Yr3PdHWHSiCTvdmgsyG3ZFM/AKIaAqJUf70wWR+5ODk8D+HX1RgS9cgJnanecbU
VTp9iDXpA8xdTOgNL3CbFmYXvv/MtBgoiND7Zw6J/tVtvBSXe+h6/K9C+Z2PQJfs
srPmY42hxXOFejaWIS91UclLQL5QFjefnBYCaTd50Gb6K07pb6dYs56KpzFdpwl1
3PdL6aFufSstfIrqrb7G4Qb4GgSYlQKc08FKU6w20RTvh3kmfAdDp1JFp1rrcP4n
1JqOnAC0Kcca2wTEcZ0ly+qjaqujTceJfAnQfg2DZKJ9CyuNDrh3xb0/uUAPYjmL
hlhdNnVBSGV4VKHAMoi/EsZqqnRqAZKAxdr/UGB56NFSZS2bulzeecR50tfGO3u+
45ApjlVNl91gFUWJK2CHyTkbjXCNQgOsYJrDzU22WSc/l66nhzFM9Lor1dXsjDdh
DepTvrxbSw46r3eCw+UmgdMYl/R0u6cZfyur+coMhZV/YgURP2v88NfOzY0M7JMM
4xA/veV5e3ld+Z/4N/w/73C4sDxbCIYFZJm6oKjPKKcz/akm0qt/iQzmXTsqoY3J
Zk/PACgCfiviPi/Usf3EF+7hJUp7hlha7H+9vuy0qJwjFVynyNDBb8mC1vC8eJIj
SS1j2+A4PoK889s/vJDWrbyxUUINA0Ir9xBvAZAEY4yrnaj6sEXmnaMZW8lTIQx4
cvYtubLfd7HYeryKWVKeZ5LjWfceEImio3dgzk9puT5ojGhWJB20UkYKF657KEXA
NghCFmZJcK26Vn7InI5WIIF8fNPiO0pHENAZU1RWcsPnmoVb8HVzzZsWFN7trDqB
uClrZvyRQxQGDOos+3c3IEuiIZSIbqgx9ApJCRw37qL7C4bbBT29P5mjHBK4xagH
F1Fzdl1Kt3PC8ghQnLPhNCMTYDl1kDNdiSqoGY4lGvG7j/qhLaY1zlzZ/9Vyagxo
pBKZ1zwSy917K0MptEY2Gph7pJqbWzbpL1HD/pxwIXn8rcjS7tcAq/5rphjeMeh1
poMRt0vMtxbEHm4Ra1vhHs+4ZYIoEWx2hlHQPgNnYSthaknetaN2AhuqhINRXCdE
jKVq39Mn3N5mnO8nqvVBxKspzT53InwYWfrxqnBMLp6upiBVtflU0RZcaRXgyaXI
Ih8Qqcb7XXOcUhseiMQQ1oP9wqmbZAoHvluPg3dMtGz7ueb1A09ogSotr0ecptvs
28DsjIQ8CiM7pHPmqEmX7R1S6G+kMp2JMCH1SPMEnuy2c3z0LVNc6SQK7q+M7k25
BI+PWfR/6arYe488mx956Klg2D883oxGGI4HafYV8RYoSOereuf18tEvk3RpSl4w
+5Zfeyw1cASe598Cik3S5kXHyhvxWwgA71xPY4s+GHwqOwxo1YqM4ThyunoVX9wB
1kK5wWaXxcBTkCHNOo2xPoRQH4FoEvk2Vyj62SazYPdz0blqw7JJ7T1midUxfEA0
i+all8Z7CiLy2x1ZLfVae3BuLKJRoubVjv7gBfWcqjRKBtSSLwR1urlM2XYcD5gu
nMvSNXECs61B8i1s9i46ONiy9Fk87lpQvRFAkEFDfPzH4b2zSQh7k4v9LLvy4geF
0bKJj87HynBnD4a+PlDnazvQAv6bZl8qTowGBxZPvQIRyJ2xZAnLu9nIaEHx+FgN
/AzcVlvxShnZfI78g2//riogB6rs/BV6lCDhAbMBKQlDB2SlM99Gnaol6x8E4YHw
T98k+9oU96VMGRb8QdkLUKgcE3ZfNpUNfkGQCwKVp1uPcNgE/AYXgLXcNoIJzK+q
Y8OU1xm1sLQXSz0jlt/3S6MwsZK2v6DVLeqCr2DuAthe16ogxRHxafSfUNuGpt8t
P84M7KueZXz3Hb5a9ueQfxSN38MhvzYljMYbsssV+RAdf1PS5aUYS8OsNPFz13GS
NQy6Kudu64+GUQYdH2VxXfYAos5gtWJENwOGTUjK6GX8AkjKvz28uBFF6E/B857Q
qcU4Kttt5HG2HAGUbof6npLkNwCPZvyQ1NHq+qCKbkl5GmCA0wJMYpuZs05L19MV
WErzs7dDFWr7isalC4MvP1Oa0tCJMRelbXjl2LS7TYfFBgVox70uOIv2fVWbL/hx
jaWCqM/wuJLJjwkkaOH8fZHUy6zi3MxeL/oaWDJkWdvwArtJTPAi0nzlBmJh3dEA
hG4/FHiB6OD0AMHuuICl5o7V+My5EDs1XbJFCHEgeCd0GAMYmqSX7mGnPPdOrS7A
VblfI6SjE6fHKYadZvgxfqFtlA97Ht28CguxjjBNAXaR2Tb4i5sZEDW1iykEq1UI
MnTVJbmRSx+hECYgguR0mKM0Bhc0lE8DFdexi4xdqf4UL+YAQvDsHmNvZMZGo3Ky
XzSqeEA+L2WvTTDxuRWgJxl7TMwpxaB/m4AW5rEpkBTtViP2yF2afuZvLdO1owuS
66pTm92R9mc3aTW8c/Y+qpG7UMbU4G3lpwfF08omFoTrrgpMFmaaYtKcw19QuNHX
hZA7thbgPQyHFoJqNPADU8EpPLnRN7qUUt8MimKAol21OauVOkAYj67UnsS0IFEt
5E1qS7ks7BRaTvWZ9CcESsa/Je+AxAOEzQL6t4BC+lTj0/wriINEvsAALZdn1qVb
aJHsQlY+nAxToMjN10kRDyvOIq2F/GiNrVywxXaxMDvol1JFtCOh5mT2oI231VWv
Jr22vMPqaHfN/bgdB8SnxOrMQvkKdSUR/ONDhiv+9SX3DduwQOrNCW028Cqka/3B
ezUWxGbvSgsjXNqDO6usdG2WHVqJZZrQnIbtW5Jo3hsLK4T+A6WYwm91JaWzSBLE
E3iNPu7Wy6q2pD+NvURPb7X7cTexDdrZKybgtDGiU1KkpPjXcK1OYapE/ZUa2WIl
YBugMh4shsRkigayFLG7CXElstqiyKl5ZgArlRIaZSAIpFMVKvpL85ZBVknHZSy4
lKUsHM93lZQeXkBNUodW0pUL88DlMjO5jGsLKwvtpRkZvoAfCc61g7rG0L90a3cq
BPDSS2O/s37Gti+/8zaN25PPqszBcOkO3R2VqrLGX31cfiz8HiSodJDBQn4iDVES
ir6mlC0nt3d189afrUMeyCKDNDgkfd+nBqcnjiZ3Y1F00WDQLMosEW83hd2JrqOq
i0B0MVTYmcBDTnhtdinE/xbC8K9+LuhLVmgfycMt7Iqi6+QnzzZRf0NxEfM6lc4Q
OT6UBv6zWcVhc8fzpMo4YAFHWW5EJOmmBZ/ApQZ9uVroeuu7xinsTDRojCPmZCTr
fFT3XafuLIVmAavlX3hwdpEHH/PIRnH4dzvoUaN5kGhkKcCV+D1NO9DCL54Efl8M
yWxX9gN9GbtGgbCis9mekDYfJnUUNrXl7NeUfrCGCOOGgpGkZbgwu7Ou0sQ2x2rd
QtGOcLZMHf3GIomcKmZIV4bFqOmGYMIYOtlvLy6yMBcU3ZjwMGcW0ghD3HnJw2Va
1wK4LzS7ijM1Wr9aIKx+RpT0wcIHeBz/k2gmpyggg2PuwVi0O005pKiSVmgSLOFS
KRpMblDO3n77lh6o6AUPAnsiHTK/PbDJQ5Q/WkoGWGyAMmzbyyXluleAaiwDXBQ3
YXoi0ljk4pcixpoqirQOQqYGDG01lEmS7r5PLFDjOfLhFWoHzL8Q213ko3K3NPeH
LqC/86uy3k3lW/jyXofOS3+3GY8tz3NmgM9FJM30xi898Sz9HmeM0MhWr5YHJPZm
gk8AAZkGXCwA0LFEibssM3rZ9pXaMlM1vmTn5cim7f78BmiZNNoxznW/Uag9fo9u
JAMFXMl1Vpr7FPnyIb8fIhxFooqOIowxIP16DAXrz0jHwntT/wW33yC8ioY1bz9a
OyFvSGHCqlfzRVT9FkGxD8pvhdWu5T87ENH9z+bfrFXMP48ggHW3oWd0M0vJD6Qh
NvxhuLkvP/RCnXP/iUyVfgxoCqCyGCgxxWW6LWTBQp5e0ntLWbhxWSssfT1ynjMn
KYyfVpmPIX6SuMLY5qJp44c6NwkPpRbjm/0CnpNcKIo9zjLHR09AkWgcXjaphqVG
QUBglnfLlyeBKxY234kA/VUTEkHAxnb+MCHnj4sYMYKvrCc9ucN/Lpq2b54kVCZv
b/UenhN0aashJYeHaQQCsN6kNTfIc2zT738XFu1Ft1poNULE/UpfjkRm8nPY+u3g
+1X49c5LtAYMgK1DBj1szNZnYZ0lszWCyFe31MJmLk5nZEUztb+9QrYyCMpk2JNe
G9fnih8TezTQCnx6I3+sa63YQQK/JlelUeEwnYqxH08dsGdctXJFl6szAw9ajTH9
AWFPQJqSdnH9/tDaOycyyY3yLQYa2Ww3Xqf0f04X2qoDfVsjYcv05ATRhWtbQLGE
LgIcz/DW42Or1ODgQBXg9Ge5Wzo0+7Hub3Mhjjc5mxDzIWbgHxCyJ5stqecc7rhT
jXik+V5wv3+pAWR5okBIRd/gcsZkAXTS8cE8ky6vR4+jMW42qRLAse506QGLijT2
s5j78F3VZeJqMC6dTugcoIPQ73Aya0DT7hzIER7yc2bsDml/UOn8iDq4OZaWfQGV
68lLeqqTmlCoG1p8csNyouGgAKScPd0/nYNHtq1pST0M+JnX6txQabtUzLCv004a
sJBo9/sK1lhrGb7bkc0zT5V9EGr5VRsLF/WDnY760CkyAQtn+GqHg6AzSaRtJ/os
wqsOdTT+oNgAfHoyNsthtbBfXQ0wdJe6+oXsO5x4uNGG9tX+RwLdkItjBXHiGgsF
zRwZ0uZX213Wr78G0g6LI2lbQ1DGNTVm/ey3rX3mzF39q0XTIhkj5XTtrLPHbDOC
nclzQxXx1xRmiVrJRZXtCPZfMg+X8qSv8xVgTSmRIoy4KHh649GW1sOjctfC6mmG
rXA0X/SLNth2nPu0iVeD3gIm4R8vUmuxWiRxvc8tiGy5ZutA3LiImlPtYK+zNkjz
UmbixFUaP59z/SQ7TUEN5e0aIZr+r09v8o31zCSjstsplTKJ5UOwssN0rrWJE3ES
efbbNhyeB7lKLU70FtWwr28IAOL9EGsgZXdig+6xGOIadZ0RHo8TYSKVz/emGwRX
n8Ivb1gV2xiwvUPMynLw94ZCsQ8+4bVY9H5hfZ83JVw0gpvcadp4zHnGK9x3JLBH
IXWvOGb86Khje/xV6N+qs6DCrzbTUgtwvK8BKdab2A3Kg14LANzDMOD6fOQtv7uu
2xYwRPhgiBKIWag8YBFu/GAVHJij1q4DrEj92ZOVdRoa/Sk5wpRssqPFSAcmsNR6
fRcNap1OYN7WuYAXr93KhDGjKFGXbSYw3q+1fyx4DamKO2+bQrbgIe5OYaRZIDHG
2hjx3nJ0nxmjnv9lqsF5dijlh1JIYL/y4/vjCJ5aIR4k2t1kIJMu0oZ8Iw7cXdEA
rkUfnSGZLUNJYWhhsYx0DlmTsJrkColus9tVtRYPcYpfQm7zZa9En6ihkvZ+VuhH
QSkne2eX1D+a1fOTXFhYqgHkI9fCeuvyDikcG7pT8002xcpS3ataKqyVkZIoeSEL
E4Fr3nnnQ51om8bJgnoJBMrtmZp9HnT3S+BIJFkmTCa8+EiM+lYMwgpiY9bqYZ/M
pcer11A7b7X3IT67BJZlF5kZKwhRr2WQANOVLlqm7rXU5oJmZnr+r70e+rzLm71T
vuuB5sC7XIUd1a7/Qo9l6dAJ0oYnhXWuWf3Az6z0haIqe3Cn29MjV+6AxaWU+R37
G7NCiyblfkBLpiaM0gDkcKZB/6+YXK+a60qxUbaM+6malMk7k6XHZtla2w/rWm6I
DvFm8dLOyr6ivHl+HUAj5xpqsjgwPXlwFbR4jlxc1WyP+dvO9ng35Vr3rtIrtEG8
cHlVfhiJ3UEmW4Lg5caY48nOPHvrWgBcwemdzJgPuOxhnSWIbWcjZur0kfELLZ7W
orak4EnrCJd1yNYAn9LXfk49mnKOP5lDAwOZYy42NF71uhZbWRCjbt2wpRXo1Uvt
80khYzP5rfNWUh+o/+gVA/6j3yk51Yola6f6WLYY3jqtd7XcIf+4m0X7Uj8cV3vA
XNpUg6tajbK1aNH8seMK2BlIQPy+LxUtLxSTPi5DNo28YV5hH85VqcAbWdxkz3FH
gHCj8HL+HyAAYrGU/yoqPEHnPTVXgI1fXp9u2nl1mBXSOggqX64i+11DX3zIQPPU
LNSuyfU4jeDMb7Mayeb6X606UpS3Nnc20N89Lo9SXKrndg0d8zA7rR/0Go8Fm/2k
j/IiQzw6URBTq/hqFQhI1mGSAFmjBkJMBDsOPHL7LT+JyBMCq9v5EJVJ8HONhSfu
mn6J17C2thXsEcObbr/991FXKeAaMMlU1bAdszl3+kk3hSmbhQGaARDBe+Fzaciv
OGdJX84v3vENMWEiQ6OBdQLZPOKmXdqizxxVNDyo1q2hhK2EcjZ/lBK1lu5j5uPg
8hmrxyEYqApXk9ar1RsEbcwB/3f1fygCoELYMDFF9rdV7T4bL5G+aKz/tw3iFIQa
Ytv4fC6FAdPT/a+/z9DtLR9kqnd669dNBDJF/3QniozmCxJWtfgsE/Qsx7X86PKF
Ya+X/Hm/9u1Wxkol3HP3+EqKrGG6M7yONCVB1FEGm1C6DwjAz+fYDgJaVt60vGsC
w1aOm+iyswWvfvTTfONB91XCyCurWCMIT6Rbqok5hMYK3GNNSo2VyEo7ur4eJv/b
TD2+ljwxdWyFhaygTBqpiyOoQODwqD9KGX5q4w9AKzaTmyfk+8PAH4YqVOXuMgNh
hCzN7kzyP4OhMm5+glEeu+BdHGjfw1VatltOwLeBmGnW2XmaQL+PH3dfcI8VEJ4a
xDnJAX6XC5JHyYl7ROydiCGy8uY3g7tAkiQGg34VxRyvoNeQg11KTuCyyP2AJjh+
R4wspTCPe/uWw8/l43d0f0SKyRN8dzU5IG5a//649g/YEcGWGHnoRlAY9/Hp9qrB
HNLe6SMrifzU56DOOKIvQrI2qHFgXH0a8WuzoUr0OGEiVy6bz5WoEaug7BmERHQx
MyMhmOKaW1Arz2zHC6566QbEEoB8ncrg7pfBYYUo1IaG1DIfrhhEMVFRZyvbrG+3
CerZf0azgW3BkAkQ2JnVxt0dDEIloZPML76q2Ngjtq+mBrG1gCkgbUMeghUY5AiD
xj+HOzHPgmGGIEsYASZOSYXAOaw6gz5lQ9vSMyhQx5Y67QfHfpX+25GlpCdRmdrb
/COmkGVI7VhpBaGqz6KtyW5LFukq+AnFpELQ54oQto5Nt48T7J8QnkXysFgCUbQV
5R3uH4eTCm9EgdZDMEqYRDBNAOu1KLLtdcKBXgEPwEa1gtAXRTkMjldxqTLLivkK
pWLMMBwV0U/vB2fVzh5j/Z7vDUQL9ks1kHk2XnFirpkJdIXlaV0wPsgz0W53jDpi
ITJ8egtDMOO6tfXSLS1h3LTfm0MGS2854hDaiEI/IeRThmsMSj8ksD5VOR7waGdh
8497jShzQeEPoEtQPYAOdLEEuec+n1zgUS7vIRB1msrQvuBCr6a2C7ujbKmxu0/D
w9//8aC9FC53jrzbw2XXnmeA4YaQCgx09qhroS3xY/X8FSqBFGpblmFq6SaBGkRX
O/AjhougI21thXHSbK0zqjSVKP+NH7V62gA2PVoEtBDFX/Z6e3wiZktl7FvoT4BO
3GizC0VxqaIONH7JI2qs0/ZPlsjfgN1TzBW+r0jfhGKCYm1G2MT+iqcR4IPPZOr6
M52EwFD4eTvFRjJhs3T2dF8GYHPizsD/kXA0DMp36DzqhRboIZZZHrgppjtWgz1p
Tf8vIEc263Yrv4v8RWfpru5BVGApZHt2FbmRyoSMboGqoLCGaiYeBoWapk+fyAbi
AG0qrLVnE7JQdTQKuVWkMgyvPSLo8UdPVch0agMOauFBy7ImosLzXag2H+RpCTCv
BVJK2UbLW3whSqYZLotoYTdc47m1BGTv4f+gsKM5IZ0N69leFAoQ1iIw1aYWWZQZ
gKjUcZS+qRxKnz6CLZ143imZ6fXgpJl7drq6VuOwN8fXEyV0B592SpFHR8YjkbY+
UhHYo9cDya/yzFr/LjjcPXn1dJvBUsJIHNXwOpNvr31tR5LgOMS66T6sPjrwFMmQ
D498azFh+onVUmyD+J4DFxYjfWU+IHaT/3EeKe+AigGClrGKCOH+WSp9FlaRlI9w
/cU67U8666TALtASowmahsuqnYRlTAHY+Fwsov5P4yNlKf1LiaMh6C8+VR6e6yLI
Qe8xI+ZLzAzdgttZuqwsJT4xk8qWXxnBvbRJ+sJYUzExV9mNwXkY8nzDLBen0r/9
ScvwcmlVX6xHltJhlk4v/8sO9jTxR7YcGG3nJ1gSuSfr2XJyHs86ZjGpDUF9V7oI
/ryFWchS4ZR79H43/nJP0R7EtQ1TsB4KLqRZLNc8xF1dM5LFob9L+9HJoBojjZ3/
OsfupUpOkZdlSP1Jeg6Ljlgq7d6F1wFdCF9Poi3qaxAOffZmUlMg5pqiCHZ5mV9a
KIuBywAwwgLjKHjCSd2weKxvrgei8eC8NwSGcqxHv+TI2u4xeLz7WiDC4KKBAVnJ
UT/gS4gLP/Zb3qeFWhPKbI2N1CiZWDziO8+wQw5dTFc4VXv0e2Ll9YLdwDj2XIHO
0mGNO9XqirniDg2SUPAvomuPsvo0lhqZDOky+zzRtuCwYH3urWJweSvFbiYoLRZ2
6tvWcmu1rhaWNek27SwKflozekNrWJozrOSTKNuGd6654wYch6a0c+RTJr8ZbF2i
O7AaPd1vjWll43cp4WkAwGOdSy0KE4c0t7QQbbNWPH5iKpXZ5OePrT98m5PzIL7/
S5C9xxBpkzGa1D41WTZD7v1J3nme/PQ5LAGfTsBYtPiipkFS4JZdAfhxxl9bPYVf
eB/+m76Su9ro2dyBbKVmxRVkIU86Qo9WYoy4JzwxoF3hrbqpxmkOrfd75QbPM9oc
xayYmkWLndvAmqD5efa7REyA29WPClCQgtxrdc87mFJzEFIlyelURKMcSFmMYFK/
RwFj0g5VeOfomgnwocd0KRBQ13rKiH0RwwGOpYCGze8XjwkBgX/ztgc2HFNhVMPm
GhzrbPGBkSA4a5fvlqiGOkDE1erYD9H/r3G4uMk3IGw1F7KjnwZQfb2NS8//JuFZ
WBkLPfAVuAPg0iQJTE/dKV1A9Z3PBxLq7dLqv7SnPOKJDhWZh0Psw2c3K+EusFhR
5au2sVE1EuN4kcIqM9S/kcWALXwLe7KGV4HWG3tW+QrFhJ0DwB1PGvMegiGYk4wP
B7XkWcIoiGYuLzMM1e9lCYPTTxhadOr1KdlAsn8x/XylzW6V7t9+F57sT2pFigKt
569JX72DmDNh+LS+5nVyGwqwDvuVPTFtlHzSzIWNJT+zivuejcm9Jxjo5TtEflWA
CO7pBTqxYjMnlm+1YUWy2LUxOwfe1B3Y4Rf/YlbWNS8OOA6cZuu3bRAsol9Fm64s
A02sfuOcuSdfof/bVrXeZi9xn9nCijtIPP4WBln19I3VHSpYQlQ8l2IdwQ5Fe8rs
9v1Dwxl5wLa8V65yb7285mKJdUar6b7ddbZz5zJwS3zc9eyqfi4lpyqyJZlmiDt3
jWqKLjyrkfsSV+k0fVGHfjRZSR8wK6gIdBsI1FZCAnQzRjKT0XhBsbGxMmBvac4Y
iV/cTDdOFir156E3u+96Imk46H7o9u1mrfWY+KaFRRz69UGniL//hF8D5GhzDYP9
VRL2hed/nT8LcfJEvmuMk1YVDw8ERRmqnPDt2y8PE12yIXWwKaFU5SqbI4oJg5Xs
VHRabqvDIZ62+bZyFtwutjNZnQXcZzJCzFfLjrEzUaehqHCqRMvwOVhiF2XGCfjx
d511SQgLzPmhcNCdEbDjLMCBSHpDIcxIk1Cb0vmCYs7jJQzFGpwWmiBPJZ2zm0il
DJaLTR3e2VhykB45yzNbYZftGIkdqEWq6mWF/OVU6gz+rdiI1SUQfOQlFpA6a0s+
aFOsyK711sI+97cbdHTS5pZsval4HGU9Nruiva2JhJ9WyyCfKVCniaI0ZVBUzCNl
t29O5hO4wiRWHfGNe2Zt4qt7BJhwNvWEI4Ro7rzNmgTfxNErfU4EmLyadSmnr+7+
NqtL1+UQFhoB+8HVbgJsdzFbQRWCWUGvHHq+4KrzmMScU3Tw720wUFQbEYXIQ66O
5kUSDU2i41sAi+z8mvXRiQ8kuSrrkgpPogdsRiSqkZbEHlLptSESKikMsp9Zuuu5
NAj2zkj5hzvqzrNv7yY+LfdjS/7535G2wFjtA88gs2/PNCj0zN5mN9xbEeqjNLij
75UmNvqZrCOTfALmhHoQA8ck3uHPvdIqMfyVRf9U66ZYCwaGR9Jjkq8gLPMaHMtD
qAo3vLs4+hNHs5PD2lMIi8jL0nKTZ6TJDQf6jGO+Ccf0jhdWXHeOZ8ENpNsxrTu7
n5nIH70e/MGFxVbjuQgmMbMWU/FZ72tuJcL4EXb+jx9w3IC3CzAc7TPBdJSBFp81
wlghGNyZP6n+1CihI7ZvVO4vOA/MFKDoSIwZYdV7ZViZrmjDfKJi29jiw1+Lb9y+
urhVcNZsV8XH7g/Gh4HNTKD3pTcQ6OZ5e2HAK2zRKfsKIRJE+aptkR/wbAGUuxNv
s6glFAQh+zaVPGAhKKHfTmVV2N7TwkxlfUzyjbjcrIrQrS+9r3Toa1pkX3xvHO5S
hm4YuElCt7zL0ahayPjZRCVZxId3R/WLeRjUvNvSOQxvZzTMArVpc3IEAmJAzg8y
mj/9XQfbp9GomD+2izVN3uTk0kh1JDaLqouGt0qu+DkYhv8gR6EZQ0l04a0PKqNR
JWl8wNfLRo6oBl4BwzG3uHAxIH5unhvdfPm1nEg8sxEHriOMD22a6hSnMHu/mB3+
8TDU1IXLZ1JZjlxzMYVBMHTMqzQnYVxZIk8UGnBg2WGJd40QX+2Saew78/YQV59R
CbkHQiJlOq48UqXWJ6pz2FB5VZbLojRYvQpaKPPxdyUt9j0Ns4k/E9J2FP2R7htb
W4m/ZFpr/T6hZ3F1LPEPQYq+kHDDLpG03BtevC3kmwopQ0RxI/MjK3/s9VItC6Qd
9YjTzHxsrMDaN2GkjEZCq6tCQyR9IdxSyxDqM3AFoL4O2I7l27+OS7Qk2pCZjWz+
LCBOQ96odjVqK0Lypvomskq1wV8s9xxx6q73XUQclyBQ5oRBdCr91Fe409W1SClx
ofhqGSsKlbImTyvAfyBDbq/lqNwGO2fJiuvhTzs5VKfdJVqxhqSnZ9y7AxmNztdG
/JjagLPzmPeud0GalMORkYthX2r+nZgR2n4/GcEYfmGSRpnmcjmI6b3YBqRZrZ9T
EJLPpPmBf9XR4VH5GEBWV6NqrH+6ty8nk45b+4E9CXZthoDxU40oo/aDdRNsKkyl
or6jRjv9jKChNMhhAArAwEGpmKsCZLg23VMzkjgNzf4krG7Dpn0LGoQHV9yqpO71
xFTyU+ELHhxozrVmPqKqWPVr5fNF+Awy3Ud4YC2LoqheO6jooTIUEn5psCOyxwjI
FPek+pUKDVW+S8TeW+DSveZCF8lXOCaO8ZFBaoZ+Lxu66Rkbe0tndyd3udheRLXv
eq0F45ItmRBbkNftmXw9+fx4jV7R8Q9H1Zm8jPtjsd0FAGXSrNyorzuiKV8o7uS9
ltZdGTk/zqWPO7cXhW4h9Do+RKkcQXFtxQyuB/YXQSHWNT9t1TH6yo6Nkpkux6Qo
KNojx7wWU3vF/77fEslc4fGzkMgKxOimzwSNqJDvOxx7UJaLioCRPzSBSx7jc+Lz
E+X2iYmWN+SpnGU/C51HxCCumKCEKTffnPa6gX5Tv4ccyaR5BXzoOG0BHha4YBaX
WFaEkrFAxo11Abl7Yx3RdazpD7ww+73QFHgJn4hDCJFXWZ3vuXuG4Woe1rC3A6zI
LzwoZTLQSTWD3FE5z90STtUg1DImIFP+K0imYpP3DA2xHD4r+ii10TQ4B4f1U2Lq
H7P3B0wXRdiXmDj9YKjUmEm3bd3Gqh/IAhBoGVgKD15JqI++ga3diW+EgwcGcbBC
xrwY9ZO95oNGawHmFMNA7UBIJXJF0TidVU3fBSGS/bvqkml+geUydYnyRtraL/uE
xfQ02n8fa/YolqFhA/e8V6uPnB5OWzoGUu1hzmTsJJuOhbmCjeZFgoj3HpW2+lm+
z/6psL2wRwT8sZ6L6+cUgBoEJLghomPTBqOjtAorzJtAzSxWN9ef6EfKrlC9w8FJ
+ZvS9YbB/PdbveqqALi/ratOqOm88Sy+1821YKiM5l5du7kpgV9qDe7HmMhVteP1
dTbAzYm5R70Ih5qRA9S9OX0X4YRIepid29xWH49cowKF0tvYPc665HGlLnuJjQbS
iPpnpX7AvsK8lkWCSlbWCQDyFQi5VsymWdaLLPISzrP64fNbthS8y/WTNSqpr0cD
NagSkMAv6X2g5HArtLQQjtkyBop/bRIEvHf0Wv9lZuO/OB5XnwEiDkPpMPgxCbn7
r+FEryE2+PA3uMyy9v7ZOeClz9o8ibesruFEnEV9TW97bUMrx3XNDpGh5JbCoZLN
mD7DJDkiUlg/1pc+Bbr1ZE99RF/p6zGWKyK9/aPoZ1boVueGd2gWsglOr16Nw7Wp
qjajI1nQBDc0xwX78HYDpuhGm5YK76iHp5ut1ZxpvZhefHdw8LYHa0iIOpUy9YUT
Ht+bCZTGEyd809y9mt0uFqcFnCaPo2ldz3h1oJaIo/XvCSbO7NBLlPm01nmOmAA7
+R9mfdXDlJfIgDkdZmYDErcTvZ3NA0B6BMtqGX9YXfqiTighK0LQ8SCAiljyUnRW
97Jq1TKfv9z8SRLln6fmQeceXJJgwPGVlD/yedLl4ncsN+SzyS+hIQeq3Cd76O58
Fzd7OIVdJzaXiPrnX+3uUcyOtjXRVNlqRr7PO+kGaGEyYmkrTnVAy/GL2T3ZWiNo
OJf6KaP4na1VtDMIgeeoQrTQ691PxZRzdyKAVVySWYhC924dKORcYnyaO4STtyHB
51nkpFZpjJp8HvpV70StbSLFwVqfiPfBHja9DPq1tawFk2peGQlimzHRSzgyhcAR
QCcypN2Rh1UzLSPOvbZ2hbdftZkYKo8olYGjiyh4KyLqDDWnTdulLJuyjDyyZvya
LOAV5Yu7detKqg+5z6c/F4qdm+pfgi7KWM3JQVRT8CI5oD7/w9AziKHiirIhEv28
74G8/WFW+G9dKvbI7CHaYM+NP/bZpsZSMAjUwa/0NdBBD8WG5YNnNx0VhqsUfoVn
X6rO322+n2PwsTUXib4I6+5XEaBMXYPJDIeKTkRh+PhtdO87Iip29lo4oA5weqeG
8syRSfEuidWW4iwgih8MedrtZZdww17iJ3r0MgH1+6WcK2sjj7hP9qydJWfz0h2Z
JTal/gBBojlPzOE+vPCUNqb+8R11yrEmjdW6aZ76grzLjwoQwXVvBwdLm7RNbOLg
5Apbdr598vL6ikVzScXoa7V7tsrtJlUqOTAPiRJVJCrlCB2w0J0XHkF1QxH7Bp6w
ZavG6scqaCg6bkOUAO760lj11s7gkY+aTUAOSRrOezdKJu7r1sC7Rdf4C9828xfU
5uh4PC2Ed63D5P+HQ7arCeF7lFT5//sATAdJMggFzXgLE2DQDTqJVVY9Bl2Ic2fG
8V7MrULOGhkbLqcsNpkzrI6hux65ifaWrpAaNjJzs/6EoaNyajg5iOv5t+MoCJNl
xdgXp9foG1gwG3Uiv83U71HRkYSUKFKUmBp+aIiFL2FO9MFllsPITqwHSROqgmIA
7+fvsgH8lVIRw5KcglFzLdiP7ErcDQMrWts4+53W38+X8lDAzGJiSTlv+Bs1idRg
hlrYhT1ibsf7SQExKUPowex3ZNye/ul5uGtLZEa5Rq7r/ihsI3DNYILay1Z/Ru2w
rNsijlsMrl3tK29pNtyv+SwCiCp/vksqwM5WJ/mQTpFgEqsfY7A2PG9hhXqwMMW4
y8QQx4oYWaUuDF5n2fGrCxPf983PKNe0NtexeV9M+hP5nSQ/xtWfzSMGTFmw/uDE
ywpQoq7Zb2Mla0MXIAAKKemi1yON10hy9niu1MjQZ9TDiKFacz9j+YR9DFWV4Ws0
KgLzOuZjTsCRzg3Us9tycNpiGXzXxDc0MwsqgQ63k2oWJB1I8qQEoR4/Tfl/6uwJ
BI0PPG1SQbLVfTnEaP4KccDjE31pFmunblUBdTGxkawmHBZ7+2fmQOuzvPhXPgBB
V7uqFGR3HNwk4GAg+o40Co7ZkqjBfKFBX1Yhga5irfO0Y0SYhvdEwcskhCjfZGVt
H6MgbJtTm1e05L+4L529LiyQM2XwN9fxnpgNbwCtRerCeL6JgR39lINWroyJ58Xs
8MqMq7djoUSo8RsVpcjnOE/AhrdmwklSwvy0U+NxWA3VjXPurwCBgozpHQmwL8px
ayPmHLDLpjaW4bjgIk66v2qUhmJHWLKNBcGdNHORva++JBLkGmCnjOPVWrqrLcJD
RuWBTSXHEXhkzoKLCPo38fShe7UbSbF8nWg+7CWSCAm9GcwolLaXV7pJulXYBDM3
W2JAIBWGwkReQsHdSyq9cIQ2vzk4HwuP+vf1nZ0ZtOGAJvYhOeyueGbIt6xd8YXI
+dHvJVkE2cBXhEEzHY7PzyXmTQR3sZAExOWbbmtZnUkHivdyqrQSNgjFfD6PiAzM
S5Pwvul+uoVpnFzbX1KlHRMUy37LTl52y4hpAtGExX6HeqMmZqv1b0v+kEExb7ul
A6iVfyVnRUOOErte8lwCJBM4KWkWtsG4JB83KndTCf8U2v4/qxmJWPHQzEd/DDoC
sSxOQ5SEvWpfIY4ZmvADVTxbcmZCk/BdjrTGiNhFt+YEwy5mESjAM85ZWnsQyOow
cUNazA1CWLdsTRzkPEBZG4/VLJQLBmJLf6IK7Ij/ajaGSPK5xURpUVtBtkB2DfuL
1MD6zpv7HiqGCx5nGX18EePjehmXAVLHHExvjsgis9UfoxnxUugWRe9Hkxe9VMYl
U0ey2S6qavwFzyN/yCgs2EmQgXbmosCmlBbGVAEskBxT4QUhfFiEvo6aUHc7anw1
GnmIqx8dLEAwh+qiqFZFxHjB1QNbKPtfo4Q1+JZnZFtuU2lrtbGUmFf/60wTy6EL
er5pm+zQVhm9WgRIWkUcJjAbsxgNGHUjPkvVNBqIE14OKqBfUU/dG652rlVWQzgg
vunAp5vCVKpW0NMWarQtsNI8VNXLgAsW1oYBA28A+ArOVGmtfVcif7jkKntHn7tj
zusfjk/zGWFC0Z6dcYhP1rJvBlBoDO10dPUKTltvKxbsvH9d7moe2Bf39m+8b2J6
vwMnffa4ttWAguDbn9W9nbAKooXhHAWxr0cKxuwogEVl+HddKIG7EsprUJsZd697
rIV3kEu8V5y5LuvpKrhH9MNPpYDvMoqkmE2GjNxzGLM9NMOp93vMupIT3Ti/iD8O
RFnjsWNtlcnpyjNAEbjEINVh++/kkh3TRGIjj6CQfLhKOHpQ4s2++NlUvMFYrkPZ
3YOpTov/k0lvV1MDj5+c2KUJiLW1eHZRZ6CYS+bM07MSCjEyRaE1+2WvmTK11v3r
vgojPX7YYV6Fa5MR7O7RoAbmth+rmrahm1aEuoW1Fj2pD5j3L/C9u39k9kd7Hhhp
3DoIalGn5FXQ1kwxlYiXVHYVZLukaXow0DeoMawXv1DESDcH89zghlHXyNuZBJew
OfMRMALnhpvAn25BTdhy2HUFf3gkQ25BPY0C6G+wYL/oP8/lBrCZSOe0qP+n4WDA
z+lk4a2WW3mrgSjKfO1aZ90uWV89MF+lCHWD3rSKykvBDa1Pd3zeUeCSh7up8z+N
XnbrG0ADL99grOmPeHbynFJWKqsjsQNn639oyLs+R3w0DyPkGHBfA+OdWHO0JPRQ
0/HqHdXFzz1j3dY4tzwYp9D95/9btresbqJLioxPLbnHwF1bouSg3JpM26nvnw6y
jkq1sZfXL4OXBAYRV9LDtjGQTCSvnmg1QePbPc92Il3aEbucnkJGoDNKy81+sEg4
gp0Izgq+7WlBif9titzsgQzzDwV+d/w99N4REJq9Sc3kH+CbVL5MuoSQYzi4+h+D
78NKCDZVIV0pJlpNISkuSwi1PL2/FpUgD1MFEKGwC6JHH1hilzt0DABfH2EPN1h6
BtdX/DW7+TdIPfRD/9FQW5+7RfgcyhaP4XlgYMd2HY0OazPWffh+CFKooN3IarXN
tG2IxdSlFXXfsI1zwLTsACGE0x+8G20hOG4I4OsWNMrjubCFw46/8zhae6oqY8fH
YbsA+tjXFPDdirtuI7Zbj1LI7xncRdv+vBMbcFreN7VtQDc/R1P5//B5F8nm7yN2
qP+4VnJIV0d0e5AHDLq3WTWE5nxtDk5umzt01/MEYUdJ+zqOSicza0Sw8fagOlOa
hMWgJlnwS0tqsV0dYxauz3DhMytjxsmzWBedKrGdXaI1KkQTC/iESDmh0MR3LD3V
zFKToKON251qdDZaPMoYf+Az1JeK2NPYhLreMjfn04mC+k7eDTqlgx69l3eNy9Df
kVAdSBraAy7xxi4HXNCTM5967DmV4YZT7+lSq7JIzgBPe+g+dRvaUSBSeb2L/cWo
7UDCe+o1WyUwd4rq7pVCJ2WyvwuigRYvKizaSPqDff+4Dxh2yBHjEgpuSI4nQnVM
FPUHj72vDpA8KpVnfvp7ETCS6KfdU9Iky0ohxOa5psHQI/ffIaOGx8GCUmasUO05
eMOohlkKoT4u8FN5ehUAtxRcQH2NdfknQHRTd3utqEd5xaHgCaq3BrDlr/c5erPg
QIOeLkrsKsuX8cmtuBCYMrWn8EScR5fLOZb2w75IkTjFT2cKoPOZyh/9bI8py+hM
AUEDVQPD1GdwPBIGYfzxH6SL1/ZlB8Gz7WOcthAeu6uUFxi6nW9a/Hk5B8Eu2FgJ
z3+kUr9gAY0W23BiTMEfoBbrK+Y1N+9sMtpZrHjetH2zDmSI0sWdt3Y++dVScYqp
F5IZaKr1iYIvAi7fYNrETEy5eMZAGehL/5QheMgVe0FqL3wdTkl/stEQGPH7+q6g
W/cII/kpyh954qdEqH3YZJJ7ta3kAaFMjD2h6xrBhMuUX8xEp0/nmoNZfR+J/nYy
qbzsZ0ny6vwChjcX6s3KlRkHf9GqXfA4Y66fJ7gIH7/iCk33dUW+WN/y6I8DFT/n
/PGuWBdIqPzBtltOUn/yH3fr9g+lKAjCizCTsvO9zIVxz8yNBHYcPzKcfVQXqFaU
ipG8HpouxqMqJJBUr+glxIEYkwqqwUij5fsfvlWJHfn9iOAy+22oAZEYgd2tbJ3Z
4IOvKKwx7d6Fdd6oXK4J4edKOzD4AiS2WbQ8O/BIJzSzl3AWMRVOY675YbkCKeho
ER/2orNIl5GQ8/rKngf14v0SPDVCcsK+67vQc1YTYlL5WhwboHUZkkYXsep+qYzJ
3RY6Yjk404jpxGuH1t62/+7FrmmEZqNDl38AzGtDIP8tpfnBUJuE9WtUXla25Kpz
CYPD40/v1EndL2fapO65Q9OGOUB1hEsa7FMcQpE/IUz9dV7wfkzZwacytlDiTkPU
LL+stizRzy3yANrRTiWLwQytneVD8f5gekFoN5p0pEIaD9nV7ZHaaCG1y2KuL4Vu
b1KltjnDuKc7eWoVYua2/RtoOltFLFwFngVhqjhWTWR7KkN9IsfEAgsFXtbqOU4J
ZkEP874HkML+TKK+zOuBktsDc/l9RqFAG5mhuoa9iiCbCzDhPdVMtmckt5aOX3eP
r87vHbcQ3GYh4lozqP0529gYJQWsRDvnT7qk4zjUl/Et/mypVk9/3UUCbZRr06sX
D0PZ0kpmKdsyy/r3AlY1BOGwL248XXLSZvtnysnNJNUigshUrHwtK0rjTFcj9cIP
0oPAu21CLCfBxGBhdkD+poknnU0ZaxRb3yVNLrIqkWZFDsEh0HjIk76uXusFsOnb
AT+an6zCXRjS5CmgELSnmk7K3ErlUE9smHeOw+j78ez8xFpC4T64bTTrVfCYJKzr
RYumIr3DF1x7Clr/EIhLyDx7BTgtPfIZCLxkrpa8INSzc/Vm+THLmYmzFeRMFuCg
Sbe6JyYQ6N4l3TS0mmaoRw==
`protect end_protected