`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
ddtXksX2+yylW5zu6QL2Lhnb2d1sD00763mmSITNX595NcHTEkwn0zB1Dry37fOW
FufOhVzEJp80NC5qZ/+F0Vk7Ik02dIR0elf3clrjeJRK85K4e3Hoo4xn7YbFUIms
l/8VZSb14+JVGURjfswrIyCUotIzlzVYZ6gzoZwDXIi5gQIBf/gI+KxNXPaKV+PQ
Ufys/12rjO6aI/pPlqSm0hCvftmBcnezN2hk1UeXgOIuKZnogjOsf0iJVX2aOOWE
6pD/psybjbnsNB6kH5uFTA5frkzIzkzl5d9+YDm9OyC+k84E83I/7/j+rk4L2dah
QJOvksSIzN867/4Qt8qYTQ==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="MvBXkzurAa5VTw+1JJ70nePUfoQXBvZOku/SMmg4TwQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
oRtzZL4VJ4iwysPsC8SXYCzXS8Fw2gtZTOskLcDV+1B9Nzn1zTyNtlo6lNICRmmK
ZRVu2BmCc2G+fmzynYlNTnSa7C0Cuel6FYpxCBlOuk3OF2tzAmLAuDyOH3Z1Yjzk
a0aHuoCdIRKv7BrZCdALt03JeUmXKPdOmIlkVGFl8yw=
`protect rights_digest_method = "sha256"
`protect end_toolblock="Jn9CQpRhJt4rnzZPRk+dOpzAubz7omckX1MrFd4p81o="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 29952 )
`protect data_block
gD6l00tciPUa6pDNTk/+tzLxvdHE2s3DQL3/JqqujQBC/Ei+vcAB8wM3doqg5vTg
mdfn9XB1bLOis2CVSfu295W2DNwHfMSTc/8BhCDRnTlLIX0UCJs9Za0+LoM0rMrV
T7EjVWppbP+Em6PkVKCwlmIQ7JKaifJ+Y+kjw9HCGboYo5074hY+K/CBbfsBQY86
AyoN0MKhsIx+eViNgnWjA6Ug86McZMSpIF0jHpZ3bCsMp4slGTgDnnyiB0TnUVTJ
QfDPj5U4P3qOVEE4G23DJnF3L3ydSMZmM1ACSiV6nxvsw7In5ok3yM7KbEdDjBkx
ZwSHbwAdXQXKYgGNC4Z7FkA88tQOEUMRGnJ10U3+Kf9zGbfKhpjtUKVAqqVq9SVF
xFutfUk4fhITAAWoT51bFq1QBPdIqgaToxlFtn/OVHQTjvpGPffHYsW8MLeJUh02
CAvjeWagjVnzdOK+6416NjUCR6+7582aSm910lIkk279pfrCOf18/Q2LM7V2nzZb
KXsJnZiRVtAn/pv4nXkOmbUPEgz1URcM30IuH3hkmI60ubIO9RdJtLTDmsuvWWKq
0+eAoCxFgi91oFi6HWUjpzIsxDHhfZf7LrXauAnWplKQhMx4kqu+AtXX4+KkzFX2
HFZH74zV+92tSjDYlt/3fiN/6Bf3X8opM8O7xseKU86+px+CjwrDka0lXatk2b5C
UmBBdWZu5bmr1IgcXWWRtWaim6sjin9hgsq9qooYZ3IKtOgfFryedSIBOW3/01yy
Iip4rNakIgPxs1GN6b3W8DknPUhtTtNfJfRvomf90357fVLABReSvq4BvPi0D29D
OUKHtjHzp6ER6o1649KgmSfSwNEKPEOd+cNXtdtfdRHzRwWOUNFktFPt85dnwKCc
SZ1TPoYoU/JO3e0ctDO8qhX9VcAYoVx/wqYqOB68i42OpSPfzpxjlBWBxMwvkH1Y
0xO0ezKIuNK1jwghyyV/V9eRDXQnC6J80g1U4iEug+lsf0AB+q9XuI9D5i0aNj8u
waFbDhREzq2+/Sb3kcRcYBX5XkdEQ8Sqh75fK4Qac7CSLttY1q0kQMmOpP0j+ORy
uXhfi2eK0zX6cabkPhwrGrW2tljXOsw3OhCtKID/MVsHvww0tEAOLX6+QVOHcfAw
8tq6NntvubimU1OO8jtU4Odd9NHpNSwygDmp4uApGWF+3fi/dEDiBQvHOWbw2bvr
W23qkHhrP2uUeBvKUDgWpUy11oljtzZdBeK0JHnOKynIZASEFzAVJDq76vNkV3lg
Yu8DmxICb/Uc/Bwzjn3CEORmPSxDszuaNmeoxklKADBRwTYf+QcPX/csmVuGSa2S
t4KxSCzEGGoK5utLH9bq7KX3TmunRD/O3Z7V9tDszabsHqWw8ygfmPGtkho+hNqL
misd7/nNRqnxWhh2WtAu4nWV0cmHRs19InDdyS8e+frK1KInYWBs3B+a3jjlkTuy
UHKEDMZp3ufNU/AfbNDeG+3/yOYkNnInpPZOMak/KnfwpCGYInBMX3vjDzQ527Qj
O8axW63ukdTBUz/0WsSeVtgOE6bjWoqqMED8/TUJTDXii+ZDljF2E6ELFhcOfv/q
aRBPfVonr1S5LlzWDxPsdiUFg/1dLO4rMtxzUcTBcHVqWIaDUyttS6ae3mLSmzUO
Se4V7UNiwYg253UJbX7WEe75t06eGHbkz+UnjXpiEsTFbDvPFnFubC64mLaFJIfp
FlfYVrzrUrvnhOz2wrNjn2FRLTvF42hchNn61oPLP64us9XxyW7gYQ3TWwpX50kL
+pEuz2ibClcufAO5xWbNI9wbt3MizJgNnrMgJPjPYW2ZOwH192ibZfJTpB/v5NiQ
Hqm5hapPynwPjLXYuI1xrwbt1Of+sA9FBeGUcgUqmuyLrT6Vs0twwoOSvJxBPwdD
r4Pa+VDu3VF52kig0DTlge85q9yW/FRQuhwEbmPEHwq8pF/fRwzIzaLcHmwRGaIR
lzWTfa5fmx2ze+mysjNpl5y2S6wEURFFQ/PP03bY+hGQ7s6l+YtpiiP3noSAubQ7
BVghf4GtLkx3Z7kTxkIbCTSEtlJdBTCQ6RmRoKGUuQv2D/NamT3DuWWVyXL3tXr4
NJ92KcsbLC7ucHf3eV3ZIXo4/pwYdjpi0AXNtfiR4uhk+q27d6MUBCAcGKwO9VGO
Sq9N0blS9VI9k2kyHlterCPxqQS47SsdkcCimLHVCX62AIJHJHVj60ZEkjRd2bPB
yGxeiI6iGUVeKOmi6uAqoJgdOeG6+1N8Y2DakG1231QAbznDpXq+PIZgQBUgSzYe
SHVCJHyHAJ8ykqpNwA7tweIeAIsV61XV42NSlMdKWJchQOe05s12MH7CCZhFvN9Z
4BCe0CNSjaLpAUyHaNDXneOSd+m9UTlHxyqhoxdHje/waA4GK7wqllT0FpLDbVp5
0fHDHCftzJVCXBXtIgBJfiOGA6vV0Ho09nGz77iGDuBrUDbQSoMBGyiNbhK878er
IWFr6Rf7VqWi0vdEmlmGvlv81JQxjqkv16Hwr3XIIbigLyuXDaSctN2i0mIOIfF+
UL0Pt4L9Xg5UGmb3hbRixJuFh6a+abH+6Zv/GpO5RbWrMy4F1QKY3gzAM6LhqZl4
kljcvEEBZZCHotwNpU8xVsAVQsUlsQiJ4cqkts5voUfGtkCsl0b3OlRI/KxAgXKS
GHGGfBxhaV4Fugh5AMwTZ1oPjIehPARHWMkyPz6RdWAFTAvSycwMl4rcjROH00EC
r6lGEaGl8tcePa46aXwMd9adynu9VqiuNsJL54Boz0uPu0Efg2B4cEoPvUtaKkjh
vnud/peanejlfYfvH3TCvwGb8jlOv0tFH0LnsozvzpCpRdr4L9rJw5hB10YpFGSE
LXhrImdEvHkpgj75xH1p9W5vbd5Tl3b3hdPHWRXU30JD1xg4Sv+h4TB7PydjLcTU
5ZvcbmA4iruWxxtPkvR8YlHQs8qumXvO8qdxXlmEdTtBxJSlHZMbp0jPPf4Ond0g
OrsBdsoIwWIdiD/+001TK8YnCVd63gHD8lF+wpGLC5xH8j3P5GlKI1a9EM5y5k8P
57OitObN+IJ+O5X7WZrjlzU9bJ1qrnBjBEaWvMcsPfGCTdm/FzUu+glwRLUk96K2
XXNAo4mGvunnyxlhyC/2tbNnhXzJs9eDWXLbW2GK6GyEhTkakbWjm2+s4IKFK/90
crCe4E3wS6z7UH8WRkB8TmYUoE0/3Cg/PeSpO7yK37A6398J+q/UVajIWWmNIa93
EFp3PK40ovyPcB6RUdAxJhmPX3NHSjk98wHoKqBysdHdskoipzw3FR/MZhhenhwC
bpJsiPVA2N7J53v44a6tNTgN1EmMPxEj6wp/VmpyabOVgBerxv/4mB9t0y4X5lvh
vHusOm3Zw/+MSe9K2ujZa/U2xdnWQ7D+ljzb0ELzabbOEB9TS5y4fOYDUW/RzWjw
bUnbDSJNpXRK7K5U5GVEd+aak38cybpu9FdM+X2F6EX/A5NNrLCwT4p/83r5RJb/
PZ/0XQOEkAr91tPI5lBcJ50L7tsfgvomdui2xSABT88C3vNva5D/cw6RjB7/vArD
481oWqWZJZUDCe6OPqhKYLKqDzmGTIeERW5/h4FR9VbTkI1q3vcx8QlRJ3xG7DMp
Q2iVkgqZ7OuQOKcVOxTTVWT6UDcmhD6zzEvEWM75u/vjBGOLnuP6fOyXWHadILJl
wZHApZCVEadToduC6zwcwoS8IBXk2ML86FGbh7PlRfqNSFLLYMfjvAAcea+8p9Re
B1d6CRb4gAMV/K1gcaO/TiXwAaeV35l49XtQdsUIcEegFrKqUdhogRvUS68tTmQn
us6qYQl+P92rbX6bfeCzDPnri5zY0zjUCwcDZu3FD0gKbVfZdNTZPCLemxOidOJV
uUp990niFSTIZOs8v6+P22Mr1NwNcCC8CgoShKGjWpAgfrDb44mI3w9b2p0CuVzS
+0iU8KRpj0w46TFgfohDG3v0cIzJldIxvxPn6la6ZhunKQKGs5Mn9f5e08hXAxbL
NzMya78HPC9lHyKGm8WrixsjGWh3z9BiVcLm9ZftUBQ6XarByNVZ8hTRgVVT7lRr
q8ik0/2xa1O3oVHS7CqyzrW1M3/MuLLaxwNEWNW0UlE99NH2051BK1TECwTj08wU
Y3tNiiIUqb6moVxqZbihwFW6FhQEzDRRS6eSmFywp0CsSpLDbLyiSf7ifKwBoJiD
EIPUZ9FmggpvrwmpCynoJrlV9wFvw6Z2Pl/fNMIwHJvxZFw1aJruLWrOKUlVr9ai
gy0KC+z9NMNAWyX+hxrxeOKsTB/2JsD11Ly7rufQttbd5Ll20vlMjKQKlPWC2En6
q39bBS/jjToCH5ZW9AH909oAzMRcWvSSNxRAJYw//EPLGST8GwjKfa5MMN7xpxGy
pWVmTd3rqS2J79s0pStXOVRGZTypuxJxeMfp7ijRt+om0/WxyfZvAArG9YFxB/nE
lPO9CKzaCeWNJnu0OHbfaf/yET88Aptu5NXRot+K0o9TNvnbr+/AXYmA0Iyp/3Td
qVnAtxilzXaoX9E/mzqO0AYdCOwVa/D8rYIqqO8CsNme01StSiagVmu90mu77CyY
EJ7hOFRvc96oRpTXNlw2hq4MsOWmI+63UWU5uCNnCwmilfKHExngRgnsCPJ4gBRq
utF+A6tahZt7UCoBVHcg3sdcc8MQfcxtidEQoPYoBvTqH5c2eH4QdJyPIirNrfbA
WFppFMJYyH+vm7SvuuxwehkMO+bDREc6nux5GOnJMIsdIelw6471JxY40DoJNG4Z
w0s9scgvQvejTXURrqwHHfrrnhApwiPeqXEpKOu78aJIBiz3pt34iTfuAlPrp6mE
wgfxy0VBxFmUjS73XXLxh0wJJC+g2/hwVA+FzsdQOKxJcGA4yp7Fk1P5Q+lWLcY0
1XTIt63DshxmQjY/UjlBuuAszu7wjFeSqx2E2Twa4F45SWSj34wD4jpCCJxRFSau
gSXW1gWUEjbmJ7lGn8s23K/ga51vdysPgawB/sbJOt8RiAOF+xu9vMgmISLbwl83
ZvTWr471I15vpIZ7rWTKQdlFvUf61Q+fUxUEJYPhSdS+J5Xb8VIsEBl/LvBf76zH
k1+iVnMW03oSHN7G/hQRMQdOHFXkGWW33yXHr+GifC+iEytk1awWzr7aO9f5KcMD
GH4Zb8V4f1dBZVQMPyG++nd0Jb5yyBhbxdk3SAMojlyqz52hxTyIx/4JWZopshUa
22zrmQLqGSPnJ+MHaAqQwYnq6GsAehBVSzeKlknclfVY3/VTVZtjugLMwYLJlY3B
ur/sGPWi9yOxqUAcbQIwOB0oBKzugGI2OHcd/7Oz6FSTsYN0GCRPpHavTtonn8L5
TFgm+FOMSR739E3l8Ogc/wzX7m8fcsslzyj6ab2RGURVX2vUpyCj9r+d6eZCEdcy
JwF2Did/y1JFzKFI9gdEJa4P2bBLrn0eQcffonybDWJz+nwhxQhKhHPLFxwB8KLg
dqlXCKL/fqiWAwt31SskK1NfxzTs+aIZ+hM12RNgA27006FR2JcNQfNev/v1vhck
SHjxR1Pt8I3ldyHWtNrM60C/vdZEkLh5O9rN0jxqoLn6s/N98PuxB/XXNKtFq4Md
sdih/iRgo5+kzFWCh0VLUjEyuZzE1syEkB4iOiIcgZgiIImm+25BELMR9Hr7Fc08
hTJ1Ip2oSRp0VD+LdlepikAiJ3WsRsoCybTOBiP9M9Q3uRifQTJk78TIuPxkylJQ
EUe6aIbeWk5ctNuGB2d9vtHdvYa5u3KMNbKI1yz6w7NZ5wanbuFIYhIeHJai2v+b
AHnxSec+GDXDVSDnjrTFDB/9o3MTphl8m9cBFqQsURWzW7ba7YN9vCPPaqO0nDDc
BE+CThPRKs7WWnQec2OTHCHMdlSdYd0xqP7WWT2+rw3Rxr0OVpY7fTAbJqYP0NOn
akBwwoZljqH6zUMNAnpjg1GQEuh5LFN9oBPZDaDMK+/kU/6fM2hCbc5tKj2pZsh5
aRuIgn4pPNZwCSpbBNuBRi2vgPoO4AI3J9A6Dg8nz3b8InBhROQTGKVHphtphNBD
QXncziyPInRwKl7im5NZzhqfdB8a9uZ/M+PWZTZiuusx62zSm0c6Kh0ZUK82o43/
dt8NrBzgG7dRz2+JdjG39ZxQeLdNPZF73/1Ocph9dDea0ROc50xzNkwivdcJ0foY
ADmwzKb81edtuR/mtdNDzT6D332ZLOoMt5T/3u5PIGiGqzoVPdZuZx3YRdjsafYX
WQ+f3n9Yn17A/TQOrdIK6dlQOCCDzp0uULdV7J9cXYOk/dRhkTc0kG3Q+q+AuMBB
vfmVfIeHHFoALfEB7ivYRHiMGQskJti2QQPZhwrPBXR5NP99K9i+IP24rfLuPHq7
RC+SJyKnXL3+Ttft/dY3kUxGBRuiZM+s+mORyWF3VvcPuuYAofPKIH0qlhJbSCDQ
NmxdyXPHH6ibtzC9LpnePBxJ57gq+lV2bPOZ/LZtOjFHqq2MiRr4Gu9ST+z2hpUb
lmGBL40DpTBlBHqfPTVqqALTctqJQy5EWJIoMAFMfEz2TNnlTy17YmgsoHen6qGd
TmteCCBmg7EOWFXZEfhcIptcMcpPCcQL7IwGbQ6wdcdNenbwcu7CztoL9n/4dwzy
JWk/wbgsuBctpAIamp7G+6aroHnn6uTRsMdgC2S/E2p0Iajme88eX2VcKVceUbE0
FvQfgE9rHJ6KEfzLS4grIu3YrvNIvyPEaPT9D+1HIrCAjS+Y6CkAj2CXdrhToQVR
FkSOGttFGMfpdmNE+zUVry5sCUHCF28Uy4+CrRx4Z5UCvSEQ8dhooregCFnHPqmG
2hwhhb3lMlRncndZWptM1W/O1IFZaeooEZ30tzRRzofPZOEXiKRxMlb2XAHhvjd4
pw1kmtROjTW+XdvqZJxbmvtst2LnJPHMSS+iXvQmkopzkY09TtJrjTnrLNu78oBk
WOyGaXeqP4GJW6OasR6/iMQTPQR2PSfZbx8Z5DwnwYZuWOukfXAvY7ZA243g6QCj
X3j3Ck+SudspE4NfEpuUMKRNMDk4aho8EqWTT5dZ6iriEdSK9YECWUSUioeE6STE
YLEU+FgmvK2ddjUf/e7qxkwtTC1bIQLlwRHMSbJ+dXDDaJEGeWcZwlFiYF1mLLto
7RbrXzTqDkClVysGUSbNBQJnTP/Rezf5nSxM7f2KZCnpn1mB7XLqSor7PphNJLJI
TBp+XJdKd1TtdO8nVKUQiLI0ZLDCQ+gzwgOIVJ1+R+pNB7hCzivff2aWFmI2Rh+s
QeNYCwNGb453XP2qLLiSclI2JFapvfpAbvRJ0jQBQeQE0HouXkORjX16u3s/jgqZ
skBL6rnqINMZQx+nLgR9HaqQOmhOWlMSocsq3jPP8FG9GcLkCBnpT7iwWhx2aeIE
HEib3t42yG5MSKqTBS1OlSqgIVWjCFlezszQmrYXaV8I1WlDhQ2tszxd4P08GK83
VJ9pt1jWqxupqUatmu6k2tp/LmFqgF4ET/ZPVpO0Umgsz69Vf2lE3p1qU8FgI19r
Pio0Sd45WLIlVGlJ4ZLBmp3dk8iFdOmta32dK6Z936saZzuYBbnwjWSZzwhWMeP7
iD2DAsvPPRtdb3kHDgNOUsXRTIfLQ3UBNGXgF+wXqZy06QiNN6kb++JNwxK7adUd
uQd5QzrAE8p9J/5wXFIFzGowqPtnoEr7ny3HwMNKeYBtIzrIsEnUL2rHTWlheD5D
tLc8n89i9Wwlq19MEAZUA0NQx5RUmySXSjJ1eTTGqJ3DBkX+8jLAl6zHsVguMUya
m+/23vjcWInfXqbxz/cxR5zOEAE5uiodYNj8JUoifvyL3IEuZXDR6B1Utf+Ta1Yq
S7gW7iowTZkqdbOozXdb1LWBf3H0aqmDlrxp5dNaAWD1Gqb1lyKjjlvf4G4SR4iM
nRyp+lTaXYq1bx/vu+kdDPa7i1QC60K6iM8iwk6Pnt+lxY+/H6gXs4DKglOwkaSh
10qZERO6IoOOknnXpYwA7kXjtHlVWr/jlbU6GFlxxU/21Cp9swQLYQ63x4N7su9a
DRH1PnNlPnedjADF0H3CXsfk7GnsPBRyhv59cHlH9hkRQrwQ2ekTqlzqvsoTG1CY
TafkQwEmdlzkEHbRo0lsEUN3xQFWAj7l1J9P8Mwp5q0YqhPrZfW1A3vfDt4m9rrE
tHT6d9vLn4anY77NI3wCXpvhgzGn/JtETfU6ifQQuzoZzOkLbvDb11xkolHUb8xL
zU2QxXrXrnnukhKM77YzWddKma6NVKkf3Jj/Khzwz79RRyMy89BejEmHm2U7aK7Y
XIh61svI/eaL8msOmI8sChruiZ3YG4yCGiWT5bI3+CQRb943Vk49gkMSbEOABbTD
kYdAhoq28h6lmv+C7i3Ip/BoloPIE+Ml1ID1Sl0CZ2lUzW42fvqZn5JS3e79CR9N
y7x8Xm+TkQuLCkRJ9Qkbxd6gzCLTGnAKwzotky0ZHqBjsWw3k3WXrvgMqX39YuZ1
KqdAj42HfeRzfK0GMbUlZJe8U1mnVw8lVYJCSYFj85Xg/FfyhD61Spo+2AOOQCRq
xgZNF9LTQDpxvwHV+Owir9GL/5r3GLXyLQlqyQ8FmfQZCsUF0W3/UwRFAcBU16ti
c1EwZqOtLk8kU0T2KVQH7XuKd4/Du29b8m/JBMF5G6CDxMvN3CFsa26Tl9kdDh6B
aNQDTvzHjiTBxrEUxQMA7aUUcNK4xiNuhIOacEcpidfvCt1UQJx0EW0T7X1hLrA7
c5DdUcjo/j8hv8cs2a36f6OxvfrMEpQSI15Q46TSiy0yOpA3zN1a8/lx99LkmCCO
ZSC2x+SUo3Un3KRyl17udT1mVUs/kIJ4u64Qkxk2i94/P8dEAtJbyCxex0TChMqX
jYM6vlYv1IcFKe8cqdPaYGJkI1tMPnXMzWMpehUDkLS+muoT5Q4JoSV0m+pEgI5Z
o3mC0bFHtnYhT+B5YM0m3bwdFYAb7zz/JFxphYcw05olYZCX14m710JzhkHemrIn
grEf1Sj+u5v7eCHNw5GkVbMW1lZ/ufpDN+pRpfrXF/66QHt+91Wq7DDQKwrQCw6r
mUV86lCK6IKqgXFH/av44HLyPAED97uBbFwZDfdpxCl+o3ZtORFOImVortDxcP7u
MxR4gCkHJJNp8OUNkFRjJryR6r9jkKiciLRYH9XAv9yZLSVx2S51SeTINTeoDxyl
4Mf1RRdQowOlCj9lkCx3JYbCCRoM5Ub4mM4orrfEhX/iH8fO2VmnSO+0QTyouEbS
QFmRQu3gjQQwmnByoc88pD8NfyX7MI+3EAF6PrmkYEaBSRATlbpAkVLuo86WeoAv
+RDvjev6hiPDVC1vOGdkNccP5716lm+GulmxtydfuDu/p7kDcRCsqw8I4rYOd+4u
89VglnzC4kV+vW2xtzm3TLBQEKNhThDwCCfwK465CPieTgWkQSgUS6sgICj8QYwN
Y5+09Pu5njUe7hXp+s+rKWWvwNIspKWg0LTucjzWr8PUgVH/kj1a+U2rIpYsBIBO
bIMj8fUNFgCb4eOGXtYWbT9jEH3Seg61sS3U3cA53AnaPzXU+AeefC79gzl2lVTy
lA1g5iG3U7xzFurzOfPKZdtTfg+7kxZXZxvKpkq2DU/3Zq+I6i8c/Hcm2dLgonZ0
069QAiAoyQ60OrkT0ShR+tch8hl6Jha6JEB7aO7gwkG6sLYW9YrgHPFom9KI7WaN
UaYr9drN89Zfv+Fp+sGtRgs3nMBjsK8EY8yLv44F09BiC5NeWSHtm/duTyDLkf4L
izKzk2DW5gFIejeB5iFcGTIWXsrGzubcZk97TMmbDHiK9z+er7bTjRgCFkFDPtg7
nOEskemetFXIWy4Ufp7XF2FdUBl+uGjKgILd5yv4NOBOqq5F84FiT6G4trAPfFzR
cQ9HPaOE6ChaVayZTMPhxf4gvpx6gDQFbDsYCJMO+Bv28OvlcFq0/NWM4N5HhyCb
CMcHlO7QCWHV7RqIwxa8ShyRMRSte+Po/t+UPddu92KYVUQcIhtR6XDg2Pg5ykRv
jl4grZmLlzlO+2828PSMF7k+PaRuJQPKiMVYx9/kxuafJdYTG66cn35vkPHtd8E/
wj191qi/4dsAdVIoil8p1W4fu0y9pjTuzuLVbYRqKTXU/qH7JQ7cIkqs7luLj+EY
6Si5sQeI4BTWN6kVUPfk5vKiKFazKp/Sr+tXBcWCOGafJoQQ4w+ftp2Ddbn97xYh
soGyg5DWItCot+WS7CfDqjE/ZJ52uoyTiLetFjMtOrtXwp3illUbnebNx5RlVr6d
gA8VZVLmy3omaubdlicdKTMuoK0SqqEOUYTehI3BGXuhqXPZxQ/WG6p+pljRBvbl
gCGZoF5HCbiyCb7Is5Az5thbqgsTRiqxwj/rBwML95T87X8gvgcWG767wN3lfdks
w+brzV+0tN9F8bOM6z8VixOpXPEm5E1lPMoSTdz8sgrdn8binhC1Z4Xxy5q9t9xt
9+DopNTctYqSTmlOoB/RTwzucTLAQoyECXGSfV9JxI1KAmwwTrkdrefAqqxp6L9I
YmIYweK3/HdAMQ5RK2qWOvcfagoq0TS1e2Gx9Jd/Ln03kB46P9wybiP9b3Kjs1yM
0EQa0ppIuLsee8w6dufMo6rIX/sDnjuFk+5OpWwp2BG2GDRLNgI8dkM5afuoHdkj
+kiUzEVW44a+xgEaqJvG4PE4I6OMLks4zjIkvZ/DoiNgtn7Xp4F1ne6WvGm1hql6
AHnihgbOXeTXG95tn08hA4xYnTUx6O+/ycZbTa7gOvU1go6jomMwgnppMiECgfjX
ivYvTW7nifDeqaZNlm+YmD3g9k7TkXR0gxqeIp5ShGuK0yAaBBzh+R7JxYxXSIiC
wgITNjOdsVtBGI4ogK73sULhWVer64bILEM69J9mW3I5SODgcw0UPEQrCaCDVP54
vRFItqbu7OJar/WEK3nW6gt+BfGEVMNIAhGZbHa5jKyzJ7OUOAN2DCw1PoHtq7Ah
63lKgZ5rgq8BT/hWOwYXrOD3vosCV7LsYbkNj6r9Dh6t7fSs4SdoMr/WkXsSvwXq
MI/t4QivP8AjBB0VG0cEYaHCC55V7GvZsPEgfrv1ekc0XgxHQPeye3N8E2iy7QIt
+gzTNwbpdNIiPyLVz02u65EJxEkJAmc5YfkiZRyUR0REJT9kZpk7h2WG+mkSu5iO
vR32RqvnJztf++K7GZ5d2bGa8xftu8kTS6Sh/awwGB+s3G46dEiJbFcved9n75s7
vE4z6u0zZwHp2wxO30/20TyOpDrNtxjDE86XqKsbz7shE9d57kzIBepBBs87axB9
zKYe+UGgxCAbUcp3r0AVPoKtnx387YGligJmQfq7k6RNfDebWgxek3l8ulXQMvfZ
mXdSbnfU5JSVGDE5qfVgLQJ292SyjDh9gHNKYuaNB+3If5JxrtYgPzbOlouYK9TX
0MZJCtIAgMIIBWVfs6eVFCDe1tWGuaobrkwMSxvjrw69UwpiNwR0VanZ+D6Z7yQr
6eGuLQTNj7tYKRJVM/ncRnLjb2hkkIwJtmSs3ZQrVSEjI47u5Z6/oerXktJLz9ge
A7LHqzNmF4EYf4CGwn1ngEl9tFKovKvrUIyv2pepH71GigpHs1wUpQMASlRgSkK4
lLpuypmcgeQAeHIuChKxTFxdufaOOH6iRwesZhn68vdT+hal2rkXHVFIjTa402Mz
DisjrvmfQiC2ffDNXbR99nRgXhasuSNu7VLssPG5+xE5fWXpm7R98wCSxnikanWC
Sn4lQA1HOlzwMC6Hebg8+kehZ9PZyAmiJXL2AdWrLC5J+zoBVeDPEP5WLZnvcUPU
sfaArLSHyjZbe1k9V+GLjnDKU7bP8STJTPg/gb+3UNcAMjdgYaTRu2YzzR1S3irG
IlKheBideE/ZPGp9+MysaFMNEByTd769QL44tFzNeiS35eMLD8Zuc819z+ooW56e
F5eQ8HJ1z0w5BViOg6Lu8GNBHXE/hdkawcnYcDBvhINR7Yb2SVWEH/+yMFg0vw9U
SfrErUJlnLe6d4j9/z8MQ2n2rMaYBYWXQ3JTV3WNbTylSvC3bYGiUlvAzZLVn3l7
RamveP6HSIFUKw7hF2RO+Omb0EUJsugVR3x00RlcgaifAZc5L/42yaS+qF9M05uz
+ciSRbZ/t0KAzKVK59EdI+yauFTHUMU6ykc39HmGF5wW8zA5ZPBlDHpLvOttjNrb
29EKDNjurKwu1GfB3K8Iah+6k2TX1ImuqGPRyHX0RhQykKpMrraUCXV4nV1+BqFl
1VNCVyElviYAbuF2E0dERS8RoqeiHo7Llwv+qn5s1fl/F4zvntEUiabEMu9Xvr1M
GD0orX45zL1SUrE/T3n2Qr9S+a2CMANCyl4aJIU9tRkZ9aLL79bBJ5wI2ZFWQd/m
jKDnva5ft5IJW2WMx7GDUXB6q265NIX+m7Zoy0gXgKeRIhH/f85T+CNAgOv9/Mkn
qIw19gAIcVV8V80RvgEBEz5dcCJaw5KWR8hJ3JNMb67YXBm2hxcmB+IUUhOwvMaP
Tr5CtLPrLfolv3uRa4qHdqyBvpTw9UG6Ir4drZVFby/fh1ewRGluB2D2FT6/yhrt
Z18BrsaKUBo3ChEudJjqvF03T+U863rjd4B0GoDD1E2ovk2Hyzo9DtLZGZ0PlO0V
6ddDIgzuLJP/s0Tr7vlZ+OtM8iF+QTd55gD0v9I68F2/YESAfBwEYy8nRi7MXsjm
kxoPjzemLFUdVj9xtCbQ/gfaPigrDHucizxZNSp+neCx9WrzWTMvBO0/mf4ZP71R
6bN+bNY634Y1zSrgs8clClHDX4hLKEIrXxbAQLOjzfnuXMGDOGeO0FnQDhyafk3t
Va42XN0Sk/NCcblRiMryHB0fPZmepGb7qtyBHn5wd8C/BiUmiAJTL7wcMKBSHwOx
QNikTKKXgZG6JjF+pcNtO0CiTN7n4hZFDyWvvICRR5IWUMlzkNTPDXtCt1jEv9xe
98OUcqgDwzeaWggJ+oIVUkcHxUYk01V7i9UqrTXX8fzpzdJYSIKwv++CwuIc+WQj
4A6MaHCVzl8rqKSs9ZwZ4LqDJcbXBSG5tI1vyaGhVV6Tfs3Dq/6nwibGnwVRmRNV
LK2H3zKaHkf1xp3rsvtMkoAyqoPYdLnd835nMxQk3EqE+9hjob3PTGLTgZ5oth4p
bu64hMZ/lszInSYDBe0P/UhXNNwzIRUgL8ojHGJ4gQkckn+mVRY/e7tW4ZKnFh39
Cpw0KyTJ7JwdVv3d9kfF2ixdEONqSgU/xMvuzxDcttmUTrIJ6oRSLDTX56g6tERR
v5CMocyOtNBEb+qs9wgjH8YJcPJb9FwB+5w6aQ47OYYCdH1+VlNJk7c3PDmbMWuO
8NPSLOVWvWlGvcgDR5AjOzmeuXVFKCLRebv/oAYHKjkynh2NwMt0CK7zEUKSeXGo
ZR1N6+twD10V9UmU8TuEMg8Z6+ryo+BwNoPplbie3aT4Xur94Ke1J68YCS3R/pCM
Fy0v63qEkgB8l7iVefNBd0QqT2r/Ml/8ZO5do1TzQTE27cw54nKUXDANOP7LH2T4
XVfmLhpvmWWpj9IcyD4CVtYIV4i6M/lWI5b6E0uX7whxMjdpjFbC2BAvE2Lh8tE2
phlE95MCQVdBDzXwUO0o8DZGcZL2hPjGARB2UAu6higqxsPxU+TTy904q46+hezw
MzysJneFfeFbm3jJ0KZ2BpmoJmG0l6ZFnQXYRlK/57VcMItdNP/4XQvK1j4609ap
W27oPRER3N/PfHm+x95Sgf3GiHm/FenrOU2gcGfUNywuQv3MXqhOr1RpyBzHbca7
tw/Mi6aY1StfwC511igRfzq0fcenv+1WRh+svU8mma7VVnJGoUfNOD2+fjY86bxY
W057uWyxngJd362/iZRjwROXBeVHSvBsF0G9aznkbYmQnEsWXglR62Do2acHXoQT
FLBcQP8h0YL8J+fmJfkzNtuvVUe7rLpuZCsw2pTMY8V2H64GXLZXw8TAVlaxqCoN
ylTl5kNrXRhQIzRiDwlowih+X67H+x+dJ/lrrgrQXoiIAOLIAn0q37d2iAvMEDTY
xt8hCRjBoH3Tfi0sc7yANcZHoLsTcSSoYiyfsGDfj2SbPL3JT3kv9e7JaE3YRoIp
fZH5g8Vvu0mZYd83NhJZ+mfKEuSJc/MBtvDvRIwdLyZ8TqFADSWhzLXUCXBNmg3Q
tKMMnjR9nWp4SmwlH+lPM+cb+HPvmYOvw4lUcyCuvSf8uJpC6gJ3Ead87xKccSX4
6ii5QtrXF0VDOwB78z9SPUPo0wlkv81GuGloZMJofkGu0LwB1UjA37yKGa2jFPgW
gvK/nfm3WTKdVS5+Cg+4RIo0V1vWp7IstgHRCsjvDnuQ9jMzNjQMbs/WMrx/rlCv
9z0zE/zVodOEcw3xvgIsvlN+2ZI+POKVNwXgd/I8nuePxkVd30no2KMXbeMLg8yM
UcWILSyZZBDQCLHNmLkAAUiidv3doZw1SGg5hXu4vzm+iO3a5zEAwlpaKpomGIc5
Xvnw11KlTF3GNbSESo8XLHLZNN7ZAPlWx3VOog4zvUyuaxhqBsVMxjKrh8KJesuY
aOTOQstSFcHDeiXI84jbz3AjAMBK1+RggApEAA+/D0KTccIRxsKNBYNF9YDo1R3F
7KhOPVi7oduyxQ15erN1ZtPhBc5+1IOfwk4lH0VycbvG0R7czP8FmzCrN8qQgXbp
XePTSNaExTHPZOUS0XtIJL4Yo4yNZQfs2q4pKWDfLuW9msTc58QAfSjPIxBCs6c9
itCR0avH3/XbJung2DE/oa/9E83ir2NiMgikxNPAqw1AQTUc20AvJ7ecvVARmCZk
rRc6t93pWJVRfQ7/xpauJ14+BUsjJrvb9RlkChVdhD7Xc+/jhe9N0X9UO47S+U6s
pO7Bd68LHz6wy8JyXaRHSQPD8y/hlSn/gVP0a0IY77TiHdlfiD4xsHbd1yOavW11
gl9q4pYtFOixe/i6sNjGX71qeTPkZimifgrYgyjEgfm3MB2ax8RpRx1givaPbHsF
WQmUaQtHAVOrnvOXuR8IHJ3A61e/IlpF4Y+316Ll8mlCCMIg4lbfiCcBN4F4LjU3
65/+X+dwrrQDSkmA+9H87YSDgaCQTK4PJisYStLAChwHAi1O7Hju5wuoSz7n8ulb
/YP0thzF2eQY3viNXU4P1zOGS4uPkasfg55idRR92KmgGXh1GGsjIAmvADCTI5Ap
a+T+xWrujXlqYvgNtMApyGtUlaaWGJVRfMACMa900iYJ2PIo30wSQFu51+RCPX5H
xWLMjw6TOaob0ox3DuhuY+cqSvkV5DEkps2rP6I2LGFVlIgnfkMSPmLnHvD2x9ro
m1FroiHVX+5SxG/tnb9586OQ8dEn8ziS2FeBMluQfv64CPDWFCYSbyLKG0YWuUh4
eckVgG1p/jpcsM5PX+vXix+ulu3gYoNG1BzCbg+9YKG8Ue7iGuRVwKGKxIaK3YpN
uTmjPbKflBuTvY5B5gAf35KoT8b2alelx5l4ehNEBsSCxWQ94s4wxZwIVNCoz6v8
Ue6J0V9VWmnd3lpowgM6koVH/Z1RzbX+OMbWw/7r7qHN7uaeKwVdHH5psC0odcmF
AFh4m+nuq1huYfArW2Qt+H8XXRRG+FRIfdX/yX8qIoVe74G7jV2pcPFwcIda1VOZ
oEHuwc1AZRXwXBgjdCLyhY5U6u7C/tUxX2593tFXZ9Xybp0Ems5ONNjfP0gLqTuW
cAlklpXjlboOkgffVVVN7qa+MaVVMOBcJ0cnD7r+vIWDRGFY6cB3eOK1GwIByddR
uBaRvjJXdYuTsoUtwAmxVnJf9+88kPBDT0gtr+lAQJJAybKpsxt5AGRTp1Igamju
kBFIHFs5It+r13VWq0yVk9tYsUCgl+fZcau8hi/OwNqMxzUSBUjqIviVsrVEEHHD
FdkLhyRfBWeyJWtFNtg0Fw4TEHb8/LPhV+DcBW55rhIjaRIYqb5tHmebqr+Z/Ovg
SMT0lSHi62DLG9NDcSM1Q7Y8gjua3EE/c5AItSDzzvby9eqiijg7etKu5S5EaP4l
IiUp4TeQ6/+lDO7KwyZUwK3mrjrhoaswj4CudzTDO0MzZnbfbpyD/fPCRIAK0X/e
G3i653DgzGPeB9PYHxkyy0++MFRjrojW6p4jYUYURFlG0QRjjjMn6m341lbmL1kd
L/4ZJUnKbHAT5X8MABmB/q2Vg6hnzyqS7LUgYshqeU54m1m2LHdOP2c6YuRNaIb+
Wvn0FXWZhnOLXDfRrzjDX/sPQ2waT++w37O9BELNSAIjjp3tljIwDiNQ34BQMZ3H
1SYuIkhOxE7dfCOtdrsEe4qsNdNE8i4qLlKWDMmqXAlyE0Zf5ygF2Dxs0FGrEoXu
kQ24G56Sovr1jyAlQ6B3evGrgXcHLKolitLSxEnrFzASF84/44khdqVPXjxP8p/I
mpzGiuSb/WGaqi9KtlwhFXQ/j/KzTZJBgz0v6ALpe5tmmolfK5mNC+hpPsRpKjPH
/Srba/k3A718zZRp9OhXOXXwuoBkxa19nQQaGz5KzGT6X8b0p68oI430pvfVcJIM
cvASPSPg8yn/Ce3L2Z2jeTOLABYMVDnxVrZH75kYopJKVsO3wBDLU6avdNfTm5EK
5sroF3cOO9nPjjznOkPjHTL/o+8Ml54wBppEAqtrlUdPbKtjGlhqNzhzfY7bP/+5
M8V3miMhkNEL4YAJqFE6+mgzcuEvHH7MmD52IylZzhJJvK83wzdkzqeK2uXRXCWv
LectHoTO0cZ23y4+iis03npCwV1+VuEmII26QLVWxyTzSEzNzuzBhWb41lUoNKK1
czPi93sHstBXsWZbGA1ZO+/hEk9HYZLuQF/jLlao62QQNehegLAL6DTMxb8ColYK
Q6fNhMBrLDxUJ/IXrh0C2Equxk9hbky3pn4xq2ij9gelQAPlExMBiY8OxW8esHuL
6JcVje1aMp+K1Nplfr6bQBEr+PJws9cCiuDzxIvsNTkH+Bd72OKCljMZ5mcnpUSH
6LmkszdwpMxdFU7hKRHUSODGB8dQgxCt4YSKXk8LSrl6xhfuy8FmXQgJoHQnFKp9
hIwbDZJSqxFry5YJyBQW7yYPoT7pDrsl+60vGKUKivLXGmYxNQvvUPlJNkd8LYo8
ofWyoPyiCum/xJufVjgM0cc0Z0po3wQD2P2URhGNvlv5d2/95C3q4Y5ayN4U0CBU
VhYC/REyn7fYiU6EgX5GgN71TNIupMCnznstez6jf4KgdOQM4ul90uUmo65VftDi
4VJWIoqjoYEAb9paj32Z7jX8+dY6yHVnfB89lpG0y+j9NGf0M1bC8eqY15OWfuZE
j37nogAryvxnl8XU1xTsldyITzzcMbPEE2BECZwTHevPOot9/eBTkkFYPcB+Y+3E
g15VqU+K/5hDEmfpSWZ3+k+R/5pLvmHdpzdeWNhlUNuhthnzyxs0ngI2awj6mU+Q
VW2DMyB1qxlAfPXDrGc7OrcNpE7miVjBmommRlvFC0DNQXF1JbmpL18zugHDPMS8
wfaKbHT0+d3MpDSzWnot/xpvgkT5EgBStqxjgzFDj9+H9jaDr7gQYMlIhQdFcMJN
mHMQVQR5ARoWHMKSSwzLny0JectN+6Uss4ppuG7Vw8nkfZJP+OwCQ/rYHDS8+dPV
VV1Afb/homKeJCufHpXjiW9Y8zembh2DZw+g9ysgnAxTFVE2u1Va1klxlm8C7QBh
EtomvmEydTFMwsQQPpDl1DSkCgAH5N9VK1/8LIi0tLDc6vV5JhdfN9cxKP5p2xgO
FcQkBhqTUXnm8xlEWiG0tBqtWOypFdXoxaXG8BHXGyEtELgJDeq02UFi+tl654y8
F3ZgApw+IvFL13LOWlBWBF7Pqr4cgFskOc7eWibsqwrGQWOwHbKCS17sRwisnIhq
3DB0ExHe3tSMAFaluG82rnUuAeBSnqXPA0umPa2A+YBRTFFMp0WVYhSBDBBYrZpf
MexdshLH4Kn0LxeLXIVnsiHCKGdvDprVWB4jpQnyJUOVghzEPAaukd5pYJt0CDWt
yAKhVzHOSm7pgzjFtOHpvxEfKzR1kC797TIHZQD9nYH58k9qBNrtrtr/dY6YEWym
4IV7KndKmJZ2763IFjEW4KtvFbxV4q0gqX2Y08rbFJW+PNgGAtAPXYIWMev471l8
7DtheXAv8F2uKjZUk1QB3wKk6+JpDVPg0lpgRqC/OA4z7w6UqElwJlOjDAATXE7G
4I5WU6zdnrnEXVfYbMxpGNwxCN0hkjD61gXVCdyUvq3Exg027b+QOl7UR2XRU8hv
QVVM8zdKghUXoXxV/CjxR/b/PACwIi5YwwxMhqyeT8/ertHqWpYlHpgVRX7Ju/aB
miYwAlTMHes6xzFbiw9jYX+JSMjv6IKzNvImg5YXf0UK+sog3IS9lynvDaaDm5JN
6WuviBJF6m7zqHy2ieVGXsNIk9+hv+213BGIbZo1L8CgSy6BrsE6gbLccpfHALPb
GupB9Q98/MMwdTjbgjb9nTaEG8qSmiQ5RelD7y9MiS3r4mgOi6QMXF/hcvIqYllY
0X+wuYX7YNE5tbrAr829KMqBQqSpIchCV20xRoi7QmO6L0uO5CfZY3DLfNb4xCHR
YWnmd/MVrKaLNec/FiJQQJv+6zqzNfrzYdmmqvZLprRfCd+fv3VN9QZ9F3XD/oJu
s8fXWYEhNbUhktlseMy9PEKF82S3oicR+q0ee4S3J4yzeVI9K/3sypSOVZPcg7xc
iGeZsv6OsMv3uE3NYk6yHCqBNwvUPrvGgzO/hC8pWVHz3JbzNjWFYITS+XAswWwJ
rL5hohuOfL225k935ZCZQyG0CW4cDh+DQN4kL6TpLvLqUgFdUFEdn1jCNBr6pXtz
v6T/jLn5jWeLkIydSFgy/5WQowDuz9QNaC7lBUUaNk6cJoAmV8ZvSOLFUICan1Eu
LrOWl/4LF8BEwtBlRKSXqgT4iNTr7ltVPkeMeUT7fjX2af6seEI7R1lls0w6FU9E
R5OIPlDcWeuTNZt5b1NRajA7P14L2q8CaHWg4Ijxc8fkcfog67l2U4jG6YtNv6eG
fmpJdu/4FjvedGjLeZahIZI6e8HJ88ODmFF2azGG8P9ZJFoLLbhuQ+UaJY6hVTV5
zL6m65D/32Uw6QI9T1QMLjhBEMYjWu85gqfFcU6BmZMYsv5+V1bACrrbQxvywgEU
83kSMtYGeVF2fXYmUeBvVLAOsFUGQgensX1IXWVwh7QociDerl1sZaxNRIf9vKYn
UtB0B33jtFoZfmkVOgyNGAH0SimxJl4+Pe80QSfKLn3EM0gdb2Ic84HtCWuLKJvC
QStJPADIiCuBKyJH++Ak8EneCFMxKJhzMiCtKD6cdP2LfXKEC+2EikSCyEC4aaci
0Xi61VGPwE9X9XE8pxTBjCbN1usTLtD43koFLwTOFMZOo5oZD0GDsupKydooe+sT
bIabLkCSlZqyZqHXZOqIH+pm1Z+1aDAbXV5SrSMsdHgBidnyzOOtpw70gVMLZSa3
GI1iC1cXGVrLcUOcbbd2OfPBU/TapQDRE3SnFu6o+GH5e7SWP8T4UhrcGFPFw8Rr
WIt3D0SQmG39jLjcDC+wfz0itobRgTvl1AEFArOvRrnb7LJc0Dza36ysIg6h+JDD
vsAMqokK8QeE2XQdQPak+fBsQjq84DOxdvBUdEaeKW1pMqqnkjPtO8qJqYKCCe4d
NV5K+QxZYEJNUSTnpOY/ugsjb2TPd61ILeiZ4vzU+DP/ZEVGdq1mEB8F+Oe/gwB2
gOHPY/xX147rDTFU4QtGplomMn6uAkXXZ2X3mQPCouivWGbE+Uosecb1/aGovqfj
W3aQsXzHUllY1JK0+xhPA/CG890T8c3vXDW9fUpOwQnOwqy9BxfU7yoUqJmolbo8
7YjLcUTelBN5wF6DmFA5VkLO8bisbGIGH9UJOaGgqipaaPGpaK6cwt3P/yIc+WxR
3nbj874thZ9vsYfDHhOx6aQ5NO+AVCVc8jBg5ZjnGKqzgeNx7z9E7AACrUY1qBMp
uLxH2yMP1NgCIi72U7+JtKqqWEt06jbzAqAqF9vRGSNi3szeH7Ei8uU7VrLghjKq
fiV9B/YLrX6nY36uOir5YRJ/PMzxZtZJSQCRbVsyWUyxEsA+Y0WDq/xezK2BxmrO
ofkKMWBmjbCX6YvTK6jSKTo4s2oZGz28f108J4MmiqwQMaXl8rHKznyy2sHF/qAB
0eid1SLG0djTugoZXOFPCrqPLHnh3LjTO/F6Xyi33U+1D1PJkGPdbkU58gWLydDQ
C1RVNkFL4ulg76Fl0D12PTZD+u9zjep2+VI6lMwEz2m4XJwVnCXgU15f7WculrxD
Fnm+yYpkFvO7t1ms+TjHYksKSPjqkHpn20NBFq87pdACGDNO+jAS/LDffkxmaH35
UgrYZa3Ncx97po/F1CNnRgDerLoMbSmmAMCWykpkxhStAHyXGnIzPFz1TJgADsLr
hUsfpmdgwLOOgAHeKVOoJ1q+b1THQwwSP8/0NYEhqfu0TfMWgw5+mhpzOtjq9Atb
EKDtgvFP0Bt9QxGPuucDoFajGogRmcjls2WQiDCnzAHLVM8xR66LPPo0OlPKG6as
0qf2PCtiAvolPPXRj3ftpzKh2OfH0bYeXMiYScAV+XqsWCwEEVJC3HFK7Q8l9Dzl
YyK3o6HGke4+SfaOnLjMd30Y9sb0KWmBG1HCFcymcOubhE5u03qSXvGHNnZfaPyh
0qlm5PyuxicjD5t4ddgAa4S8UOAUCG7vUbrhaooJmnJoknaU4vP2HSl3JwzEOnDW
sDG5NE0tUfzbejlfi4V89iGaVcsqYlp6XMEgVgyHzveDzle8u+tP5Kjog+bzS0Ax
OMt/+tOCB6zS5+T8SSpszvmie/G+M1+5CRp/N8Gzwex+AJIeZqcKEja8Kg6xuuJs
Zf/HCKkbJNJmX4ryEzvMXBfWjWKofFmtC9bQFZQIwPjO2/kTuwf6QHyJJeXizo22
BMvlIYvGoyGfrh+0UvLePANlZ5j1qshPR3aVaSiFY3bElgO78Y2OKsKQtHNokqat
6EnC8f+ntAwQsGCbLTc+Y0apj9p6RQA0N2R++l6rPneQz9E42wqnvMxu1B5NGC5y
3CdQz8UHWzw2ze6RAJx0lAc81TgOU2I0TunpgK6+pWonxJeBkdmT9L9jneO1NfPL
/encfZV71I90ZxEkHSAPGPhJgwkxYEkK4h1axgvKYmFO5eWyTeYWqHMRxk7/GQJV
Md0ESjk6xlDtM7JsKqGs4Mr/+nQx+T/KX1jRGO3Evin2XD00Ruw/va1I3CdmbYeW
JABbrFIf8BdTMaTOvs38JBveT0gwI2abn8rkhNiQjvfU69WVhgaEbTQZXIG0QjIc
tBQ2QdjRz8pJwyEjRiX7jrxLXQVurlJ6DhX8bGFIRXnOWe/53hw+7GnL6Eo+gyNV
5tKn8hJ9cOI3mOZ4QZoOZb4U47Wt1p47nmh5Ub4ZTmv9ukpdg1Wi5iAsPsaeT2i8
C7Zob3rBa1vfyPNx1fN6j5utrJmlQpvgGgO1O6lepa2It88dCZry3M46GVY/rR1T
JeqzzV4YpiYcCh9bn2WGlymf+Y0Sg98HyO3ERs01G0f3dWmJHInUq9HNcqBlySAo
wbe3/STuZ2D2Dt1LmdmX2lC96lytYrJSoY9POf+pFsUbk6aJHdzjNXqFN/IExPQS
cxY8H9v6pa1bzxTjG0d/9BOJwWd45zfJM0wP295+Jg6jOkagvqMcjVrPFegcuOnN
mjPK8bdrLUmWr14YmjAMfyOM9JGNnMYCuYTLkVfKhOMsPGshTdPQ259clwtkgjx4
KhUgTrB994oDzhWGAuXMiCv0Kgu1r11/6TSxkn6jVM0bOnH/uwCAPK/HnYfOhSdF
7z+LL645O0ql3KrCq6qilJJdk+MrJJ8pvV8lhRGiOUioeQOuy3mPNIkk9EoSozn1
10chmgRwvscS4xkho7JSKyA9Uzi5sa5/z276pw4uiDkUH5IlNobpyHdTx3xIcYji
OvQ3MxyaEhQKfpCvRqE0Yb20VyCFNA8uuH/ui4Mqws8Y/pCpBRmMAJTmgXRgJ7+3
IF2ea/rLktHluhaekK9+K9sWISQF3Eqk5TBBbUrHMJ+tomxEpp1zW/hniynhs6Kk
qmVTra35wlQDwuI4FWW0R2PLkVZuVmG4gCala+yCDn3xZM0k+NRZCU/ATtu6FwAA
g0CIIhgZszJK6qeNpQHsM0xGb19M1V57LWxSyU+3I20Ot5MmZvY3ayVALZFcOLfE
zewf+skBeBi5ceqOsRF6Xmse4mz/BSa76HoTyTHau1XIIBKKrE+OMFlsvoyPUTn2
cdiz4uFdSkCJxTR9BBjsJa45PYipVz4XeLnNCaix5a7KToCPZOby+K8mOuKouay4
kbJF/n49XshYrFcksLiPVKTmQeDdHoRlcVYpiqKpRi0+PoZJ+5s9MCE/zkEGTq0E
ZipgKY7WrGOMsnsIfeIlCDTPzFLl5oy0XK4pPKC845dzUbC2XEdkS2bH8TsTJlHy
oaiBlilRodyvpfoitrv0mFMniip8gizYgoxmw2gtf0GeqOKvJLMEFhekrgIkFLpV
+MNEoRVssHhT1waw8hsJdCOV01aszYp2wWXI3jrZqkafq0ZNiOJPuB6D2/HdEtXv
OwmhjqyRZouD/NNH/kKCwlOdDk14Yd+0WTvxSC5ONVfsr8gpyLbhS1CIrTwcA043
gmBvo0lKt3nAdHIei6lcPQfbdOZeu4YE9o8j7Cx4XEDgYGVy/A1OCU1ojLZnYN9B
jS8Af4lxO7fVEP+/J8FOicu1GlmFZeUR/VkFHrs9s3S65LO2kr6mscrajO2BMQn6
B/nUZb3Uj9dZK/5uJ2umlK3JsVLN43e71wCkMlg8cm4BjJnoUJO9azZTwicz/8Nf
qXsNAd0QzWcezyzgZ1JAGjdz+DAMHH91QUpOa6s5AMGpKq2LzhzV6/wkvirSQb7J
nrTMm6yNnr7hTksqGXsDXt2XRRuOGaax5sL2eRAN8kBaDyjV3WRwtFVmYTdn2lOG
JfN5rCx1znxSke/K+TBjZDGemSKDti6mfmPgyqKNl8uN4QVSm1x8jpMRLc5lRyPY
uBFE3B532Pgqoy67abm0gQgNLI9GNyHOdQ8LLg7IUYJGelTeoktcgYEBXp8unP5H
Fr2cAw3YiCKN0zLV7sIE4nhCthU0Q6YwIUrCJr8bLF8TeT5E17L2/lupTl34FuU4
8gXzNK67b+wk0ZbTELEw12xj6g8tbuOADgOHNtcpn0csy08KOMx5EfOV3V5pAyBR
hwB0vaZ88b5DBecDZsCNCq/zZfI7gzPm/vZlg8BYenk4PbhB+QjnmXrhf2m+RXIl
RFBnTXqNJGxSIpD9L8baDDBmZsBWS2Jp/Q6DElZVohHPo7itFdIrT6rcpJ3h7zEf
/4MO7/gmNdvAy0Ab6ndXBPkaQPrH+Unuw3i/9VsQQ7F9lX6mVuzN2gpm0g5kWfFu
El9Zqy0MIV2JYocyUVaWXVm2uzReoJUOPm/18AHJItH+DRB4ym9cB7efxjcYd/18
Gow8Mxw6Z6tunlvLEM1Q6KXZNLHbLtapmPPoLku7D4+aazhhX5OfZCHH09qcIgz5
9Pa7guyhCqbQQWq1OZOam/NmknXmbg1X+4TzrKIB0486lU+F4tG80pZaUghgcA2k
bIPTV3xrUzNDM2q0TgLjrQPftLwW+E11xkdemoTDhoJk+Ibecyq34i9Dzui0nlmr
TnmEavdRjGFHXtEaB4qOd20ImBYMhgm0WbHM81y+uSg2Eq7lA1kcbPC5f6MQoNkH
7H9lcldL/UeWt5/P5HahqMklWbfqOUu+gcrO/Y5LI/Wg0eO45u8T9cw/cLJzD5G7
Q/guBjhIcxDERdYJF+45dtGrmVycBe4CcdrS6Vk39bbjzByccpwWFO9I1w2uyN5K
4eTx8JRqpt2aPEr3+MnOC3dRn9U3MFsPYiNrKMOFWp7avcyNNs3rTIag9yKywOG1
topgcvvVgVE5NWWwnQze1LrmnUpiEeiHIw6N0dhu8pe7VdqZyhegBvuhCHPs2ae4
8Ci/Qfmgoxa64GwWME7GKbrzsLWUVqx2vGUPD2A94iSEI4Q+q2tP3If2g1YfqUTI
aPtwFJR/9tVSRrGDhV2SNKoaskxmNxtlGsFABceq38BxX/+Sfp/gF9skV+DPYCnt
2SJIf2wJlXnY1zBQQdUrWtksuX57AAzQc1qOh8Kz6rJqp7HtuSDQeYoNtRDHAasK
n5jOYD+P1N7l/4pwqPaSGR+dWuuNqx7bSV9Ys8J7fvY4ictycrPhg7UYIfEuQmFQ
zJeXDuN3u9HCYfUZS+4/HUHp20K+aHOG7n9Wpj6601qOcrU3suJBae1MEaIVBDYP
r+CenStF7cgKJ0xpqWfKVIQXeSRfNlsqNK1r4Gar+fjAkTOrm9SANgbaIOnOCQU8
wfStMSgn6L/kfKVHa+oPedBjtumROTOvSTKExeG3oj95NOk+6C7T6zOSpcBgC0hK
2UakYgSAOrMvks2apZ6HhKMYEYgBrHsfGARDAysybyJ9mWVVpwcyR/ItUMcaqNWE
mtlbNpKPH9fzpUyXQD+TYuaY9IYbxw1OdQyPb5aEDNsVMNo9QK33ilE81TJCxwsq
cR/5TSkwtUbCt7HsACqxV5Le8dmgR8GiFiuLN97fqWLbPJs1W+0T0GHjxoWFUuTy
y2BzhGZfb8Dx8Sm5M4oK+go5H8JGHxluQVyeCkVQhN8KCtXm/UCQG9wYPpghvBTj
MQRxZYh8RHDjBug0m/vIhGK3b8hLj+rjQ8qRgAW4fFAuzcWh8Ka+zEP611/OMJT9
8im3mihQ3ZfFGaRndqQzJiCe7mmmeoOiHN7EtUjJZ2jeVF8QBJgDeK8++xucBDS2
FdYyXCCEXPb6M+ekx9W+1/5he5JYgZk1uQAMPFj+fSv42pt+RgIwA1sdoOPwGwhy
lTLrmceBPXERVWEPLILxihM019vEY/2zXCghrgK6orNYCurASRX0VDpSUn9bvrEG
NdnI/iP+6Q1ugUoBJ0SXPUXbt7C3g5lZy04L/NdUdJ98QLVl2dkF4nmYdHpftCzB
jSvmmmdZVAkr3qCRKGYTOlt+AkNIAw8ncHsmJtDjRmlgj1bbYgdOULg04w8V9sIK
YApC4pOSpWmomELhmnFn6sNWqcFsy2ygYdeulonYgGrg8Pha2DjMJjLwM0kewDnB
ii8kHMC7i5OjYs/MWYlmp0jENXBuwKqc2BCYilYJj2WFIkc975vioB7lEmvuw4HS
9JhPAS7GH+nNQc9b8QrGaZ+DNvemwrELkz/oWsNn5HJ99S8l2Nm6UE0CbhceiFQ9
cfbjb/tu9NTVGWS/H4ApDmhHFG+zrIyQ4ta3RXTFw+zbKcKh6oRQQSstJHGUmBmQ
tNUxMwF3QbdLBljlxpgMAhYBwFrLU01qEFiKXVvjHg1ZRWYyqXc4kw4NEFlmQLmD
3/y6N9sNRr/h4CxHzy9+CuPUrElCWoDLwBqrcwEh9SK3LJSt6UoD38ULiorAzULy
wB+fqFHWfLkLtu5jwOpreSBwc7SqFHDV3k/nqYYaW4daL0dBpmdbQuG9BdeOqrEq
iqcmgX+pFPPFT37BdxlQirgetBp4R4XULKwcCna28qbnBSOS8sQDNP0gdv5OfEw7
dTkk8QQwpFFdyhoW/CG55UyIvlsuKYjgW+EjqlVbvLFBRjlrMXHPN8vR+xeA1oeP
g288Tp5mYFSPoyOcsyQ0l2XFlvob4bD2oSJIanleWA1BQ1gAjCxSgv6GUof9dnVh
SokBxUsiojHq3qBdYeObdB6g5/tkIoYMe5a0O3ZW0cbxpfCmFxoI6jSNlYci0MX5
IGEgh0yFuV2rxsgGjY0/jryi7LrvO7I7PHZ4IomBl4iA7JY/sggh7aO8SBXyhls/
lwgNw2ytkVJh0W4wODQtudh0MMRL09oYO1bUbPYyEmaue0y+Lw2BgGMeNUxd4Whk
Rxnqsm7F5V0WtKWL8YKa50v51AReoOY60NbnhjV6sx/WQttIja57c4kwSBsQt+zE
AtJNRlaxz6pq194VtW5frDhdeRs5PWFeoUeSh/lmwaAdiydebfmUUL/hchGqcXti
dXf9FDnvH+ksUjli1eXRKNmuHEI7ZeHKRuFd1hmPZj85xhnXIBFvKmHpPlK8Akq4
7gDFsBlAZH+bQfRABCsu3lcvnF6OGXq/5wDd4XBGNYeW9kGoIDCj7TlH6GjfQzvf
7tPS6DlQ/292GV4SF+lD26DtGwzI9smCAhrB/nJAhj2wan79ZioqMtdDEzvC0qDa
rdD8OM9gIAQKFwWZWA826S6jFdXXxum5W/bokQvWzyAgMFqv+xcDZOADVj49L8EX
WCK8TxP0YpC3bRmPenhHgVC046+J/RZX+UFrtJkD4DGEJkWPS6wuHdkFqKb4xwnx
Yt0wb/OXyUAEjVvVBaBVSuD1TlpoEn08pLrFY0n8eK8R7Cy3+Gwp+Y2A3qecr7L3
B8VmFrB3pbkTlqDdsuuUB9ESdM78yhSFOPgsnkaiW6viiqi8VR6RH2f+HovWg/NP
sHBnJY/gJf+z1R+aFx+hm2jBIZDaiynC+KZrBKym9xdXO2dcVNWp5vLFF9wYk+EX
ixqvMe/MCSZQrSxFtPxpo5bEpogb2+2h8ryFuIQu4yH42YOtLi7Jn9+EwhdSX3Cw
Su3VvK1b1px317hno/7ug6g0/+9V0IySf4387B5tUGsgcVFDtB6aEvj2ywDaYh21
pihg6lvkz+XCnl2Sfue9MaOuk9TqjBodmNz21rKsEusezGhbbj7pKwQysV28p3Sh
l7aIcCwhpLFid1X6+tkXfpXms0bg3CL2SGjUx61z4c1K0A5AKVbDOWQToNEXXfVg
EodimE0sm64wq9QFBH+0YPhG9b5SBndqgF2jSrR/I5uuH9fkpH4nESUW4/9BRJQP
ETOjS5AEovSbUR3TaF3r8DxfItC8SU+GDfcTGW77ebUdeK7Pv1HUS6dVXxAwCwm/
kSjvdeICp+NXu2c5Lu97BSHsJmSxwI3RarXE0suD7SO604JEghflUpyuYJ1QQ6+P
O6FjcTYcEhE1uaRNjL7ksVYr2C005yUOhH8Z9QmLkncy6IbaK0r8q+pfeU/N9ekg
3Jc0YXyOrJkT1BAUqVH9GPJv/BoGjeF4dYhlwyM8M/rUfUhv+RWPuQqo8m4jKOL2
Owi5H9Z6erXZFQGTh9/Y8JFOFUDIiwg88EbPw2QZwx0bFgqFczmHkMCJRx/IctxF
mymcZ+G467Wbj8+hNEXKmu3jBzU74BreHtMytrAYPsxJ7vtRuahmypGR7BxrLcb6
+rOjbwgeUpofHMRwJiJSE6bcB+CUinn6QPSZ9H/Gfjiwku9YIGOTiUigYnMpKxPq
ITWrzsOj+MvTtoF7qjzbRv2wqT0m72bh273NH2c+1uxZrK+vpaMz4iws17mwhtD1
p40GYUX4t+9hTUL2puM3SBWcVIsr8ahZSBiD/tvI3OEQqtmlai6HNsmWR4Zln/lD
j+nylChQ2VRTvL4TYSuAAYhy7JwtnPO/fnWLAd8Soh+aphXTI4n6khSRSpXUlMIq
TxD9K/YY2M0JEOwZWzEJlixtnME/oGmyuV0Gf+IO5jGjzBzvGMZx89csc0LcekGs
S2uCZRZz8hGApk3aCN52KE4iicQrDNMp/7EX8MABAandE5mPf+dmH2mNFy6Hc3TA
HNtUUabvr0ut/R3yl+8Q38DovNf9GDLSlQJQr++rfgSOf5wgMMKS2tRBbXPx7jrw
Bn3Og3NEq678oQHV31Ve4T6UsC5n1AGWC6V4NppHVhUOz8JkABDcWQ7ClSDZ9hTg
Eu/p8ZfFrH+SwlzAmIas4r9hgKCdTYtl0ym6ThrScVBw6WMJEZLWrnv5+gLvLgf+
fAEzDRIIBmq/2j++6wiG1AS5CCg12Phi56vBrQDSlO6TJ5YccQEZ8T17krQgeEuw
bKubYwSp9ZhSk3e16uW+VBA+Or6lIdOncB2p9wAiLCAqg4ZQVrAMBF4A6PLsJ0AF
yKaLkXusZu4HkkcJ9OEgz9FN9BVv/htRR3nVWGAEYxog8fmWr/6drZLju5ga+8cA
zf/O+HdjVq0DNxaHot2+PC8FWD5TAPyI9eGR6fp03zpJqHGUE6rRR8XCjZ+4K6XB
6vHWtldwAuw9rrNgv2BXNhc0WO1pdeIdcXvE1kdMCPFKYZA9+ogfNJS3oUQORd2A
o7mHHYYVd4oeqwN+lflgkUPzWzR8XB8Rnaa/3391Ncg1Pg5Z4kiiMfLu5aaZxPRu
RIboStKhhAMkRsvgWJIFKx+OVg5UrXKyJ9J4IKBWno1fn0NpOCYpUVcbunwwEFfT
5lyVGIW/zJnpKryndm11b2uygxrbpA9Df44C2VReJIbRZd2SfvngXUa26uGT50Tv
sDaFPG3Ra16ZcbGJXqik3LdwJgpv8Cpc8CN5NJPvkE08RyxZ7okRdVFeetDCMMoT
SunwoVojg/Chy9lVf7ht0NlwYlCsPg0DAb11IA/cUQrE3r6kA/OIQWbG6WgAUvo1
O+D+e1M9Ks6LAawJaM59CfxH6x/A0b7Xuj/Pog+qNymBw+fi+TJF5qlgdQQsJImP
zZu8F/eaUrdoK3/92usmHy7ysWEXqROfEhoSanFz3Whh4bJ6M7O6cDesxoJc8/qn
WTmFrfpJIQn719QM2ChEcW5eXwlOToiAPCQSKL8FsJwCfb7B4RV42Vb1Ur5O0Ec5
EMIsjw7kS5XPdfOJnpB4ksZksJW1SiMmwekP1vQxlsj5SKr0FS9MpOPyw7DhUzXz
TkO3XChZXcp5y24w+I5N1X5W64ASeFW8Hj+3lIve3zF83bt3r1ZoLBW6j+lYEbvS
D/fa1luiUfsxrjubgn/ZgZ9GBhWnKz1v0UVJp5st1nHSyNApfHAsEjADYVSo+9/l
f1UYTa57guuXwJ0JL5+yLbHlCSl8ia1aHxinzyc8iCNKvfdVIOs8KlZ/U+Lmq7rG
aEa8fSNAVP8tkviIF7KPVw4hV2ttqVbAGB4aYfXtXqd6lfFDBtJz09epD6GlVr6H
EhXNT9ZFRigqZOUs18qlW2e8UNiMzuS2ao3R2ox/kswG95mUjUXvaXMYoWL0rWDQ
hnMIsPPYvDJvvPWIyaNCHp8d7kkhOfNN6MnhYR8DoKUSiFVcKbiJKMFr0C6gKyFB
rrPfz0SBx2k9eHK16XVkccIlFQmc0bUfKFyTgi4AaG7vsWTGnL/BbOFDWTyVFKIm
PL82uozED8+3yDIniIfsLGEmM1LUDiozF8cowZgdf6kEDQgqjkQIxn/sHj2RjPaC
TED2ZYXBhs00pCCWG8cBSm1ANzK4PwD5dizLh08vF4jWpZ8ilxH0vuK/egRTyTE+
RICDFu0waPwiTTvY0W6PapfWiPpF2vdePKZZlYhJct9FdpBbqxPVysQGhgMR/wMY
24Z268tagPfKW6UUkS96PQGYCdSsU2H2qeqJVbAgkmL2nIBbe7fxravkxhsiERMX
8nAtLirAXda88z50zj49Et0O9aSeBJiOMo6u4N2Q0n9o928kMLaIe3Gyy6WIEd9+
eIiCPQOSbpqWP+7spnWg3fHzW9Tzlq+RsaORMpa1IzYYMNDLocOKOk473Q+MQjTw
/SqVEIYsNNcZg4jxrw/GoheRi+xfv8oPNY6lLdaVK0qs0x9rdwySStUCq7LqbEVF
BINfYFe9Oct4D5jFuV41m52t3kskGC+XT5e/J1bAhjce9gTmnoP61BPUEXJTIlk8
rd5upWvI3N2CbHpz/KZiAMTLZ1FcI6kxU8e9ek7AEgWzJt9X4fksigWLtbYfoimr
pF3UEvzD6a8AIUbLS3/+fAVJqHAUN3dMK73gPWEK3bJyQA5Ti13H+BODQCGc4RNT
to0W2oM7ZkKrEhaFvD+vohleHl/uDqz7iBVRaSy7XJ9JfUD0Ahr8U7whtV/RJpjR
yXW4p1jmYgmqeK1684npyE1NfbtH0RiRxW0rVBmch1i/EmcTYBlVKc88PtxrcZia
SFpDy1fQ0PJBKwxmO/9VHoEiqNulypjljmMPRa8hfYc416wBZbKgWrKWlsWg+Hme
J0g07Fiu/7T0WLZWuCDVRbE0waBK01eoDlQf74uloDKd2JOm0zInuEwL5rzJ3gcU
2UHOEFEL2dbBLOmSB5h4tpw+5Fb/hMTscFjbgyyRRkOtNZOzS1j+CCS14Le+Lv6o
quWi7J0VYbaP7/c7OmJzum7JG7LMyHGc3p2eg01pBKrUdQ9MT7M/jJmvNHcj89aK
oqv828lTCmFsKoQ87j/bCGadXfcU8z+TdzPmnrtz2zfiKY9Eow4lquI+3NyeWlgx
nW/jusP40b7T39GX6CpzYPqPq/itLCwJwCOrSz32pBuZa3B++yoinXqZTSHKnGp4
IBY/+KY813TYeU2i4NL3ZH79bWN1KZq6hEqJsW2QnJKAR5pEKUvSysT9v/XnEG7E
y4mjSWBoajBak+P2NrPpdU2c6zroKJNbW9s3gFy2zuUxHhkQ4uOPVRU/J48Lznap
99MO+z9T9NlaVRxjJm77VbSu4HwgFf80zAm68/3C+NQK/evG2Ph3vQ2amUUHflIg
di4rScg2ddR0Hbw0/hzE6i6L07XxP4ek0aT7vdtUv4OMsEvcbE9J8rBclZxLWSsw
1k60Lrw0D/g9iSEIEFM83mZOOf1QGo+B7qdGBvabX9wAUP7vBPU3+aRTwheIKPCI
cDhEuVpXrfBwhBsNtUKSBU0KK0mPKP3X0SH3tsGcQXqPc0pJx2ird6OsDWHK2C6R
8jrLJeM/JLtjY4Hw1z/fhfhmLdr8z0nWozJnIq3QdIYAq1jbhgQNc3KMVc0pNeYK
T/kzXSfJQ2rsrMJ8Sd4n1YJbUF4b7jOPgDF6YL8LKb4dN3FjnpEh3C6UKKBSmfbq
bgTNH2kB2imlpx0dzdH6j5rr1qYwxyDQ6QALiZr9jEbhzDyGpOOHrx+JEwgm4Z1H
LtiQgaBJ69k4k9T2HPBDPgQFmXYkfisTWZWFuVmHVipftHPHMBPBZovNRZSSy7LE
JkHQCLhYIkUa9feEsGc/A1ZmIqbWYNDEJtOkiXI0tn9Im3YUfg5DQIQMiC5aHAMz
lYchH2HOokVMz84g6bmHYGopM1EP6yAMeZWsx+LwiFbkyFgNOK1+lN3OKY9PL1tJ
t+V0682lr3GgBbq2di6TvYuIjm0Mc2GF6OHTw906PnYJE5McHOfNjUJ8iRYuR/f9
MmUPGUD9btEFXH4bQcduuMPlpIhoEWdfL46rHAslWnjC2zzeZKQdGrvpuEUMp1Ez
h/AauM78qe3NyM9s/OsblLgezl1/HpPNMrIzJ9JGu69fL5fF7UIHNuvxDkcaGxJk
D2oBNvPcOVzCgausKussjNyPezJ/5dVNUDAG7ThBJWiYHOWVjRjpAxBhwOFYAXtX
VazwLVQ6CJ/g7FNLz3KyTKpXoISnpV6ZcLQ/Y2w+Xa/FKk1zILO40/EGjvZpQRTl
B7STDeTgTo2Ds277bo9mF2kNVHHiX6Yc1gsK1fDl3fews5CzWI3JjEMh0/1xMje6
K5fZvYUHyzC0XUGp9qy4KrgeOK8rQl9kGjgksR6+8RXbXHk3wxtxf/rElkJtRjfK
9+G7L4lQUNrlMbdZ2836BioZvZBTvwfoIr08/XS8KVuMk3FGUUuKgn3P1xWJgQgk
iPCm6AcrV6KWbxc3MqPGvzXIdgcT95kQ9Z3rtYm43x7KKrLH+rxOZqoQSryPiReF
HfBLbCp8tqEMDZaYYv3ZGMpWhODzSqdPagVAaQgx/itdgJaXeKkRXR8WRdGU4PNK
D0UcKSK/JozD3Z70XU63LzJxhLv/8shNQQLzhTSY+lPlZnJDe6Ls5bQZf6GBTuZ1
RxoeP3FrRupJuFJzsZfZrC1gkv2TRlVw7ogqPWlC5X/7CQxxl1x7PllUMr3toQ/C
BBWbzjCuZM4LEqE0+HQ4HgwJQLdDouiLfZ/+HsxiGntDTwkLoGn6KZ02ANsKFTqO
wRYIlB8lyRLp4pWV+Wg+LptZPsncxMxiXdL3AO03hxg13HymNJBKeTThO6XjBfyS
jiAJAkHnhyQSnNAi61VOuJSwMmN0JfOhEJ9Anh1jOS9i461eQ7LdsoHhN+4bjyj5
q9Sf1AxxX020R0Ui1tf0koVxjCKj6TS9aDRMcmZj3xIyoXACjlX0sWgvVa6+cpeg
u3/B6tOjpxykbyPydImzWcCKD6XlGC8w+EdGH32rEzQ8zKLAwbB/VLfcW9upRDEN
dlpPXL+vhOpUrYOZ0Amckxv2dJuBgiMLs5tn0DfPO7fCQaERInkkmTXWck2p7nMY
QRINiSrlmZDkvxx4o/FS/5A+ND3EZYSAmnQ5qvXziIBh4JCImSCo8luIoUukHLuP
Uaf96e5jtInvSOxXGvqmFJ6j1uer94Sj1KIAHdhp7O79UWdSpIrSthOvqkcpHAZL
hizYlyQCOT8cPPV5SNhsYTWce+7iGEH/paJ7W1POxyQ1W2bYbAPAtV0Lru6JaEJn
8sY/cCx4fpo9lycudt38ObdavnQidF/xjuGgaZ6tDJVgbfXBz90mSwqWY0D9937f
q+KTcjpbcBNGBszstu2MMkG5Db9zYDf+5ntj7AqGEbK0TBKH+RpQ7tkguHsdlQr4
7Se9xrIKBln3w1IqJHJuq8oF+0ksGNBhq9ziHpObCCRmi54qQ0q6gZ4iHUshQpkg
2SqlKyOmgtjFF7CZEu+DUngAJPppBa8GFVgIJ90SAhQhpdZ/abg2CYifLrXIOaXa
r+5qUUJT4cy1okJyZMGANJch9GJcMPNsn7rV2V1hVTnNbor41Lyz6NO1u/dJ3jCx
uMmAVXyiwJBmTrYBQt/6f8ERWQ70hVx4fQqIjoNlBlbDgFZiFjP3pATR/oybRJN8
1oMWxiQZFUmbCDrSIrWOZ4NFiOsr7/Oa7NqJxbOBgOS0JIZSR8EgzvLrrflftSJO
5PBMQ53/Van1gB6TyAkhQ4iOIKEZlFFKGBlIqf2SzvYNnqApr1ZN+Yxyaifpc9+6
yOKWG9gStU/bul8HpB/9sxlskgYRvUBiRNJZelJZqOHD5axHQftlxLU0IDI6PCc1
vHqqG6DQv4bs5TbB1Oj1BvxPgeVWC3w8f8fL6gVTxJVXQIDV3D76l4fDQEVrwmrG
+hNZ0EL0dkp9GpDNBX23z5ENoK9arboggSWkvzU/KY0g8zdLf4HN95aC+WvpDy/8
HS/oHJE0CB6VWYCVlrcgQliL5V90a+yAD279dO+wjx9iM3WPAHWj1R/Bd66W4gUo
6S4VpHr5mAAn28DC21GP1lD0xWARGo4ZvynrSxduR0xtSIi0Shi9f82hzZFi3tQM
0ndcYD5aVPliu0VB4jxJ7J4xL78/d+ZyxIxInG0OXzTDZeUEEw6f5EvGYIcPj4Nw
kJGhy/HY9DfadPf+0OsNWqbOf1jlIKJ6Kc9PsxUAZRrX7VmTn5m2rs9skIiXZz1q
etwN2kFRJ/OcE2k+JEfcgaOQAKoJn2Ipgzs3okWTebUCKl76ix70ex3cexTTtM7f
LZjn4Sq0z0P4HJlCFWMPoQ0wRcTWv7sfjFFRBPdL3VKoFpK1CBRdWT1sqpVrG8BZ
eCxDRto6CyhbbmGBuwG+4M2zcsf0k52xLtkQ6kJPX5ns6iy9+KvyEWGTQiocz1ZF
SPHp3ZOnXCCdaahpqKparf8+xYphy53DeG5FF166VjExofbrsjHBnMJWmdeOg6e4
SJq//3ep/7CV9hT2x5nV5RQiY4l26H6uajbkeDVXwo3R9WXp8H2A5kWTE/MfXfrx
bzS4B0l76hl9zCltLkZTJZ1aG69cdj7uCVcyl2I+2wHGGidEGmJBciDDa9vUvaus
IywxH5r21iLFhselVNiYr3k8J+MrlbBkgdBYvQfAduFYUD+sukb/5rhYpDa+Dt+r
cvD58no98IhZoRaSNNgVG+iy2EzjzmOckMBY1PZqXJHCLpsH2Nin0cwfEdH1MXmL
bzpyB5/Frq14B/pRtE0xti24GklKnGWpH5j+uy6rTnhH5TUzim2vn79zDSGUQMFe
+/jZgrGCTfOBp5DiUzYwd8DBcrppxUAaeZilobPC8sVMtL6NNdrpCiCBoS2GwBvY
GCmFM0mWZHtZ5IPG/sSQHIvwU/YBkl+pMMILYKMlBQt3tEPCKDMKiHxItcPgG0y9
LeTquYJTcR4QhFjHoh8EzV6Bw+Mgf+fWIc5CAGEVNPV/g5A7O0fbl1XJkMSFomMU
6hwqRsDoUZNOtKqCkl0L6s+8OdlHDUOTZfb6FgWOUlXzO1PZS6bNI6Hva1U+oUdw
KkQecDdxHycskw1Jl/L42YEGGWH6SqY/HhP6N+Ar07Z3fYqdT0+MZnec1s1I8Hbn
qE0aLE2J1rlLyjzbrgzLlHQ5egqq6KabNstaMunuAT8fLZ5oAlFz1ByrkZcfV+9v
PqWxwFCdoeOhYYJTBhEgoUYhDonvtZWe30w3D9eRJcX1YEyQiiYONAgyD6xVhZRp
Zwo9rfjtLHt2VRFfvwikWJ1ASamyxeliJoCXKBBSr6be8yppnrEypb/7XCTWHIU3
MMnBjPUsRjdjeJcp3GlGHcXnd0WVZIkRNFT82UbrA3W+Zl9L9x7lTouL1FVwuiAc
ZK6SctPB7gcHd+uY8B3bTpOQV5YZBqmwCyQvFaoX9/XsgmYzrWZ/B5W3svNL6bml
s67mYW/XOMf1FEZ3FjWf5y2drWcgJt7fpD3mbQTpWMgV4hGnV3WXgr5SvdiTZe1G
CgpG/pwWJrcJ+8Z3JhdUEgGHbbmGYbAA2nYjfGMnpw5qbndo/VdpGUctxuMQ0lwH
tj3IdObeyu36kdZLkw9QCM+9rWIcRA54BhDpZ3Oot1P5r0HBUBx0fdHrBE8koLH0
W54j3/SDxAm+j2HZ96arlsIO9GLTvqCy0+uMy9J+SHeW/+pQgTkvlhuyeH2v0c2p
trr+JJ+DCd5dQ6kIlhhsfJvDjBOpQsG1TAtMMtI+g6qZ0n7mgGq9YFxIF7XV73Oj
QIj1t8su65/j2BdR3cWD6pGbGldBw/Y+yk99zR+l9WERcLQ07dYBA2cb1rQOiW9r
2QuN8SxjXjHRR0zPcyYhYaKfQ1d+3boIjhobzhmaxnHGIf8tL9vBh4rUZHLWQ2KR
0z8PdNsJjQWOk9WV/3OeT7pS9cl2nGtB7V2Q7/fjguymeENvN0XWl4q+3bttJvdd
B4mFgbY0LDnCyyXhTDakJV+97PaR4WPzNjWN/uJmziutJ6foRcO4tAjMqzj/dFtL
MFRAOoWD7hgl9s6P9Fn4rcjU4Nd8rKd5EgEJiLdcMtr6n/Zbbjfb+p2HnHuB17pr
4IKEmd51ITw2KHR0tOhsSxIlmczn0II63z93tafsrauo+ZxQddTqLF7SOKUiqGUm
pGXsfq5bdZxZwmbQctHtWOp/x3yIHwrrveGZr88rMus+sm8pjltKUoA6NY6ntYMI
AgtMNgGJfj9LSc8lCwMUH0zEZmVW6TxV+J50I5Gc4ogWre3yhyrThDTCNszC9uSq
aO9qYwB0DgXmJPVOzOrIqBDngw/qHFAuNrBItaZbkOzvOFuHZ0a097CXeeRvh5D6
5mVFkPAbxm8fOJVwC+UgObXl0PUFeVpMj3fIbVukxs8lddo6jYTi3ZiAw1JCDVvN
/USH7KGtrxgK1gVurJFmofRowKHtxLLttVf8DgU+/hqWDqha0N5Da0sjrX8bOD3X
yEFYd3xQrl8Pl8EWxRCWSBhc/xfkgw97CbNGdP3HV+rCOaE0dKgZ2WifF1vzn9Iz
xBZCB2A0As4tcpwgSF2I2/1h8a4RxWV5soSO9oJ2Ray7xUxq5Wr7KDb8hp55xZ7V
VvvMZYoLbGNbsxRml5yxXFMEbuFDsv5norm1lehQJzmjuH42wjn0kjOaCtybO8k7
oZMrbbUNs6A8IfdUkxjXbZKGmx7pqksZKnnAaFlc42hk3ZKWqXIGekeJ1GivbDmz
eQqzVdsyZVAdLPbwxBuawe/hy/Qj3CJgbxxZ9vkLHkqHaFhkuU38Z1DpRM6D51GT
aoLhra2temAJVYYwiVJNSEefQ5V0qiP3DCMC7X3PKVZ/dzz2LGvcRK/Ny4wn4d0Z
73gZlbhQawLEQp08u4CiMwa7jJWDaKSix8XYVMqzGwd7LpEshEf1EUK2kkyFTXA5
HSHSdjyLhrAdYGwW6LAu5r3XJ1FL/nkxyGNS3jioeHyO/IRk7IhXKJ8RNNudoT0k
+2opnqwINa3lMKL/+NclLCZXn+BS11vMWt1yIX/kV+HNqDOmm95J4p/jSgMVZFfC
lhcHMCyfUZRU4xwKQK76BB/svBnpgkW+jq8pkk9vdUX1Wvl44DGi4UUe+YCtHP3G
GV1mlN8MTwcBJjJlvZ+sA64D+N5SJWIVg4EliUm+p19Iaizd3Jt9whlKPofXedag
6HupZZ6mVXscXkwsQSJYd1D/7lTuZ7oazki9lszk+crTPer2N4oGvxeU4G+fUIzj
pxGVl4nUiB9lcsFNtEifhXJgLg+FXIQXevnybTPVh4PFcTl3M6hEstxGyjoDSq81
AV7jjGJzDPCjSy7eQFATAK8gO5/J39O07d3X5XipgPCC4bEB+UuZNNXmEvPbmeN6
lfjILdEDAyooHPukhjjmI66K9mchIlcQb6yDSJunULUHDWIJSkSfiRfspqr0kEc5
3ok/joEXfog4s8uDZrD1KGj+cmSFo2q3js9Cbae66oNkvK+60BB0viWVycZ1Q8rO
6lmnSccM/gOSbng0YOw0lDBg2LMvp39ZvhBkN2rrABun8cZ27DBH/UX25Ecmv8gi
Re5YMdywSXSQK0fbP4jR5hlscbbPZ7WylIP4QTnNzqxgHlhuJ3xKP+eJ/dROdtD/
2xvaUsKj2Bi9Mahxzgy3HrvRrt3tHUGYOwTw7lnBdgRXccEa7sqmv0x2gIL5f624
WCjevmbZfF5qe/zpYp2HxTifq1sUpev5FthkHUJt+3PvGf2iGNsIaKGblkZTNr+K
2ro1cAsY3D5EwxvAL/psBfyt+4PALBxRIy4UsP9tKSrvbCHeQR3f5o31sBXSSME0
UjZoZkRdsTkOhT3A0zLZf9knI4uclynyMfpd34c8dNQHECBGObgN6dYYFoAh1aSX
2RnLtmU1XoXQqhsxBAb+WCCI5zwhGZbUl/jp+r5Fqs7WqykDSC2u6dehsp0k7WSl
VYKiFdd+QoGy3RyBJObJ3h3/QvNzMYk9ILLlY3W1a0et2KDhXdPtKQt+AOfkWCkf
FJq1dQTcJqox00jgauK5OCEHxL2yV6MOiuKpvsBR+Fwj5M8ADmIF4Q0f9M3CAcNU
WLBZqwj9cTGowOiCM95BGpP18H3CclbTr8jusShBKlX0F6GjXqeFGN5bSg5sWDMb
OoYnxATOixSo4O7F/8lIP7kY95vnPRXLbhiuSuLnvqDtvVIc/MK+QzTNBK8kUcJe
gjWhzB7570lcM94Roc61pGE5cEjVlP6CCqpdaxlLx06GqWGk6aKE0N6SAaQREhBr
Yu48iBfbC8JpPBOfIl3uyHDD8mej3mKrA5UW7Q/0nWH2fisUUFbL9iGJ9fKIAYaE
pElk2ctx5TjoZ4/rgg7e/3M30Lq2oNW80zUW6aZ2DUm/qnRdOeT+WnWA1WouRjhB
hoGjnB1Soz1eqDmXuBOn4wjg2DrFoP/ZFII4ESipC3VZvJ/e12/Smpv1VT9ItIII
9j3BBH1XhSm85sxtRaerWvSFB67X1/HNAg09GObN/3MbWR8xdkeY3lN1mGC7Q7kE
08wUmFIEucPpr5PPLvFAoimloh6xoqkt6VsPPlNE+PiaQa2Z8Z47owSV8F3jZD7h
RBzGcNocAXNM1QoEX67iw6OvdQWC9qY1QyVj95vDclTkEQ+r0+Pib8SadKkE2abg
qpLTZSYJn18MNh9TdhCZPN6UyTd/nSaaFfMbYDqQSd53dIn485FWrXaA7Gbt4VlJ
zJkteD0cf0MO4rLDY3vdXpxL12yDaXV/DD01CNpRrLsX/dZ462pIT7LoByJeXfFv
AyWYS6IOb4ERAVOPHm0i2RwjbB3o71eQAkWTHPO5yJkc/Sr1ngu/XEVEMRLL3rzj
0cVgw0nc5zKLggZbgrAVHpvtBSxCEAtYi/YKDQyy6wbQ5mclnsaRScrMBzkugl/H
/WAndMqwxB090B2r873Deml8oMJ59cmN1WKLtagrQSto2Y0ycY/SUiK/pOcbWdQF
ti0QwRwtsaEut9TJAuq2KO/F7pmb5ajNoLuPHrY/8MctMmMsYE8+6WWtflcKUyHp
9/m+5dzNu0Mmcy/YvdzMF0SMclBF1tZyFjFHvZiRSaSZmVCZXTy28Of2j+I/XqlD
dKdILi7zxxzrOEtbcgRrDPJSD/rS2/xCVWUqcPAHw/tQ7ama7seCdJGAI+GxcqJB
v7+Dbh3EBI1u2SBtZqWK6x80HKgU2t6oN0EVNBLmWFJtEdRO1kP2zfCXKMjNNLnV
s42FGZlS1vNVmalhHYRGSGvU9ePT+A1BmJVfSr4eZpOuN1mjdYxaWKmfYGgQcNcU
j52LZkl6yXzL3CtAIQu0lkMF8KXhEZUlj71whm2fR5mfCqzUzNRCoLD8Ak3AjaMq
P1cZlS/HOe85zgdpNnGblTk/XDRfDCXD73mxADjw6MJmpggnNV5uoaGB21nL315/
34+kVKwbVHEBFSs1pkN41/fzUeddkFwKiaHWmSFnZwj1fKqPu3IB6bSAGL/iinGi
DkietUyVvtuoxWlwvkvExuKJEVIvcbHJGr7Euj2hStrWIf79x2ISFrjm4emELHkZ
R+BBdruRt44mvUA6AwxNOFTovRPM8z1vRznWrbdNT2ANM7jSU7C685hTz3wrZxkl
HQJ9oWnh5FmtvC9SgXSXwqzsD/jtTQWgeL3jkTJ6dy2Uut68TRbgIguTQakc43qk
+e84s1QY1DsDT62xstmYwLL0KTWf+XlJPBFxU9CK48WtdjuylOtETSVSlwt1Z3W4
SUHAjMXi44Gd9kkkB/K72ucd/NGHiZKyBKnrPVoK8N22oshLF8egYUHfI+dBIjM4
LCwPVs1lHvwRB9F1spe5HU/9dQaMkPeSlMZRgSvo5EUA/53AWRf7PyijS8Z8vDhD
9u/sezXsc+liwfj7JU/5hTzo77jebuu6Gr04LFTcaNXPp+KWTO7q/SOQ9y8VcK5C
FtfbbaT5ygLDvRvLooY/d0gCWoLZ2y92uq1lvXm+A7OApwjfBT6WyfJbYEJQqs5Q
Ei5jN/vK5o3xcZX2jnC9QnBIzjB2ZFA47J/b3+slJIsMkKbThWNIiao9ZJNFlFtu
NAAICznEbQNAWZsJP0WSdlkKG2iVa08aEN3eNt1OmdYOjOyheuSzvx2mSUburaaz
DVk6ltEyzmL/Mbph/nesaHqoX/W2EzFt3gEbWhj5x2tMjgfMRYegJLbGUocvtepF
2A2a04dzB+Mwvuav2QzFRtAvZi0B9LtJ5o54Vtc+x+r8bE0zNHQZ6Z6RldsENAw+
Gew6Y8ifbjBd4H1PdIc7kMqWlvVs+S5fp64tuSEoZUUJZoW7IcZlUKnmyfc1+KmV
Pe3SaazeR1JFyJlpoBk2tl1FFJ0PK8Hi0FO+ce7GFOTOWMNSjMSh+b+QCxEqgvOc
2oMsfBrRoHV1pocNLKzs3aeEBE258vEMwDjyAq9EXlXJIgH61gJ/t5iEhJo+i8pL
sFfT+qtrCxxHTemHeNTiHe5RgloQsYpFX1rogkIJ1Q/ve9FBz4hWklycjksEXD47
//ENp3lGw3YhfqNKnq7B1fEQmn88N1fI0+5Mtg4zkNrhxMJ2AKXiooGZGuGSGp+L
7QnWFDBVBo3TqNx3+rLKEQWbK7hGXg/n11ytHWEqyodGCfg2A5MYdevEuoxlQq0W
BGUK/q0f3tyWrZYWh8GU13cuV+HEqLaw9466hrIKw/t7jdwlvuwpR4aguMgY30D4
`protect end_protected