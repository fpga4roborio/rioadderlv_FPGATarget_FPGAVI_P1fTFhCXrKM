`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
ddtXksX2+yylW5zu6QL2Lhnb2d1sD00763mmSITNX595NcHTEkwn0zB1Dry37fOW
FufOhVzEJp80NC5qZ/+F0Vk7Ik02dIR0elf3clrjeJRK85K4e3Hoo4xn7YbFUIms
l/8VZSb14+JVGURjfswrIyCUotIzlzVYZ6gzoZwDXIi5gQIBf/gI+KxNXPaKV+PQ
Ufys/12rjO6aI/pPlqSm0hCvftmBcnezN2hk1UeXgOIuKZnogjOsf0iJVX2aOOWE
6pD/psybjbnsNB6kH5uFTA5frkzIzkzl5d9+YDm9OyC+k84E83I/7/j+rk4L2dah
QJOvksSIzN867/4Qt8qYTQ==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="MvBXkzurAa5VTw+1JJ70nePUfoQXBvZOku/SMmg4TwQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
oRtzZL4VJ4iwysPsC8SXYCzXS8Fw2gtZTOskLcDV+1B9Nzn1zTyNtlo6lNICRmmK
ZRVu2BmCc2G+fmzynYlNTnSa7C0Cuel6FYpxCBlOuk3OF2tzAmLAuDyOH3Z1Yjzk
a0aHuoCdIRKv7BrZCdALt03JeUmXKPdOmIlkVGFl8yw=
`protect rights_digest_method = "sha256"
`protect end_toolblock="Jn9CQpRhJt4rnzZPRk+dOpzAubz7omckX1MrFd4p81o="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 9472 )
`protect data_block
gD6l00tciPUa6pDNTk/+t0OO0nC/UTtBwLB41d4inuAUA3i/ALrNyoJVcBnAmEQW
ptbcNp5fxEUJjnOxnedyZEuEBxWRieZFQnkRdF269oPO2ZQWeuzMW/sUdfEP8jmH
KMyp4gSGV181GFW7ngVZBHABAiLmgDGXw4b18vI/W9bxEJ8RMqOWXttsTFhMxp/U
DXZUZ599msFgSAKx0DddCsotXJ0TKYTv9ysQ3it6Agsgbsu2CczvCeVKUpOfPz9p
STYEEPsc21QyJMssYo//httjISvr50zFXE5MS+wkNKZJSucUPoXubY+ELYJuQj7m
5giO0He8LPIGqI7y4aUG/XyK+w1rZGcCd5XEDJy2b2Ftkg5DqympwrkILQkZ6WNw
36bmWF3lUpaYM3P4op/Qgfco1ba276PJ1HYb6JlxkSrsBAeOYDWM1AmLM3SjmnqY
ddENVa3V7IwsmenitF5j2Zti+JRhvLRcDduzjKcA8pX9tmXzOdqBLe8BIcy9IuRk
GoAnDlN2RxKkEorwmrGFdggF/70aLgEu4JiSadupuXw1+bx4/s2JTSD2lB3yaaGr
vzqp/AXUL0BjtJwgikReu1GKTSxQDjkIb/Iolvx1sia6Ak4H6E0Wb14b8qoDXvfo
hqAw3jWuBVvdH1SP4gTvKREO1iytmF1/z+SA6tRKQWz3mMDj+3i28fjPeFG9ujfG
YfIiPT1mVdGJ/LayUHobd0HPPRZBU1R4FIY1DfjU0WaGBu6ybepHCyRY2zOHBFIH
9RCNpsklZrsldT08XCDAXzlH30/c5OzNr7G89MIHj+9Ny90On7GN+WufHTvWINPu
4c68M1TsU61Fa89Xlt3BO6UNh+CEE87pdIAnY/MEJOr84mpFLa07IOEb5thcszMR
ffo8eplIW82wc5UH0HpKB2Dpkdh+s1j6T3aT73Ehw3DweENclgs7MXKHZC939SGK
YMs0XfmXe5Bbi+OnpvCeH0lBiGDslXPrgMovgpB3sPn2LSDo6GaFV7BIJV0SyelS
dN10RhKM6PlUKbbqnxPXF22mWJ8FzHhVESX1JIoUgAaYrG0TjcuwtJZCeTX3jO/u
HdBwSb7mPKnvUG4PoLPv6Fp7fydCSbFpKaHRBDT2DrbK38ocd5F4dcn6FE9ef80q
85jjmCWSOzbmQ3yz+Ak+atdIvnRmT3g9/TGs4Ad9QEPZdjr2Ho7eDDJvbLzsCzde
AF39VRj/4U+jPfBtOL4J2ikxhBShpapmMzJ0v0JF7FKUCTPlhrMtV3I/sfSfkr5U
SdLJG4gINpgH1CUxqnghrwskqO2t60SWeDdPHjVcxBDOgEmyR5ZhRUh+wZ+aQDE4
w6D1SZSN4Q01Jytwfwq5ABYwQArl/An5Luxh7pWzIa8ImlFJuVp1TSS31Mx4Huo6
jV8Pr5yuQfg+HfPN0oENeOdlYNvTLfV3UKZeEVapvoG2ZMNeXDzzRmdpRHQttWX/
q3YDC9dqLSe93x9av/C0MiDurpQnpKiCRmzp8JQ6xJ+d0gyI/JRMHEgtC9Tm2vFf
zb3w6H2fj2MZx+po+v+btLnNl7bGjXm2n1+WDW938dXKlZTms062jwdorhSU+6aX
Szt5pYC39C5Rbz/zzVTVb8WiSOwSDs2JWfXN36amz+imRmlOR6owMYAtbK0MWxK4
xEHomlyoQ8NXJeb4TjXBn2ZLyYJhFsIRRxEc0vSQe1f1fF1Tvf92sjlXVLYv6Rt9
QHfqqEsdlAD9YlgYBxxZ0Ca2ixVbEQLjbFok94pHGQOgv0wcYfMj4HIqlG5M1Tp9
S8COHPNj2SuWHnnLTFJPP1J72OUt+91zfrIlP/IU2h7riQX7k5OyIRS/xoHrXdBD
v+Al5Ot/4J98gYx8GFLX+ecVUnYHYElX8c+xiSG/o4nwm36cmWm4oFmXfoqBK36C
hyTDiSQnoigoZgVv4dmhx/o7XEk79tJWh1q9a0W/KHz3VzAdIjwnte29USIY9nGF
ZgRW3Bs0b5faWLrGk/BQ5wKyxW8sg4JhUh6Onpsm0Je2WuEN/TGeJOP86/CbHF3L
zffUQeFt9q0XZ1h7OKMWqiGV3wQc1kllBw/dxsRG85OY3MxnsIdDQZah1pjBoe/d
gGqnqueVme8FdEafH/bEwvqzsDa5A4MF8iVps7phceLi2Eu1pgX/ml/n7lnQ+rbO
7y3rsvFMoJO0NaXOwD/Y0Yz4+9mXskvlOs3LuCejUyIyzDFjK9UeVG0PD5FSNTn7
vd7cGyIfbyrge/FqQQt5dRHVAoHNOP6anJGZnPvnhsqaLI+c2V/cbbS949iiXNPV
cGtOf7uXDD2q5tn19nfBgWwUCMfNRl4Ej2TJ84VuVkhBSSN01BrNKFspRICaAjjW
ONWWtYvHFbKYpDh0wOH76uI0wSH9pdB4jn8Cv3/7KJj9GsJKT9R0hoa7e/ITI2gY
ckspVBl/hnM/NT1TORtaYRqgA15O2HPa3IIprocOpW78nDHaMYGE/IL79oanDNka
cgMwYHFW/bB0ArvxFNyk+8HlMNI/q4PMoKsORgDpqE6viAnxF+e0cj0W0MaUZD/l
6n7SbJO/ymkCQ617TnDkhTG1Q+k+PHkkGV4XrVP3QEEEJlXqFvQA257B4oevDsPv
7r6bLk77mqVtbYpr09tlMhEitHSQms70hgy+Nv3oG4QGW1w7+lyf9ADC4NiCdTuU
8S04PEMLaCcOoPRg5pgydH15FvdFNRPlje7Oir2i0Ms/Tnks5MiUx0BE6odvbvKJ
jywVr0iVQPzqg0+xspCtQsf5GNR9t1DtXPnLhhCxOQFInWs/qT+IteBr+1LmWmJ8
v+jlBtNZ/BV955HjtCt/9UwzxdMrdC1h+UMYlErzdmT5raIRDjVq2PQbPA4ZCGsB
ODKIsiX1oIIfTdPwaqGHDgsdJvoa3S/mo3XKgB95yqNtBILmlJoGeoGWhkhyDQaH
KAOtDLIFWg/WDPxZPewJWutL0pifqnHNn5Q20CBEv6gumxy1Ti1ouJhCNYWELV13
doT+xH+El9wYd4TpkXsbQFDShicN/6qX3gQbaUUNxq6EAVdNdkL9zFuGRnLXqBes
5UQ+gdjc1nKht8G6GHLd4Bw1c4UQF8klcwIDsqtYFxQ7KwFeXOEMOWl7ehODpkP1
8baP+Z5oVVo8vHWcv7E5MKl2zSqamLTBkS+WUBDwLeBiJKXtS2hKunyvg+tDB6HF
jaGEOr5aqJFQCuc5I4jzY5FWgBNaCslcXZf0MempVUWFi3EBuzms+ayX9q5O7Y5W
qkORQSFEDcst2RouRjc8ow75xOqecAaXD0pOQSdlV7jQDAYNMbmLuP3lnaBS3kFZ
HvV6PwmVt8vYrzH3Xb5w6+5Luxvu8+SnWNNjaI7kPkUL70CTcnAca9lZ0F/cKZIr
2WISHFr23Vir8gkd+sLLfWDzY3OnoqAeUrJNOtVK+xdEZBa/pRPVk/IbFgeATRSO
mOOiHy9Dk9T0iqBldVs476rc7EZXcMz8TgEiryFRCxLsJpkQ1H5XQVmrArFIfYzt
u+h4KL6zWpokpOOmS9carml7P5MxXWEmFLK1sfpgttOF/qIDpymk5k1ANRnuHXJB
BdiiNizEUnMQOynq2Tu23fGqaDYAM1grsQhalbFReZVuDgVM/4GozSp2JV4XTaH2
AGBtLJZPmzjTzCUnjcUZl7e5vl3akCl9gywwmmT2Bn5M/Lx4XS23BVj7XWCR87Ql
G5iCxy7uyUq5awXAntesXF1ScSbegEKxdyLYNuuj7ikobjrWG8i9QvDlmoqPBlFm
sKJ2bhI9oMn3bX6kfngb4Gnzi+Q9NDW3foDsHQY+C/Cx15ZZEhDDf3Lwti3JOJiK
JgHjOnFS018kbKdJdLdd7fvx86aNKtvqwWV2AqN//D1DUVKb2rB0/ukt7fU1a4Gq
ccyvFUG50PCidOr71Q/OQa43IyRzZTqrMojb3c+BvL3FkzRqDESrGF+mZz9zAntZ
JRq7oU7TD1lF4SFR9cntDjheM+Onap5jhG4GAAW35qKOSrE758y/tmY4bZtWmjSB
8SRXH+uZCLiaUjNcK5+bYNWZe+nRVMk3CukeS7o2QJZUpnOME9QiC2hOl5nxw/dI
fKYpsEy5oG5CAx+Ao915XatF2FKDI8wi8w+evKh1Rue1khs81KdJrEA3pmIllhXg
XJi7GVndFcFWB1t+KNrAQY9o85IcZpqKTAZz7ELJNtWdMTWofypzXFrzenNtg0my
A2LJCMdsQGVVw/HD7IxvoQj1Podaz8pxtW/tQDQJwEciFVRY3kdESq3bK90gYVAm
8bA3YRjFqf0QeLEh7OLZDLnTAc/ygi1UEI+jr9SYghEk4fnHFhQ9SxbJP1Tj6Svc
y9dYEd/6pDTIyAXk31FFjvUsXkqjJsFaNJBm6kmaRq0CuLvdSqhuohzkMlJddJ8L
CBrGcxxf1MBFQ+wl1lhuPxtX45X79SZJ5nT3IvTx9whmtYjuFvty8d9G8Nesd20g
fVpuCEHwetfbVo6s/uBdAOPFSSPyHKMoin0zia43wYO78V9j5/Itn53lYsexejwd
W4AdQLyd94XtTHTsXeIggk1oVLZSDq4RsZuUhcmv5GVT/S1h9Gf/09kYPsk7Aljt
ZAoKUArqXhAx41QJwdvJMXqO4UPEWAiBa8oC9FKj8THt1KUJYLz1ZNUO3LmmoMyo
ba//gVz7thfVGFZDsmxbRuNLVac3rGFqd32tWYMzw1aZnqVOZN936gLOvtAG4iIY
5dcytBaSvn607A2HwLkMFr90fvCJZB+MXZRIgs7MqyUTowQoWqeG1IDhS7AA2kbv
LAnRbfoTXZwv9uNiEOkq4eCxjowhY03G74FQvSz3eTaZ+wR5V7D+amkSbmLoCBwK
eIk9dGFJ3uNucqnpCrqzUtsaRLlW2aGuuWZjtVQTsXdqHNpY1DYmyayUcc0PbyRL
54hocoYKZbplfPe4LFCbrHsDuQpiiYKxhosfnxEEszYRw6cndfiSqEF0T8AIwrHE
2FGAeYN8Mjhfb1vtcGTMZZh6nWXngPtagYWEBmaK12AU5H5wKLZUdxeMNvFArUz+
2Vbb4eilhFqyOYa4WGNqh62wKkoIjeJdhNXtQlvqCI5EvOgVbOIV+FeEPwJWOnsg
GMmjPLxYN97sIy6rFC6tCX7SM1oLZAzI9SuXcW71ycSWP2fzQFm5DKV+2h6je+Z7
nV/spsMOaXVIB7Hwldvmyem333McZDMEAb3BKzK6zjxb33oFzxgkWxQpHXE5v600
CIr7Jv4Ss9eSxOfQsvas0TN7K9dv6kg6QsCf4HxNrSY4zlUKFe9gPArjmk2js3Ih
gWv9KB/KhdSmSwIoK8Ju8LBKDtye/FTTcHri8LxY5Aww8vJYcu5jxksCHNDvdTNg
UQX0qTRXYcinpm9xfvMR4ZxdR49A2Afhs+67aDGuFiCcfKsY9Ee/ucCF4NrhkpHU
1CTj+IVDzyWQuboW9Ao1x1mrNieux6ajxanuiW+s4+SmeDjGzkRPQ1m20ZI8zmoL
4EpF0/bp8MdIV4bWOuCaPvqfPQdhGDRS7e8LDzu/hmg6Wx/VKjmct6+pd8TT78TR
6v31nNXpLXI50aKOIH/Q/bNAjKDNqun0okaC1kOO/AvZRsLbTPRywhByAnNM/d8O
n3LGVPa/tS0aftrhRLKsm62d3vp2jM4y4xGirXg87N3cL38RqoyBA+no44atQ1c5
Y2TdLvgS6mK4ZhOPzIKbu8YJSZO7LTz4oSahDj/9Ee9g4nnMZdXxyvcUbu3ipM9K
4KtF44hHOkU8OboNt+DPVXrP6Z+GmmaNuv+fFm8DOI0B/0t0c15JX9HCaszU9X0l
AaISxOz8KbabLVddNO5ZinfAWJM9uRoYR9Ypin1dH+zunfmo1PpBB93BA9eC4i0e
V6XaDXqblX76gFwkqqVuJTJIeXELYy3+89dQGEOKiMvBwLecAKAoq2LI8zhZJm7O
+hJzcW6NuQctIpriQ2GH5iVEddwsxEj6yJvDoa8qs/RJ4HcNcnu4Qlv8x/YtDJWe
IHu/Fln8ZitOW3Zkdji40TQSswJ5dTcF6Okldii+aunCGDvWvf2e3HtAEZfyA5hU
kK33cZ1wl7ZvUZT0mcYIpJ2haT6/E0/3NxWAd8JAtcPAyXzA8uxJ/O6m+FIpjxXJ
Uzq85KaIH9jgB6ix2TPub/NnpJXaRYCx4G2xrNfW8gCEIXKMsBO8UplrVdFsJVuH
JdjsoLtr2aN3MtXTsx0Wrpr2CaEDvAQwM8TNQZaiaZ8YVkIWBicXSdSyOQeXr1Ru
44KnsokQT3jTayWu/30FnF9/4pExx8xwawdWO4Bq9+FeYFpWdit8OaWCRkVBQRY8
MdKh686sVzakqPOwsquYrC+TrZC9WpatPMG3SXddrqyGPodqxhayzg1UfNwxCsct
69Huq0v/ByjUwMvbeHGYbaGIUCZ0ycZUi+4ltIg/Ewy9wRoXanTU+VX2SsRmlFm3
DDk4AbwltG2tSR22IWBfZqossnrSK1NwQOan7306okTEPG68RK5Pj1tx1yKIK9PI
i5AMo0dxOdj2dXwbUXYdwq7bvt7gUSvrx1e/Ep1p2Aq4mDBLSHkr3xsXFoLTTZu2
JyD+r+V12MYjGEMebjcWEuo2EHNvQ+ckboB6gIW8Av6sI3q+HsbUBtAFspsD0VXY
KextSxB09Hi5jKSPPIM3W14Xlrj8tjDj+tIIU3zGJdDKqLqiW1xzjrJPHR+e6vE+
Pm7NoFobYYNcO3adjEXQkdsxOON+YWbxjNgRCMRKZ1BCU6TIRA8YVI6tx8hfvGIz
MKqAS2xYXZUpHmQb4gBC78sgev0CHFY2ar6DpI45MUS6HUOVZDzgYu5XHREVzvJ4
FEpS6VU1noxPHm2w4CUBKsGaYd0kIoGnGt/zdvl03r3VbPzHnhWHeZtl1afmvAqJ
kJKTAJ6BDwFiWpW4xG2QAJemk8rnPmIo28XYZlqEqJipug2srl9+GExPzOe9juA4
zjKBTF7P7JNdbtoCojDySSJt0PYRyKYVQC2tAywO0Wzo8i6YlTtFWoNTWQAUQFxx
OfQv/vZK166GPYZAmOAo9hOlepf0ZsAEsE8Mr9lrI+IrMHe0g+S5D+4YXkzszHQP
0HaVGBnzGwQrJsyJR5GOe4WuIWtD3lmwTl86ikhM4EJckgHF/BFMwLxd0V/3l7B9
9HF+kAshoaj/13Kry8M8qwRDUyVUK8nl7MermrtlFK4kkz6x72XbxWY2uDeL/P8u
9AR/Vb48zmvWzdXIQi3unyT73SMXWonTzaC0u1QtH32I+UMPWgLO4pZXfizROdVX
EJEGzWbP9r9B17eToVjvKLctQ0lxJQNKyktbyVTXo/agQhdQBwRpUS0WrYagikWf
PlBc3MIKII+Ig+tZITvxZXJ6pdXmbjGVN4sktjGwsBE55QJgRcbMfNITMq6xOqD+
y0J02MTtNwoksYponBbzqlZugchH1LfxF4zIwhPQZfNfRrKTR0Ox6/yJOfvtpnjZ
jiq2NoFpzXeCSIqtoaCZXEDMrlvq758FTmlY/+T9AJvnM2GCUfDl81Jk3LV/f9Gh
OZ07P2mhmnnt7S/GNiNWSizTY4tCTc8a0O1AEErnBmsdiLgeI0jiGXd+73ej7hnB
r6FZ8sjj3muKBvVu2khjwVoK0WH/o1Bn8PPKXD73HJOr2gMsB6YbnBflFmunUunr
re4Zx8BIg3Ycsnkr1suJ67XIPhxmqOz6y8ZvhZ+diKy32bdxY2XBb0Ea9kUGAUfO
ISAy2HR2miodYnAZroFDSv4TzO3goEiJtwSSWk/KNHOZdApwirgWJMpF9R9dTVPt
NCt5nNNBdqpu5ito00jeFFX46qUbb/mkvWyCwUvC2lH2I5U1DUPwZ6gE60NeLqVg
r402W4IzpTk+vGO89N00qHpOyKYGhtwfiSPC9PvSnyuLFPYDK6Lm55seQSeRMDGv
1SSFSy1bVU1sXV4aSheLy58QnxZ6ZxRrqa2I8xVNfa1Fh9sQtyZmgA137D/jcE2E
SyAykrRgF4P1Jn+BhtWjQQfJxT/aJSsxW4BE/MDiwmpAo1YzsOx8woRhyp2G1E3M
G3JfB4poPIXFFNYIeR47l5Mz3Vvy7GiiKV2Jb1zCSlbHM3j7+sU1B52aDaF9nHjK
17gP0UJxQX0KXJYmzzpLz252JHgtCpGrQaQlfJQ+qvlm/QAUDZxmY7wM1SZC+Dtt
txxBnSLliJP/zBlXlGrvRClyaKAUO+XBfXIOdqVcyh405LNlZSguM/yojgRb5aKH
pMGF9LHHXL7nmTt/0FZKACpgOBzmOZ5ahEumSLEbbcTYJ6cDusUvZlWRXR/nd9JM
HEMfVgAzXjYSKs1SAX+0IfbUY3+MshthjayJaS3jBru53XjqwSAhPgIeyjt9oGxs
XQdOscYOht6sl1I6KdMncs0OlAkihcSnUJ6Evm1jUWd2XHYD5ieQFKaeAD8WcIG4
24Of9cnX6UTO29mN6eUP39ILbDVxRGhBQqASI17YNriVDhzca9MdHjRvOhPkOXvt
ovgXDYGIEpH2ilColy+lQzkqlfrMWSIaavl36MnMIeZMLN/HdcrW6Q6LUMuRsThx
0VbfXu0kLSwMs8e5fHOUeibM4zU8c2XaHptI+Ul+4z/V4E5Zi3r/XeqbBSsAP2q0
bCzED6neUL5/yvRxsct9GtsZ4PcnHHKg9vN4lnyMTbQljvb+l8CTUGtN+L3qzEGk
JAXrMHDqzkCcZrCPKZ4ky9lLprDzMbWzqZTzb2AGwbgUelVkzylxZtAxwmfygeKC
7TjH+xBfrTsliuN9lIFKfcanTUNgZU6IIaF1On58hUsWY5B8/5YYhj/9dsdKwzXF
GIyvPf27Hy86D1au8pEbNb61sTD5YzYEHzNfC5V6wZdP6Wi7gtv4rwD8civhYjMi
nm84PSg+h4mznQFUcnblACqPWLGrI9GQ5RvmrcG04ENXfqiYMpc2vm2GOJpkHdrq
X5u8qjtYuGXCiiswqlmpNH8UJACiDb6EUdZ2BIKRNYoSKktkQHDJf5BEJ0qldoM3
N9+XuimgmUSv+4/DGaFyDG14ZZoYOFOS2/GE9PH4/v61ew9kj6kGk0ix5o/2mF8R
wrh9l9qtcFnPQdqUksjrf9H2WPZ95+PifETHbrMuNRdQ3QRt3IK6RRWqvMeKpso4
8UQ+Xm4+eI89/WKkpYeZW2K3/w5ns2m+5SXaq7FJYoOw8r9xYcfefaP2oSc6l2aK
e4i05qDkrQMwS0po+dB3bE305jLVW0x+fGGuOJ6wAtUrNfsKLUZAklOrVW/5WXyU
KluzYnZeDZs086r2ZWcx+Pesv8Nf4FsxIjzDqAO8SFn6nt8sGmSQuk5ITG+9cbjG
VWTU3qdW2EsvKD2R9+5J46L9FulbwYgwAgCfC8EcsltiRATedeGuGl4t98xaxO8I
SfanLrPzPwNm8Y0VCbp8+Gz/G5qmZqIhUvNB1EC1cB8TkGDvAE6cgDr1r3Nd1zFp
RSXCrrlZdexMPAz+uHnnMV3tl8aKRtU7otA8zoZIK07h/FLEA2t81ZVixnPhfLGf
thUrY1wP5RCR4E67Si5yaQ5scHPqGab+v51071Zw16t4VMKDNXkGER7zR4AFeiWY
ORUw74KEg9oLgQreXHSrHj4InUNKAwxIr2GSpV2POmufC4djhES6IVDzfLlLARNQ
vtb/8ENQ8TTfXBmbmkWHoQQNoWBGmN/ee+Bhm0xLB/lUEuhGzn9TxrNU8VKJIpU+
6aU+CNt7ZGUkNSGPNTb8YL/t5jHPyGhirTpAF5i39SW4qAmtDcgfyEbFh4+ykAzz
dkO1lHIMGHMoo2nn+fvTiMNoQA7OrfMRSLBevnsb47GyhNw57nrp/LtAiv4cVAb7
thxGvUkgqMO+VF9EF1J/g2JFS3h9/87CYZz90+aFJMlo9LkYAgYnwAUhum/PksqS
zGgLRNV0biLgQRWHzMVfHgURSKkR9EqN179S+tIC/WJaJcU3YIot7Gs+xojoEqzE
i9RfZMBxuhBcGq4lAZfd1sW0YFHkvRwUDthgaat5MGCHoZSlHUhOihLIhNBcQV4t
vtyUfxW/3V3py4W6M3cOvD56glzRgdL9e3IQkLcrF1HJvkHBRyIKKWzfA6ZQafRh
6D/5+L7oXJ1SFfPc9G6NrMjTmaNbde78csytcfqnHrEdPF4rNPN/bfZnObkrvYPW
xd4QIWwu3fQFVLbKQQSqUQiwq9DGUTl1qvl6xOS3ejglaqmpDlAGtuTY5kwhe5XE
AobvVJ44D/7/X9u9Zzqi9zxox2f+YSnvX7xZGfJNNiQXuOt94eG8tr86CT/0tC+g
OCRJjGW3F/9ovVcIOLg3bJ9Hg41Z/CTAfqZLdgb9eXsxkRSUUm6/aQ9GgMJj15Pl
WRKth/GnMPB+azrtUH/dOT/aqNGitM5u5r4Fy7vNJVaQ9+drF5Xb3CPz3RUUiVT4
lLfXnIMm0wLCDIwd2nNyGlkMZUn4hEqp50rsWEsiOxZ6xCn3H1NfyTWaiift3Qu7
ZOjLVOKuDtkTxsXU2HAW/6OqaBEUpgsKAaw8r+E6kn8QSnuW1nknvAc4zzgbUX58
QBzcLROQqry4vcZDLebbGPtpJnSo/SMMTgKDFT/RDuJXUy0FXQyPjgovneS4NZat
CPIzqpEeZp1b2MtjTP/MPytNAOsYzo4wddbWiWubLm9jmkWC3CuyWJnMMx+UTSeW
by3gLLoCi1xqkS/5k3bEwhf2KHKyGF6K/NgjRIEg1SviIWCxZbNuFR0VedQa6aRh
1Jp8n99V6NrfXib9Ag6sgYkOjoiAap2gwAOhVlESYeFcHuP6Pw+TDFcL+6mV1SVC
sbnaaHAKnNdwehTDCLWer8+C/U/Tx4yoBHs6uHhDzXUFJXdHyP0eOseKUwhvUmMW
SrcmcYTGS8TTkMj6fe1BjzB6Vu5JgTMc+de6hWL5k8vBMsOHWOqzEiwtmENLVt3h
6cjWiogWJqp2Ik6I66IOgpOd3wz7LlSgFDNO5V+mFHOiQ01A7WjPCkZr57LovNxH
geNXhp3y46oLpJbeigJ5RpkX488db1qDju9qwv2kgrOvobNXrx05y/Mi0eStjV9F
XbPQDrJxb1AEwkCACpvrKjelZQenlQT42wMVaZrwe+4t1oGWSmFIHDhmOVkfsQOp
V+OGNzW7QnYrNQYSXHHFY3f+Q3RJYO+p/80gq26+aaXzk2KZzNAr9nOTAyzevKjM
bmtWAamLTo2Crm91hs0P+aACNG+ip7XQuomEy3Fd5YseGcy9ai+s5LMIlaEfRN5m
HbM2fjrxCKiGK6swb95AX/xV2zoO+kXlyaYmuWN72SjAhOAaMoGwQpSnWfGNSdTY
gBXn7eCvB9p+fkCm2IkDYfjOq4sadFLjZ1SpZQ8lVkmbpR/jc5YrHXnIYCURzxL2
slZo46Mibe6lDLFKhCDucI2sHI620PI87649WDL+oMqfqq2gv7mxOHKb8OB83Ujc
LfvHe7YOHpQrYcKGthMJkQ9C1wBaHF7fhynWahj8y9AUsDX5ucO7WQh6UhcZGCYz
sBnF8/Al6ElklHmNTIgyd4rMY4RUeOqllYXE7PBBygysBNTN8YbVgWPRy0KfWusT
GhG7jH+V6/NXRJVh0Vne68Df5i3ePLROsPkZGJx6y3vGM1s6omw9d23WCrnIi5DV
YmK6qsqYFp/LPVUjXheb8ohIo1W4l8bQssZFYGt8B1sFnJIqi3yUuIcZFRcDaVB/
Y/93FIlBGtyFWemBeuzgZxw6cFKcnGHS00bjyD472xrhHeEAzERHD1xvVbwMAhlG
cfndbjok0HExkUKZ4/QjlrnTUpjQ6oN1KHIcF/yjZtkQ5xtepiAQSmQSvIZomXlG
GPdJrJar0CVCpHlrCQtlE6XdAnxGP8Ke2DAm4RNppP/yQnLan/L5WOMCevzqU7ZZ
PUMZx0cnrBETepmP5B2L1aQYui6IpdKr3/gkfrMi8VweuzJ9cGyHuvit3DjNuGbI
XWV90h+nl8h2SmU0Dv5p1Zwb5p12XUS7CoIcj7aOsZPNYytlyJvbf0UooTqDJkn9
4sMo5HqskqWCfPFkBiZJjlln9xCSpFx39pbjnRwLYMwb49JNZNKlcVPRL7XwdkRJ
qL+zT1ZNqR2IrIdNEgcJUt3edkI7GAaVQO672hptqcXGyzUkbEQv1kZybw/oUENm
4kim9sVW0IDyl40cYM/nYwNRC4kApnWpO0MC4ysYH/DEv1GHTFLImQaDhr1Ce6vx
cHUYrHAVaLJRn2THuEQUnEYANspmOlTQBeIGpY7t4jvPSoHJlAbkh72/2l/53E47
Am2cJ/fcxcjONH7XNkwiVz4LvrcsmziBY2cxY6qieOupTEMuOixIsSel5eVpsKTz
R7wUHF1IcpOYy+bEoLhOv99iPNdmXGQqUzB7KL3pDBTq5/ZTBmCnHCINwKXKQgji
DgjRmej261SJlGagNKdcbjreBtk6DUiLrYw2T+vFo3Xz2LTiFFxXkIt46J/4rLlZ
FODC993Wv8fBuZ8D0sXYOUoPvoT3hrQCWER1Gn+/6cQMOl2LfZhvST06Y/P+DTG3
nlp+KY3hgDIUw129vEPd4WV4uU7t93wH3vA6ISpzvryhDa4fd0LWHzVeJQa8wMyF
0wkQgjK7P25prOkQeJNxxQ==
`protect end_protected