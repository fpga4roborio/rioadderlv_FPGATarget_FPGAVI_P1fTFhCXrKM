`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
ddtXksX2+yylW5zu6QL2Lhnb2d1sD00763mmSITNX595NcHTEkwn0zB1Dry37fOW
FufOhVzEJp80NC5qZ/+F0Vk7Ik02dIR0elf3clrjeJRK85K4e3Hoo4xn7YbFUIms
l/8VZSb14+JVGURjfswrIyCUotIzlzVYZ6gzoZwDXIi5gQIBf/gI+KxNXPaKV+PQ
Ufys/12rjO6aI/pPlqSm0hCvftmBcnezN2hk1UeXgOIuKZnogjOsf0iJVX2aOOWE
6pD/psybjbnsNB6kH5uFTA5frkzIzkzl5d9+YDm9OyC+k84E83I/7/j+rk4L2dah
QJOvksSIzN867/4Qt8qYTQ==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="MvBXkzurAa5VTw+1JJ70nePUfoQXBvZOku/SMmg4TwQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
oRtzZL4VJ4iwysPsC8SXYCzXS8Fw2gtZTOskLcDV+1B9Nzn1zTyNtlo6lNICRmmK
ZRVu2BmCc2G+fmzynYlNTnSa7C0Cuel6FYpxCBlOuk3OF2tzAmLAuDyOH3Z1Yjzk
a0aHuoCdIRKv7BrZCdALt03JeUmXKPdOmIlkVGFl8yw=
`protect rights_digest_method = "sha256"
`protect end_toolblock="Jn9CQpRhJt4rnzZPRk+dOpzAubz7omckX1MrFd4p81o="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 19984 )
`protect data_block
gD6l00tciPUa6pDNTk/+t0OO0nC/UTtBwLB41d4inuAUA3i/ALrNyoJVcBnAmEQW
ptbcNp5fxEUJjnOxnedyZEuEBxWRieZFQnkRdF269oP88vF6xePoTnu3jnkaw9LV
GUj53Ro+hZem+lG5G9DGc0PmDbxMOL7kVCeCUnIH3TrPoLcvUU64CB7LqD2jlorn
XdvWTTO8Kf13vC2xNWnh6Z8HlVl9Z8QJl8sQO9wuSSbYIoAXvcubmv+eAM5oABHf
QbgLsWR5rf4QY451cvjcpb3BTeYcraqxw+fqmXiOlzSPpVRkepk7iyjgb6/AbwMH
VFuRiouWSbWB9rrDfXjulW8SWzGszE+boef08/8vSVqSua7d37DXpI1Xew7cxTyL
h0a3A35Fhh/3hiRRUSZoVP5ExBbWLwzFvCMzdMRYP50cDb3jHzg3LYRaGJm14QyQ
fde1tGVoyTsHLYnVGd+eVU9O1K+4F/Z0BOocdHpORzdrTg+X8dQivqkl1lSKl+zV
rrboQ4hw1R7Nm1DTan0+STGa6LxZmzRpI/2yN3oE4OG4kjJjX/VfLHc6Mb1N/s/f
7IWcINzlZA/aeDqcowaRfQVw3ar148/NKYv+J2Tboa8lsCD7QW3shOA11KJV9ZAD
St31snT/D88lR4rt4lJ2cpCD4jxxkE0Cbw/e8PY5W7ZlDMAmgeoUvGmLkXbZHJk6
9MeVIdcqrdm/aqRUOGvj9dQ4Jn0DDkV6Bjv4iYAuVlU9NqZQzu+WUzRelOFf2/jx
swOxwRUqUQrIkp2c9Imq0jMw4dzmtxDnXSfkjMiyBwJYsJ+O7yLOWVnYSWZFqlUe
9shazUqN6RqruTSrQTGjEXHiJdu4CTT+6t+YYaVn9RGUfEQU1ncjeHG9bnZpfRBP
+3/Hz1X/aXVO8odjy0fuUgEhyORCIs18fvOZf+q14ZQEWYNZFZdomjKTUeHduYrg
EcW8z0gPuYeC62kVI9Q66ORU1e5UeG2S8bL8XVf4IqKivKKBk7+nVcJwZ/4y+y8S
xggktQ+xeFMW9b9NDN7s3wT5NlLRmGgr/XGkZJUDCyqmb37VG+KjFoMyKAhylN20
v+4PHVHeUOAM944LnoqYrxc62wkj5dAF/pOB4svYz0wZ2odG9A8LGHVL9OLqqTLG
8MMeFK9O4ckfaNrhVccodyd06W5or1lna7F6hveGu2sdRjM49S4/MG6WMPMP7aXV
j3H1kiLdSbJGs2dos44V/k2tzxg9y29rBkiPqqYkn7OFadd/ACZ+DxmASz/zRxRL
Mi3z2EvVAL8qHT5URb+OgRuBgHGrhzDde67PRFXaEG+fqO+liY3cK9/Za3ZVsMQU
17QgDNvixk/5Wf1hG7wISPLUScyoqOayj7P6l3H2+REnwJL1sNQ8mTeLfExidm3q
4SyVBN+hBWX9aBjPiR3JqC7UQ0Ge3C2ifqg0eZ+hEvTHXohwqDYL8rrQpn1BIlc5
XNXQlEor0CCFDYQ7ztWhlhydoWwoF0oPN7Zzxg03CrihlEkTcud78EDWPnL0SYbC
T8byoW6Ii9UPZAP6ykJo/nglDtTzWQe8jWxI6SiW43yksJqGdixXEJkGKbxS1oOa
LGRBvZBubI6kQiJavGeDWtj7YanWNWd0KubCV61z4lphg65vLvq5KdzrHZkJDtw7
wj54euM8oswcnlvHbL82hXXHiqgRnC2ivosn/SC756KpS1upKs0dht7y9uniD4NC
gBH2BwWPV0twPHHVRpXPsJFm394YdhCLZz3/lbwizU4qBSpDIYR4ofZCA0u81MCf
YMTvkXn5xyb59lUhYrqCyd3QdLFDXZQc5agojnP27hKmgPpSXEy+VGqx1necS4u9
kIwR63o7/ayyZVaEiV6DgT7YNOpzzRhoYnwudbIOu5qJXNpYNNcdwrfzwKw4BIvF
HfnQiP43KNkP3ZtspT8x1ltWx2SkjLjOMDwnaJSS+8F05TM/a1tCW6fatYsqPk6w
c9asTXU4LHqNHqxHzNQ/KBWwM/l5OauatXiIZmjEfT7pyWYKitkKhF3uLivkdtDQ
WLQwqdnESPRCgR1BTfMiJKqmEwrm5WzMHtQM78yFo1Z9OWvcIA4RtZbo0WMZguDN
A05TOj+zfkOnsH5yfXm63ympARYG4Crdyq+4jXgCKv2mW5qv091DocUbyi35LqG0
79T8ldb7J/1p+Sa83eR1gNIt9+LCIloBEfB8dN7daJvpA+QJWWu9NadGLgmIguTw
FWZylGwBo63uqmtCLL07hzBpvqGF6wNN0gPA8gMqIMmANNMNIHO2+L9VuouW+IDj
EE+d4CMNOrL/gf9kcvePMdp4Gwn72e0uedj2KXcIaGWD4pXwX/gyRxqg3122jDJR
nSNtgGBjqqS4q0hD/4fY6/0C4Og7Nm+05I2VOKGRIi2cXEvEdXcbufLxkbsp8cSW
irFJbGEXV3J2Oe4Ig6ce7TGIAsVdVs4npeX/PyeYIoycDLWfpfK44v2gDh/jv+gf
b9B03F6rrKx1hEqLVrDO0aRiiPZZkiCfvB5cLNRejI01R/OvxaeMmutkIAfAxmoo
WwkS+2G2dIosuenpVjRy96vitITL0UXrey9qC7JhoYgdIzqL9otQK+tqvZ+zrIRP
Q9n0cvCJcMudh8V9jNLGgs2sS7ZqwnwA9pN7EUJ+rq2BuBbk9p8Nb2YNf84XRER6
pw6GT5JXrL/Dg2u1P6bfnHWrBqOHNwM8nsph5N/jRGAbthOeIlWl7uVKP1MAwqmF
qkXw7gckYsrpcTJYgjqfdoMBo/MiRzRWf1CNvBECrNwwov9uuMZR12lo/jznWBQq
fgg1b9f7uG6ATvvgW7LsBvRB2IDT0HZkC8SDlvD5QW7JenMf+EItbgk2tT+8vw5S
zLIj3KlhzirMbnPubgHG6bU2RjJiUd2EUdi/gd6hlTj8aD9GoasfzYCLQvXI4I13
dAmWI8xHo4Anx7H7bW2Vyfc3MwAjhXivw1ewAoh9lX4HWTiFY2eBSnih47ffRBzg
HSRKWfCZqtTfNJyTvcJ2CylxdiwEMPAfkMbe/t4ed6hULxCFAiwecMoDUVlT95Hl
AfSlu9bm6CQYEbv2VQoHECvWaPO7BfovIyEJZfXHfDiEuUS6xGrVuJvevdePsrd5
PYkP3HEAWs4uRz6cBugfQC64DKC3VIwm55CnsUXvdOZSSkG9vDOljIOTbi6KLDNt
Ox+IWcXSbl8uMJHj82us9OXdskPjsSyrKvWv+m6BdIsgC2LZAmcv4IZPqBbjZRpY
3Rlckt7eR0zJnP5ixTk7aSBeRZly+C4DiXMkymkg/aEYydejBWOB3oUQwhykoJtj
gSDQDJIfR5PpCPoAtJZOjM1NOThC1WVIsdRqGr1FS0zDkst7eJm3Wl+RyLeamVqN
MdmUwkr7w8GqWFqyhiHBqbwHlHxm4wc92eMbaquP9KHFeMUc8KlsCFlufBJH+CvJ
OD5THJV19s3H/Bl2l7iRjPKrOmkTj7p1swd10Z62KKOLCxfK5LgGYR2+iauxI5fn
0Jya4m/cQzEWFgYyBosmGf+dp+/7R2yWNPDbiSd2WtL9Ps7Dq4RUlBhD+JoOY7qh
fk4vya/Dgjw3dpfB1qYqH+ZfyUsVQLKlJy1W93XJ2oIs2RFqEZgZx2kLepDrS4Zd
lkAXzBpyMlyCqSERp05UHFMJ+rZce7Al7WAo/XX3bLpUyEUxdmZ6h09bSl62WskT
9ByOl3/EEOUBttumGXaLN9XwrEldcP+U7nrqReEfNcyAmRCYKyicbNulRVoQb301
PR9gZoU8VzEy3W+YuQi9N17oABB8DGV7A4Gi4OVwGqp2vJnayVF7QeXDbpsCpFzG
TEhuDriXl47foD/MA8aL/1OCE1/r3YfKkGpoAUs4QNOFdcS0QZim5a1LK0N7MBG6
AC6qQHyg6t9PPU6XBJ0+SOPqCvVt6glUX5rbTPgme4x5bAgXWu+8JHMEKMqzrzD3
YqBsQpQdA1fbSzPwjndz6Z86sxIQwaeTlPYV/eXh75J7EW009wcAGdFO4K8pTBcR
iaLaB+0QDOzzvaiVcvflSbPzvPC65mVsQwq349ugnapN3rIHK3HCScxhIdRY8LDv
UvWLu2tzYWeI7Vz/6QIrtANWnvuggYFVexfwRCfB5Air8ai0dRqLbHwW7b00T9Ia
vp2yjgd2IG+QNGq5V8844CL3ARrN0pY3VTKJfuSJmrNkLIPGLNkFkFzVw49IAw2k
JDzykFWqQ/9TPUy1Blb+i7NSbCYp+Of55Z5TMn3xCfncPxj2Oak25QJ/EMd4uxnQ
xWw77ZL2i16GeoL7wal4+wmf4XPJYVFV6Ux1sFAtai0G2H52iIpO9EyNfr1o646c
69LHXepYlDxPxpA6BT3S66cILv82gTYvyxoXrfUeWurYXj/QLgd76KWjlaAYbNoA
XkEfvxgLoXeHt6RM/urkUZessslWf2qeeEaMVs8VJBFQYK3hlzk2D/0S4VjKqkxj
Ivgzpxsu8YurQwKGMzdwMHlyZdmc9X7Ffo7ZEjTWvj1wKs6yzQfB2jeN8vhDh2L1
NujX9l062Mzlb7cq+BY0tda+m7QAjuj/X5qlvzFaE7svSiTgSt/ROULYaANMcMhJ
2LMOT3dQ/0yGV+vwX3nDuSfkI0Qnnm/msbeuW0FmOGpgUWRuWHAR74a5YBGfFTg+
/27hAITr2N9eT3rrqFoII1Qw6IX8VRyf/B5N4L1v25dIXYMy3DF47x5Bfn5boQpx
vzvL757B3E6JrN12NDrLuMhKsSA0QSxxiwNbQBrQCESAeN5AdNwNSK1zkK45JFRz
sT180feMO0KsZWiCbXLyqYB0yErPD4GJrbnYkZTA+DsZDXQk8OCPK4iEYfvc+rii
bNhh7yUetjiFhCpIESx1mapySh4EZ4WkfmzWqzlSNi76/RqFv+g6MOSUZ+b3x3V8
XrRV9846QANooAuMVqiSE5BJhCB99C96Rj979vyWujvsNDeselweWaCJVZDvl+Ew
ktQ0h8nlsf5iFHNzvQh1PRftJo4gI+NMc9HUgVvAipMi3V5IjVc9wUXjhush9pRh
r86aDisNHYZj9G97EDhWzX1p2QJIiVlDNWa/WmJ+6C/nSgn+8cX5pxSe8OJkwnro
MquSuIccnQJ7UIlEWOVGR7/gpCIMIEDmzRvrQvbZ2Z6r8V8cubmM9O1uZgr5EJn6
gby9CsdHpiHle1O4qHnCntxWkvtQuNy/7LYxphkpd0BWAPgYC3GN/Bei3SjoJ065
pp1xBlisO8du5z40hVkI5SpgTzaQ872dUAubLXZZ9Oa8JbB61H2zBRlaYGBjot0L
/KMLICF0USm2teumjaPfgVO1bYnesqSEiTV+ws7Vx1r8GJfjgR8UQQUdiBPP/QGF
3igoc7BSSj/hJ+EZ5z0rmhslVyoG9GPrJMCzCMrrU+cS56Icql8CEnVU68+hgMJF
TgSpL1T8FhVizc9IfI3yNcjtTC200Qij23gsZoTv6rJ4D5G7i3DXrvA73hnKFMb0
IZ6pye9a1nyNNO4MdjZjr7Vq1zgD0W3jZiSOAxTVqb+fhlTizVMiGpdbPKNqAfD7
FIYTfyagctVnp7Scym/Y7lTECFodJb8MYuVNZ5x/IF05DAj8b200kkaWH+tSwvKF
aznLjSxVqQX1pPySqH13tC4HTZfqwBStRNXJPdCIGqVkj4p0suucY4Hfh5kER5uE
Cn7LhEr/giEPbc6NMxGF42V42RatRj/U6zIsLTEoOiNdq2L8OAg0GWONgq8pGJgg
1PwR8+KCxNWn5iAT2n5qXXDcxt1aFg2pASlil2w2Pzd3fS3/pWBKq2RDZdpPCl2E
5JhLlinXn1ypXQX79mqrH9ZkHTzATvxoXoWQqTklhceFO2q3TsLiAREAMKbv5FS8
5oJRZBk5pT2HhiW/C0SwYmdjMTphC+FW6JdQ5mswKGUUBYoe/ymD5WmoDF2o4FIy
nebJldjEV/FTWkh9XYBQDka6t5/XWWtOiEMBx3mJt8KlsDrKaIYJxXawge3I+yj+
pfyTI2A5wr4w+f5dpnp8XkeX+VRvnzB6McbxOhRGPBHwt3eYF4n09PCt09Utgh2A
SrN73vHSAt8WbF2i2vwBmdeLYOKSq61r09llBEy0ahjFfTBADPrlklYqzvtjRHRX
RNwLlAjD9VBsitioX/uqw9PVIKb5aWsGz6OV1Y05nRLDm6Cu4H0DQqFfklccZyM0
P17ig3RRM/hKHcFDUG7/aHju1MLRDZ3wciqnk7aYiwgxYDbw2JkiJY1GeJ7JDaMI
eFMAKDRc6oiCjU903hkka5noVVY2dZ0LVTcFlzjcui/dDp+b4JAEXeJ/LH6uOFzu
3Ln+ctbxbKVEaYU/UUjAv8n0aqZe4udYJkBowchF+jXqKEduzgvLhX4GV+G6gh+Z
xdTuHLxvF+HxuAwRBAE6qJ/ar+Ax1ta0EBvQCEP9Skm2jlpvY+QmZfI25PL65Zdt
MjN/OUj/HXMnPBm22G1NqLgIJSom07uj0I4OpalhVntTIGqjREqyFE2PChivj89j
N8zsHGWo1yy+XcbWoeq9TBObAg5Gg4RlCU231gh6D3ZuEWAgIns26Hj9c0D0KmQV
jQoO8vdkI2qKUiU6sWyCHlEHZSfHOlj+drlKTwBXW3Bh1OdaCQNmiJtXktCEXS0I
Jm8JiDjswn1XXqR5mduhbuPBMG58rkJlZmlBdTpi9k+NLZDdfqNZhgSE7FMc7qR+
3DFI1BDbl775IssTb9p0Kgq92M5rb1t1ZPvwCaq7x5rWeHT1nV4h892TJGaXTAF+
u2z3Hq8spa4JNY+8GtiKPL7OjyV/bI/mTSaeya43yDmp/JlQq1FmHZCDbWXrCN/L
zj7Ib9WBWyxV3cBJmejnmkircULM0wkpBw5KO2avgs/8PdTQ3yPeslsYrnwRgEKL
Xm+BFVj+dbfqFmz6/uj5Vjz7lyTWYmyO56V3gqJ3Qb+Kg2QiJ4iDD8fbP9BV4Du9
VRfxz8it9ZiEZH8D/PmgcQ+OsZBIhvmZneFs74hQ2eOHnTUJAuBJkeNstuiNUIn8
eCaqTl0yAzNbRhwqmgzkRVZRIVRQlLiiQ2gm+8DPw4HcOyqf6XLVXgAHMz5wHkJv
LNnkD4nvao76fGYhITSd5N5WMI1ZCcJF6P4oA0DbmbLFWAs1MF9CX8uqYSA40Tdt
lxlG49CibhVHOSLRJEnVrG2jar2nNlG6B1dY8SmOhk9doiPsXGYFkg2j+HD//CTu
e7YlK5Ja/P3CNth/V9i1ma7vbPCY2lTV8KH+V25FeuwTHrBu5EQHG6Tpbvoliztc
hE+bCaBdKTuLYX/mTrizgx6OIn9G/cSKi+abfd7ypigOd0z4sz1W8rwBKt8JJTUe
c8DTh+5rJ8vXEPoNcfrXMCSdkKAffPCtjVgVsS4Ia1Juh9Vi35vUopqYvzW8Movx
gzohbBFND3lIn1A9eKJKqlutt7iU1FIo0SqtRUo6wqPsrGf+7vGkk+RfC829o/ZZ
Kc5jRgwpjKMsA33Xzj6pDsc26LD+lSNxysmNQTlZKJN/xmMN7vk0hEw8RWOHRrpg
dJUqGjSCSvXOyI/O1FXSyJUc9UGEABrZL/DY+PDZPOr6A6X2QSlkzz+8QqFNQx7U
+V/PFVexIagDk+hAFxqWQLhS/prQd20CTlpEXDSWDzT6PjsVLr4RYtwk/XjeDBUn
oUiUGwPZ5uaS6HtwhbWSFe+9/RMgb721hS3k6Qf08R4V9syyyKspwFvca+0103Mz
dve5VgYqJLrBv+LmgFe5sIgnsqNYD+QQQl+5O803S6R+nqcfeIThCfpVnLlU4pTi
MQt7SC3+PH+sXdh5smiHb0J0zgQdP0Uj4i7PH64Re5rZVCZMUMNZT0HdVkM/FeUQ
ciM0qCdiIWnvajat+Lr0GdAGmNr1iyyyK54kY/MSWKMRWpfNctAb7aKcydyhIwOP
YcN7sfZmBwPUtVqoZagFcgN6G5e2EoTKTNojH8gv84IOnj8WhEKPlNtTLiybqUAv
Vs/yzLhMZhsVIE7683QzS7n5EgI3vV31z6GRN1BNbEW19+efUbC+QvNn4VLwadbn
Fj09/Qi1RP+lWzFuuYUEKqIaZOFVJ2EwrH2k1u8h1309iCq1Nb81W1xifo8Awktb
zuOm+hAVKWfnZKrQEhHo7I6WsA9zg+haWbeIqQC7TrCq0vY5j66/g4h4rM0u50CS
t69+sHGU7d7nypu14od9YKviIcDi+DwRfVRcTA/ywdD0A1+R0WHi/y9GIz30X0Yh
bhfhmomNEf/oOao3vWi18hfyy+K2F/gA+2qSglKHgKLsfLAiFhk6vSeEZUgERfmE
fjJCMcm9wX6nqoSJzT1/3va7eGNSaJjeG/e/Pu9Bxx6ucI/eMH32CrUYlPMGRBGg
IcFZGkawfU37Z87Zox0sM3L1wRGKybzeyEG9sunE1lYO85/XXWbqu3iilO6cVGxf
U4phNg/JV8O9Py1ysgX6wApiJ6asH+BrguiGZD5biU8whDtZX5iKNZUWWfdrrx2L
8Sc+3xPEaCQXxVxU+mgmbpyG7lDPTDgRthP9E3PlY7QEZfvGR5pGhAHHMQVrk/3N
w42sStubBOGVg8u7LTQ68JZ80pZ/Phw41S3lYgItlJGaS9WhVypxhY97OINemma8
aXHxxDZ9ZjIOF9M/6juAa1kjKMHPfjnt73b8DapHM7njzqaYSTJBNEf4UcbyEtdU
Pd6raB7kX5LfShUBn7nTWjBuarDS/cBDYGEuMd2oSuu+0uo6vV3lW69T5kPiZpDr
BKOm4j7RmbyVANmoQ2pvJeOHyi6ljFsjNl50ByqhX187RCiAZX1btizq2QCiG6nq
klwjDPuj6hrQ9o8SR3OKjXmv4deowhxP2r9KrCBFKMIOuZaRvZcNonD1x98+nTTG
L2EChsBRs1VuVM3Ow4ggkwDTM0Ef8PRTjyCY2qB8WccrX86+CtfHX9Zi54FfspO7
vPFXrHmyvltAMIYO5ph1HfRiyQv6Lxh4icCkHijNUJvGrw7vLIk6Ax9CoDr6thki
1G2ERjoFP398nL7mP6V0hvW0XxewuoH9QSX0wKVT0EcQ4zBs2O0tRArptpPOPYEM
P4hYr0NGxmGpP5KEqXjyYCboApVA9xzx8UCGG0pCQYvu56/fZVW4R+6LNw992Nbq
PbyIPd7hfJLMNykNv0sDTXFAKp8vdkd/pxmls6wGbN+vWOR1uezedN6KVQE+TTGq
nBHEMHqo0ku+quNMTsE0K9XCW7l7LLm+kNukjrBFWaPQkQQ4REtUp62wJZ7UMI1/
ghcKDQSCy21huHvH3UKejIH7OLojp/Z8trpzB6xd/twx9KAqfCP2dD3XlmPsRzmU
25+EawNZXSj51wkQF+g+BtbqzjNNBUZQTOURYUGLzVcvhOisq4/85tk2zuUTx2Tp
NCOwzII1cDvECY5A/70H0U5RgaUaqjlkt2+gG5bvSo4Gl617+fXmPqGz4UEWgUVQ
vD6gOCWbwaNK1SUN+o3rNHg1BQXiQKqCe/R16nEbkINkSZUuXLDL0+gnxCZZbBPc
55fPun62x8aDHIeZAPK4tOQhbifr8rQS5ISV64XWq6W/oyGLSKRbzvlEHPHs83Yj
DxY2isOP0OyYgnjg+h5VQTTJSbHfLkEyRTEZDciDW5xWJ3ZJDkEO4IbXxniTCm27
JAi5puLDEozqkQQ9oKn6qW8T/U/OgK7NTOHBv2FljsYf0wFse8v2d6DLstXl2cyS
P7+Z0ka6lZmNZsCAAek+HrdbdoNED1ZAm42tVAg8knl/bmB66nk1Bb+umhc9ptCH
qfV5QyXevyA5rCS0VUqr7ZdiWeOvoZx0PBm51frr1ajb/nrqhfoJ9Ydgc6jLK7jr
RkHrd33Nc/FPqqdvjWzLW49tQgAtdsAScRNBpqtEbu6JRQ5bPvtkdvl1MsGIvagW
Q42KpfADUlDQr0SiFVfxIkf/Yh+7ziExRRyjOQpXguVGCy/T2p6WZ7cmOyMp2XU3
+2rndkB00vHodq86jv13Z5Lu84J5X0QkFgistotkZksNYcUxblcpKtG9tK/64VWA
oi1HP1YMmkkIqvCK9Q3Hzks+W3CUzA6npsMNmVpI/g2KuWhCrUPOyXW88BNItrow
8eduFfyxEvGHsnZ9E4xxJ8SD29Ymf7biaknaG3fW+m/vL9TaQZYFEEYAN+x0Jz7c
lPCh0pq3GdipM13pHTJZov2x3y/5TYEpxJn2oDt0G1K/6R7VRZgQherZGktcgy3u
CWCJC+jaLBL/o5czGTKqnUQQ2TX2CzwEmo3ffZjgRfxS1cW8kQ7bt6fP8YqFJiNZ
Atn+RD//uww8kaMZ7uWWrg/F4hmgWqsZj1aP2MVuDPLUyBBMPewlBvYGoPWE+uZF
srSmzX2qxCfTIGgnQDGzDSC+qpSLPj8SAW5vFqjKBwCqX1AoA0C5fbXgjZs7Ohat
+sH2jtjPm0AkmLCnGTr3tJl/a1+8dj6v/skw/IOwaFCVmM+z7a+rUD0HiFYI6Ub1
0HHxO3U025iwokHPC7RIFSO9d3MVZiFbUzQV8MU3//f+3p4CgsO3gh0+HUq/MN+K
3pQMamRgcPGFxubI1Pd/IPCOE4fFaWaf0yfC3ZnzuXvZmoYxLFKFY6gCaglGahB5
gaUaNp9KzdyFoknrVgbZJdl4AVp/zY8mCDCyJNuup6NIQNJFEnMQ1q9XvNuLlNr2
m7MDVLki/+8//zca4z42c3JH/QiknKO1jI7OTjiRLVG7eQW2lgoy+DSBIk2zwLQU
8hRZFERg3w80H1hPD4rFQauyBKHCiklKq8nvFKH5brw2IZtSRMr8ZRGjOuXM+QVu
r7Y5T1/2EnfkoeokgljOBuOXtv1of8Ntsp7EcKsLSQypj5bbgF3bMJNDOqvEeu0V
GfMjKs+Pt67Ef8DPhjsQUH5yL9UwAmiSUAJq0/+ilU5BQB9fJbtwQS66kymUVw6y
ZAPL3XS0g2gITNcRQCMtObO4rtSUFcvFv1ZtDSBsH5QOWPXbC5XD3b0Qc31GOBCz
8sS0bnKahcBXXmmg34YT+WTwLzuGik9g0EMlbaLj3lXhQYp0iGpw6t1e0RaBg9s9
AKsvi4lPU6gt6BqSlJvzGgc9oBW25cN1MQCheUaSBR75AAUUQFx2NGThwOhVk/5T
6wnchaOCWwKUucbqFZ7qoUr1fF690PBF86TaLy6h2xyeyeCX3t/3iB0VNdMUoY3F
94NH2wS4otYDMEmCFRAM675YKsYrHUKgOwC7MzyfAv3eE8KMrECsyorS20Rh7QLh
Hm544D1Nj2fKDfHP/RbN0dUoB6NnC3xQcBnaAaBpDma1jzofDTVYUD8QGdi7Iqj/
NdzLj9S5lOcRiHSOk+y2c2dZIrfd3ELOVuWc+JvyZlMpatuf4zAzC0N17CyY9ird
jutJH9zAfZKxNE1bGCQsrJNRMTFIlKSiS8MwYUI8kRLvwk1QajV6tz86k5OLpQ6Y
NBkMkh1lsc5YT8auZENq4g+UKY0qQwxRGHIuvcvnOzSp23Scp4B1Zbo6B+YGDC48
GreY92gMNYhgSi/rrtDDB8Cuh2Hpe6fCwOIxG4gNWy64OQzs72OsiWI0RHlkgK33
ShSwvGrMd2QZPfTx5icVyz5EEcl5zJNqdV/SE3DluIPI1RayewGcSFfiNjGvOi4d
1JjyJuQra6wg4EDfxNzaOaU2pUwJ0tFyrDdZHzRou0Sz0asEeP6vMtplmgNw4tg7
qJI7U2ra2oHf9WzRjkgCuEyyg80NBNzlTj75FJaqX3DGmiwoiLmlZ3C84KJC5hFc
jEKRgdWgMuVHBiR6W5ZPl1+/G8fSDIxwbYtfnajXN0RP0yjaVJnpIbc+hmKrVhWZ
aLLf4roy9WFVijuIpff1PmLF7aHoKCuilM8kgLj3RzmkS8jk5ovNcDOhFW7EdDgF
OqdjsVnSWbV8A8Y4PXrB7HPc+qNg6uckqJGAlL4Rbg3vD2zyLuVK0f8RF7GbBuKc
vJHw2eCApxcCe+R+9wDhwPC39rnwu8rCRMwSezpZNtuak0xJXgqHjrZIzU3DxNQu
XVseg7MeDNbp8IJ1XPtIuWJzFq+7Ul8XAJSdfoFItQLSjtx/R0yEGwJe/4LOCdYX
JuS3UfcP8cLSpKOwSvzsT//BgvvWlQkP5v9WctBzV2avW7BDHV9rCgbOKp/s7uEs
fqMbPLPq7sBNdAxhWvTBiAD/ufcy5KteaqtKCZCBF7CPPYZPlZ+QJS0USz0zra0w
BYJ32glxFQmNOL/lqUSwC23hLuwjIFhTT85gMj9+SbVK/YVgrne2c7uegwFlUFt1
2J+fsbOUJcaD18shrNylscji8jOZOcXkmoue1nhwcx1U/OpAMHB4lvTowX42xJl8
joalX1gLJydtwrE+NNO5iVkcBofBMUSaJQC3ta7NX/4TjweTzeZFFq1j2u3xNL7T
PM59kIDaEe3uLX8oPrkpLkLsCOl1E3JQ4dG5ief2zrndicMvoQtS7Zs3PYCwDdue
UoT/DjwVQ5FLN1BwTvYQk2aBsSwb4Pim+IJ2n7YiNdBdwWCO6HhihpS18TEoOk9Z
y3bqZ6qE7AUVCl2t58/rp5w7py9sE3A5zdg0FULMOAdp9+dRofjRqp7ud5lOq5HD
PYJjKfAWZ58w0JGQDNU6qXd4xpi532OPaaxIHgsZXVKyKut6HLKA7leKLSxnFw1y
RLSc95Apvsr/zpw5dynts93SJbXjuPs3H8W72pp5gGotJ1/tuiVTBN3n/8QSKIqA
rsZCqcW97DO8l04RoIE8OMz2VjlNpZAZ3MznbDfErWtaLYz7S65TIEFaHo2wgIGO
EPx8mIcg2pnEjCxTNfxwGMI8T/DNJqaz/YVgfDEEsdnecWgduCRu7AhnZDTrBOfi
DCwoZLzggfN720+3zTu/v/W0ryH98amJeq1t28MF31M/bfSCNzbL9dPrYzJ++yW+
7EJupt0EMOur3knOAFRoOj5iR9b8g31mvk2eTFfH7pmk/UrCNsvbG9fM1YzpTtvP
gFVPSjKkB41Y9wJmoPVn6m9/zMn72/IvHDC69zNDOfpVKV1OpDMck09J2W29W4x4
RcpqKHd2fmAxJcNAcEJSw03Wb+KBHrndd4W1LCxsAJn4JuP4KRrGhnoy29DzDDmJ
JjZ9MkHTCU6GuxEUGc7s0YtDcrKqpeClGCFpH1qb+Jz3Q1Es4kzxG4ExzJwlHOqj
v/IpxFO5WTgErFYz5I0EQ6Ipxf2AIXi1rD/UvviVGErftXvPUP7o1OEeI+gkGru5
KUpo9z8yVodVFN+6QOgpRbO9roWx3UxS0sq0sGBVsK6PwCy4TYtiyKryiW+XWYna
oyj2tEXs1KCd6oQ8Mii7EghNpHj1MKgO1klVYzmj4NtHT2r+2GZT3ALC0UdOFGOk
bLQrpOUy0EKh1KF2DPTOYtbOjkBrjBvS7OW1G+srHjlJn6EYNP+H5DqUE4wB4VEo
fGo1mkVmCxIdnZ1Gv3AkdjVnncVUNNuLZyU61vmgVS+KkKih0mag1br7hCYEIg3k
rFfVmqNPGWaVfL4QfExqd+1Nt1POKRVjQmKcR7rfTl4Y99ZjQaPw+Ic9tfsQ4x/A
WLMhWYYJK3e8gTHx5umhFXT0DSqcEHN8LAfVKKQ4torP5wO+zYSrH2+crc1P3GXa
DcJBvz+8UY6ZEhE7SyfEsVgmCmlloGFlfrEr7uJAcyAaKDguEeaeAGTHQr3dR3S7
ZW1maHcHetg0W4IvZwDVD3PlBxWz5iVxj2AsSIMrtrhtvG9VwjDmkFr5pUwclbtY
hT/BmJsMYJ1LC7OOmBr8d0Fkml75RmEd85hNM6gAZy/WsRa6jCC3/5ASPsfuQOb5
d4jFSOkqFpzpiJEXRvQ0hsmKjB/FMS4fIH+UMBCHijKZ1WiTM+oNhwkVFx4x7IKw
reZu9+gDPmyjvsMT435GQNHWFCYPxfPiapCKR4Q1XCGrWj3vTgXGnxRMVW0bcozy
kUS2j2NdrvzWjmUosJr6DAoJ551t4C1LWW7aMZEWd/rzXJlhYJhowqy5a+4gYuLZ
KoQImDzrlWSLv97WdY+VTlZWFyR2ldfzsPShT4Fxv5liZk5OUGio4U/Lbb28Yy2V
Dv14Dt//TAAPYsKM8UyGzz0Euwr6BtTWts+QNIM5bOyN7GZPKOdbJSu/nqvZE1dv
ZRuM7PABz4J/fHgX9x9yFzaBRGy0kKpRoXd1ohlE42J7i50ybOYnvXTRxEGMTNYa
60JOnQ7LoPPoxdlRlCSNXKE5V1SMu1iQzUziWlz80JwOVyet2uuzGpFcSu887T+W
MQvYBFjZB09GdkIhJbcbxtGjf9Mf9rleSLAsxXVerm8gfrhY34te7XRbjMilUjYd
vgtRLt/k1xaNoaTritAfqQRzx7YBX+hl26OuobmQlSgtztQ4AM/HC6g1KZ8OXo1B
k9UqzcApGxOHVBJbeUgVgSnNqjRQtiE8ONOn7ie+FyOwqJ4vu59+QZlWTVRVqplJ
OK6g5HMT92b3ElVDHpZ79S4eaQ/eeMYjJGEbYnjm73GCDeqM42Rl8E8p3RaAR6hE
3XnmJs30+lxoxgziAdFNg0ALV3YKE7emFFaWGrNRT0zJXDACcq5cvyqzu4YT4Xow
GrjUQPMkZH1fwj5Bpgv/cveccdMgzLBe3UnbHmaNq2NGDvkpVnT1D/awGBq3AOmY
hLV8ZYnNNVtgsTHVRXD7mld310u+pN4UIYwVngFN4yzFhd5m2nco4fvaGVAWlJ07
XDjRsWg3OGpvrtJJ45QjiCo4NUF6BIRB40JhH3ufvQPsH+9SRICeTEqN4/ScfEnt
PvI+sSSYow1feP4YyV4sIxZ6NdNzcBIrD4DFteqnuzAdyiMWLq8lrKfLmLaXZFkk
5BwVIL+/cBH3S1zu5XeTSppT8BSBqY2dIJWQozSWBOI8FBHD7M7kgQPyd/rY6AsU
qD09gu8/o1JIClkm+C3W/ZP/QZFczR+U/sXA7Z8cOE1/1r3KIc1gfUdJojn8kqql
JcPqkN+W6EX0ZNgphZUyQN1eDF8TMaZw5d1KmtzEYnwi2cmw9kl+LvMapR3hRqDd
BiktO2M9tyJqzJVd2yreawXQyUXb6dupflEi/OGrWoVDQZGqBqaWUT6/NHPlCDxS
DLewoFGISBlKUrYqRlNLYOcf4eyWQadkhJDEgd0ZH1e5Po6dR0uovotv5Q1mcqOo
UxiVjtmUCpYPw2lIbiru1KTky6S9cY+KBXSoPCOfGvqXaT2TAH85F3/fTJQUXiVH
5jNcihe2EJmy7muxS3VBFJ1GLUv5T4QQR3m/VLKjUZHLlQMUEA4XhLdgW2CJUO2z
4zAU5fncSfxwwA7RJtXsP+aoqqdcUCRz95LbN+JFDbvG4ZRN3UwPm5lqZP+R5f06
2eaFD8+PRl/HKtT1PXg8Q7LgdSG8UnnWWdVKSYPrtOeFtPfaQjcIZx214pcI1okc
7REBI9jxOflOamnIK8nQfeH4C5f0p/5nB8pORoC4Tq7G8o6sj4neqGV6Arr9EOg6
WIzfOeP46UWR2hEUk4OZUgx1jbCkL9OPnOSkjuyQSAtKX4EX+LimgNBNpCZWjbBu
TyFBNSjMHd2hlZ9aPxke7R5fJNco8pEQWwK0wqiflOqKMFAm078MtyuVc2c10hUw
KN6GbcAXB0dm1XEqeBHgy/ZUOBGkemAdC99KS3+ilHNQE1+SnfUWHBLthQPnYFrQ
Z70g80qkvbmeT+2zPsJ60gOfa1CLCcfeu+Nso/PW5RZyMyNbkZnyHuURMIz8RjcV
X7U68N+VBTw9sRkrx0MDBrkIvMW0ku7J9fUbkFC4Lx14l9Z2OX2qJPMpr0VBzBTf
BPKdFc0FItyF7UgEGP1kyczoSq3sNFDuABMh0POXhacmeCWER9Cb1LLSZWHU/K39
srdxxFBTkoZhW4MHig+cWNWGXLqKJQY3lWfVANGPO8INILh+KSHAalIpCxumFsh1
+jL5fh0mrxvXmojjHJvYN0AnC3K/A/ujRYQI+ohMmTFwRFzV9GVqz8ZhUApg8AJ1
Pppc//pLTRFdteHXN6wc1j9XFHG9cmJk/tpY6RbqWT3QD+Eo6sV19mjI+Tpvj+b4
vPiu7+qpE63Ecohu0hKegG9UmyBXJYejt1jTZHnmbWZ0TtHFKzHAcVQHvMU8nKw2
prhqQBifOsue1Ushn36+7HMcJTfif8LPKqBXqgaMcES/i4/Uk8mrHeZBd0IT68bf
M6GGSuQKLozjf47OKpn6PB1d1hFq+GifMO0hVTtrBPMwk/VgG8hu0njI2dDP1pv2
Dr4kscWT93ZNXV/NUK4GLu74HTZAljPbQ0ACBUB/g0xisZrOI470/E7yNtDhfc7V
0RiZnmyEu78Dmeb+44bw+MtABOFm5NX8lmO+DAq7RES5snoGedzBAkHBGa6jAStr
gQmJthe11YGCzEAb+k1rq0i35LJT+jCXVWW5wMY8OOXfVlLjC5Dk9LCUr3j5sdVH
YB+th6d3tfcN4AB2MYHUEtihc/rCRQ5OaamrMbTU2ENi2VeQk2JoG2RMZz5X5EsM
8AFf1cIO0m/nvR9TSAx0kx4VI+JtiiN+fuVBWMX5Gpq5biQ7v53pWtD1lSXP2TEA
vtGxc4LL8ot0opzrQq009Vb/PgLokeTiKtRo3FKjkSVb8txOHqA00LbQLWQqwcPN
Ef4xtIp1aWjzOQGLDdK1LlptZxRzF/HeOYm7wLAhrHw4bxMem+xVnKVRYaGLmWFR
OiEciLJ90heNGduEoFltl+VKQyQhof/sTLnMSQyC1zAcXPPzsfrOS0caLNo8zmhX
2o8gMXP2ZW9ySxHCEiZcytju4vNAMCCsxdA3/ebTuB1t8S/2GkhHyIm2RCA531TM
buHQZBAPw0F0nTBfksf9tw9/qkAyAuUIsYAFRpeU/y4csGC9WeFff7/sq0kqX36R
DiiLM/QWe+DhtPJK6T+2Hn2/sYSa6Jb/TlN7w0dQYobHQ936YjXY7Ao4BExV19Tt
M/K4CZJ7zJyK26wJ5wR3EN1AHX+apQeP3iW0ykHWCg/6ot2kuDdgLp/139/QLKyV
GyCKQJJ+tv3YjiEbLWH9WEC2lmRwYcjyHmXvQ8tInD1LsY/T4vCwtnoFKwePSkSD
LAhrmAMh76ABpXH4iiSwShVzKk5IW7ysdYEZbj6Q3bN1yuA2X5bSgQKYdd0vYgGc
WQx8aX6NkslEyFszm6cqoTQjoTrvSvxH9BhkEJ7ic3OM2jRVpoJIEu9ikmzSuSzX
NlGGmEDBxT7HI83yJWroXs1/sArJsVhPW+jmOV0FNANDoevjD55gMxNcOu66JaPA
DQmp2AcFae1A+WHesjsAwjiUTM2vSQTFJHCB0gH+nktI5wqz1XPucCyTAYkIg6Wo
5M5bIq5bmDq28UC1dEOyssFU7J6N++4DiV2NAoWmLezrhhhW6xDVypdy7+0iIr4W
4/+9rCD9QiWXEnCnuDSVqN992hy9SGJmPgalouJuEjw5k1039aW43CzTlP0cBwII
PYSmUJVbCFtrcQtExW41+tpCvz+84kUGOYUbm59y04XZMbRf3enqaAAXfBtf6iBf
1Kby2yrEVZ+S3let7nYaA0Ra5gKfb/4ZM+vsDq27fqnPVmpofOlyNjw06soADUTj
vbuqwO0ivX8hWtKWlPDJnRjyttepXV4IINGNlTajmAks3VlV1kJL7LBq5iH2lazf
Z8mQletkijd4PeiMNuiAwSdmqJOpKMrLpdJo+hpUoUmd+97PlNkYkqpGJIWK/Q8a
317E67d8ZFvr9uYi1uA+e9HO5xS/KmFPNH97CcxubMlahbg9xl3VasjcCrJWYMG3
yZW8N2QCgSJVbaDfnRnu2Yy8+ROGGO/twue2kFx/xAL5VAnaWxlT7BvS6b6Rs1GL
lHLLrJBlc+pG5ukJ4zPxEBFY5vPjX/S9P4isAtbPmol3gZvlrylnz04RhMcAEKt+
NKo3ybmjoljNN4lV8y7x4Rp206KrJwuhnntysyFIpF/H3zh7pzDNcYpjhg3wqgDe
eOD7FeTWuOiaLd2pQefD7UhdzHvFXirDxPt4px64SX8wd9wvQetVeH4kJavS5T3U
0TQwirf+oLZw8WFwbie3+87xLABEeoyX8kW6WseXBMmuVpEkUgaq4dsx69sO/Mgn
vG3Hkko9xtXJKVsAB3cJKJCbLe4bsjC1YLTqQnJ9GFYkndVnKexd0VfnIoCKV63D
fgmFU15rOtEdlvRa4stoPb9/qhGh809Z/uMnZuN8Aw9Lr8mORERj1s9sxLB/SwO2
Bn6kYZVMp6Cxu6KBVgzMokEuO7Qw089gBhbhzfZJpzGBhu9eRS88Nnx96hYZNlcI
4we+2oJ0m57EqMfRcSwioHvCS17V6H6yTI8U4/NDSp/KXisaYDA6/14lnpD2qP8D
aZiIoG1iAe4oJ0y2fIQQmq+bsWcy6lFQBT+EwJsyTgQ4I36t6WM3GHpwtek0UOCQ
hfxr5RBasCivAUD3fsotM8/WhcSUq2nLX+vXLT+/Qjt/BDKdc+5IyIpuL/M7qVdX
GXqwJDIntN9M8h5V4PT3dgj4Y5k5xQFiHu/cAPhocsXMUrd69oUe8W5e1b1qrY+z
uIUmKt0jKvm1adXW8k3foBgMbtth1065VRxPnvw/FEKVaot9DY/Ydt2F/jMbCaQ4
qXirUFCWPWchF2DRY8hVZSjdJD6ctbTeKKHX3K9kvS5L9f5AoldAV2FDwr6wh484
WqAlbrrOUuYcEdjFoMPlZTKCMndpPG8oxkRA6pl4LBsBR8XlvxoD5GIVYS5FyLk6
QHzdS10UTcvQzrxK6dB6dbNtVih4MRqGSHjfq98c4ZppCWTMqAkMoVX9GVrUIyDj
2tsgog20aA45nJO26P/7THJhKOVPD0AZT+bZ+F5NBJdojXfq0pXoDGrtsDNLHu38
WrycDBZtqIT4g30PQb4vHtOvItAFU/ff3ZFgTMEOLc19zRSvqdJFz/EupLL4uQqe
SNmXPzTSZjuakz/ObJu1xIAi6ldnhCyr66/4B71x/CvvS9Na/kzKn2LC0/8wzobN
TrQVWGNGAFWzFvb5E38nO/E33eciTIO/MPrVPjYEdwIKVwxa2oeCGiSktQv8m0z+
d5yUyqEybAlpw0xfQBVJtX3b6utDccc/wueiuANqLj1XeAPr38lmA3mKratrAQur
lkXS1gmzpvA4guBWGxyiDpG3MkM/PpNeVSOXvKZeL8QGqTMQ2Mk7vxuA1mS8qZo7
I/McdNV1+JgFuW2gMjFTc7VGuu9XrcJWtKBbfah6sEt8Hyo59i4lk128Ty0PDnCR
HId36Se0yOZpOCbhOG1DQdaAGyS0eX9RMTEDjD/xVDH5JNrpvwtndufn4TN6LaJ/
uQsuCn1i1YESuMIfBm3eOQVCpo3EFRLA6isB6+0bXutSjf8//5YQa7a+TYwW8DtH
GJNWNg5nXunSb/Se1F/YgYJLFmU+Fs2NUXmjWxRxdAuFy6DP76zmQ5vsFOddWqpo
Cm+oNitzSIG3sjqxA+zGTga1RG1sR6DeFlHMW0j+zwA1+taE7UmYD/jsceWKjpjk
rzIU+Y5pVYcKClDoHmgHFGktGqJXFSj4ovjDtjlWpTQoakvKvpTCCKkSHcMkok1S
/m4s6CFeUfxlyxd70OyXY3MYIEQskFAUuHYXotfH8ILf/MRBROd1LYUbofkn3FSH
3GjyDB/g7gSp6PHzpn5eYWvvpmHJl4E6r1EMAn/+iXLCQQSOzFde7GPfkX/niJr1
HlhZ3ZVQ7eEua+0BxPfDCRs3Lwp4rsW9NS8IANQW6HuduBwOLcLtH7Gz9KPB4z7l
V9wYdDZtgarD/Xfpem9VqtOFuYev/Qt1u18H2pn0iDFhbLryYIuEhSZQP25395oD
3F2gm+4rY7GUe4mp6Za9Fgejs9uOknV72jaYU+DSrubZA+3X2huTj+raMBH5g3fS
jHijQBxlk/iUes1mrv2jwh38L7+Vyltra8SOUvZfRvh0dC0QfETzmtgFMQ0upwRn
0asg1qx+Ir5/J7Y2gZAUjiTTNXYFFc/ZYaveCi0+jpwXGXTex/PryGgRoGcByVX6
dsO4vYvF5EOpXqZgfA/NI6tZTe1eBMVtI9xoh57XpeVKHwg0Hnfdoxo7TkyQHuIW
rPkLDrGebwTtW1G1OBlaPORwp3mSHKwojCZtg06W+RSjgk1m26Qi089TKkKRBQd5
8wQprOgLKBA0aUz6taZYEBWJAz5QK5M4YhgO8FddJLAN89sBD31emUVCuOEuF9P9
IrA10MNUfhBx+wgEmwFQQDyN6P9SfkcJXWVIhrqQr1xLgOebv9XnEEIYQKnHadMY
/juLN2+Yq+etc/wILIGXUr9rNE3mbqcJyS6wAcH9KyxUe6ZOVYkckVV5JzCZV0oX
AJD7lBAizb7q+bsFCMhOSYMnhoCbk/kuLjMg7M3bp3OBr1sZnxOV1+np4YW+qEAu
Xa3TdWxZisgXE9Gu/Qur0JdEgK03Wuf6cmS3rYkOmIVoYCJThV8klmv4GVg4WIG8
F8dL/02s9bR0qLXLJY+dzfKxkBD//KucImhN/chDpeTVjd74/k5nakYhkoU4Zhow
Yd3e0Yaw1UqJWi2CzxvImS0GTMMNELkMaD1s3zOW/Riy+RYwSAASU3Yq7LBnneA4
ga33eDquLJBy2eok5+mhF/2grXlt2T/Ep2E6Lajj6dL7lrwm2C6YNADg9bOKJvRp
7tpIYZBM90wIHiMqFybM0wcfI07NFwV9IjjTOCwWVNfqg/+TI/W5lHUtC2dMxscD
Dkr+z2RYa2X1r+Ap3SlC/OmXi/+1feZkjOONR5jm2AhF5hf21Nj2Yi4dauAAAHAF
h1c9YHfaRtnJ4auxpTNdkg41YDdUsh3NWyfQppw4wmpxeIDT+VszqFL8q79H3sH/
nxb+jDY/PUrYgPOZ+m+ZBf7iYFxRDIN+qfVGxO5Z4RwMW4QSoiAmbkLrVs2MaNiS
QqNcttZaQQI/7a74UcHmWvGdyRZkmisXqzCeTmFLWeH08XEcEKLswaaLjVG8zTTE
0s2wNn5A8m7Lz22ssFjnMXJKgsNrzoGUsbIb6C42E1oKKKrwbOf8wfRXya1pnmJm
1cXDsqucYkCp7O867+fBqzW4nvsG0QQ5pNxu0lAIf973LhPZCJ1Vsii451xJmKeP
ArXNxrIDIfXTYYPi0L5JKaXkkE8wF+kf7BzHOSN2IVlTcTxgI5A4aj9AGGmu8AOv
lAmGa0lOOCF7c/uJdcYt6bnQvnATsWByXzQ8ef/Jn3ythvpaJYXIs6ltnckiddFD
HjOLUe3+GMXebvbT31zZASytykO8kFOeUaUV1wS7JUA2wlLN2p4M1DsMueeD1Hoc
QWxzj7+VxTu04NSFwjRdhs49aBDJLYIbPYKMG9KqQgXHHtQgMmm6fH83ZKI36Z1C
fsc3jhabc7NicEq7yIxI05MhYjNbHnjguUbHtf5No2OuBmK6SpgEbSYq6FWuxn0b
wYqU7uWeze87cH1X59oBie+fo4Y5ya5glIjRNH70Djgilf8rmlqBMBo4SM2Z4Wrl
Pb9iGPPbvKgcMRRTC0b14V3xQfOHX1nLJDHP3R24P8k9GgwZqqdsKf/czDSP5FzN
+NsuMcdUqP/VMDWWjxsHe/84UPBhRb0yU7kzd80BcwWKDHZga2KDi2w51vNkj1bR
AdXj94ra5XiHmIo2z/l0qxSG/jmDu4XvafxjQhIrCaP73t7V0IYh0AWCUY56OJh6
VXZXTRS//UJnnrkQP63OlE9Q+VRdn8+Mp195i0inUGj49i9geWv9DzUjfPZgtlR8
tfvDoZYEgUsWCc/Iicq1tIjdZHNw5I3/5Wvkye0uXgTg+OVG9YGWGO6MGJPZemO7
iAfSX0aiuuuyGgjHrBxCv0rfsZIrYF3t+9L/iwaOBwNBpLtK/KZamG2OAvgnvJYm
Bu6pE4Im+HUqzq/0+qDAa5AhWtLRcGj74PfEw+MGM/uOIXlW+KV1vkOI4fkm7iuy
27O3F3woO17vLMIBEIuD1hBxFBLWOEQs96bk1RDJ9w2I89wKXk7aTQS9vjWii7E2
YbbDdYidw+LXVe694dU3MNjKytlL2jc48GM3UcB5l7c0OUMROyxbRSneaJHOmfP2
xHPbNtw/ppwoNxxwcGIGnPz2nB+vi+trcYi/zKVj/M5/DQvI6r0YK9Ljdm3Gfzlq
EADsHEJbywCLDlIpSUbGWOhM+fPYf19bV0LKhIp6bDf9z/lvumcB9TvCwkakNYDp
DC+SicVSDIYd7rHJNO1u1yxtJRTVgR/7a3Z2UEkcGobCH4uHLvIwfOIUJT/32FS6
8cR6hw2vIluPwAmyIk6xL6x/uBDDmBOe4bitpoiWV9cq9h4oQjDE9fubPPaW8JxG
ElDf+IaAKNTY+Q4+jRJFEmIuZRRq9fcnFN5Za9Gfcqx2AahQ3VpnhZnRvDKF9nYT
MhAARnbkEcdzIozREwpqoMWfa+Wk/kVcWLd6AWRfTmk/3vRRjR1Ta4O98f0pXRis
8L7P6Lgdn1Plvr0V1uOVQ/t+4unJH70KbAVlmnhcmBBez0upMWZLi9/GmI9GyZMC
OEboHwffAFGKzz2DfcfWCyUwAI38eggVhAOdLfqB+7nH0EKbd3YdhTIDQHYz0I6T
zPxAvjjlYJwW6oO3OXb9+i8cmPK9RYxEdLj4mw9O7jDcKCVWMlLL37FFkURwgT43
0YRoYqVbvKB/RTP9Eh9o+es1FYvQ2fgvq7F0tAwpV5VtE9xRG8sHUyZI9sUKYkdc
m2ugs0MfBLHALHTBxdz2wbWJFkcepvhl44DcXbT0O/FYz6vFEi3lss+lYZuEICUw
brN13qOl4OA/XfW/b53RcbdEsIG73w/V4Gy1SboLmZypCTAEDFNFc+GMMnxTq480
TMrcwQHQllu0oXsCdB8RBnfYdgc7KkZHX5cTxe2bQLmWbK2d2lAXWosUhEJmXsrI
6hybNUMf3VgrX3KSaPJdmO+2TbwTXN2plYpOeV0FRLBq+hxad933cWuOmCOew8dz
V2WlxbUWfI7Ohof8N2RX1wzbEZcOX3zBwUWARUaVS4zSW2Q/EGo0J+VyGh+KGIex
NIVnZlyr2vjdx+a3/pAr3WHK/0O3eT2pqFUtRJ7dK/7VmMlnE8/4eYRzd/M0nmd5
uq2BQfUgww3TJ3LuAoNKL7UfXVukOF0Oi7IwF4T2hr03moqxlRGurytiQxGaew7D
QoonuJvlG5CCdz1cFuFR022KqcBG1XAKCZakaH2+60oKwX5GTo5zsgxIPhlh6fy4
YwV8FLoClQGEzPnDqsz7kJgE7xSzyvHa/1wSWLB+XeNpOJGc9ufoZfcZIZRXqNEZ
1YJQ7eX3zJ5BdqtatXe7dRdfaRiuMfCDy5XIwrj59QpAwtnN6EJYsrH0EfV89Qcb
YsNTBFW0jsT2D6hjkvX4CWuYyi5w1mfUpcoFufbaEvd5THKWw4vL7FyDD/qYgdcw
heI0U3L0yme00byKkDHrO58vFNhrOvisckaZVOpMlWWDT9YOxTEmws0buNZsY9f9
mAqX4yfTHVdiBRZxUF7gC51sGvjZx023vt/NFt1APJ7fao544Jc7UfV5+TnRqR1B
PqKbhpz6fvcGciiwLFfv59gM3A/Ai+dcP1boWPNKYD2dHox54zHmf1BnhZHUuRza
0Apz80i5Han7CxY7PNYtR/GMPIc0lqYePO0DM3ZzE0CpSL1U/rOoNfRGCrtvw9O2
TL+HN2mpnez6iU2B35+Q6kTf62TZa+PDqxpnSkUdOjbeCarqeUa84WfidqUyWiVV
H70bQoKOgZtkgVxSoTNVYmF6GV3d6tm2FNKRy9iaKHYPATf7ril2/S8292si5rFh
ZgChPFpvZtCV1QtOj3FOlpGCNAeyE4dlAsRgtm/fYxqTVzJ+rSFC24L5C9L/WRh6
Cb/v7W5ENIVAmq9vxiBOfLmr1N0xxpBYm4stcZh6I2PX2+BybpqzR0hF4ZtXujsS
I/SukOMLit2AVNECk2kWwGijK8x2QpIICscn1nHzepXiv+kKLWwwH85DT0818XnE
U1V/+u4Ni1RNP7qRiWKoPaabBB93/szjhrs1ryTfjmgkOHCmoER/VY9w2L3Q9ed4
lEHYw0ZNDh2VbhrsQfHRQPreCliDHfwQQ5xao9CLJG4mLvkWRaldUgd+cMnWsEtZ
segjrfM4ZgHanBgKhcswACGQMleNAhqSbCZM5Oppvto23bBstbd4lJIR9WKLRc0J
BMJhP5SrYzIuIgVwyyYFE+Qm69dClBlzKLSilJQW05pfja3BMUK4v39r3nhq+tme
6hstG6nMpE2+J2/jyxWUlNEecgG/YRRxi6BLe8rnhORmwhoqoj8no85NG8DHWX0L
j0brkUc88lQJEKUOjfdQAPCFy17m9vM24RbWg8k9qhquhdgNN+j5uKyv8UdAX6kM
UeCURBeDjJDI8qqvM6j6REAeLiuVm1wXDuUTtxNE94G94Gwson5eo+wQc+23zrhX
0+yt69RMlhiZtIAPs0uRjCn4fy7nk7dHaqwiyG9xwtdvdJmWFlRkdjuLCXY+PNPD
9wwEKGuEtAZM4T2er3EChLmERtiLsvb+/Aajdh8JAhQWuFTYj42NUmBNi/77p1SO
ZwqvAaO3qyb/7S9R99wmwwnSo8OpoqsnLVKTmIHMAIKhLZ/H3TFDeuDV2HrrKgZU
JLt9FwouZSALfIQ0mfEdar53ULHagLt4VJjASCnGuebB/E8XSjNyMo+Bg/ZlP9kA
OHtBBh4dECUHuW3tBbIs4vXt7ICa9dh5lpnAqFa09sl51J8i52bk5KT+iqeR2VBr
qTGrxfkWjQV5OGl4NPKYWHRxDPV0AINkum3EfX9jpqmVcl98dM0YZSN+rXR1dP5T
uk9Y2UaC2Zw8VdObaMsnP2HnTuIXxcrxh5Oi1RlA0aQDhev0Rl4yLLSrltLTtprk
nOW5pSI7wP+93Ja6Jsi7DhkFOwLnzRHgZMU/qAqYVQDQNBlIyQE8l7VwyKAjJ+yM
0Q09bpcWQE43BPJqy5ENzXoA7ki8NVq2N71beP8a9HmPyDihe97L8ViStkQCGfW0
VQ/jOSgnDR+bxH007yMBSL8oDYlMPcz0d8F4i5Ug2uckbrHnT3ireSYtee9j/7OR
GHz3ATVh3jpYCw9Drae9SjAflwq9IztFswXPmyW9QVmaLz+zwPSev2LEaDG4S+X7
rGIJuG836s8MCmvHZyOKDea0c00g3Dfb70zMbqd77ps2ah9JdyAl6ikLvs2DDeda
M+j1h1+Q+khmgexTnPvEVJ5N1oT3gilNNTq2xSEX3KHVc3jcE2VvhkR3PiCMXIXk
SDcTan2wv3U9hwYEkqokVPvnjqGxxh0ong66e/kN2t3yQSUJvyt7vj7A9eyhs+a/
8VEhEfMc3QCJ+8k8IxIFPIqhBJQL//+ZbiSM0bnZCI3lpJqwshB/djqlkDvQAK5s
NnjJIezAhOw/+HP5it/AgE3PYB9AX1BgIbsdPub8XhGMW35O9XxBoLSQPydf5h9f
Ck/E1woplfxmykou5ZSyxOailtk1If7hTiWuSB0anD8N7OZFdT8Ye5yCSRffgl7p
3sqGV0R3axJ1/Lb8AbMTBR9j3hogBIQyRGRMZesA98CsRKh7mTtkjhoZCD9tURjU
rwc9TPzyqfpeDp06LuJz8bqJJrWkuHYU82mKXL/qnxzpaAPt8e9DOc4nQnaiE3o1
sSvZxwRNADRot/20bsgymkXeqDByVxqwLXWmyHzLWppTrz+Kfxl2Gw49o9W/06qb
k6Nve5KoZuaJr0GZ0uePnisT1Gbj3ODFUX2ERDzFs2isARVIXE6mOkmB+sIKj1X5
U1SgId4/ukUbxgWWBzO2BFevwpbD7NHLbVmMHvs2YeWxYSF6hjB037o2aSew/VlG
FF2/5+PSeqry8sm/diQe1Pu3mShXBD5emnMb3zSPSvXnL6hTnHiOIfIzMd6RbiyC
B0fCl5YLFZW/pDRnkO0cRYvoj5p9kBGl6az3gdgWS+fgxMjwDfaAJ3VQz76dwWMW
/Tip8v5RKTV/JmLueefc0sGrZ/YIoq1L17/eI46L4BgcQyNcWSmljkoRLsoeaGU+
WtHni+iDfQIzw+XabEC/MAms4n/je+XVFLsY2TcWhU7OEVLK3N0/8yrr/fjJDRcH
Eo8WZ4s4DYYPzhi+WXePVqjb1VCQeV5yuTO+m+eJDisgon2r5QKBfw5SIJ7UROGn
N5m8/Jkcu73pX6yMeHyXZisyjBRc2VCLggNwiKRxWSl+F8D+TRuoc6F6yKIR3fsa
wSwPt+P3yY7c2vumi96Gp2J6jNBK6J1l5TI+Nm1+/d2Mu0dZKOMlsTHpfZaMbJPp
gBwOaIyGu6AfcQ29o9i0yM89Z8Riqq2ag68pCPnARPwgj2i1TwVQ6Hel+wIXBx7R
6CtPZ2lsT4264zoTnIdZ5lhxJRMxHDWu+T06Ge3PYbzkgmqUaY7jsRH/jK2358dK
31vK0AiZTlK9YT4gn2LMDBD3zU/r1r9+X93aSf1rLt2qzUkGKHdDkU7UiFLG1nL4
OWH5nZSA05QBESQvpj7m4kWhg3Tp6KI0UhCLuUHYMDBX87R/GAeZqZT4VJ+Pyl7e
Kj8baQXdrmCV3xSkjlVKnkxKgnTOBCF8xB9aaz6MfYRwnCEdgDaSR03hWNM6fvIl
bkbdoDv6sQbtvkTnmGTQ6Q==
`protect end_protected