`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
ddtXksX2+yylW5zu6QL2Lhnb2d1sD00763mmSITNX595NcHTEkwn0zB1Dry37fOW
FufOhVzEJp80NC5qZ/+F0Vk7Ik02dIR0elf3clrjeJRK85K4e3Hoo4xn7YbFUIms
l/8VZSb14+JVGURjfswrIyCUotIzlzVYZ6gzoZwDXIi5gQIBf/gI+KxNXPaKV+PQ
Ufys/12rjO6aI/pPlqSm0hCvftmBcnezN2hk1UeXgOIuKZnogjOsf0iJVX2aOOWE
6pD/psybjbnsNB6kH5uFTA5frkzIzkzl5d9+YDm9OyC+k84E83I/7/j+rk4L2dah
QJOvksSIzN867/4Qt8qYTQ==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="MvBXkzurAa5VTw+1JJ70nePUfoQXBvZOku/SMmg4TwQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
oRtzZL4VJ4iwysPsC8SXYCzXS8Fw2gtZTOskLcDV+1B9Nzn1zTyNtlo6lNICRmmK
ZRVu2BmCc2G+fmzynYlNTnSa7C0Cuel6FYpxCBlOuk3OF2tzAmLAuDyOH3Z1Yjzk
a0aHuoCdIRKv7BrZCdALt03JeUmXKPdOmIlkVGFl8yw=
`protect rights_digest_method = "sha256"
`protect end_toolblock="Jn9CQpRhJt4rnzZPRk+dOpzAubz7omckX1MrFd4p81o="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 9472 )
`protect data_block
gD6l00tciPUa6pDNTk/+t0OO0nC/UTtBwLB41d4inuAUA3i/ALrNyoJVcBnAmEQW
ptbcNp5fxEUJjnOxnedyZEuEBxWRieZFQnkRdF269oNy3EtIftV8eTvMbAlInmpf
A2yL9rKDcparWP9gc129++q9fgPRxNm0TjePNoW+I3uX0/nG0GGPb+s0z/iw151y
0WCFUN1QwnzaE8aDSOTxEpDq0WWGdFCT7GaGq/wtNbhJxjIKHdguHWRvw5KWnOOp
UuDvdu9PCu/kzMHM9C5aCindlCNpR630AXRu9Dccv03He5qebbADNECH+ndpAkJN
/+WFN6QFWTmZkg5GWqDfCGnR9kxGS5/zFg6uIiq5qpYbgh7PVTBDGK0/iMkVT02w
b7qvtK6a8DE1G7RAW1AF9FGzOlRBbHJ0iSBC3ToZjx27mZa59f+8bvhwqkOsozlu
Bqrxc/14WIFy33Hq8vBS99siL72JV9pSSPIaLgapkITdTJ0GngGV62ZOMsXq7hr+
HfiNAPEiOyYWxgELi0FIfR00+bkl2sbOL3NbblOxQDZfoXV3MdtMdRufAhnF+ub+
8b6RxxgvtbqUcwAnvhINbPlvqor1PMvnZkSLmV707BoWU/22BQrdqwmeGDxn6eko
M3TdFBLlLm6EJEKEZKqkS/e9KUW3thlbhuT4RcBh+AhmqJHsRMVGOSe9rIdhAFxZ
xeQcqr15M8wyGCXqhLng25TzQyZYIQridyRAfVYhX6qHdCHfSC9+DdrGf1dgxZax
38b8I8kyz1F68SY4eRYkNZyr+GdifYDhXjiba0pRy5oAjZxmxT4CE311tnb2xcKl
dpkqxvpEyGHRNmcATzeQCsC9aCxulK3TEeqba++0L2wbMNlnKcdr5C6Yi+3WvkzC
m/hGXTDD5U00hpGOJz8Gb+UQSNL973cpVol3+qMSCdmtayUaK3F7hj9IHtM46kZ+
88a4qnw+qkNCSCHi97h+cE5CO8WGWzxJM6mHIkapTlAl7JorSTmutp2VEukLuNWt
IQmlTDyWKJXZwoSSAVPxgtICfiTj9AriV7wiye3CzWcZrPlA5VHU/KkBUCsqkD8G
m6QYYmKuANCbUASsIXqAMhnO5KS8SAJwGmMZBd5sjkVAth0MS2pPW0X1rmWTA5aB
KOrma5owznCsj1+hMgF7jfYmdI6DoJOPBSxQINQeDi5DEChEWm23O+eArwM1W6F4
E8t80Z467547vbx02jTsdX7eic0xsRKLcXfpdRRXW/cQnd32y+eMAVqXdS7FtYcM
75qyQCy6BypH6aoOJ5Lz45A6SDUFySQo0Ohwd4w6Zh++K+9DFDxhLC4wqDsjrW94
kQVlK4HDSVBS/Mph+fZPuqAQuBnqCvwPIBnTqJA2LCryun2xfYPXVZO1H0xG4yxU
u4lxRELbltVgl3bg3toTqGfaoPdM1S3eGheOBYkBWl/OIq8FTy53j5qzjSf4VKBH
L6pOBuV8upHRuZf3mzRb27Sw4zQmKxKgWN2FRIdafSPb3cSFF740gtXWj5BbvY6A
M+Ip3lOJP9t6PCokjWoHhWs5LFd9THBpX2X+e3Z/hcjZSiwv+GzF0AKDfxoRiPTA
PIqGBrhPH6a55hhzcfKA5QTLOKcwsDISnJzZOhSTEzmoWZI0XNauh7HFvLEDKntf
mXTPAqYapACc59X5s3ycyamlZF9CPTnzBSUmmPdqqlHsTD2mta6gjRP9AyCuu3kx
EB/Sn7+KsqmV0ANtoC2YLSr16r9aQhvfrt1Ug1cCoJtiLE7L4NOEVJLTlyS3LjV5
jRp1Jk0oTBslrPmnHYysJpKR5PpwtTm4qwwLLf15LoSYe2wIMEj6q8dPfiuJWsRG
ZIQW8KRPd38zSLu8hw80mJKJbmVa6Fb2jKmfkklxLOzyOzHYuvbmaHxMN4t35rOG
3GHpUoWgUes/ajIRyS4+RZ013+TXX58iiMvI9p7J/4nnno2fWfBq2OPKiUmV/qo/
h3uLlKzeBgUNIAD4iylYFzPYYOmvrugSaFULzLWT1hY7r3l9h9vpgcYOYIo/CqHi
GSjqFngur+1PC4ptN9sqDmijp3MWkjmYoNPqATBAMuzp6gwo1OPtBcxpYcPd0S0z
/tLwjo0qDxn0D3RgWE/kq2GEA7Gj3WhS/pmaFv04OBAO+yVPQkSrNLEDwXj5MZRk
GzOU8TFKj7e34LBq4VYauzVA9MdrhGCRjBhzALg0FwWeMS2YrizxZ9z4q8ch7Pk5
A4NOXumJFS+EGNCQwPVos48lIKsU844aQuLkPH9qhyJCeHyslhkMZyleKxkJubz+
Py+Az47HM7COH17Zv6r0C+FQwk2hVWLre7p/p//aaOhe+P9cdRrLK6W6vVY7YQRo
9KkU4MX/dgbOnN7CZ6c7BjjxBcE/C8D1A2k1EYWhrvt6ELWj76mWYBr/euKctJUv
8WQXrhbjjHY/0WBGQ6n0hAfxIz4xye+k3IOs495PhHlbzSrx2RNzt1Qer/6G2lKd
UCihW2ReIPmvLzx8xPTNce4tRpidgGyJWxIk1/dZMhstISu9Zkacol5R/DO3OLkV
/kucSLY9OG1bChJoMqrAA7Otpptjm1seZ3Nl6rB6GGU7OA5HAnruFRXjDohMxl/t
54F6zjeEk3jj8gwdknjKEEbF100XPpZtwlc49t9EkahG3nXfK2sBu/uF/zGs4X7z
TVI8Xml/EPJqXili6ajzT52XHVT06OLxi3QB4eQ0URzcuBqwq1EnAljHLxELeNxo
wjLh+UetBPE6Q7V4Smo9UC6TieTmfiO3LiRHAo3lP4w3n0ik3A1ecr/nTE26th28
GESpS9hFf9MLlvmPYm26tvDoLPhQBau0l9kcD8yq98G2X4WiHmx+Pzb0IZkjNySu
ZgSGvJA0WaQzVJdoUUKNF0/rxrz/m+vUPw/S3Ril1Ud3oRhUKeuhfx3Nf18liK+Q
XPcZPsMVuL02BcxT255D1e04//i7bTZevQd7YRN2nVS0xEnw5XnP4WaRH9Rj204X
wE+Ozrf1KetitovWzlVga1Npt+FYAITogUiaATMhTovCQjsCUzUOjwkELlWxsypY
nzF+jC8xUTUh5GsBvrQRwiWNykiaD+kifY9foYbKP1LjAEivDQxNF4FLQj5+wJEQ
cgrjznxXcoWZK+DJIBJt7+vg0+ked5eQUYoysEPyVnfTxkv9PD4kfjS7Y3tDz57L
KT2MXDMZiN0OMo3v27SmKtcH2sR7g2gVTGOTaKw253FxikYxkQsJMOgeK/iY2pag
VzHROK7SjFsyIVJCsxhPqB2zmRhf84zCv8zuTGMk/jpaOp5rYMH5MhO0cLZOvBAY
QnsJ+ll1GewBt8kH58JpEemhVQ+r+W9/GfP+y7InGuq8zLaw5f3AXfBncv3RyXY/
Ad2i56ag0vH3BUskb8GotTj/W52GSxpFMoB0oqyK5gGJxV/uf31pC2BOqtRq8lbA
ZWspLF9g6jcCeAqlCIMTx1rwAGldGJujpBAcL5cc/gOL3QLvyXrcDGdYBR2GVbFj
JS4vX4NWRRsauzMTss/aGnTJekAXKBevc9JNSDfRiPdSotx2cgtrdUD/mVs6fdPN
NkKAVx9QC7Jswej84D5xYo0AptW1PmDuY/F8wEfePwxzCcqQ6tTc4tNyF2zaNpIs
38P48M+p8+wgdDF80By/egarYFC4aPRcbf2UrNuArJcKLLU2HlxVPgLNmVZ/vV1M
pjWqkCirkq1ue6+jjplz9z/MOqsizzmyHFmPQIqwKIrHSWT1n7VXx70P9cAMTNIB
968My48mmHI/JyROE288bIsOfteZXNEVJ99ctiuP5Dz/+p+Umjuq5wwN5f5mnXMw
N3qFtC5rZTp9YqycNki2v4c4SHDFgv7QNq9V3o2tqyQjPPTv3zm8m+YR4WYckPM4
mcoNxt31U3CmBgGCGU63Zm1pbfqphQpwXRtv/4+832e/eua+el5M1lSxACFw+tuv
re3o/sgEli1eehr+ZM6Hs9tyIcsOhtAMxmSkllVM6jlYwemEs/6I+TBFj11k9BAz
ja3cTJI0KOmMofehtndv08uOnRejIo+snZAOwcRutdO2AXMorJ6srP/MXtQmpJnP
mk39GIVY2QbTXNZtXQ6oGMpDjdfrgPIb4xU63qBVT341newRsi9JplwJvzep5Erg
VTqcUzgxmC/u7FQneXKoFkDzYz9Hpt4TIdij7woGAYvDs3T4HMjh9yc2F1lFp+Gi
bgO+rqdYFnroAN6IlaJzn4octv28+btH86ClbWxK8MUJkfrbCHe5tcCyRih7UXzf
WkURTtueE8NVESwSvfmMYuRO17yPLoIzbYisH2JkxyF5F3zQzj2cbkgFAsfVWEvi
XRMwrIbPCEZhogSwDyOpXH2aHwJK/MxxA1RPolnUYf6kvoQncvF7oFmisgjalhcc
xd3Fu5/5QvuyTND9qcMdBxpI4M3Tf4Sc9W1VRk3+Cb0hBmqNtzVPbzEfBrV51h9d
re1lVPzk/0nJ7VNL51zHNlmDHxVJRIjqYG7j6zyeG5B2wG1qG+iF49BNJXIfMSjq
dQIRuylhwYg4sPE0hJK+hpabhen11UMvEiafwL9VeCjVfUND6qbPU3y98/+PqPsv
FTZVsiOGBL+tG2OfzQgCmXGQ7jgXgZ0d2/4roV8n7GGL2xtxPclIU+dfKZuP0CwW
uBYYBjVRBq/cl2eMwCSGJ0twD9TjVoe7I6/NcUpkHlZ18SrtvMb/rJrwRWVyXn84
2SwVkNWH1i8Xbd0TKh9w0saS1DfxF+aHCUTpiawdMKf8gMZ0ISxRK3EQ0H45wcB+
mBBJxxhVMn7U13KLZE+ubz5bKrgP26/hqr0+6wSFRDfRGNhCm3Vrt2LPz2GJ1Erk
DlUT3zMtgA2YvYdw5SvZjbH6A5+rLZXGpxmQJ6jK5qcQKfcVXr56yB2lQVbjQcLN
AdkwnUScLx6xSPC5dLZwPFjOo6b6hYD+r8QEWnldt0uSHldnuN2/v81rKaYezTF2
R27lEh6wgYoDfzyrGZzyxqBYDDHoI1TplvdwhBm5k4YipJNb+msSthkQQkIM85xA
MX4qmrwl8GmTrTd/SwazC3dhURKlzC/F5NoppB1raQL7WCjzoYEEpxACI2gFx7vE
HaD9YgIlF9HiTbkH6hh3rnrxU3sURb1cTFRqhBuX6Q56GlMkPDahgo7pD4qqQO+7
onCuoYp6I1pc+YsXFbKeK0R7z9aZEXWJ1UYAFh3DmEdVZrBSt3oKR+V/qpHaXOa+
D/G3HX0WxFZzUuaO7avlOPNLFduDkNw36eiR0WO8Vp+KthcO8aWc73gkhqCLhloo
A2+Gu7DHAIseCGTGTkTjQN+1bB0zvGJH7TQ5eG63GkK7KZyMZfCvwy591lDUMAxd
NsxESJGnjTPf1rJCsZQc9+ZyFG2LsZQPTIFS0pcCnSCySgNxmNyxKohlypY+x602
++E6cAZHbMpWDOXYmD5UNkcvP7MkWUFVy9QnpgSBllLOQ0LD477Xz73QzPqW3VZ2
5WEojDNPcXoDKNDSADnyPkUsY6vwqi3CfvoB82JvI6Vdxq+ZPLmzYjTjKHHUVnpF
hGCRDFVKA8IWPUXgRVUtZUfyIFIIXH/MoHqDKe6T3KYVXaOEiGpT6PwcDdkKmmkr
kp77hUdXIBPKaSn7GnyKbsqybJkwMhiiVoRYyRxP32R6l2TWguIFNTqSJc3pou2h
v3o+q+rF5JT4lRxmLSc1epZm/GRGxHklbYfFitSHNCKlu0/aOGIdaPq7de+LzJJb
PhKgqR3shdWmzfEAOaCc3gV9uT6TlEz4QBZjUg79O2FHzBSKiePz4+u/FbBVfsgP
UNqy4QMA9JYcEX9GXX3cMeKjuj8vdHF4dWtMHiaDj0/TyFS2w3NXDULTcf/0A3Zx
iuqhKGfdPSYmFpVuqIdHyBxzEpCdqoDp/GQ7PnBDXz4uAPViFTRaKJEq+qVJuA5U
d5QYF6Xsh28m2f0iDU4d/NmtpzDaXQtAaYhyKy0bHBAH2rmuu7hDC3u8QMYu8Slj
zEUc3YsbYquijeixYT6XUOfRKey94xHzc2hBg4QzLyeUcZIdXoH5qKGrLEF5dtrt
4Jh1CJx1ifOqGpT+kSIzWQpuHFL/oeAdw+G8TZQCDqFLbDcb6uwpXUVRxkdjdHSa
geHF2uPAsYedEpJGuudZrrOMGs2nyP8U9twQpQfMxt2vuvyB2dHkVi32k83z3a38
oPlc2R1oe3SeITSde6wybbbM/hXbZm/WAvNX8dL3hOcc+p0IBuS9zWHZQs5Kx/hi
Bz/H1CYgXISCXZk2nYacwzatwZ+IQ9FEa3vUlKyOAmMySzeEuYgmDx56RnePtZww
VdNxa2GefEa2rIwhm1oEBHPfnVkjq1Ejc+bVIkMyTaNPUWe2jXnUDtCAk5vCwcl4
A6mkPtLl/N0h4PfK7og66Kzy6FGgaWd9vK154dX3QB0/SgaNmbgOKYvSD0JAxpVG
kl+XT3mpkLMmXW1oHogBz5ms1/ufSArpE7uRfF3TXNikhbTAGdT4gJ58v1m0NDot
rXZQdJID1WYU8ytbdiziv5dR+MspxPnfc4lNRKMK2FJLBpvx+XZDbyuFSquQdI3T
mRHw2RFS5tVPrnvSjalIDCERpndZ4wB9d07QSaKlcBXwHlEPfJ3EPxU/wDVEjr2E
ZrNB0SQosaSiEnz/qa+jN01oOg5ZCWrm+eJxlSIgVdvUhiKmFKTXZwKcH/z6I0tL
SlwjFKV7hjMNDBvCquLJv9KF0SOaJbUzlDKooXdRWmmPP4f4voBteht6phcMBNX5
L9O6i6xb2IvbHQVEmPBomz0MUi96gK2LDdDUpepzuDaYxCgWllsdB4g0pFsKpMSF
QTxhNKYbyD9Pzq2F6MRvz2DmV136hjBSlL1yfSfvSFRltx6oX1HZx/691IdXsOQl
/LKsVTfpRusERsjuBwR2UCNulhUNhTGY04+pc+6a1qXS9OeTiKBlob1rL5YV0eWt
TEROsuNdUPdf/15gptBva+SBI3+JqAEBatc4xApB2v+pX3LTwPyjdWWRsFBSGc+w
tcCegTHBYEbck7MIOK6rmWx8yL5jRr4v5V0tEnMSru9bH95zebfnXYbqHPRZVadF
xiaxfvlZ++jEmH4YM8sKgbwTeyyOv7PZmW8w9ykxB99YuPgmuLRrHT7/Z/Sp1gZH
U8YGTYSnhZhfj+58XN9/QhqKXhws1qIyw+C06/iYOROWqUYdEzLfDaSB89JKxs2o
4NPwnXI31mzNnGx0pF0o+MESlYXsEYG2NpC7iNO1d5CEAIALvC5qhjOGHba3yYLx
J36MsUofEeAxLb+bgoGPnxyu71xYM1sF/sdsp9d5tbcLPKrfMTuFbMx3shafu59z
kbboF0uqeOZY4OLTEyXUP7Es145fn6H77x3oMOwYIZpsycAU3mehx86ZH4h8gdQY
XZnqJYJDhaUab46o8YHA3nTb5sAI3OO1Ug03n8kDSFZ2WR3fYnYhSwPAuo3zqGsj
jA6N3G8Autl7f0kpNCEJDUwFJphNA9Ryc/xTpGQWo5Vt4IB1QCufQGB29JkHRXwS
v3b4XltOHMjs2SgoH9lv5OYUxBP8fXjMlXk337pbT3EOxUGmqRGFMZ8hCYpCe+hM
XtnA3ceInjMFVsr4M7KcHQ+W/7oDAXD77ZNzYdlYT6uSED8nivNKPpz6UOehCKAa
ip+CbW/b6yjZRadTEELOdUhpJ0AvDmyuZltFeXC6/PLQHn77Hj60cXx1DPpTGFHD
J/FIhAZaTn3uhLKSXxcHoyCRdqEykIGX66REsKT6lHiWFX3il+6UIJ7daTjZlsPU
jDKcR+ED/R5/zdmlqbtVvNKo0KJMZnZOHFA1jFhT3H7DMcCWSgyZLKSnVur3CiAL
oJ7r0MjQ0p32foPsfJMvFFgOFca6l9vlDUCekzk/uMDMJOL0pF+zSvQs6/4LPRDs
tgVnDW0M7guJDRarvViZhr8XIViOo2IADHQJxkNvZLO7XEZxkKcHGMhAl7B057va
WL2cWxK3ZkDsto86zgQChtFYejQq4vC2xDkiVbbuSzUgODjH5afeEDLaT79DEwAg
locFbKn46lu0GblJwjB9YBat+I9Ty5M3+fRnF8gdwDf2N2Uh1c2uddKya+LywQ4K
RkN2AiYXKmpD/7H+wCkCt9E1uu5KEKymSVlwX2/xrrv46m3gXXja/4UIl4QKMXxg
rChSMcahiFwV8MwX0AiXhlur1veNV9YWLrfBzjaKUSt8d0a+7L9YarDXALnZOYxM
Q8aL2woHuQEP1icT20yFKslyp7RTLtX1dexx47LFRdo1Su81ExN76U6sQuDFddnJ
g5uVoGD1A9hJ/iNeF6TlGIF1cWLi6Ka7yOWVwuBqUyciTBYOC/fLYWstJU2wqf/0
OSS7vyN3+BfOtD08rU4jVX2/RDDZK7dJ7esKQb9qvGze2THw/kSfRb0z/nEAJ1KV
U9aJqG06jxKRrVBO+cp1gRft/xSh0Ewkg017jqLxrreNTZBvcR27JUJlA/3FnU9r
1kIBs0cpqyHoOjXaF4GJ2uF7SQ5sHBsoC86Pyn8F0zWiGASV5+iWGg8JDIdLJTma
FQIrBMjXmeQCtT+27I0JPsnaIQen+taJ8poT+/T60pUPFN6Sq+vNcJw/+fSfqeKX
s1ttBDJZUFiJQJM9Kt7R5q5r+s6XM9qgGwGlgQMRdkqo4wElIod/DebE4b8yLy1B
rGBvY0stfF2CEhqULVU7tgfa7ERs0TsGJpkhR9yU+g75vDHdBEixeThA/R4SNPPE
nXOY7zkjNdeXYsZniQqx2USYtoT6g42lOwnlVisEQ774H/Gtx/EZYxSyRA2br2Sw
GwgPK7s2AVqPoBW13FgAz2a91wWcl83Ui/DCjkoL92uzq4giG2nDbPrKgeWaKqJB
fFEx7HknCqHwg3bLX5v6sj4UtxyLz479d9kwdmAMJ2yfwFSa4sNrp4k3G5MGvpRT
WoiwrA9oZ1oKcr4GyuBdeaI9dyvunp+ej1w91M/rxNASnU8O84hOc4E1fSl1GgjB
SIM5haVBrlCabgzfXMgzz4AY5k1KrvBp56z1lPkiPb/JReftQNqEgojBvgliuYGP
cXBxkdDtTSyMWevHLE1s0kK5rKdXfJ5esLZy5q978PrL8HSCq6zNVuEZbakt/D2M
TQujsTPitT1D/hhNfY72lZRPapUueNr+aOLyIRgBNUaklOcidavpkJaWvzZTclcp
HvnPlO1Scobzt6ug4oLGQShZS3KVRBqNVR+O2ZOX6AZVDKoGfTS4zliyx88WKAkA
xavB+NZ8wPMRKrYpSwjtfJzo+OxSmZhWAMpqBF+rEsgKN5VAoz15MFNRxDXMC0bg
4b7P/iELoM5OyulXeoP72YR4mlgNHI1AACa+wMakkzVFChgAkgDOahYMcOJ0H+Io
biahGwMIzcwN4hrG/eGe+Mx4Qf+dpXi8mUWDdvsFDltiOelJyKK+vCMwR9fNxCV9
119HNRzlGP3KCyHdHZkv/ZdxN1D/Ao6Q0xt/N12Dcefrt6tsHO+IiLroUtuqW56N
AZZA5e7GTgosHPrrp/0gDZoxQCB3recf1QmDLSfYDSj4tl1d2IqruVtyFR9sTPpl
9ZX9XsptMt0wH3TL8n6nGxwZ783jaCHYSDZaB2RySCaVtfKOY9rmFfJqCDFl7ZYQ
mxUROMCJu7A78iKzItmN+pPOt2jovPmvZrOP8vswYqAQykIAlcu+tY7fQBj44DZ6
Q6S0YzcqoD9x0tb+HLKEu3WjgNUqQbDTBxZLmgH1Pcc9HORmdwgRkLyKj/KtOk3s
cD4yMUqmWw4AYyELgQeHQq5tvocW1/uqCoFpJ1dN2Vt2W9sfQfcIgf6NLNfGEKo+
UlZYLHOZrx3Xa1xcIaKwKoIJjRyx9hOHJO2HNupQMjVA2DIJaIKXceE4fseWNLNv
86waqLsdu16A95LwKolsw0wl8Qh+bJiWbRM1VdgQMvehQvibkB5Q10qK0NtNoTGr
0zf3Z32JW2LhLBvD1Usx1e/gz9G30YmLG2OmzyOlGJgLc/n6UunqRR3VEurhiAVI
BJMCeB8MJ1nPU5bBVPRHklDmFZJ0HE5d2sutGqj7sAmkO1mJBR3bIXcgnCzNmMbC
8h2wG1bZcRgrf0VeGWB0fX2s4RSmDnIj7oOFAGzd9eAFTnRgcaggTgDur3F5EvCf
pMQNWnnJh1cU2yWYvIzY85ywCQrw4SHkjUAGjaaSYvApiwLO5/KIJztn7aZK8elf
ZZZ/z1to7cL64yLnQtPyYsa2Q/uudDmQrwAzlS6AxmGlpmmzVIEEdysBpm5jBQ9j
QaGt2AkNtTlUCOdBObik8set2iiLgcBFN/NSxXWBWQvpHwwoUm2oHtLDx9uUnN4A
tTHIBbZGKHWPiJ5+9teMenhDK2CMroxEc3sBJujyAHJ5rWvo85jJKqWVabDKn9SN
MmPQesDpCoOjAnQMZ6O504i+sC4Sx5fpCM2Q5ijpnjAGslbZFzPOqtzkxEAacdfA
Uz2jc3nQ3Crh60SDtdJpx2EU7GCDvgg92X40y/Z1K4P6LlyRgtverPWXlwC/xCvl
SMvGTeQWjf2ZImRPtXDC7JncFVQNTxh1g8qCIqKmPxAKAft8sMptkZ1WH9Nhl1jn
4SKXi4kNOn3O62mBxicAyrJC1uK0N7i8MsdnfXVbUPb3TS/m1SQZlRgcjNBmWg3g
annJZgtj2jvH7foSp6wBZH+ttj0Lp6Az1IBb1/YOlrqmMoD/eTIIHSgfNmqyG1vF
DcfyW7gyglD8prjO4Z/Bw/4F+JzHl/sp47hyozegLkMrHhgFcvya/goDBmmsia+3
4CHzSnagDPGq3KH7Ruk/VMKk4flPUGgMapZ2KOYlwtvSj74r07OnA0UgEJ37InZd
0zGv3QQaclp94OUqUBDJseWrYOfD5FX+aWfUkjuunW0DnCkPxi4nE0fPbYYdrQaT
DwzL56R1Q7yqwD1P0yLSL6CCM/biS59YJIOAc5Ygd8ppYlNr0utKg7xBUQRa+RsR
eFBaT7S2KuqXnx1xQrHavv6As+M447egMRuDf0MNUb1BM5cpd/3aK5J9eY/iqdAz
0x9n1Ik9nuCTmsN7AowdpL7k9a+wsVcGnj00zUrvap9PZgqXPKi14Q/HVp9mskdG
vL81cF5aTS2F2N4YOVcD+cX1kc6qscbb4f7EfEANzxOhsPtOy5sLtpVN90LhGx/F
4MG31HMuCQo8IJFzbud0Ag+qGjzVZf15qqoCuI3MPoOa+6x+Oy+bWknnFLfVJLKh
Pg7f0l+4jb+f6UafpFhPmYeU6ouMX5zwg7VpQF21BeNubd9L/MXU0uH2i7m23Tne
vopwDEseuuHKjbrmzImXz0Sq2Xom/vfAlsE6jUl0cYLqVWz5f41ExTgE7nDywbzd
p5JmYXwN4pX3vRbYSlopXMbGl56+NeMAcz8BtTjzk/5RBAlDpRCdQowQFrGo2v61
lG0sdaxvjZYnRxAjF85ObGSdwpCHz/7XPKOuBYe0JXA30guKxxQkLDxQjdSBdrcy
O6tdbwqAE7QP55SJBnAcCZJA2wVnZYbDmxCptgl5LW4Qz76CI/lfTGWs/NEBikVm
4/nWcG3zEX4MirW7RBJPVUzVcHph3dc/YZ80tBt8XA0zulLwR3txfC7Bsd6NwgX0
GqnvosWgmkS3GjTtZNXt6ZCX2OD3Kf60/k1EqJ2qBKo17K+kjG84c84XNvYvcP+q
DAkaYk7+pPPFlX6bFqqcEldInywyi/qaODNsRjr8kGcv+Qk97B7L/+buyClPfW7G
PnK1h1dWn7dksMP4SW7joOPopdrSwn/7e7ZjWE70DUGFpMZaDFwyYeXCiC3lP41f
XuOhsvcWQgYqCeOfbw8JfFKhFOA0+4+e2lWtfPW+E1ayhANMRyrunufkgA+fWw+h
MHWONDID3TKbo5/zbBkVPPAMH2aLoiDbDVtH4b7UTx0M1pa30/hb9S9mmtdceBRt
ZeQ2iG6PdztIwTPKNIfgQuIO+SR+wap1sV1suIuec3StSiRyuipqgfJDDqb3LBpE
uJZoGfgyhaANHlFKlQhXPJKkQsUNEdNlrq+umE+77stBG6c/qo3uD02k86o5pZaP
a/xeCB1DdhR5k4vS+eVH6eFaM0njXKiIEklLSOAqC31Vw1JwZAUwsEQZyvmqk9a0
8ftiMhrAdRjtNETdXyUvQyJ8b5Q9qcAn4iZ2iDURQnno8pMWHWiBb9VRP59lxbQ0
giIsZQTR4lK1Iyii+v9i5XMFjQk7cZ7DqYQYmWm7bD2jkqLgBn4pyBP8FfSP+51M
XxnnCAd09RVVugPLg2CYvj0keDCLrtB7pY+wzVlOxioVxDYT2FVlxB/5SmyReej7
f6rNjZgDJ3o8VXSgn/wzA1q7Qu+wbwdHdJ7hoKyrJx0Y7i3r5GuOBMproCNgIlOl
sRyjRycqfsvf4o88fAkSms0jBSK3jGb8Fo+PM4K9+MBbCKIoEHPZbjUls3S/N3Ai
ZG1Z1fL6xSOJL7waZQD1cqo4n/OtSfUBzjqT8T/lOazQXmsZ4dEVwP7iGvfEITjW
/dIf1nfRlb78YQ1G6/RpHgMRSbK6ekCVluqnfK16HG6nIskscV6PwVxeGQMXdmK1
GwcXBrYhWx+le77x9gKWnQ==
`protect end_protected