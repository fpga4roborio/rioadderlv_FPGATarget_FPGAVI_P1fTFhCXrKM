`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
ddtXksX2+yylW5zu6QL2Lhnb2d1sD00763mmSITNX595NcHTEkwn0zB1Dry37fOW
FufOhVzEJp80NC5qZ/+F0Vk7Ik02dIR0elf3clrjeJRK85K4e3Hoo4xn7YbFUIms
l/8VZSb14+JVGURjfswrIyCUotIzlzVYZ6gzoZwDXIi5gQIBf/gI+KxNXPaKV+PQ
Ufys/12rjO6aI/pPlqSm0hCvftmBcnezN2hk1UeXgOIuKZnogjOsf0iJVX2aOOWE
6pD/psybjbnsNB6kH5uFTA5frkzIzkzl5d9+YDm9OyC+k84E83I/7/j+rk4L2dah
QJOvksSIzN867/4Qt8qYTQ==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="MvBXkzurAa5VTw+1JJ70nePUfoQXBvZOku/SMmg4TwQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
oRtzZL4VJ4iwysPsC8SXYCzXS8Fw2gtZTOskLcDV+1B9Nzn1zTyNtlo6lNICRmmK
ZRVu2BmCc2G+fmzynYlNTnSa7C0Cuel6FYpxCBlOuk3OF2tzAmLAuDyOH3Z1Yjzk
a0aHuoCdIRKv7BrZCdALt03JeUmXKPdOmIlkVGFl8yw=
`protect rights_digest_method = "sha256"
`protect end_toolblock="Jn9CQpRhJt4rnzZPRk+dOpzAubz7omckX1MrFd4p81o="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 4544 )
`protect data_block
gD6l00tciPUa6pDNTk/+t0OO0nC/UTtBwLB41d4inuAUA3i/ALrNyoJVcBnAmEQW
ptbcNp5fxEUJjnOxnedyZEuEBxWRieZFQnkRdF269oMy5NrI2dcqrODe6q9cwki0
9ErWYRcAyOLixabjP7gnEOivOziw39ec3Dj+cFIfv0Ri60Qk/q2pkiDolQ+beW/F
0lbpVJysHt2d2O6V3Ck2V08/5+tbGK2pdNXenjS8UALaixe52PwiH6+TurWpaA3J
2tHxSdOtzSeULvhIyHUY1YIG/2ErtC201Ast+ceDoqLPhRwh2JUVsandqvC7NdnP
ye/5ZAcuW2xubJ0eQvJPvlxK1pVCSp+Hk0Ug9K1Ci2Yj6ttFLZWSP9eH/r+CRvf6
ACmrGyqMCD76wIgO6MmwCgQG+foOUjwNMuWp1Gdd0ruzUGxMdpgImDt6DRYOVW3s
aXzsudCmFk1MqMsMs2zD5v2/WXJGs82zCaqd2kOYklEhsEWbvqIBzwPh9ji7ZUeI
+32/IIxAz3QTBiZMNrOoGXovjAdJl6KMtWdyUJzy5sCkCHGguyz1aVlRrKzDeLM7
GTnzgtmlFUEK00hJF7aWwcbNh02VVwrqA/wZZVtzL/b3QXQ0MRbA18n6m7yIEMO1
SByp74yp8N8FK193ivGjbTWk+3NF3OYHEmA3tS+GZI850wXDpo1d4xO7RQUrtmNw
vgvs6gdJA1yS9Da1eRFR9qKbBqHObtYO7D1HC0B3+3ZgRL1ISYsuqKhq9Q1i471M
xziGb6EBWe2lmyVP3V4LNPVbOVtvSHNjsd6pcNRduYfAKRC5uIau+JJlMKTvyDKD
k9fw8E/QrA4Q0Pb44E7bzzeRV+whtjb8DDGpffNpSABbJyYfV8/TjtOjX0r10TMr
rRg14/nMiOw5IzgrRtqLs8UcAKd5WzE5dZjeojK6o/5NrN5oVIsa2FTadccAVlT0
LRMVPJw8yrNb8LyszbW+/KRhgyfhkYWzNE4ETQcUmokjPHplipP01CYF+iCXnmNk
BMJ8sKlMrDJpcBa4bdVghbiFvUs2zNqGVOYPr083yIabWCrU4dT4GqCaAid4UMOK
34xcLhgb4Es9ux8JEo1PMu1pSfD8ARWZOnZkxo7D5p0M+Ae5Cn+PucrRpUk3GTKX
UihZ300bX/jxB0bIyxELklcH7QhdwEEfEnk/sE082A/Rr0y0Ia+tIdXyFo5o9cqG
ic+puZoE7Dk7n8lHzWBYBHnbyIQ9coFb5LDT7PobX8vE6Q9B3sPZcWQ/yv+q7Yr3
INatCJNf7oMFwhRDSuz52PncJgOhDyWu2jd0hGdZj1Saj51fEsYTP9gQE2cmDljb
SZT4K26+cbBFtsCeO266D8brWGlPDESC1zY6h8q50/RFJHqI5mWV/6d35RUZ90TM
iRuUbRWhNzXK02GAnwHe4cW3YiK7InpNf9nbBgH0Zds60oln/BxtopkUmkk/RPnP
1gWdXIKqV5MTS2HReiUvuoEAO2GbW/IX7EtUl9IBHn9FV0zAzeKZvLi1QRrv0wR8
m5TVBs7lGWT8MeElymIincKomtjQIk4ijpTBoXSSYhyvawW0tVbMP3CQwGf1otPU
mwUq4HSyufrAuQuVXG727fWNi5vLwloixKSJ4MT5LWHESzp85saMQTUQ2wBrBlsd
S2WI1wPFBhr6nNv8DsEGw3rOjat2RHtrFDnvxlMPSQ8GBnPCh10kxMkGj6CjLpv9
nqPYEODbyoIKe3ml4DVNT0rbeutYKX2rzCEYjmor8uhcIQxAiQ8vh0hV9YlpPanJ
hCFII6JjcwqvBRDV1RE5Lj6CJ9rmAZQow7QThAd7KB6DWl7EG56upTEzq2jDFdX7
jQNfD0xXAhpUYbhMmGchU2HfWdAxhB1I5Ojx8zC1O82PrgYAqxzLHqg44K4ui+7C
uhTNHveM+1iCCOZBvBjFxpiiHPvSni1aVyzbkXrOpHmRn+5jLkCEE9G6+KwxZp7H
4LP7i2sLukJOFNd4FHnJPwKsNKbdQaeWz47Iwae77zhjD1XKUKdJwiyjI8rVBZzz
ysBZFPwO8bPO7NUNjASiEsb7gvFtQF5jqAI3lKT+aVOFDEGZQb0vavqFPCTfzrO/
2ZRu9tNbNsuVuUCdUbivz7/xbMLp9Hg7erldlorRSLzPpDnGo2Ey7ApGbkU/Av4K
fZOYyXV3L9NRVevWvjz5CZeC+FV9sUarBZ/xihEMC2l7CEVbChJHjKAdGx9liNNt
tuh+snIINpvRCjmXqsnwwB0QWqC1rDAidc2b9+3+uOUrR4GxrwaFNVK/pEEAB/bC
Xwl5SMD2yaDDAUKO6O3l+BC6drCqFcHwLqdEzk8prWyQsYVActqauUmIpjyS7TUb
MMQeKYNHw8+PWa+mYqmGOkcTFxixkRdRMHO5jNwyqJsHIsWHVrs5bA7H+l/X7+96
BKd/R13GCvURyb8meQxlH0fBy4VzJr4XmaO0AZ3X0mtncXNYx18fFgR237XAg74k
QMUpKF0l3htCCspNTq99XoJuM31Eke8SO3CuE6xpUXJwrccTMgPgozub64b/+YlH
SBHsqaspg7l5gH0/pOAvi0gRLngz6X8xWPXVhmjAZyTK4TCvQC96Zoy4mS5fZ4b4
cu7pWvp0Wb+RY9qcRKJ42C1irZzQWA8Lij6SjY9J3e5+6QhCW9/J5XcAUde6dt3T
Kz3mVBNUH78V47NcF4jpt6zPJ0lhFPUnL/8NjAWYwDwHcLcTo0LwGf16r/mXem2J
HjMVQ8HjcD5B+MyGyU8WP+HwzuJ7BGpQAhkg7SjSUZiBN3wtT133pfQs5mIvlOMT
/DiQ35O3/53aA9nb3NuSM2Bo3eqtrNrLC9BbWxnehDPowWeCR5go9hZPFJwDwk3M
hegP9Vnb3XAGcowvQOdAuc6/BhABMqDkFGPpCLaAWrqM6tV70BKay0nxwV3s5K1h
JKRV/O1oZWyLOLxIsELJYx+seQENfCR/jExmbGvIWYUmnJpwBGbv7stopEePQz8Q
XwNr8M+BBQpgFzSwGO7uRjvfmsgveF03wDsntp9GGw0uxgmNnF+Upb6noPF2NIjs
NyN13AxBO8+GJJpTIYWjeN8P3ioRN3EL0Ow/bt/1qk5DKTN7snKaGXX5rkEdrkV1
QP2A6G4bpfD0GEpAxh8Zkmgm99yYR3Sc1hUsB4i5uYoOpYn3O/I598B4Vri1Ifi0
Ih7nIJoZeEaTKsEzcTqbGoZxfmW+17OpHxH2lZ7IPLRsGNbcLFFMTrA3fNSkbt34
9UItFjf9a+X54bqqyeqCWF32nGLdLbQLKEFwac4MBK1tkHDomCpEYjtDInplA1KR
Kt2cVWVXtQAePxei3AyXPrX+7lsKWHxn4sZadJYAvyRq+IiFCid2RrFtRrtuSYac
pOsxiqbtytrbDTnD154RMQnYFJPsgrRqoe/NOGQWU9KCEaI88r5jzmjCWwzGfRzw
hzJxWgM67MgoHn9Um0TsfwtdfM41MOx051m/CsRoERmt7e7Cxq7PC219b6XDMQt0
qi5fFe9Q5fDl1aKq/LkeXdSA7Rm5/j0szhxWVP+mn7A2wkZjOkxjTzCsDPOqYtlw
XagxTa0ktPVjANt6OBZ47CDzL0KkyjNTYcbZyKsPbiFp5eTztY5LuSTz2LbfRyCx
0ZzW0XY2R3u1ww9POAzOg3aXhNmBNa7FV+oePBdjJNljKvzLrRNtUy4C4TaD6HLa
f+rGfGSNVrGTk2fh7lZ4pETiwc7/SFwkrhNmlhS/Tf1UNDGvrkAAvmcU3tO5SOWE
/834oojPOUFI3Ox7wXMu0SGxIHtxizmdIbyc71UpCao9lFpATKGpb3yEFMkRbIRJ
AT3uaxbtPjQlv8TpDmZ9vS7etbwgC0I16eQdkKc0sBrdXJw/NSmSI5XEjzGHL60Y
+zTreTn3u8i1/guFj+9L0l0c4mQWIl/47xEMJEhz7qBasKjUdH+eme553Mc/MBzd
I+xM4RfRA+3ZnKophZZ363AMWOG3pLK445Q53O+yy9GeB7iEIo+IQLmGXXUOS8z8
1GBRgQhMq9GfTvprq22pLAVGjm6Qs72PWk7da6B2R9YjuVbHAu9zSUlv20JXUWwu
Ddsu6/aPSuIwpuU2nqfmG3FnfELKsiIWPfQIUcBmiyy4CM270gceaFdyVRQe2xGn
4rc9SXevAw2j/75C3yaMyKetmEoPc2uSowcoIjz113uV26412o+070uRn9hEy0uU
YduLgKuVWPRF2P474R73G+iMnXBLSEoonVF6U6+UveHqwMRoM+3hRInUrs5Wpz6+
IVt064MnDkYWf9Pb7tijhtJZDGNBVe06qwC2DcP21YFcKVR8BJT5QIa06KQjfIAS
8a89witkucvySYTNnYk8w+NYWfj/eEq3aFiHlTopsz2QZM2pevowW4UKNN7l77fl
iua5A9c7+KeHLwp39OkLADoJvVlxf6GqYdjXqDKA0OnQpkaDBYMIPq3nYgWWhN4T
5APvcoX7dz4BM3gJ9/bsa5wD4+chN61OUHUZr/6oF5H/Y8rEYrNg9c0LnfeXA+g2
0l+GzqrTsp9+QnLbV/BwApzO1Nk6iVINzexGJCxUVRA1CPKpo91gv0Wp69fEMne/
UMZhOsmvyPXZXRbMeZPN/CKtC0FAU4+Bkl1Enc1Lb4qkusTGMKjKrCSACbQWCgim
MfsDYhJgpAS1Uj2wnZzpSW2znLLF2JFQSWdczwDbWl8VKf8u6ivzvU0TzBboaCFA
F1itYLjPC0J31d/WzQ71S0a2wu3x6tnFj5Y04eozPxNj9xmE+ew74NqIkKX+qKme
U9cn5APavTOSZX0ImAbMeN0vt3oKMc3OPYiwzDD7tzJ4cfJ2BbDyql0Y0wIWAxh6
ERc2XyeM9Q5wEJ/KYnNIkXmWQHdLO1Q+/7ohrq3ziixKQeAnjzorPUk0O5KL7Ror
fBw7fTmqxagmrFFZ2MxJOLEviCBPZFHvTg2YkXOZJXGLIe0iI/1Rfl7SwRpVSmwn
gPUgC682RAeR4+wmoVpequQdrdhWiaFF3mFIfqSRC2+rXuogVHuhVfxK/crVel/b
Zd5dfOyOfIbf7llwjKzn94/XBX5rfaWK7B2MWeV9mUUPnF6nD/pjJDJKHpTbxryQ
pEqf241L8Wp9wN9YrbIid3ZF+D1tKUhV+lYIY5Oab8Z38AC4fm+Ux5m9H8O/Zk0b
y6KLv+lvxl7u5a9GgvXymmU5zLr0TdbR7qOTIacCga+4puEDE6OvHJqZSIULxlaL
vHzFEnxcyVTL/PDRMox7ed4X9WtUVyXbpRFUn4UPYwTQPKGp4rF3X9cG5D0BM+9Z
N+FUrh8CxwWnql7MaGCzOaG1tCQFl1DE/aJlvyR757Mv5nsSGm3YFzP4x+yXsdfN
TQXMn68tDnTAkMXLluDplAqE9v3UDkNbIYtrQOlkeIj1/7hhgl9Wcm+Izs2yZHbO
S41vVTVtUmOP8c/FBSNkPf6MPYxGOueUJdB9TbMSrqqbw/k2+6bjjo7PEHes6Uho
/wtpelXdgGV2KIz0Y3qtdITqtjf66enX7UyncDajJe4eshjYhqpiOCwJ8LwRIUJ3
N+YSY6ya0uzO03VpLHDs2qZ9hqmBdbKt/jrhSX8IHhf0eFRF8jVZdppOXE0RBLpf
tQOOhVGoasAArlAHO/iY76e7d5Hbzg8pskgo3aZn7ZhusNMQhsfSY/aQqByBrOOf
Lx2S0E0kzxS3HhzMXCQxjd3a5vnhKg3uwVW9AnC8xOKi7jFd8PEr0gxYMkMWP3PB
+9ff305ZADpvxXAHJsQC5lg1rXspk9PcltbQ45jX/57hZLLY8HpkGS9gGbpRnEOb
1t6fAmVOCtVs8R0Tj/gX3uB3ff1V+a0NZ43QPtl509RO8NdvCkn7hpzv8apnq68N
Uj7hCt6XhZN45HQU1IRlMrI0vw4DgDzmq4XLdT4aSdCaHMR+6w6WVfEnXWrJWNzk
0AyziaMyXHmG7XtWSroz/DZr27+S33QuHc+vjLjp6O1jykETvVsocsTVbCA4s1WZ
ylLz3P0rWJaT9gjqQynjmwGHtYmc0pouANe6bHpxcyE=
`protect end_protected