`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
ddtXksX2+yylW5zu6QL2Lhnb2d1sD00763mmSITNX595NcHTEkwn0zB1Dry37fOW
FufOhVzEJp80NC5qZ/+F0Vk7Ik02dIR0elf3clrjeJRK85K4e3Hoo4xn7YbFUIms
l/8VZSb14+JVGURjfswrIyCUotIzlzVYZ6gzoZwDXIi5gQIBf/gI+KxNXPaKV+PQ
Ufys/12rjO6aI/pPlqSm0hCvftmBcnezN2hk1UeXgOIuKZnogjOsf0iJVX2aOOWE
6pD/psybjbnsNB6kH5uFTA5frkzIzkzl5d9+YDm9OyC+k84E83I/7/j+rk4L2dah
QJOvksSIzN867/4Qt8qYTQ==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="MvBXkzurAa5VTw+1JJ70nePUfoQXBvZOku/SMmg4TwQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
oRtzZL4VJ4iwysPsC8SXYCzXS8Fw2gtZTOskLcDV+1B9Nzn1zTyNtlo6lNICRmmK
ZRVu2BmCc2G+fmzynYlNTnSa7C0Cuel6FYpxCBlOuk3OF2tzAmLAuDyOH3Z1Yjzk
a0aHuoCdIRKv7BrZCdALt03JeUmXKPdOmIlkVGFl8yw=
`protect rights_digest_method = "sha256"
`protect end_toolblock="Jn9CQpRhJt4rnzZPRk+dOpzAubz7omckX1MrFd4p81o="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 25952 )
`protect data_block
gD6l00tciPUa6pDNTk/+tzLxvdHE2s3DQL3/JqqujQBC/Ei+vcAB8wM3doqg5vTg
mdfn9XB1bLOis2CVSfu295W2DNwHfMSTc/8BhCDRnTlLIX0UCJs9Za0+LoM0rMrV
T7EjVWppbP+Em6PkVKCwlmIQ7JKaifJ+Y+kjw9HCGboYo5074hY+K/CBbfsBQY86
XpZyvRDWHldynRDiChLubVfGjzO7PwT4nLR/HBiyWz/IjAyBqJbfDK71AaW1pD0R
wmVG1ks7W4+9BeRPEEQb8vQf9qMLQzIiyHa9NHPVUUGSKrvcmlOhirM3TDZNMtuW
A++6/UpG3ffUNwOHgkQeq5tKIy3UExuIqlPSWfYVtpnY+pj+x4ZrVPvEkE3SnFTy
S/An0WQQy2ro7a8W5NZKjWGn0Mzj6jxfNpPR1iAWg5J40thNXU8NYnGI0nuql4rb
fquXn22Yf0NrLnkRKwFCG8xtDURNLVgp7GdkE1WJW6HLu9BUY8rk7f2OWozBGben
Rh18pJ0enUNW0MncDnKx68+2/uuNdXJau5v7sKvc7R5ocBOs4eCRt6wqfvdqpAE8
009rSbTj8Di11F+d5fRA3DYccTun01Qts5Zv4bMeTlIW8TuJIwOKwtwr56EqFMYv
U7uI0+y0LTyV3JXXNI1ML6vQtlbAuecauRwk9n0z5cP4UrgX3sB91EfuZKEEQuIo
IL/RA5OpMTERHisSZtsm33dTjYwObSVuvv4mExXXYdRBmFFxgLAZ3keYfNs/oNbg
O1S5xR0p/zw4XE41bLq+RJBXtPC2Khyek0a49llBtzNm+P6Mo3oaYZS034eG4doa
UqFeV9WUKgCRsZPYitkPubVfwR9wHal7Y2FMOJy2+UHIOiAejqt88ycmMMCrWxsd
rpk4PR1zzv366xUgcec9xVys1PxCuT5s6bU87JRVvFUryXJs04koubEyMRSD5SZ4
70UrKSjCp76gnTRV+CTYnMGyu4qTtdqZo5ZmDFixYLVxvpMLz+1q+LdNP4jV5+OT
drRESK5vCghks5XpJKQtvyS1Gdmqkx17+KOOaHRG5lns4EdRPzwbiufA2F5UfLXv
JtRqsVXFVsQlvnBUcfFuF9yecBMmmV+/p3Pk52Q+/vsn4p5E3zrkxC4JD9/bSkOd
iyPqlhlyUVnikT8AvW8suNO1tP7iWlnpPQf1SJfp7r5pnu/vX9FCfrdFt7YCBVeW
mobHrTEqwqdihtjANjUPsN+/0r9td5EtG7FRyRsfPxql9DKPQmpLsvAwknzR2NnN
aEbb7P5I0d7Ev7geBHSKPsXiMMDVfkuDZjXIamSHjB/l1CxApd3QTKqvIWaL2bOI
PuARU7CqICp0svdFfMfrto78zl8HIF0mS3mu0la4zD9W4Ok28fr2e0EJ/Bn68VPw
YIVo9i9SkSluIOfajdunplKQv6NvnU6zuKd+/vTtF2Gnm6P4zr6XrodnxyC3CAXT
myc+FPs1quHOjwfw1pD62hKKbZrBJ23BTDLiL2NrAJN29S/533iVA8tvmbpM4jVn
Hn/QtFl4ne0iN4WRYzZknJpIMzhMgqvm5UDsDZwzJ2TM2NkmUEPZ56+FpG0me8xC
bgPIwSwdhJ9nDYfhmAn+xNGSMustJUW2BtLxLDzDEZLbehql/jDmFkafJpwv1EUn
xT6EXiG5V8MDcmFYmUsuwGFya294WE5FEyM8oqw+12CEu0gw7mjN8o9svBsuqRB0
Hx4qYR5EiPL54oEWSjxjTld+WuSBipyzxJiLTAyhfOwL5KCgPc6AptECYuFqUi+u
kEDEbOUS9+H3Ps4iLWlUbDkA4R3pmKXb3RaVCGBm9dpl+9w+8ekoI+mhPqHFqdmP
tZFfqhaGmMMxZvn1Fz8kPjb//sNgkHKj9pRr+fUkXAEARwebLm5J29aM497pzoXz
GbQVdAOg6fq71IA1uqaF+N2dfeguLwmN7JDceCPKpUEAMO99AAsRfKUcEQ9/QNla
e4UblMokFWPojtzs0bHwKE0Y+iTkr03QzAPxKgWiPXgT3cxynivLFfwolET8zUqa
TmJ+cVrng6jkYRWWasINyoSJOfFu8Wlg+zdXLdKzErF9xX1zgo462UUAEELz599o
4eOcMMSzq0Hr5BUUAvh8uTzMl2NBauCHNa4m8zkvQhGEMV1f4y/BZJHfSHcwwOVn
0M6/xBQcZVggUNNS+w48tKop90P0wBABJspNXGmQXHLtOQJlLOX9On9/LzoAexnn
mi5RTmhdqpTwEHUjRUpCKmr4hfi0xJu+r7IiSNSclieOW9Ir5V39+n2D+OcHKA/V
8S/mfFhpj9qFcLFc1nt0WSv70E3ob9fQZluoQmzKnM+Lu+4W4JUupW9r5iCJbkm3
s+e6I3Nn7OSHcVZTrr1TxOKyvJARYxemnJDINq0X/jfGugxL80LvxHZ+75hQGk7l
odmGGqCtFl6CIbPFbsIkFYHUA0N/04jPywnRqiiQn06qihXHYJex7UW924LeXAeR
dElRWWRxST7lJOPWslOFEkukHwnfuGsl8koOrdoiZuYn8MdJC0BYTnk9Uh0fLOFx
66N6i5+4bx8VclAlOvgVGBHn4NYrZ1RFoU+1OsovsMwZU9Wi4EJTQ3az8c/I6Pgk
2q5IL3VIgGhcNjmz6q0FD4MGAYmDnj3tNDen55/Hctup5+V25XBTILAPmjztnhnj
ES7zzKF4PL21IXEYkoUFOlzTd5pzs3dkkST0ZndPFGgDWcBMzCSUPauK+JKooFDD
6PfUcpnABoVVitQRQG+vmusgXqT3LAK4FW/gHflFaMitgkO/f6tvkIsB/kXquU1a
pMQa4voDqEwvnkTOZdZ9fAAUufSO6IovC1xrePir5Db6YnLvOUOwiRWXVF0kVvjo
xC6PN2Yn+dC/peE/KxAKn6gp2/D2Q49VlWCj/e5XVQQx2Pv63vJMgBE/cvrOVnQu
YFokHImiqv2Bg7D3nuRADcMy/dL21EmhVcDUzhrjEJuWlNJ+QgAuhAAruMTZnBgK
xHYMeW6K4YoAfRH2QRNfN4/6hcqTtJSSvuOyJPAAu06XWDqC6R3PA1Ct2CwKz4+6
dzgMy5TlcxLw+2JMkZtLHvaCnU5U6hNr2B/NlYTyFV0ULqaIfiBOzh5v6eD0zV0g
oI2Ip30uo2b535ds0iNqpzrV5ttODZnftGhsacA11w2EK/NgobiT+5smhd31xoJA
o2AqWMypR61NnMp9OFxpZMqOjAgqH3QL59MzVmCZxblMM1fV32epwBDcNu7I+pKE
VD99TxRIDPdoeuP/hPdn4QPUvgIbLOA297WBOULEKTbzu155H7hHIfln8A85PKql
dVn1vQaRoSJrcMq5nL7DHGLZbZ3AGvYBvBaqjCp132DF2NI7xqczwF/GnodZ2stP
TEbx1/dsAkZjGXy1LrKLBfDdzKDv8HXNp+jFZ83wUQTfFzxNXRRV56r9kVmL1ECu
GfRDift7nKs5GpmwdiTdJNHAjcoJcfc7S9OLo+2nN0DgzKUsJ+bvA7UH2y4nEgkl
PKkjq2RUV2+UNEGbguBHQTlRaSfvzRwPotstn6xWkwkMNOTUHoHRVA44CqnAqN4d
fHxJHVYHrkTxPKLRs4cw0wtemFF6YyUtoCV6mkgsxqd15ouSvlD+7B0IPJxNvPiF
HxTDzQhMicZZYJo4FeMMCbOARCC9T/FhTOsTbSJxHJMLtig18KFEL5Bl49PRCrhP
4LdcX2TVaQm7FeqzBr8or2p/8GSPpjjZQkIsX/n8EYVMW2rGSgm9tLhCJwHSsApa
UTQhbMctrRJs0AOGigOMyYX3ql/Yy9ZLqXQCieDu7mnDzAWL8rj2K5VSZupD6nek
UdlPV1tHWt7sxZeFgfCZbuwmGkUXvBPWR4iS4y4/mEQh3naXe2zhCDdKrkeCzBia
yfsuxBVJDsAlpMk5Az0xVfvcFjl50fhHurxLFVckmOX7cHC8MVGyAsCRVO4jry4Z
SAiY2qNyrxIG5Pff34mRPwZX0dRuLtkzvY2SegWEpVnGvAsvHHxSg5T4+ysx6gPg
V8QrBy5ECaU1L/gZQazm1fnO8D6SKIN71HCQMjOIWYxkMg3c01um/dK2iIp48SrZ
4ZzRRVMa1kCvvBG+POYrc5ZhPY0moun3aMcjYVS6qrU7PcP/z5zRXSByV+651JGx
id0zFfCRghdAzSQkxOAj9MvzMc/5hcOkrvU+zxD1IXBDZliUPK9uPoPvzAqvrWsE
PjKbcCO2sZ8db5WgknmGdr1sHDQvybcdnnDDc307yOQaGFDQax8nFTtZsA/gvIbk
etQDOSmlI1RWAOiQhjEr7Vc3eUTa7sAnuGTUqYts12MLbLD8FY9k2ipM0lH5+KIw
d/559hlPXhpWGRL8f6vW3A7JDmf8+Ofp1VmQZtaAcNG01YInFj3qzMnfUuiNpbN3
J9pF+GUtbXWp9OVY19d3v6JqoSyoJb0bmal98vWo/oHnfW9TfAd36BLGOgTHh5nH
nmRNW1eu/tk+oUdM7t4niTiHa6SJsWhLnMAt6Qh974t4rHSuREX/JD6UtcA1g3jD
NuRr8xCBIOmihdYSQcUgzeH/0Yy16e4IFmOIyjE20iWio3oGCj5UQ5MDqYbkoX1m
UZ5ns591H15kwakT1Sx728VTK8bcHbHgaZ+V/lb2mLBNgOJQOlqiQiVNYo+D4sFI
nlqn1esbDeSwihiVjgAF7D6yQQdTe8cE+8ExMXl60CTnLtq//LeecSlsDSiYyyIV
D+uEuQF95z49dz3o4rCv3UyhL0SN71RkKWtwqmIPIUwXd88V2C/f+gq9K66A+65r
y7bt42R0pgdsBECIaSBY8wqLy8o5B9f8QoKkIHte7iUCRltGpSHcG41qJI0mKi/O
x00Hij6T6TYdlBP+LNdsxgguScsBpl7rDsn3Z9+fmn4WWS/IaOMLO2tsruGmiOTW
Xu+ySxnVkIaFWtW/VSFlg8zpevVodZOImGvechX98qzG1Xylwol3hH+fV5tl2Ucv
KkCcxCt0zAPp7KIol4XlHNKCPSIHll5IOk8M6ow3ZOdQqwJ67yELeFksGFFmp892
089ouqD98XDS1MrVh7XaQIZ9cljLaQw6rfsUBpLR/3Mr53amVYg8WlVV+XFL2z8h
wfoz8T3tPYVDY8EICm9OErl709wUpety3sq9jfmfYGAZ12D6GFoc6ey8noqXOtr0
CTZEXaT2vuOrP+uroffL9usqiRSChl7PWBaS6b3O8HYvGFYtlOaGtpHSsDi9ySnz
dkeLdTxviIHiCt8THctFhehN3gZpYWN/o5MiBBw0icWWPNDW7Ub5z0xdMzXQIWCx
qZXOtYPEJaIw4Xu8v2JHc42bNm/iO8K4Dtv9xZb+6ZSURNfIiJWDnL8d2SnH9HCC
/lXiV6LCZ3qekuzankAkjBgNh4xczVzwhgExiztdiiKiq9gNHG52pS6BejRx+0VS
baAPMOPZqozf/aIiY1M28s+9h6kG5VCqFs5hCg9ZxNgWoTqgQp6Ft3+3pea5ddMx
QkP0Eaiw5GyMs59Hgs/g9bHugX8aqMeHzNmNmV3v++qB769QQXojEYohZte8JgHS
iuWOmr8JxgVeDJI8LIpyS9T5Il4UZgk0/K79UwWu8ib/VAzgbXmeB2Yr3Xd3p/U2
BeaXXZrHv+WhJ3GIUkFTdpGHd7csTe4sBhpD++8hAw3+0nhrH7TZ99s4AOayOFZ7
tpHiMGJXN54DHnzEIWvJ+mvcm7Ob8PpH5y52KqBiJ+vdTJDYDB4flXHhcU5WpJ23
f2s0VUsbb4mFNFtaSax/jx38JsS4kVqA5yiQhz1Y4rXkk9aLRb1hi6ONwLg4u1bW
8ZxxykLhNh2LS9cllkn2Xq/eythxlsbeMT7AoVxSNnvZAla7iJBLft19rFH1j/2T
5c3mMvg7wAwJlto2tEw2Jh4NLnrFX4iDdUelwslA7oad/VDrs/yowqMxOAHYeEKA
1ifVVjY4Se4eFWLGnfh3LK4GT9hGSpzNrYu30ZJhOaukatAVUrkzefXppz2QRUEx
GqgFSfmn76LVQq1ufVC9L7xTDjQnmtXd0BN6t19geXz5EXK529K2zE0yrr1qS0FG
K/GCI47tQfD1iFfC3rayNB2ME9dhCgeF+ZS2u/lpgz84VeDiq4eogmBFlnsU81mS
6UrFovCNiAKI2Dz5b2h3PGBPhwm3O+PIeqnfJ5GKdh9Dq6UhALUoLqxYMqPxG9iN
AOiyWFpjgeTVLIg7p44yYbjOsX9KmDa4WNT+QwyAspXQ6yOYaknXm7nnI9qssd9u
t7dwxrDyYWq08FzO1ND9REeBcH5uStgzkQFVAe2A46iqgT1hl4rAyYDckyxJjrot
iQdxM1IXtbMevQ6LEs22Pxvst1Hi86rJ5EHWvWQOWl+YwTyPhOkSNF04uV/Lryn3
lLIxa5Ksslr9Cj1X+HB6xYkAKkrXT6gYvnLLbszK8iCcofqWdF1HAM9ObOouuZ+g
0GvyU0ECft4HKb3LjqObxdH7OY9fJpQgN2LBfQ8s9u4xDr8AFzBkDt67IUufDUOP
1JOXxzOp440Z6S8YiLMag9RiC+douHCWikUd4jYfZHuan6jXKUSOhxuKJjY1H+tW
qv2MeBKX9dHjJC35fpgxn8w7sHoXw7XgwWYxYAhOtZ2PqXSfcB0rBPSxCfxuW+w2
U3TQZc/WAlqrn/fXwJsyje3tVb+eRi1XAgOVqeAlqFYPKOn4wORAG+UTeYqR02Gx
25FIPdxelgnKzhmCSREo9PuDl3lvKDEcdEoFWg3I9iJPY/Djs97J80mF5riu52gl
tXjnDtZqIYEAvlbCQ5712+ip7H+4fDJpKk1+F7l3+LbKPJW7sCLnhxiTHNkL9hT1
KYRRZQU7eN4omjTyB2vosw/ARhzLBb6kFFNcYUUN2RPBAG8/wevb1HJsyEWAhlIh
kJmjxFN4LZLt6Hth5L21zcOu8PPjcOZ+SacC5fMOWZEQD1LQSPEXL5Ksk7Epyrjc
5yslGeXe528fMq0Z4zvJou+lwhzQH1UosyBBesNXml1le6XsLdGDvUCfzTuLs2NM
LKPGoLsR2tScYnAGOonS2sXLcqIO0IR7LTpcYSq2r1Gtve/4tTCngjQQSGcftsXu
w2Y44VjCwdb4Kjol4P8Pr+mYYW/tsJzLIS5xADmVTvDr7hf8tdPTwvpTFu4+qxFY
PdVI8ZnvQfXmyLMMSXV14GbV5JUme47k8mVla5zW6MhKmXaAzcVRHkiMAJYBX8nN
PFLsFJJhTufad1cZM5gN8jCcaZ8BEqY2Gagle6PwE+bJTMwFc4yAZXStJkdBB2/X
V5IeUhFdRAohyEORXtKLL7ehKHqDcj7GKGLpHN2iQtjZhf2gFv2X/WKYiRF2Hrlk
pLmOwKFUqgBad3j3PoHZ9b5gy2CvQKLRiz5mKob0Sswm4ZF6v26fn2P5b5iIbExR
VA46Ap/OwjoZYNiUhNe5qRK1ItbLHCqCRzcYfGIicYIlUTt/3wClKuTiaicZKLSC
l8hFSfUiTKS+pyTekxySY4sq0ROvwkWFfV1Z5UO7tTP7+aCZfepP65v8/vJkTLkK
MayOvPVOxkIpi31k1U3Mt+aNbaCdeVafBewyWXBAr8L0F0aT7IRTAKbpNk6n2uhB
Jh862SBWEJEAMdxeAJkBneCfOicx210TRtfQwqMAjvcHu7XnqfcYYcU70121K+Yb
+bI6DPaoGEN15IJ736pnfSTJp6f6P2JhHdLMpR9jXoSvv09VgF2eMZKvzbSnBGfw
HOpQlfWiPCI7md0tUpc/v9j4Mtj5sCgKuDCQwfK/oHmkvxTugj6mRC4PwLeLGFyj
NPldHTy7G35vLfbinDRlmNmAU995YTZvYz5dfwc/vmupikHXP0PCCLZNUWpcZZKL
aST/J2Gd+ppqmr7EnMUZhsztkBhU9mcjFNe3o7NNiPoUnPcEY/5gIRoUtEnd0Huy
ZYxOSDqkZy+Rh8fLqqwkeCd/ZDMnos2jDi+SCIlpHEHHc5FmmQOHlw6XzUpHRabq
mYOjzCcrd3Ks84UL3Dv6mZCMBEqlxh4yiFfGrhAICvGZkcvZFvSO5F4Y4+MLzitx
j/bYGa/NKm65kXKFZzGNK97yPSYon9iE1eQ15g95qHtLn2dlaggHOH01ZcnCjgjU
xoOJH79P771bEIGXNfDxK40C2HPboIsSP3/WCM7HZGQJqzPHzdWZC61stcm6gLUB
H8FWRzzAU32rEeFvaYyf+rbBY6juI9AqkFBQGwecskb/n0HRHkd30X24ybDjM1SL
pp0BJduPHNoD3C4cFZs9+GB9AoJhCoHwevgty0XZpErUwhSa9BkXFgohXyVo53Dl
cgXFk1pWRMplT7Xrcd4NQJaUU3J1x00l8ROS7rDeyHB8+ccSaiv6/OllXRBfs1xC
QI28J2gSE/+ktlI+rubLReTvl2nTKVjutlX6ev2tXgf920/TwkGLt5yBXD/qFuxd
ZbDIUza9Re/3bzOHsC04By62Y6yPmnqNwLIgUtifWCLSIdbzG2uwut8lRI4+4gaO
Q/eyBr013N68TfiasU291VKxMedvBGNzcTyQ6RUdgcKLcgirOC4/4yUmMbLGXyO1
bBjn8Ulvq1AHZEOGYJkamAYxZYvskXdwKjPFASu1ptF/2RsnHh4jGSE5S83H4H7P
4EHhHh79dCK2lLWGHcV8ArUAFqXc4ZVpN/7SheB3I/U1/LezHTV8hxQPdWlJUrnx
UMcbaWUNUWDgooXLUecBMSYfP9M7ZLUj+ct/nJ03v3dTl7mDk11qyVVDXslh5WDP
UkLl/jt/ZGoXFDp51kfNP8NPa1gVLDw10BxOKAf9bas6WTvnPSmXAPgoDI8CeTdu
QtuFeVCL0AX9GzMLdITefq5tR4w9JmZpEh2UvGId9ZMptTTowLI9PKPVI+N5h5+k
ZpCkAwpC7kk1XG/rpI+smMebzqrHz+bmMHqBH2KEu8Cnl9azIQJmtDLOm6Y3ErMv
TLBRsiUDAzkLVeaCdsxChoaIvQxsOvmWJYhyj+qii8740NJVD4P+qodu8dp0p4jk
hwkFcpIyqNSzyJMGwAZGL//4JbWu+QXND0P4dqCfAPvUJAUdRZq1hJqYGwiJdh2a
+NGYgSc1f8zle53MzV8MSw542LDmMVU+NrEe5N4NjIv1yO0jw9zBua5rODlzbllB
1KH4YSnT2QcTcT8HDPOzxxu12ZjmA20+U+rPoUkcvV90C5M9DrZY947kNOdk7+JV
A8FN1+R0/Bz34nvWJ4PGgfwdCPN10xFb7NKezOel7+tCwzhvRgrwQZSVYJ2ATlY5
kYlRALZQkftErFNN0Lyqowzdvwm5IcIoBUx15xDd0uFxrZLgZQVnV1NHiuaxfs5v
yqheBNX1hhcRv0k0X21qD6UsuEeuDNLpNxGpBp6uZaEOSwVhwEQs4Br5BgT1ZTnK
QFo0QSkIxqfVCm0gL3ZAFLllwL4CrSSAfIXI0FX8Jvk7CVrvrMAs+TsnciN7e7CZ
tb5exvnaAuhNXThT08lwpbfPIUBvk2Sgj9XgZJ88NpZqhsVJ8UQgiiuFs33SFGJZ
32xKHIAzZD+1PMlHd2ZDwP6lZeX/2kdOpJYjoJcTwAZ0cf/R4+BWdW8Mp4pqOLNu
8oBGRywX6wvcashjlJ1xVmcfv03RLZ82V4eG7ZfzYA2HImX5YEtxbVwQ5ChjEHpt
G3vlv8DPzFRs9ulnGqESS0RVYEXLTAprMMZZPMX5UMTQ6w0ePOlVLzpGEFSqA+t5
wBcG3r8wuoKF+sr0mKV0JVHMk9OP9X94m3SqDg9HQ3sEESBQKl7IJAwlxHXkgD9N
GtOZ5FKlZMQHZ6jb4RRIaxJ+M3T8lMtaRVF4aEzbK/w66d2JtNJY3HbINhvSoyRW
72EXC7MYvo3zpL+TV9umLpzHtog39aC9XPI5BoM5gXwAM7gA6RFcvW+Z/rNiHV+i
vDGRSy+MS61x5+SzaKHSk2IYBB8Zo11PS6JPYFreRWT5BRTjYXaz3UJvMTDnAOb1
3V6V5TKb1QgiQZgyrVO0a7RCM1OmZ07UV2ceUzativvShq+BstMyayLj+3vcSqFo
KYaA/ExYhv8XBJfs2xb3DPe61knKBs1fKmUAYqlZ9XQwncAgLf8YsC8sA058LWW3
hRZqtSiIJJehErDuQIlQpXCWxdXjyXFeNInFQehAV8bG6lRL/W6p3hsfYBkA5Rwl
n9MPcei9wm2IuEvjGfJwVViZIByTjj8WBUlXUOQkdRGi9cg3rhge3FSVK55kxNYi
c7KlW3axLQwO6d4cO8a8rQy+bA3OEDBYh01yDrhNcYaLFx1NgFtGsNg3E+g6icWI
bf5JmFZJ5FBH5wFWKha1ZWp0h1/ynEl7NGxL0aY/mGWNHBDoeVR+1rGbkUd57TNi
DkDOv+ZtLSpYYKs5tfvB49esnGKm28myF/NMfzzXqfr9QOgbxb2JOtvKOCx43jdZ
9i6JpjWCffa4h4Vo+ktWs3MBMMgj+XFLQrir2S3eXbcLsghvYly3D/npdrYdSXsE
PUpImt81XAfnSRVM5BpTj/u1lOS7tvNwb5e6XuQ9/BxqoeVqYNtkyRIYJ3yno/yU
FO0uBvjmyLK+TkWOO2k7NJB/Ssy4SbYpLhHmvlrAoZXjcKSW30Dcl5Vd4EVtD1Vy
+EwMjbLT1RSYdVa3bsf5RPXRx1ZQY9izC7QAkYYien4zOUBZVeH7yB9T9q+9vkdv
WXVi8MGgvGnA07VjuTT6CCPD/tJ3QiI/ToXidiiVVv/Q1GKaU/Lv1kEVGj1QW42S
sWzeF4IqH0Z3MWtuRS2NSiv6Og5hPLfRO9rEZ5z1zGnOQm5W6LhPsCDrwgx0rfh5
sTu++46CtQqY6jk5fefTQwZDPiQ1q/C04yoXc9M4zLVXugZ0BpODn0s5Etq3HQ52
OgQJGuKUunct83dKHzjnJXM8u7MnwmrDVz952ztKmdalNYA7nG6PTycMcx9sVtcs
DGI/6Uxzsyco5/oAfIkdjt3Gh7K0YvQHkAJGiuWW8ADWcc1JgmSgdiIkYkzuA9Jj
3RVTqN5JOGYfn9L+kRC05bH4HKDiHDFTDtu24PEijDHwH3fdijyB95EjWbC46MbK
dfSwjEJL1jdnR411dO+y/Blrbx+FCRe8GTdFPfhOfvlaE21EenwJ8hV8NKUcu1v7
A+BzdTovCHAB0pdhnEY+7jpXjOhHm72nf+ellsmgaDBpi72NdOyvfTeot0aJVbG1
gew/EwWnPK8vnghXnWGXgHTZ6Ajj0FoEIDRdHMlujpdKc7UMtZuHJns3GhHMQq5w
2TBEP0A3uF+0adcVLD81AZxWU5OjP8ZHsdCiBErbAfep8nB+9jBKu4ot3quX0YYP
5bkdS3zdaDQLjI0Qc5dw0jFgfZpdTew4cRNP7f6UG8CYPY3TjNOqrJGLRyKvETuu
QLIuFi3k9/sXLaBYP3UHQoqkIxrThuJUKOe1rsMixnR12je7amPwpl57bbLFtH+q
9MJo5NXisHyXUGiIE1K+dkjpX/YgUDRnzTmpY9JV4yQ2Kuq06T64g0PNvztPzM1X
jmm3x2HHfw7jMxkaEmfj+XkDLfOfY1xrHlkiZO5vJcJlY5QnRxqweV13N31Vrv5O
NB8Hx2rwMGbmJeop49ishe+n/oUT2eQT+PJDCpuEwU1Mlg9UP6YnbuVrF/7x+WCh
G6SwGg7mtbWf60gHvhvbICuxSmk0ryX9bk3uqzkgOSMLuadpxyoNK7Kq77RR1TPl
CO56pnWZm4bl7E+BZe1KQ5d8hQkmEKeFsQOfUq+X6R5Gaa3ep/sEzfZdJjL68BV7
I7zGUmLMf1hQ0Ml0NIE9T9q4hf6rvFO0XXtpZImf1L/IlgW5ECIKxPOw5wm5429s
0r4trPQD9cKZNFLcwQyz+GiAhQQ4hIPfF6ILrLv/wqqO3KDV2qNYxHeXTr9aVc4e
TZy7n2lEYg3k3MwS5giYoKbCt+1Tf8ipYQWMLvB58O0N8/oivlvaWOzzq7iGDZGR
xn4x7f1xdqlL+VqzHwmjUTLL/LB7yc1frHailHMBODwH2xitq41xHcM7C9Q1FuHP
o6hKljID9H79RcBMx5mmk4rawsinXwzRxpLDBASnKMYMeslafO+OilGVNFFSr2ry
IBN2mKQhXxcMb7NPZLJhLaSqV/UBdrlwe5PwEtARM3lycSSKoPr7d9Cg2Gd2R9jf
dk2YVkXd50kDdi8+Ksx3VBkcz82PkdFhfuoI0czXEGwnKuYBXJg1DmeNHdtV5DVA
diHHA1i4yNYiWoCg9bd+QTCQ4WZsH4s5GOS7XSsTKjrNOh2O2onVspchIAG692sh
8uM0iwDqVLVG7/cMWhR/wtIexydrRdKS/BoJDmQHVsAv/fsQl/rV7EaxK0mnDwfd
iR0pu2GiISNej3YKB+Ap1GQ0WYEWGtrFDpq1dZlCNHh0+cO3EFLvMJCIbud/e+Hm
9EXPNBOv3dFxhZi17CaAPQY6sDwcfHz7QYbKfgaL9c/xd0OYt2SchyEYrNeCt/Kd
Ig0iDO0OxOLVBpYLgwhYK6Yvzylv4h94OHXLOWO3uxUTaUodm+UC58pD/1b6I/zD
QjfPdi3O7Gw00V8aadtYLctci4wnImA0JB6G1723dAmao4v7TqD2hRLaJNzC13lC
kOtmr+I2SXsi2B5aG4jsZIrrOOhkGNUaK9kZAZDivU7O45SuQivCwADFtiIFVJTO
UAA2VAIkDfZk8WbtM/rZRnKyzCsFP4XLOBg4BJRFPGFuf62oq7x66Imf8UEuPUvu
D4YUGnm8Zbk2ZZtyIIXfJIivDuliZirX+WMtHVxqHpoCVCIpNPsyObMSxY/1VU0z
RQRn7fShI0GyCzepXHx8oqMD3K7ssQlnTiOlxzIJJnvNldx0dEFK80thUznbG3EN
rid8B1SdpxHaq0I4qilipcAdxXzrtT8F5Pmiy1NJ2cBhbJYQ0mwXdIoMPkBfOYDO
iNXsDPDR0rsFPjNV4Qb218x54BvwF6cHh2nQBu/SgCWC6kdinNYeFAO9lXbueG8C
bhkUWkbX/kFNYy4pwfI23cw5UdEa1/OfCakSrxhA447u7ffG0XT6j3eusZiOXYnT
EEeQdM3V5Y9Ygabv7+GY/c5BEZg6JT1oRWMCHbRjBjSf4XC7goa5LFf6+clxm2YD
xjIm3F+4WbAlfaEMFUv/285kQuPTH1RE7Reg2D657AIKMvNKJWIZg0TAKI6X1AcP
ojujg9xENUpro8WpMENuAnGuxPfMKus+3dPAjVFKr8z6ZFyM1COg2HLhLn+T23hs
HZjha51Re20AybNIDOr2V3lLV+N1YPoWPSYjpurLOLtt7owWXZ15dpnBJWT64U5F
HZXKQFy7XFljIH0K43CqsmTngdQWJJrBxTk/KKUJDEN8Zv9KED9zTe0v8L5ZZniH
dO7cWGkPnxhDU2StgHr0oTxd6/tpXjBs7nI5r56xQ9zr0aUlVA0ivpDZwQkcI8Go
C7b75ClBQ+DBLB9uYjyTo2C7dgvu6Fgin82Jc98vd8DvoRn/HLkSZZK8rVmo62sj
oV2aMaJCrIGPP1hJnDhN4Q+0Lt9wpfI3PAPCcUs2r/uC5OpX+b4J6E7l7V5pCLjl
nSVX1hIVInPNYrRduJP8o3bcCjrPTUVyxP4cs+0vPX/CzxqBI52TPvVKy30szbAd
c9mwA/t2X7MkF5VAl5Esi6MBtOT6sE4eeO/r94lVBQ7uX23EquPHiLJZ+jAVbgf1
lekul2jq/tWk9TBDvmBtaf0GBUBgjvachtPA3FkHz63z8s4nUCaqYLG5vODZ7RQc
y9sBZ8+QQFMDnXiSN8bmApkqCrs2JSIR7+877pMPmbzPpgI2wQ05GwAzjbc8Uy4m
SXXSMCRsQ8xeUon8fsAl63JvJxBMoYCuyFAvHYuGEnrHIh45ZEICk3FMkjbTqCTL
PcmuTMguGCQj9oZ1j5AoxhIdf2JfiN58xuVzN1L7IcXqu9RnxbQ4dyaUBAtFpNJI
SQYdlvhNWzIM/mknweL+F5OGs+bV1IZvwKVVvZifTxmDf7ImU+M6cDmqiBROA7a6
Sw2luVOcMIeuoMwfoumBI+0cRtE7zVI1pSa0wpmJ7knPasW/yEco+mXnPSSElppP
DjoY4Lfivg4ham0sFHtO6qVVm+IZzOdXspozMFGsJ1pPlajdcicxI9uPCuZi7SWr
L8Xk2zXWQP9G9RNvgQHawMUJTG3M1cRKtjvrzMXzmO5Yp/fXO44dhnxSozdRV695
oyJyvFMvRVBBltA2ChcaVY/DboQm+f1DrZSJH++rWIMqOYL1+ZjH4iE/OklDedTv
iWMDeuCm3uVuohV0Oen7fkFgSUVCl2tp3V9cBc7MGdRP1Hxfq3758mhYJ2b5tcmD
PnKOsswpGDKjOTa+8ZSh853qbAEX9b4T4wrL67IGjSfqWFxX3rj+havuZtMmvioC
59b3d6uAF7taBP6yEHyC+yE1dH94AEBuUFg048cKgZWaOVL91TpPvDdldLkHipLL
dfO7Xo+6FCBSZb3dsolnnYK4Wl/N8FaBBsg7RaF056CJ5ps1XU+4HVO0ZPNTcWry
lgtQfYyDGamZhrvk7eSulCzYClR7TNxZVT5Umt/pW6wuXBVv4a5QOPsy1cIlwvTc
JtqoJ8SoQaOJvDqDIbpUFrORoe4W+c4P2sLzfpX0zGs2pRCD+5UmcD3WpIxzvLQh
Y5CBWUdr6kEQMQHm4ezGszp/6kQxeQps/ZQVefj4sTJ2B54TgjRxSVJhSy750ct8
7cqYJNVc5Bw+LcmnDR2y5VX5EarSHUnedXI36Vo/f/MXNc5VitQB9ynSiqTDlPal
vP2YWYgxGN5ImB2YbjaZDI5L9XF67TMMDAu/8Pt2XTOdyr0ESQnpcuLLeyLcC4zF
MuGBabiIgz821wEcV4o+lLf9q/wMj2APBArmbE4KnEXVEk4VdHfx6+r+6Bo8Bxd5
WYHYgNQzISkUqdd314RlaIS+jWkOMxsCDU8gYcK0mUYo38FWHvSRDa21zyh2WgDb
n4XSgEeWvmuDRCtK9cifM3QdFitJ4oOQZ1pIp2dkyB+lsrd5mIsM80TqrW0YNPCA
KDMbs7CI5zzRjGu9pYrug1MYxa4DhhvaaUWsPhARuLa0b5ug0Lfesn9JHBZh3KDs
lKmzYxkolD3uJgQtZtk96lzPI1L4nEIKIiW4Y+4kYWHtLX2GEHRUipvFbSvulLGs
wV5qN2PC5D+XWtEsn0Jri7RKl1bJvbiGD+2q4xKmAVnd7VzAYzU6oRRDMwJyqWbf
KI52jhWYZoirCIE78nqPuE357+FLdVDfzIgDEQyXWrtNC2PQAFhoKfzVT/Q+TNIP
f/3xlMiUWXsqs4d7APyUZRkd0qtM+bPHAu5pG6IykMtpNJVMMe4d/T3IJJsd1xGm
CU0+E6FsXbzeXoOFidzX99FlPBVhNc5YyKaplQ+DB9pred2WTGDWDjOr3XgMbv64
eVxlqC+YnPaDKJSkD1rRllw97bde0yg8LTiKYLVSLlqoRxdK46ORoEGpLlXEGlDS
EH5c1zpqLA1pYAkhFwybP1bhNs4ws7LQCCrUkoFpkMKLGNvvasL+iSBbHf0fABJK
S+LIXugCOIb9pBecD8Bd0lcHBs7GAcJgdQFFW9MOKHr5IqAVfuXAUO0YmqsRzlpi
uCc7Euh2d2pysExZEV9Blq1pP1v50jEaHrA9Ixf+xn8uGKi0ltIHDZBB9QHeqBK8
9P5NSwiy4OYT66/TVqKTEp59KeAy4q1bVGMKimUfCODzzcEL7F5juJShc7lRJ9K/
qjTUM7C9/uJCaCz5Cg4U+T3jWdam2sxpZwYES0DZFy6L651cWVM17Ja3OAZYiFvr
txpM5PSZdaumzWVWExVTvv5XcnJYiHKglB+opuoJHUF8cYTEYMyv3+osBcayaOwC
N7uGMJDwXdZYOZk1BezuF0SCsG/EYXI9ku6JPw6p3I3faetU3m2sSKfICejsy42R
BW+AQhQk9T809k222KI+bDqUClm01yVr8GqokPl88yRBO/YgKWw8PHOU2nwEh8WI
ZHxLv2zx2SS3Yb30lLHquchIM190XcaF/RFI6bkxd6xnOKmNgxiv6M1fdf4QJMXn
iEV9BClqsG7uTUbHg4l0L+3CSK5c3YxSWANBFZSL1rPtXFJJ8YXnisgMznxGY9eR
A7VGw9rxlOyGdut1NabBVClaGmAQ9uK+5KF/JLQAUCnO3zB9D0i7LmTcYCGIugiP
GJo8EXcLAWQbYTFQObwJRp3ZgZnv7NMxt2kM8YhwHiwVK88nT/huEQ/hI5wwt7ei
P2bqeA+C9DVP57Lac2Lc7C3kgbYxoAjzJrB59x3F3vvyxegjAUfVOPYABYMYMn3c
ePS00XTJimEVxfsRK4cbqLchd34h2fEJCi00TuA40sZrJt4Wp6BxLJoxMqAreQnl
BzPWvBmAIsvGvVDzPR5wRMGivJy+mDyZMymEsK5zuk5XHgQXMLePoCn0pyICCTya
Ni3LI8KtHRBzv9Jz9qB4Wu6NjF4YbEMb410PCRwd6m5gLQKjiFr9683TbFzLik+9
tBevNlsKCOw10mirde/UUWPJTygkx8bhDDoWVKH03bgWmSUBVx0QHnz9Sgbtxkew
yWGIRjfUuYRdTI5BhNlfKckQmvJ1vniNfxxBOZ211xb4RzA4bducAX4gXpVu4wC9
uSQUFZiQfulajU3Eo7jRS0Gk/sRChKJE+3titVt6BUxVmeFxSi/WzXfTPWYfJOGn
d22wzdfJ4FGHYkUsQpSX4DXldlv+wZ/aRKbf0GOC17XGpuPhRBj2l3zV2SszH0rQ
xqltdV/XqnjfzDLKT7PdWbvFxe7oFZ/xP49SCTbeko+TL2bhspVu5PQOCDyWbMUe
mJTas1wykzOrApFK3Vh7BmHXy02v8MjsALpZuF7AHRdDd8QsLvbd6xlIRpn+TYCG
dlYB0gO+j3Z3zg6f6uAvlhWmhPAYWPIgRGIsLHnWfcyINRVvtH2WYbO2qnRlOp4/
WQTjzmFn+0Jtnul//YzCzwj3fre1Ykw2I1MB743qtq8GiknDvyQkK2Bc72WbuCLq
mGsMpIcuGbWEnFRPkIL4O0aRy1U6kovCDsuk/hccc20NJuxd/RCpeJqOs1x+v+kB
KK1rGOZ5o55lRSPR1t95D0VwXeCtuDMeS9ewI/G3KKLIvPRIuWJzg+WSuHZ1Up6G
eEdwOX10oIrCGIsqnCvSH9+Fu0nDP3MrG5j8ZF3lOZ3NfLsJXS3HLYoTAbnwNx8h
o8KAjZkM6L9lsRtCPTKAWwfyCw1wi8aLRl+L+VHWJVPf68Zyq1SN9dvzxbV2Mqgf
OYNeQ1l8wI4Ks1RDvVYc6GMDo8nwPKcmUPC6e+FzxR31sTN3PYIx44InlDUpnZKy
crIemRXZ91QO0yunO7/3damjcuG1ieDUmFZUUOkni/akFxZwWcSfKhzY60mDnVcv
bvimxPBYj6Bfx/1forhAYS8EYS9brkrUWE9apBPw2Wqwr2Ie61YlNx6qNT4pngOQ
2Ok4AGtty6MGAuPdv7FusbmObeAAnzDH95PLd3vUdjx2hQSQOCv9ZRmeAMHDHnVA
dDnWjsI74XXUKtC0Yh1+RDjSKfqhHe2aRRyY4O6TLWrUomIIlMts5QnoWpYzJir7
cbU7GdV/qixG3w/4cWhxgi+QrtvL46pL+dMqP5xn99xbDMnKpICtT9wxpdIHBBHO
nSsIfwPV98M7WMPoPUCA+MmJlb4AINzVAMHg5DvDphMTywRAqQKtt9dm5i4XCHpk
9+9+7oKvu7TIyGfMvnqtN73feadlM7LacYBO090eUrKh5qSnvxMeDaILF3+cFDRG
A/dtufQT/FtftBynQtWlHO8F8EcxVQiEAVRqMMEFdsslyNxttHGzwFYGteYM3lH1
nKWP0/AoBuD3v7YNmrUEbpJkwdDq/Se1t/04E2lCgDZ89vbl7qi8vcBjSiD0nMMw
zB1FhI8M0NQHQwxKsH1DufjrIulaVrwsm+RgTms9F/OnOsKoSnvNDb8hDq45UL/Q
61MameFsB7tGDC3TBrINR8+g6cgtPoxw7BGGXgZfJw8Mnl1FTy4S0f71eqKKcSXX
d4++5E1twIduFv7cPlElheqXmJGs9vfr2Ef93Ahwg7ZaPo05WVeHqLrmvlkRjs2/
WMONhZzS4BBu2rzrsfcx//47l+J6gphFvFCcnkVSo0bCedMJPzemndprKTyD0kC0
kY5gCL/Ep3QETwBSd0vylkpP9q6E0bDsT7/db2bzKZrjhrxhtHsfBQt7Xn7dtEE0
W70PjhmW32OC/n3vYe/J9BVEN8lTX3qcAC4iWd0aub7ruALbXbAgd7gt57cHdquv
Ztx52PanLNVfg6mfGRBP3Vd36e6+WLzncwzW9KrE9j90CyXH0cuCuSxJt0szTHRL
EshgwCs4erMFrO0oG8TbNgBA+qA3p/AN22mg2fVB6mmgeDLmFcoTtNhXVDhaw/ZU
zSg1prn3tHUXt6VAbPrRG+V6bh93bZCikRc3IT39TBh7OBhrPos84Wr2F6Y0szjp
SpEzZXTkB3txzKkmbCG3niRAenhvXYDL4tBjW/IoLp8lSpof7fJk1XngeiQEKB/t
Yf52GA4OVayhpdgLNIgwAovax1DtCGQuFunzgDkQ3SbAOlHL0a3UArX96t1YQckj
NMkQdfAyGVY8Ax/14g8ZH+cZCqawfDBQIytu5XUqQjb3dD3CNohmC7xaIPZFufbW
c1EC1Hx6Zkx1m0qpRG3Nyd1uFxZ/qo48bO4IDZw1p3wmlJ1AjMKq605fDNkzwCQt
mjowLLu1yoNbnBQR0h47tnHjSrDabl59emAy752lOyIqqO8iAOhph81J3bO0j6N+
tadYk7ia3gHzXSzsvkkfujTUYQlMGGpbWUrkwQNrDm7x/5u8i//rifMcDOwl8Law
fYz8c8AvnnF6kQAWMMR9w812USEG3p6hXFE7b8BEbTTaclH0VjcpvuOCj/YZ0biN
SLFfqBzg4mu+hxIriTyJhZ1VC/3V5O8ArYyIkOubFGmGSyt07HtyoZ9mu32ee8Se
BKr7o9w3e1CqNbYhV9qmisLpT3iGaQi1xpyAOI1PNdEhfKKpEmSUhU9BIvIA1FLc
keAo38wgMzyBBta7u4ESEZLjDgdNmd42rKrr6hLaOGVIbuLMWB2W8Hb6SZAq+Xml
2kbt1udHBDqoD8gZ4tUGzjeX08JX8c7nepBfJpwG/yBpOof/40pVNAVhD6G5TlC1
UhIlsQEMFMLEcs6JXvM6oEwVs0FlWkvT+21Gpd2RBsrjTFp/Dt7DKuKBBtJXSWs0
GgECBff+zkdD/xdxc+u2I/Yl5kNVCi1LIzTZneD7lYnioVZ6IrNYjkIbgQ4o6US4
CzakfF7h9Y2FB6BaGvJ5ghOXMg88IsaOAvStUilRHS7wNnpnyZK+rhx13pm3wJHT
oGLI6GSuTZD3qzUNcldJUlAcbMRg/HcEhEYAHcM/HEss8jx0CbCBBYECF1MrpxKV
ukuEMk1Se8p24M+6/Qnw+XCS+q2juOEW5olKJRGxJ+WJFhSZtunyo8B8JyUZ9WjI
4V8/DHnGYeVyoY1ZbWk6p5FrEYE4R7d58sw1N+Rn6dCaU7z+DzFZ6NmeLk0qrE1C
l64FZ385xyfNol3HfGGE/JpMBLAD4WLfQjrLugaMrYxvxWNWN8wLM7gx9DvYi9+D
vTPcGcMsmMueXGZyTYqMmCuE1kxbepi9pK2YOq2zIPSd+ZxbiyPw5nH66yhOPNLy
AJ9w3jefWhMBAFCgslVIEhcxYhzBVuc5Ksqq3wD90IvJakJiG/988JFDi5n4DlUp
xKbebqXnSA2wloGf1Tt6aalZTiSaQ6cF5DEhlBfdMBHebLtcUSBGcWjb1O6sg4MS
SYRzbaUDXXaEyzXotfdbLitrC8NDzbQd5hJFiwVNIZRokGnbgQWRCTt/EzslcNvX
aN/kIDnK4/J8U881Fyz+ptmKzOL5aiEuvsfjnUckyJ9xaU3Qs1mfLTbUzJcIxDlK
G4QqXGZst5qbXppknHtzJF1yJoHcr8v8zowtsMLPitQpj/Z+MsKyuzV3McZLVnot
1vBhu8DkTp3iH7DJBtLCemf/p0bZjiwFEiVrJ7BA+/F2nWXIdIsgQjM4dNrZ37Lg
Nr0H91DPPrJuRy5xYzs/B+9pfYKI7E+iIKRhoucPUKm8WMd5T9XgHx4Bte0GGQ5z
kqq9xlxodC1ggFDHsshv+Sn+6J9X1l4pVUTYuNhjS3ptak1j9t+NvfWYSFmfpLfq
Nzwh/V2XUXxU4hYlBTdErwx/9gRCp0BRp1AqDLf6b6opfQHa7eLrdPejO7bwoTK0
IknY6dUpyfLPJy1k69XiWzOOhhiB1muFQ24fER+4vRGf1ZzqL+axQ313PQvKHJ6i
d6MFQnSCXygbVsyP/YyHHhyHq6Vp3CKXBq9joorO+PE0TG8k/yzPvucxzkIewX1b
CL2zoxRXAoOYtVVFjQRbq4QvSsalbJAvGKrrU09Cl9nYy2P37OxwIs4sX4Xz7BZ4
rIsIP6O+PmJZnaoEflmEyCt2THGD8Y2/zmsZoe7X9ZrrNecUm8ZpO6lHQXTu+zV6
DJkvxmaw65vCK/CX7fPERBGqrjq6KJjUzMClvkvUQYn7OVWzjxDkfkzmi81Lt+nC
9HB7NfsfZ06wRQe9EQlQAH1CHUc4Yx9L4X45RvmTEQYFiFrcNUX7KyNLjDBy3dmt
7NBMEWAJcrf1V0bCNOW/X9OGrq5SVM/U2GD+3QDECHIDAnXfb9oUQki7BPpV8BHr
HVyHTLNOy9EQdmcpXcA96EV4+LTRi7icoxzn1b02IomwBTGMUNuIJKjxl4WvwgN7
fbf/aBCqJ/zGaALxUSJYx0fWcz0xV/mzrqhaeIyIubL9EDz5mgCKkcnt9H2kp8v9
cR4Q7XwBm7W7/2KWXdFnjRT0M6oq6vLAYJbC1uCLgnnbGpS97Sj/SQu8vO/JvWil
k8IjCE3UjwC3cBuohKSlS78zvOAHejDy9ZEl7Y1IAR7RcgRs7gRwCq92LLgtmrQv
Aeq3cNsWV3CU1Pl/YO0Ho9B5pCIJ2nYLawY45xUlEKL800A27Lt3k0WWKOuwmdHV
ijbruBUAVsCY/X7ZxGnsP6WP2Jpn6ZYmtF+2jGNAvCol0B0c8dAA1XqdUu57c8VT
zX/gHXPARZu2KHZu85usPGI3IsXJbRKSZ8Jo3dFeT99aMOiPNnTvDxIUTh54/Hz/
/992Yqe6PpQvodyyPq4Wxp9yQ0ZBaU5N+YLnAN0OdT5fJtLcSE4lg4F/3tRQG4O0
AvP8M5IIQDOgJcdY+gC12pSiUJqqvSvq+POeJfkIaXQVTegtl30wnpI7Fvs8INIR
8Ro3Lz4VcYFxalQ3fr9COzdMzLqCvB3AfkrdvUEF9V1uNySh1+2EXUYWf2709G9q
7Tiy7/K/St+woZ3biSBNomkhB1Z5cyDcxoPgsgjrFee4eiIOo6pseFFR/szIcpsn
DdiIP/6XqcyMwwK71o5PRcdquiUXouyGX+10R+rEQJ3yhOeB9WQEsnp2iTeNpABJ
Zf9td64O3vaMDF/tiy4zZDj1F+qoE3ctLBvOyZtPZE6qYzS2q90iRwvnff8svYUh
1+uxzN0Jz1WsviYqLlckM+RJwpcTd7XUznBNSEjGygS8NZ82ycUV02r84NzZYg/a
FjKZe979Tno6YHTFrSB37qBSE+cl90xLt05GOSqS65C8Yz7chnipnePlAPSiKbux
LzJPl//iAU85O1cbhh6sbqA4fm3kN49p7lEUdlfQNChdahMIrbkKJtbY6pYH3esL
wwhr+P5hCLDbktxpN8zjiTghvomSJWcNYR8LmOaLpikYo8rsQZ9ehTWknttzcGse
Q5QNMKZGpypTAW7EpUlngky84rmSG1wGST5pZoHhbcnLv3TVK5rCnUJjCKNsjhfG
+kycZDzWw7mb1JqW3k2MCw358QBBwdckaRR7y3GLIbsW3VUAA8SJvVsAQ6wk2tcE
z5LEGLszWCgdoE2RZ60R7T040ZO2mEHUkxqdAVxv0LH6vcUd+FET0S0d8bQF2O0I
d49Ip/0YnlAo4B4DWjOHC/XcSs/JftgbzTMdkF1nshhjhT6xDIVJCXYcSnIFhffA
NYfdymzWXj4xDsGQYWqrt7ffXxjBhDTRXVFMNM3rYsjf/Zz530ugK45nD95+if3z
hwfnHH1ZkTRnaKJPU3JiNLhV3/m3+4cpZX+VOYYmHolPwfjt9edG9VIoBDi+k7jY
jrB1msQmI47bkpe3QaMQ7PqIWy1x1bDsiH7endFtLr3oBTXuFnAEhevirNzMUGD5
iPSpd8gcLqi9U0gzyEQp9qWCH4VGaVlfk89ySlX6KL3gAgOpxcCxC2RPxO0WF0il
QSkkCikoxIHJrdbruo9RB72FPAtkCBuhFCHwFf/AJlCTpfc94Ffl/xHkoxPbEzOp
iNNUiwQ0bCT5fJrfq7jxrBjgAFi6H3IrcvwXPM0wI9Rud6bhJZCb4LrQgKL4qaWd
c/oXxNVHZspeyI2MJoqiFUv2pJVzK5RvYvdiFu2JAFEBF7CmCcMs9ptzNNxRY96Q
P5KDoNYLqLalOK95wmHKFyc5RUfzkjPdg6OD7os/vYCG/1oxeFk08BlqHJEE/E0/
ZaBGiOuO8Nkz7AlmhiAdzqPjYkyEPwGr0HV2m6hXL/7KIwP9VipfVee2zJUIiD4F
7+CR/bVrUNV4j1o6kxf89bz2EDRVpnKt3XmMDlnQYW3U+RLHdkJbMFLKodciOy3t
IhJXqzHQ7SCkgnXz6NMRxOHY845yGK/xmMdfSapo/Skpuh857OxXl8hEk8LMEBBi
yPvxDUnRgJ8iioVYAA92FQ64ABFODpxwIIj4UWHJw1nzEOytYp9HlO/lLp+6C5dU
PjriBTGBO2KMP5P3bUtXq5Ddl0LH2l55lE14XVp47uZVPbotvBnNoAnokgAM0MBt
6dh9Ms9CYzhcycfukDwnBr0SC43YDF/vkG2LRVEvvUguj2w/DElezC5qJQ4iptrd
Mz4QldeZPWUWR/wSaP+19KxEU7IwkUMeBL2NEIeLEAkRJ3L3pJGKIUbAWGu3yXXP
GzRvn5OxMdDufd49pcmham/QDZzcSWfanvK2m2tTdjEfPkz7AEap5AZcaODmjqan
nEH5KzyWXZGNYa4CLzob4GerddE3HEOpVJ/WISLecNBbtgKP1bzrZK/8E1ymW2ws
MmsRUVv5SjmT58kgMsMX8WFk3cH7sSXYMQjBRcU33YXwT9FGnP51cUwRsO6GJjnJ
A6idZxYGTU1MVymy27YfZfGQxeOxNGdlXhb+hpclC9GCvrAF1mWZbyksoShJD4qk
lQLXoCc59EAbhOR9LigAKRD8kjqBNRyohucD7f3/+G9N14iGUIy/hrbBxqeZUrc7
0s05cjD6KcxjlOmn02DwGqhlcj/O2+KRshRNJVPLvbsV0J0j52lCCtFG0AGwnZ1X
T2UiGGAXQUtwsETmf9TOjQ207/DH467AZoPPlaomCbIj36xFOXRtVJsd2FYxaXCh
MiUzwZ79nNjFkxy9PS9q/4F8k9/uyugasEP8GO1L1hfoQrfuqYcO5xfWqIdyK2qN
Bz/+PxyadlrBGzkOTTnJuoJ0hfih+BycTEziJxDkc9glvgnnjw2/tPjISqc50MvX
RpnM27Q3N5mIPd8d+glGpTS+zmoiAozEXAK/XCVxDdPAGkSwcBPhsz0UDLRHfbXS
0pTUdqPbkNNthXMeNuI2cdGBu9NlCWyXsBX3EmgyvZYTl6ptPQUu/gy39VvXOIZ1
I+/LSv/b0+p6kUZUsm6iA2p/tq49+hPwlVMxCiAX9J/deTanDAYCy4d7MmYE/ACC
sBDaYclya/fyUNTiqrn0KibJ55B03Hg+R6GsCmlfQJLnhPRN20VeUKFULQRJO1mE
7NbCrU5hthME6W2JNpuqmZMSv7R2PTESpo9Uq/BrURL9RunMbkfckFlx8S/g+BMT
eSAaraDGzOVFnFgLEt2asBTuTACjD/bb1UHHztSJTlgeGPRCrTbZxWskmm0pU/Kc
GLyCoJFDEiXtDzYrgCpbK/b2wpjXGUOuaqlcD4NCVZiRDOwlVm6AXENFLunkPo1B
tvu2slyUNijtuKPZ+mWbSJHltn1Q7XOhADMGXg1otv1sZxMeWSpTBaSrNzgoiD+a
zqB4nx4YmacNtvaebFbdV8a6NdPqSFEhOyVFJqAvjjhtA14BwT+j4YYed9Cf/kdR
ZlNJhgRUh3wyzRUYqqrGQM1brKuwf+arVL0Iovn6HtAm8fCkjQsivDGdWPX2hYWc
VsDyrVj9C1Okre+jYpGXrTTbjE/5Cq9/cMds3CIU9oU+dQa5r7k0lac/5ZjqyQC0
2mYEwft/tF6pRAUptzFy5FwhuevKDGJO81V4TdTt6zBWijFO8upiobX2HIw5WjyQ
GumqNPQxPJTre648q35PidtJX3bqGcXxQMuFXbFhsvU1oEBbuf1ILRGRXKmKmBwC
DS9m/aySnb50BUA6UMCVM/WxZ1dEoQcGKvJjmkAVNCMn5JhrA+4cd+6I9W0Kkold
JcySQxOor0v/kmvgw8hfN8LGY0KxBdzsDQAfGlBW7TSdv0ppaMitFgFdrasmD7VT
+TXMTy1sweQnwewkVpmdIfGIld0S9/e5QiEPsqzIySFzAgo5Wr/lWv0pF+htVAlh
RQWaK6AKnYnqzxh1L5Nh9AydahrhFbaNqss/RA8VDd37pv0Z3ZGDSl8FRJuPa+pk
t57jav2id6p9rNJknYvC0Xhu4WZNXoYOUA35rRzB7+cYf+fi1VPeMjtCxtCyCk+n
SD4jps7UmOz+S0sO/6pDQ1cRpfhqiL4V5j/I6SJolaO2HXn+o21oXjX4oVOQjU53
fbMUkWEK+GLH0/0QkM7o0CKx3gmPF4uwsir3CfzyUXeWg6q7tMlcRlUiM8gWaANy
ZO9IpcXJQHie1K3z00ONSa1tteOF/MIiLjTCrTMaaX4siymgVT+e1gx9zBKsQSIU
BAxKMALPDr0dIcxcFFcKozpOzkfDpYgDsG1TpBHeZWWDShipseWJAwmFdygubrCB
yWV+QcEzyaaVBvprayONFKwSS2T0eh7sH4XkL6T2ciMJo7BtWcSMPz/7tNytZQo5
i22tv/yn0W1I8MlgUM7NWv08hhPNrGezABHpLRMRyoLy6vgPGfPfd+H2jXFKrJP2
75r9dU+GGz+yx6PAyhVZShlwIumMT4kFA+KHngpsSHQIy2fPY05JUg3GXGbLIvNb
YFQ7XlxiH5EAlmqfnSCyxTYE9RQf3kECONtuirxbmmeoWb7SNP0xQQyHhuBRw+8p
iDtz+aUqz7hVuMz3Uz6tvb/e9lSwBEUs1+Zqg40K9hhI9DINokSU7ZwKB4eu6Va0
lpcWbQ/PPthcqOU1s3Ddyff/JOwmjZ1e/uELoKNhr28aVDFnoIWpVr9Xk3cq5G61
1DsprJMGkxpm4FBFNdNZEJNqXfrlraGquBIhmTY0/o7BUZmO8TSirBwp7XmnZpiM
Q1yrldeuXhLWz8dvHyeFqEWYJScgC74pFyximw0dRcRy/2iiR4slF4pOt0NYOP62
8OiIRFb0qw+7tUFhIUXIrzusNJKz0x1YkwtliRJ4ncbk4AszKH297tMkF/XoRr1c
fwfEdd0EhzJBfb63sOLVnO1D1zvIfGF1/syaEiB1xvJGBGrQRSgfI6c8iU7qZa4f
FH8ARFZSNfeLwmbwKpHqtCFLhz7fV6x/ZP6pgaMaGpYo4fCHwTOge/VpdJ4FEAa2
cT7t20+UjeQjXOXQy4LmAo/PmoOnMt7g2XIgCpDbhfysYUVphE1zyRV85Zlgyubg
LFpBo2jXyx1URnO5Bm0LFhOPLO++dlRrYFHzEs6YQVW5OZTmEoyF3FYcwyefuoRr
u50D+T//6kR55iYDXrS/YrNwkO5BA6Z2hoD3kB9bXcArT5bW/mz/sLjrY6AZ+P61
vrJ7vma7s+Y7yErHRFM/fRg1XWYB2l6Ecqm+xyQIYCIcciF3RieQII3b2DOD4I7E
6Zt1DQIW/2S4goCtsvNWAipD9d8hA5tmFmUgE50rCHa/pdD0xuXoLaDbCvrPCGAZ
2u+iWsoOLm42xOmFIfLEvfwsMcmfgljU0o0+Bloc2+oquzoED9pmwsXtTVa1WlOg
afsRNmQReBr3SAzSxXXgBgsyGN0XDZdnGn/tKbKoWQjHnCVYrpDqPDDCERbuSmSG
d7YqszMXGQwDjgZ3e10NSgCik7lCnWsP/QGTGMWwoPkdbqcu8j4rZ0o5Hlb6Q1Fg
IZ0ik6b2xOiYsdgSR8vf8rumJqY6olkyC0RpRZZEGz5qlTbURTu4GSpc2QFyk59C
+5LOb5D9pW+kIgKsN1evFZRqevPV/5eM4SIaWOrpMeN0fQr0jYXtay2hcBdtjPIb
Ab65hZJ9f7Yw2m/LeguG9fcavv20KVE2WtkreOT6qLk9y78/PKacb7mFBCs13o1o
Zp6qVLjpJH8owUFiNdhnyYoJC/rG6yYcfSQKPfn4tjc1NfJTMh0kRfm5sMDJ1yw+
8B3dGHCUZUd+rES4YR8T5f1KzWBnMA0VmUqbwLy/2rBZLIEQRuXf5RqWkgNZe8Ir
0hEhi8a2LjZWMmUkwxySDjQhP2wvGt/YwKqGgFwPAl4ScUlRs75WNOkKC+4qtqWu
tIgrTE2F1N76S+w4VzsxG2Wolhrp16eWlbs8mjTfCCn1Yo+nN5B+6jzrwf1romIP
+e156NocZY/L/su+87zGYQrJQKcKL7c8mSzZT8PI7qbQ4yTYheomCqVzxdOojJVx
omG+UvyHZpnSDp7IqGy2pL0cpb4H6rRXPIS3aaMf/gFuXjsaX23pv5JhuAmxBcc3
i4+5gF2obvx8gno1gd5booqBr3TM9iOwlo+74bA/Y48IG1cEIhFq/y7pxNKe0Z11
GR/M0CIGo6XrxIVZVLgizqEst5rry+6Z0xPoAzhxbsM5TXACOKfKoTgx+Wh1/JeG
48RAoPqnlS2ova2k/9Bi65NjtacBKfMSNyASsYx9L5xx1+VwDprYZiBcEYAy3S5S
d//xKobSxjEj9GM5t4Sg75g/n/OEIHgQqSQDwisV3RWz31naFuPv618IbsfwS9zV
4vg9v/fmF98lWOA+5NF4FrSXujcqYEi/ElZ3Zj5vI91evj4BcmdnxOPVZRkzv3n7
5SiT4UEVxilM5xg/oy+prG07FGgEy1TEdxLOyBTCjGlkhLia6VWaO8x0ST3e22/v
VyH0WvsYfRfqBNBNIQ5BrYRC6oRVWfI2bSwxotGytfSc9pv5CIOCf7uLQkMSBqXl
uSvvgdYx0zzh05q8CzimmercMZskvEJI0YJc/0SHIO1kY1QXaAx3p2dA9quDrCcL
kUpdkyrBueOcEMx4XU9Bn4JEqMYjkVyVGsVyUSA2GGJ6HhK7f4iEcd+PLT4g1anl
YwQ3CbKR0A5ZWok7aRHlMyJq5mEY8dWSlyp1oiydVvsHrzV6tJ4cf5j24G8Li4Tt
56hwDF6OwlWhVc8o0STleu0T6trD72uCuk6G92Srn3MXLxf3H//i7p/B+5As3FCH
hMq0ES2WEHZ1Uvb6+/lyp0ADn3DqKZCHQZKP49DlFHDBxfAoolwE7momIU/nB7Bb
WlVZstId4ufqbPr6mCQy75iycdebvA/TF8SJeAIiPaSKSvUVBjOG6nn7yc1OrpYR
DywYRs78J01W09EGC5G4YA+jNQirqcMD5TLW0xiLiRgdovvYIgN/dSZTOkGQ1bwD
FqgfKe0Y6jyn97ZxlPQKiebUGt4hED+SiNTeQDFPmbN6GuUnomRqqvXDP4S0kgog
120aYHldVmST9rhJHPe1nT7URuxU8oigB/ETxCiIQTNU6Xhph34ZhyIWcNo31uZS
1xScLq4b7Q8urRQ58yNoEsasviVpFCNVBLunn6UjToLhqNBQcfvsfJ0d/f58KjNL
GC7CMqYEZpComXYeW3v/1w/AyN2drSVxo15SRpzPtPpILBlBpLArhnV7cVXD5Xkj
IqNExSVLL29JmtpiJN9Jjn+uD7nqh7mJhSPEghWcTt9aetZG8JLYz8aEq7dGujjK
2yfjMWHu1M6pwZPrkSbgMyUx5iE+CqjqXc0qUuk78DBRJd1xluuxLP6TOoNCUu6p
nPD1oJ/iY9Ccm0PGx/o8UOiMKh1LgJdaP10u35nZzkkIxHtcDlvzMiRnRRpnTjnJ
JuLVAd+WSmH9JDuULHXw7/uC+9zCJJA+wiQpJ/+ANF3BNqOE7pAQQ980L5YgzSNG
sTyGgSqXA3Cp69wXwfj57wogIzIcYCUTMY9SPoAYJzy5li+M2kzV6ir7R2qtGnps
uezjoxPB0cqV7w0ge6bBTLHIwqfEc8jSnmdRAiV0bk6UDFa1v3vM8g5Kk1NK5SRa
5YzpZbomZdGmGVLi6pXwrtVtSjPcn7qB2iBi81gl50g8Qmu8AAeNx6ony+T+/tct
jMoocc8QGrOeu95Qg5GbGtUh4Wq+493Zq9Lb4Pt0a0p+7ADGpLNY8YcgSc0FWpRx
DEA2XaOUWCqhtkwzt8fVYuXSsLozRF64P4TYJbMsMW/GlOETyXuCQoXrWBh4sZL1
EEwxeJieYjkLvKNwz6mnl0xByFC1Eo5tOUZH3DQZ8sRr49Kk0a4E0fySAx7c9zoR
9dhrDr3TWOZeiSuKDSmQl0vPrEOpnLRJ8uUfQDA5Xz6sE8e3Tl/Y5yNoRHaxHt56
1GDKYyolz0P+SzvTIKzz6xgaqY7h4yClErSi0YP+Cvb4JfY9yoh2ipyu5r+C7n3D
sdmZXHA4258GmLxJK4tBeUd/L2X67Ya1QD1ZVWXlDnse1zTr4LE2xHutryvp7TfY
UA5e52v9Gw/y0JRkhqLxmxGMX5KbJ2dSmnrlxkcdTodRU2yKjQNx5bnf9UgFYxJJ
BG1J1k6XsAgoGwKSemvOewtf9luBrGOhv6Lg1dWYywfM/jr2FXqZCt5CpYEq8+uU
MqE3kLBg5BUP7A46Eb3y9qRECgu5pbnCejwMEy6xUFfrgEyByEiRcaQola7CHNi6
IeJALFQT73/xAXdCtqUHz0KXqboPbttAhCXCgUOoWOUoDptOG5gwSrlLb3CBSrGH
sYjVlSDse7RbEcWiMJU7CaOyEWLbj8IuYKOH5K7jEDcV/Gz3CHfSNePR0kvqvvMI
znQU0JJRRSWNU0ZVs0XMuhKX+22OkhWPqwE9RUzYjQ/1zCLXjO/Pm8HIshtsHw3A
VW6A15viZAo5RI7toHNzbguwBgcD1PkIccTHF4glg5/2M1HaQvg2LZzxIYz81ddl
+ZTY0VMfo0Erb4IitZYXvsswiBfxGhquZX+kFg1lZMR37/bk+yXUiu2EMgI0SESc
34CKWNNhGEbnu41gEc4FuwUNttg/Yc2VmU+zxFm9jGr08Tn5uZzda1sDCYVq1Vyg
VxuZmHejnV7ARrz0FPtsA4n3Wtu+sgm6YMtDRISu2CYoReA9SgE9n6w2J6U5doBM
8rVYuDVS+0kzEcMxDEB0gnZuXIkjk6If/AD56OzYpu252HuPtnQQwIcNcLmOhDOT
vdgMV+8OENpwzs0Q02r7qAKg0n6srwa7L60MuBNn93ndDdCIxJiJY24MknRGTgIm
2xvJRq+LNc0y/LPyAEc0L+JOBHNv1strBfq16k+zSRCDnVpaoITUN53XQHAxSdSc
u5k7ZeYSr4AwDGE6L5es78vjDrG6xzGKPbxc5N5lj8LR4r7G8a5OScX11HiR+5ze
JDp0QPTYy0Z2t3JMUGXKbqNRjtc+gQ0LeE6sXnOujIkf9nh+hhkiwbaCGO121Phd
0AaBDZBgLl6w2nri1rooPiM6DuW3y1jozSfzzErBgkPKR+adC5vXBX7B6JiUJFQI
UDpEr4PLzCTPyayElZV1g0j2ISOkO1EpLEmYlwsjNkd+Ieqprukmgylhh54xreSq
J82kNbVoWUjjEs3Mwkfbhs8uDoi/lBOruExBpNQ1cKgQIgROhgXHpbeE8U1G0UkB
YNm4+cnTUBr54a5zOhlBR/12qF8WKFbtjDmynSoREkg7C4MPcVsrhHYnrK7AkJwq
HK/epPFLs2Lc7gA2ivL5FUeEISYrZHhGTEFgVGIvK/Gqfv+0nQBknKK04FmaX6rz
mgl20JaE0bIWMh4dh1lLIgnR4Og/mVAOqTyRoDURpdwmUNM77sya9ifzYqsvYYrF
+hnKV/ohgEudb462JXUNpb2wosztXYGSeoOcrZR75sOSB0SY/Tv7zH8JsT+LVoDq
N6kY9VY2472+NHQuGv6HGwkuWuyi6nuYjzglRXekNzpWC0ll7dluytydonjLctM0
OZDRsLybvvMKqJHXgBi4mi0LcvRGpY1F0mxw/AKgOgwd/4cQgQTWk8zrcvdTqq68
cY/VHi7HPWnGxIFxxPC6sBhXgXXHCo7+YOdPeQVLw+HkzodZedESA9pN0jYto4Y7
NBc5P8Vz442iCz9Nw/ZkFeHV5mc9y6GqNqo3ejVKbbeN+sBK5okE6SHZW1UNsWW/
+naP/0RNM65CDV+j2U0ntFsQzs9rtOWt6zXCBWyGVwoPy+EmLDNpq47wEvgxH4zt
5oifxbiS9P0ouBpA3p9jlDAbB5MHO4m2A/fW1YhzKWKsS3jeBYdsY/G8wyhqCB06
JfM7LKszIrMqEA2oUd2vDM+yPc5bJLP1OVLG8Jx6B3Nc5lV3jfZzcqMrNlgIg8FK
qMhvJN/Tkf/p4pAfjFqm8ajUd8+gN4yW9l5ggtL1U7d9a2Vsms+ejX+GBrFYKUmM
T1PpFhGTHy9EPnFlAhgaGcDqQPMde0WW2mF6IDFniYDNDxNp/B98+8/7D5lxUOkM
/KTBZegbODADghMlXQgR8dKMfK4G2luIYwr0sam2gHsK3yl5lob6UkY0Re7px3/R
SaFSXKEosF5sx+iAI2/qW9xD3znmpu9KjjkX/eD8yT+J0TExQMNkHLlHZSam4ov2
Ho3l07qM1B3KgvqUaafK0GzlxlogDUFJ91TdeVM/w2xzIBpNJKh8B1lRAu2VmJ46
X3aa1ulmQ+cfXz8tfnlDr6M6982QVoA+6cXYWWiEDprG86tQAWLF6+f0blhvff0t
EngWCDDOcl7TRZgzuHQHPAu5jDStJTwOPlWjCCRUvi569kNhz7j2yOVoX8llimIn
qnMtKzp8EhRrk/nYo7Jk19Z3ConMJ/fiqHATgdGfG+37Ilk4/5IvcECLFCnTQ1Cb
8QbCeymsEu2xbbUawXreLXkrj/qajoIiBbHrfRGK1GZC0rzm8Im6WMckIZ4jshiy
plbB6aaIhWpWH8DIdIUucnLEeX6kjglHDf1vxb+67tFW5VStbhI/+d+yDmfHl80A
+qr1rg4L70vvqcZCzAMh0ysvZQBKjdIs9eyOylKpUzh61dvc3TMhk/91UnD65EWh
o3LOoN8IyPHG0dzSYmzXsMmYnqFg+W/z2TSGegcokMNSkZCnijPy5u1I95GS+Iff
TxviAnqOlYlccPLR43652atP0yj2YspkH6QVT2sZA4wE16u3AgTcBg+pU3qOPZLk
gcZMO8+h59VbB69J44Gk/WmacPlPnbb4p4ootFEuCJzuORcbGmHrM0HWDLRogd+d
eafqEoAOBRqqMAiva7oDQ5/KSVLMISjThETQM2tjSDgSSyrMsY/BuxMNE7OyIjmW
xf7z6zkSX+tln6XL+pnweYZ2XSZb9YPw2z3RA8r8OEZFgotsRvamlYH4MN4jsuMf
HyniuHg1fR4FbUm447FrgqRSH8YPkPHcJ8M/FS2cKzBiZp/BysyaqwHaIufizskZ
IVwMZGtEh82rsA5u1xLrQOHK8TA9qxObSfhg8n2ZC/rchm4jatf7x2P4bsRnS0iX
ZXNTRp3e3CCGyCG3kpZ7Xdr5XFIjGmi7Vc+dfw8hTSaX+h7A+RV5cPx47Fs+Dcga
j274WyEJhAczMATzbZZNvsInIPUdU6T46An5HnNY7ma8AdzBLAZeW6Jppigu8XQE
Xf8rXyPZzVsqHgnD0YdcBfHvZLQfU76Rb1kVWgZfOzMtF0odTjuEv29kMy7ED4Rv
e9qPmG5c2mzpl+EATBy4/l8jeokpwB7opdPxiv+jizHFBYkuauqU2dxu8HTZgVKi
3CJB4/Y8wJqH5G/kNv5D/p3FQfzwRWvrsUpSX622Wq9IswO3E6bJ8u5Cs21iJm+X
VCiJDIzreW45O3Ij4zQP1+FETfTiAGXqG/kqbgNZ58UE0peOxmkkd+8AxhqXVhIg
u1iYNmGMs2DeHXZcZPN9wdqocjEN0SpPGH7VfAyguM0CckFUj4q8c5wfWK11VMNs
q+cqM2u7iU6xFIGzQTW1u7DCA/iqYGFWVxctQk9+ymgAibsP/fRLmVv9sELNfkvM
X2xO7cH4A9lxOsjqjzO6Aq6WBeL8V3V9kJQe6RBHHNaYPAVBa1Bvf68RXnfc1A87
uCQZA81qY3Ord9Ka5ds1LzBYMQ2gDrZaUyKnsFxsTaXbDsqShKoSEbODJZdJNEal
Zyg7TJ85Pka+bqdDQDiZGs4yP/qiXoCuktyRACHOoa+UIz/ZAJut2GTqLdbDMvOd
iwnq0Fh4a5f2iuOBTvH0gWivvPG1Csm9GGUL9d13zSbNCGD/cyaqDQzF1CjVSCDo
W+109JGBdSqTJzmz/bZ1vxHKgMdcK6aypvsqi4FTgjcmoXzvtHerYN+yJOpNBuZd
Ew//3Lnh6R5iEkQkgEBilq24of4B8iljFIznO6dShf0Jx+23wydSDD6vYO0G/GtI
cVF+a7IQdA5gu6q+vCB4y/Ko0squSPIO8UJ/5GKE0pmp1HiSauS7G78NTbqoFIkI
KHs/2aOCkvfaeo5eZ4Xt+oqd8TMRchGoKMqSioKZ5qABzll2PTyRDQjBTVRkqwfC
v1ZBF9FXeenznH5FUk6dQzafC6byT/ByYTZr7yd8qg8TNuwQixOv+rq674+7JoL+
zo9HTB/PNJSQQh2xR9DfshpOJIPVGguKMAaadQ/C9lz6LV71er54hP9vkBu0/kSq
/2KI+0AYp/EtiAjCLHT+PJ5ErquRFRFKfj6qq9WDyPtI6c0cjGwh5+AS8SGwJ012
H3TPQu+z6wVezk6uK903e1DMGf5UkmiokQluN268UABS88h7UBvbLBaQq+lHf+oW
pLKvNBLTwtCeIvOgngm5JjDCV/mwxY/24gLFRTlnimkvIsIBxTJfNqyApwgPE7qV
AkqvxNDZyUGZZPK7r1f9X25eLTGqMfkcdm2EGD68DGgmGn4DrHB1PyqulaEGUd+u
GwyC1Nm9/MJCSYISEnfhQmn+opL7u47uPWYIj/L4PpLfhcvu0gVrERfIMwh6VAbb
Vo70+kyADMh2QowDapem9+oXeR3PqfyL1rLrKKw5u/mBwM4AuZUcj6hXO8AMCHF2
3fH5k+rxXz1wTsHhfAB3WXIrIefNC2FNpwfD5nRIBOhiiLp/DAeOMovsPXoXx5wf
n9EwuBZTRqcIqiKTFCfeBWrIxA0Mpg6b7UsG6XWDeTtf1/7813OZaTk7HEW4zRTD
uwxUXiilLvtkbhmT5V1YFOhtjzA4wwAi3rlzf1z6psMKXi6k2gHTF6QaojyXEOuz
zvPRWioXu+k4EtK5hvssdGrld+wksr+C33djYriZPEsmi9zi1PRhMo+ScO2EhA/j
aCR0M7vokAc+bUShKx2XFht7kOG5HH08Roq/hs6AG1qozHYtBhdExzYm+Ly89hFj
M7ZCeBvNGcTUdXVBpE5pQXIxXdUHBll/WZM88mhBiVtxw/XxUj0cVTyhrW83g5xz
TwetauGm4EAna8N/CukIn8apeOvHu9z3BqT3aKN1NvtwLqSn1WQQzeBi40RtPYxX
m9YoAIsYCSnUntgzDUpjnaNQ0NZi5UfsyFyWbGiAicba3Gmx2HjMaN1u791CakbY
k9v6rGrkdH7eV0dMVu7gZGDd11z0ZTAHns8pdThVU7IJONJGCKRme9t59GYKzo4F
73v5/7FiBUab5YTNdnyW9l3aZh84EDO7UuuW26ZV2/+tKLOZuGB/9NdpKPV4XspM
zfVrp4JimVAYwkrjObXviJ3yXKznTjpff1xssuCWW4iTF237grR6TWiqilUleF+v
e+y9hVvrpKvJI9suvTTEJ1aRui7zE6r0j1TepZ12BE/ET82+nqBTfymAJty/hc5x
Wd4eu2E8U1a7jey8oAVygJGL2cSHF/Np2vO4fK3neQ/qFdORkjiQrTe70tHpi8jz
38CTK3gVYb3XbZga9XmHToJ2s4xtWKiPi6h0KXWz/wmL3WR5M3eDW/+gmAiElN2D
+WFSdeBXXfrwfHAlWIQBWwFLND25lD1Wzgb0sowiABw7U0p0ZL8wR+vzfxBo5C2b
QhxXygQZjlOFga6avRdRqmKViCDDyoj5q5csvDazXUfiS+SOcT9a7iwfZZOax2D1
C3G+DyHehfAUDcKhMZc9lGj/6lLYgW7L4X4oaAN+M9pG0x/3OruhCnau8YWY0Ziw
9TjOrzBAHGtqXsgC+dkdZmt8Vf2sf5NrCUbRmwE1g9W6tW5ENhgtQ9L+CuDhIPK0
uG0DyQhkKzG/q0XsXNU6QcUrXqrAtGwolNz8fQ4T0dDA/a2mFSrbi7e2OxZBhNh+
hLwp8FeJSx+MUcI+BHhPGM6W2xJPIjN0euAOoNtApDw=
`protect end_protected