`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
ddtXksX2+yylW5zu6QL2Lhnb2d1sD00763mmSITNX595NcHTEkwn0zB1Dry37fOW
FufOhVzEJp80NC5qZ/+F0Vk7Ik02dIR0elf3clrjeJRK85K4e3Hoo4xn7YbFUIms
l/8VZSb14+JVGURjfswrIyCUotIzlzVYZ6gzoZwDXIi5gQIBf/gI+KxNXPaKV+PQ
Ufys/12rjO6aI/pPlqSm0hCvftmBcnezN2hk1UeXgOIuKZnogjOsf0iJVX2aOOWE
6pD/psybjbnsNB6kH5uFTA5frkzIzkzl5d9+YDm9OyC+k84E83I/7/j+rk4L2dah
QJOvksSIzN867/4Qt8qYTQ==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="MvBXkzurAa5VTw+1JJ70nePUfoQXBvZOku/SMmg4TwQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
oRtzZL4VJ4iwysPsC8SXYCzXS8Fw2gtZTOskLcDV+1B9Nzn1zTyNtlo6lNICRmmK
ZRVu2BmCc2G+fmzynYlNTnSa7C0Cuel6FYpxCBlOuk3OF2tzAmLAuDyOH3Z1Yjzk
a0aHuoCdIRKv7BrZCdALt03JeUmXKPdOmIlkVGFl8yw=
`protect rights_digest_method = "sha256"
`protect end_toolblock="Jn9CQpRhJt4rnzZPRk+dOpzAubz7omckX1MrFd4p81o="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 3888 )
`protect data_block
gD6l00tciPUa6pDNTk/+txp9YJ6lFS7W7YO7BrMYAvj6x5dueVnllZWesGWXkK4/
dR7lrgJAmoiN6kmqMp1E6aEVmrJicH8bcGscpAs8Z1+fv0Hk4cMZH2GJ2LLS2yHY
95vJzfFkvuYT6HEA1+lf7h8VwS5FaFPgywxicaMihnRXx+jMEg1lgPjVq8GdbJ/P
a9qf8kusnqPTrJi4Ep4zfE5/R7UAeQbU8jf72yE0C6w0l7WrTaJkrEXrcWndzLUP
DVReRc5cMT8kL9Tix2gioBTDH2T31t/wth8up6VlmN8KE5rzFGn5pSolEa2O5SIt
So28L6jo+kBFky4W65Es5dGxkWtNEFcyD3ZDXlzMMmxMQ1vSRC4ajgJA9xzPyb0E
31bZDlkqtZPcij8LvvoRLrqmYRpCV3n/T3PNAMj6JnUTJxZeAVoMZDQmsopFalCH
qqjcrJLgDMlVF9NSyYIlhSaEOGI3A3gI/VRNMiRw7QUVtVBZ3uMIeDXe9I9FNe0D
P6YKoXNXWGVnZrnMpdMsAvPz5JT5vK6yvylGBLa/htvTlLP/RWEnLM0vcpYVR20X
uCPkvPyKSgzR0VavwVRQgUl/TZ0Ik9raE3o4WsgNSteK1szCJn0geCKllm/BKxAE
JEVBNOjpt6z+wzzJPzJCu/ilfni36/vXcqaD0ikDl465MdkTKLUAKb+WcRS30F6F
psJPiosEOXFhmmK6JCDDHP0TKB6rAE6muZKJ8jgiDs6DBwMeHa0OMxWxserKb+Fh
KUUSHdW6JaNnFbbSXfF+Bwj4VGjek/R11vssiPnVfzhs65kgG0+awTCVYUbif8Dy
wt2boYaInakrZsgjgzWkEZt00RyGuGOOsOjPstNc1ifM67fFasmRGnnpuWLXpOT+
JhcvKz1jvDZcQCA2vlwiOSMaxD5fdjJ/Ibm/Q5ZUQrTijmTIZHb+9o5fFpqtEYli
pYf6Z6u43Xcz3R60n02dY4uewV4Bi4Nd63nazXw3nvFYUdnoNgr5KZpMAaqYBPUl
rnl4is+9N8XY/7SwZPoFmebN9JmOehgVwkRkqv56iS+vGkTmSQJb0OydFTCQP0O5
YrPhgtuCGqi/C2NsoIr1vWAvw5V7EDjocZZVocgjarCsDHcSDnars3er/cI5xlyb
UgLjOoNeUuQjXxYgrlVKVCMnzXLaO6R1RbYKEtr3aGhwLEw6mOemXfJOkebp5G53
39biXygV1VSajndw8qBDngXYpe6Sv8dOl3RKUIx6U0NyKvOtt81mfeanW5rVotDv
kPR5hstXk2gIRIH4dUVh1MFhz5BnujbbFSvxPyNH+VKNZ8MV31BDh7b8gcCPMAKI
3jVrSMUHwBL8s1+lRmpkr3E0T0fyoblaGQqm8mrU5VFtpEtD4oKNUrHMGZvfvbdG
bYrZH400ds+CEYPdkMdIldMfNqWki434i1s++qNFMcJxNPVOvEBXtl2Z61BdBbMo
5KlJwDG4tlJR8L8jkI975UmD00ex7enEMOkaYCJ1GwWLwd96Dz/1gsRfqx9Gu4bv
v0St4jMMBS4Jfawxi3gDcCJlIPychZysYWawB9Rs7Bfvvi7XS5CDEmyFcdlJd0JI
RZSWeqbJj2Do8sDUnwv+amUj8ahY0rBcY/6Un+0rVqJWHWUH1fPcN1dPVjKkBDGX
nyyBTRhjaZAgSsZ+s6UIB/vFOx8m6mm4eAPo6qKu23DhW/QI5HjBrZ4gdvYyJBLw
meTDlrsGzRJHjGRAvK2VW3NLZvEUkqcJZaen+21G79xiIPXshq5ktrBCE2kT1LDI
WYYn/osNEWBFlrMG1I2lRh3xUfJ56fbvSaN4nuERpSoQNK1ChNDZj8cxNonTLrzF
0abrUSHFelrX3P0rQ6Oflg2pIFaMsvKqG77PnXm8LGqV1ufAAVcn9mzsKAOCoSMV
DpixmG5rnm3lxKpVQWyIWqpBRoEI7tIxW7IUT7ETTf4ZpVE51QA/d8eu8/YoWcv7
zJ1GgFeIvDNI5dPTGZWZWAKW53Q2UpGE6ErD0yK0vkLg1qHGFSJ5HW3gEH8NN9bp
X6X1wAludGJDVD6bs9xFLADDCkN8ZrmGA5V+HojTRvzMbC5lvprnBkLesRLcMore
2F7ADFtK2/7up2T5GDcQZO2eH+DSllX8N8lEAdluAyx8Prqtl5zSPxvwNweceFLx
ZuW1XEygX2kTlbWTHfUScUeW5we/Zp7ErIK94XhYtcixw3KBlFlykClV4gt+rd9T
rtaYpTCDl3FZ7Q9BHKwV7jzupxsRiLCvXY0TeIdEspCIToEA8/uYFZXSOXR0Cj0I
I22UMdRWDzLfmZZc4ybMar8y0Ks08ddpp+tqt5YwIuCo8x5LOsBdATxq2W83YG15
QLFHMhAnvualQn4wgCV4PVPabI0fV6U6idVvysTaCwMjAEB1DwaU5IP9GPPYEg4z
hNIWCY9//gR0IetCCErCSDcq5EPav+BO9qhD8DdQ5YngMvJg/FTvOUjw3/Bueow/
Aij1/1g9IgMCoqzp/41VJVTksu+WNAV7iMrdHS9aNAS9Dl6h5Tu6sJty1RXTmrgk
uXdqL33u5bDID50M7xzcntTsE+7GQpuKFgdUtPx/26daM0NtSAzbmg2EttEG5qYq
cmVUAMxCaecLTkrouPC8vDv3nw9zl5RMdLu4BtzEVRdc0OD1USXBkqbETsQbS1kj
oUQTqYWPYUzSZUNBZaCbrrONVXisDW3ggoHM5ANsdkzZkTqT538nR99CsmN+rxXH
w5atMH4NEuybIFa6IUlpCOY7fOB2xoaVmAtGYqLNBrVbaVQqob23mqmvjQVJPm+3
0CRrME9staXLeHIDoTtmML9yCB5dm9prUzVSj1/1WthgOqjAvjdn31qJVwbFQew/
TA+cHPCDiClqxGN1VUMyM333JpGV019drNBp+EQkdLqQeFH5CQvw5rQegFNJd6ux
0XsGQz2n/cWM//bEmMnpAJTq5Zmf/6kZvGmN/oDhnGDbIkr+77GWsj3aYjaWt+J9
6A6MLWSe4V61uPikQ+jKCFFTBhMi++Js4Y9ePbfGUNmp13WR6soh6FFvFG0g5auI
jsljSHH/ZqaVLysPSr9Qzl7THvdCtgfYfli0wGwEUwDNleFRxSkB5SRUfCXFh44p
HcSDjN3CpGe5v0J76m0iSSw4VvGjSBWvYpZzEqmyjMpevXewqUozeZ0ecUS4xsiR
XhaHlnpiINJ/USEreJw5/XGc1mTmvPfE0ouXqUruD5Aj6DLaag/WB17YO95KOcp6
jnxo8TrEsP626c8epAY6ahvWB13m/yzcX9xDI4Ag56Yz33cKvQ0GV1ODlHL6M8EB
3Hx8e8DKbEKs365mPdyW0OW/eBhcmd0UXC5uZ14Gtz+I6VLFN8g8AQhiUzwhAIhg
eZjl0BfcO4+peV2W+xqKUOp07yshz2EEha/85FDHDl3QUlkorpTKjdU3eCb2JUzV
3MAfwjKTg0LP/n4AlAVFiIXlhEBw7OmOeiWBm/jP3NFdeJISikdsHP3UrUEJD4KF
KviuFyy+SAljGEHXYjJtLBR8DCEPTHZl5lAXiQfAS6FJiC2kpBQwcEgu0D60m8xN
6WP3Y7AAtJJCNo/7kKRHPLoCReRhuSXXmowCazknj6VICFGomDLMRbzXL6WNJqao
grzRbJfSTWGgTQx7YxsOmQnlRdb+S9cSwzcB1tyrfUHPAtVJMnEEn7eE+Pku0w4B
oA/O0C0X5o9aPfR2Mb32wcetTknnmkHZLjloTjFy3sl34CI7KGVWlyoY5gtLEHAH
RT7y5aXbW4fRSgSgWe0IwEo6uofaLmtE+8vfOCw2YnPK5Yw48sti7gvEqjOLIYPS
O5LW2bx+ir0jAclJr/SL6RsIAbXEriMeI6y9bj4iRXENEDTi2+5llLXKS9nqmiA2
SddZKWUDAFGPFuSJMQTWKRyZCGPA67vt6VmVOOQ2fkipMLFRaePg1uuicdrdKL0r
sW/qmHElIwmtgFJQZ1xNahKWhg9Gw214ROTvz4hBM9jgnsPl+fbgSZXRA1lzvGAj
IqcwO8bLpggjX8STSOJ5q14BfjVVIO4hW/wd0KvLrw/t4Xis2rEowG2Gxxs/MEkx
kwESuvEC/grMmY4D1kb0jFiGZ46XDnj7q+HbaEXpf8uU2jQ4OQ/kmpoil07xaVZc
xABorp4iFjCYby3vHD3lzA3W5rntN5CLhW3CuZ+G1DJtqr8Ph19F7KJmFUypvcQf
RiCxv5Ep2IZEKjrKvEJoLRv0Gc4kM9soqRlazmCsm2KctVebH78SuX5KGpZhFOQP
f+TB/KIvIAOU6CTrchu7bx5juMFSgjREUFR/GK1P28ZeOD5M3OAkLRpcIciWX/TB
cpoSTsqsrcRIOgW5xNp3CLGXzKQQSAN5P03T5faw72o9yHAixmSK8v86tZu/+7hc
+yloP6QeTYSMhtNnjuizAJXuapk/XouC35UInjJPRSqarmiZ1XkYn1e0TWlpxL2G
lOCPVV5XQD1P6kIZVqA5zHzs9RgmPTGZs0y6bpE0oY2VQtQiFn3LouHjhZbvNdZk
8GgDLtgezighlvaN+noqTddJWg+UKOQ3TpFf6VyjaWqhYls4LfTupayN1QONhnWW
FYHDvzmpOVsB9tZ/H8TJFNPAE5nqL3hdVkfyKLi7Y/90ZQD9eGSzPVthpQADTmwU
5enontA+VYvxvo9UcpfCxPskUembGuv0BauPtW3V/rf5+fjHIf8P+D8LN8VThe35
Ql4Zi8jALNZ7MkzhM6FnZ1GeV4Ny5gCuFX/5i0dIC19TyeJOYe9jsteDtN0ixeQn
W/yI6QBMVwtmS2/6Rdle5XQcrlffj9H9g0++YCXMsoVhddLeB7XkD07QOW0Z81Ic
0XyIeRmCjBY9kkDCarmOlYEjqdv0I+aJtCH8wkXl50rz87qy3ThXcnBLj1/lDfG5
gdLa6fwP9PbvRzW8eVOy4OIiQifP4G+xwp7fS/KCk9GFVCFQGMRoo3A/4Jd27AKm
6M5jXZwJSUqilGssGJXoDLC8Ai2thPHvF/Zp9tkRfyR43U+5gYg3fMnmUYbr62ax
475uuSEyU4I0rvyNDh8rttTowYHz/Ki2/yoADz7FVW9S1Aoc8u9ceFy5xrrAQPWQ
aBmMF/mXdvfeco3f2pGhK+nkwB56IAF3zcW++XRj03X7VpMMSHRZmAYcRqWZ36Q/
`protect end_protected