`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
ddtXksX2+yylW5zu6QL2Lhnb2d1sD00763mmSITNX595NcHTEkwn0zB1Dry37fOW
FufOhVzEJp80NC5qZ/+F0Vk7Ik02dIR0elf3clrjeJRK85K4e3Hoo4xn7YbFUIms
l/8VZSb14+JVGURjfswrIyCUotIzlzVYZ6gzoZwDXIi5gQIBf/gI+KxNXPaKV+PQ
Ufys/12rjO6aI/pPlqSm0hCvftmBcnezN2hk1UeXgOIuKZnogjOsf0iJVX2aOOWE
6pD/psybjbnsNB6kH5uFTA5frkzIzkzl5d9+YDm9OyC+k84E83I/7/j+rk4L2dah
QJOvksSIzN867/4Qt8qYTQ==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="MvBXkzurAa5VTw+1JJ70nePUfoQXBvZOku/SMmg4TwQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
oRtzZL4VJ4iwysPsC8SXYCzXS8Fw2gtZTOskLcDV+1B9Nzn1zTyNtlo6lNICRmmK
ZRVu2BmCc2G+fmzynYlNTnSa7C0Cuel6FYpxCBlOuk3OF2tzAmLAuDyOH3Z1Yjzk
a0aHuoCdIRKv7BrZCdALt03JeUmXKPdOmIlkVGFl8yw=
`protect rights_digest_method = "sha256"
`protect end_toolblock="Jn9CQpRhJt4rnzZPRk+dOpzAubz7omckX1MrFd4p81o="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 49408 )
`protect data_block
gD6l00tciPUa6pDNTk/+t0OO0nC/UTtBwLB41d4inuAUA3i/ALrNyoJVcBnAmEQW
ptbcNp5fxEUJjnOxnedyZEuEBxWRieZFQnkRdF269oMokHpEI1sEQyXzq8+V+pKA
qA9E+zOQ4B35sl9a+/Wm7Se06xdCBFob1Jcxk9Gyf+lyC1rtxdSO5Nc06UFrpLaw
L2KHFz67iajYIT9RYxWc+674BSf4VKQCoPgUe/DhAOOaveaAGkGczhBbfvdG8x21
jSl1RRYRvQePY/OqmFrQcrgTiGdrd5taLLKg4wikxqeJ3gIJuHcIpC/oSmZvKHfj
i6eRhV1SFYimVIBvEIMalXp9/4LrR1vr06IZdml8T4ZJcDWoW0x23nE/PXtDSojc
Xjf8kJtC7ThPx/yqhePEjPHBIw+bE2Ks8bHkHMp2UMmeMu4lNsTZORUk9vvdbDrN
n65NN4WRZttjxrSXxDapLkBxwIftGcT8xPMw1A1NpxtV0s1KdGfLNF3kI9fCZMdA
RLta17hT0Czf+DUqBYfqaTq6qGxbLAMEEIP598eRdeUipP/F6Roe5m+dwBMyyrfl
ZE4PgpHR3U841KbALydniJefIv5l/ekH/9m4NMI4enQN1U6aCUMIVAhXuiyPatiq
HaaYvESyrgHjF4aaYkjLh+vQKRfHoibGOn4oZa84LfCZNDGf+8wXZybb5YQhrniH
KCqNxUWoLeHKeSkcvT4hcoXD1S8WnE0EXiHnJ2mRIj+I1vQvmoFjHBVxR9N/5kRm
Xp4YpvW2bdDJeXG7gIkET/GqVC0WKSUO5ORsdqeV9GxSMEHrqU1wBmQSGrmfeVcN
CXTBHewx/mIS7OIuFzJU8bKvTrupqRsZql8YU3yA8PqOZSsn4tcmiX4QFoC4fhd7
/cPZJ2TlDygIV01Yq0YbtyjMj/gHP2dHuX0/G+gHns3/Wj8g1sJYh71ROo/+IXXt
aufHG2gZkl7v3hcY+pPIyop9AbJNBlb/PnA9AAENYCnPn4CYqWjfnOglltR/9M6B
aWblKdeWGd4NJXMzBYVwOW6Qd12uF9EqSsIgi06UDCTuzpjqtai3IVcjMsNIPEAG
FaSS5XkGfLVp0SHNmWtS2gX7Ni6JNWR72auiOg+br8f98vME8SvbpU1m0XP1nlSY
Z9+RtCwlkiNsOdlrlm+iZYw+/A2sZ4VYB/O/FaQ5ieMZTNd+NxKbRhzfNb97XfyM
RWzm2IKeUw5LvuhD3hcyBKWTTJhciOpGKoL5wh+BbsJ7OLGRrf0ZmP782iUIuX4n
DLWbQlmfEinIH/CXO7mzYHi2pM778mapPJASIk+vHvtEXR9swqmgmxI7eJ5gm8bb
i0clBM4g5NXq26h4XepVf1HHBuNU+YdFT1xqQEOfs0rDKUzYKm+AzMvSS3mNHCa/
/GzZfPeTmPcmrCNsF7Dh3TMf6U4yHZzLbsQDkquuo9WSJ87qryGSvuXpjT1Of9xO
3e8jnF0sz4LtrWoustEA+yw3onZFtTwPlUfhBgjcysZWbv/SiujT7T7qyrT4RxJn
kJFibF1mMvue6kL1LrYJcvqlIimh4i7PluIdV8yB1SI19XLVk5m0uvDgzBKA2RLi
222QALZtg/NWpjBsUqX7wOeUsVo8lMiWX8/oFDNUTck8A3RjvWARN6Uz2jSQ3gQY
xvL2evD4MgWiwzsaAjE+Mzn7TvmCUNqacAacWTxGV7LeptehLtQg3El2PYvfAkO6
mwh97ZtqYjRWZIynsYVGImyf4/Ee/L5INBCbD3Zc9kPNTRatyoWo/upvl4rMOCQL
KDHXSgKb8GOxX6LPvQvvbcTPBmNHTXfFy3n+YfvnfKtz0TEDazPdqGqhSJRrolLY
0JrjuzmzA1UjArzsK5FhaR6UX+yDG2Nf5EBefCorE37rt1zwsQV4tXnSYd7vevVR
CkIwzsXH781r39RF1EY3xEPKk9Ae5JFOTQVqRcVCG8BPW9Q9eYMFr7bb2Zn5biuL
1lNnHJvSU9Yq15GvXQiq98FSXIYhlWYbddQn9XNQ7GYffDw8QG1Ec6cuVdThG32o
P6vUb/DbKgq2qzHw1okT/WRXDKBqQ6ZVW9CZk1LxI+JVno3EHzLjc+lj5yKCX+vK
r2K67SW9xm4eR7WDpigHMn4B+1KqBhSzddugPbUPTS6XXa+3A0E7KDY3oVBOhHCU
46WDnjj2sdhBlIzEpL4xL7XBaeKCb3I53dCrEffWFcXZreBb03x2N2JxMlwyzcxI
RZDbUKr/vvBO9J36j4O0FjWE/EFMNjG2VkAp5PpxafJhUwzVPtvdx3NqHh2Dr2e5
NYRUFBpdIo0Juznlaszcvs2LwnujA22uvgd5A9qrp1n2IdEGOzZthMsHTOdN6gpp
OcYBWzTbStRb48FBI18bMEPeUq7db2UnmNwS2S1ydwxycw9bop/p9soZfyWkFEg9
QSzfqDSvfoqczyJnw33K2BcmRYjpwt2raRrS8PeaNwRokRVWenhXxNXZfloFv4P9
7PtdpL30JkT3IB7FZw13iya4ugHzoypIWdsMw1CdTc1IsppSexuZFF9MVpQ1YWnx
lUYvtdQjYErL4IKV/p6G/cL3Tm1MhA2uB/BtOaBfHXhcApAYIUHK3BjoJO6J5pXN
lKGIxgvV5gp25X7p+Fj7AQL6jRyKky5hUNkxrXKHJEACDPe2S/4GS4KifiQqHU5S
qa3QSvYRmYhYqCztPe6xOrjD7n0++pldqhTEtbcRM6QY46rFrbuHq0M69VBVZ9LL
GUDwxN7GOV7OnGuRjixrSCjt/D+oy4S1Hp5WFRrsdeKTazISG/F05p6EHlsLNZzM
Z2zG8nosBq3DTkhBLH6X1AGJmyUMUsd6mxXF0J0I/NIGsYZ5ebsrebs5JKVpxow7
AuSEeBxiHHFgoHa9NF4C8oiabIjbkEalt/8aKreA3NNQfqM7afls7Gu67kwOcHFz
K7YGFDEC9MTc0iyjrYy3QcMbTSDMeu8XqU35MICJRPjhuB/P1mCJB9vWEZ7EGHYE
NFszUTPFVHvbXwSLbxZBqrA6wdyzltZ1or4+4pIkELUfUvWN+VY3LYMhad9bLJCo
R2kidL8UCmcmoARBuf/VIpWETptfLtbotjL+N1SJDWeQI8JTzNfjbtjBFsguagJX
9mvwPm1r2ZX8EwRNd0YG0OfspzTP/s8vlR4jyH6CJDTOBX5n1XTKI/PLXPRrMNnp
+NBXQBXBtYvBIXjN0UMMiJgmlqalVdJsTRZ2pkWmhBy3RRmrUnCrFxEDF60JHVpe
0462pWJsrPARkImumdzrtxT9D4vBR3rmcrh6e4IE8K5Qx79e94OfVGoaedSuQVI2
cKq3pTtj/sD2aE60Jdjip2u/M1sniryUgrtNRFhn7wT4qoBHiV1wzNeSvjXc44vR
QedeLGdpb/CNCqtqFgL/GnXjmmFs4T3xazGVTgFNVKzCTLuv/dauytjVQRRN8IpH
RsnxonqQlTjax5zqwkksZRuJF90+efTGzLEeA1Xe+1D4UTvgCLK89JpcgGL/9SZn
vG0hA2LIx5JA9wR92uxE5MPrOkXfbbwpiShMtu09q0rH6mDOSxJaLR0moM6m2nOX
UPdZRnTieoNE4x8K5iEGDy7/33RKfYKya5xrjXd7RRA0Ky6kdG6uy0xkNTBPzfgr
h8JJKM/QBKj2pPfZ1LKXEw7ZgRo1s/byEGNJiq7UQLMFP115mh8LQ96M3+mLeCMB
Vw0ulCO8zJR6/v0eztfn9VydpitrS0+IWXbEl9QmzUrPy/nmFPgqO9j/k/2emC4k
oQdJzviXsPqys7LkTdB9TGn1CIrUPRNZHVjsdhYoauWWBUHskTrzJwNCJAwF0m/2
+bOnESwSTYKLSFL3k40KDW6c8w3Cx2xLvH1BGIqEFSI0Eqw/aL0Bsx1/ZlBHT7Ey
1NGghKoKpqk8we0KQoztwCdF3ySIvKJUy7cvDrPfvmbsWFiTM45/+bVFYMmPVvqX
YtFn3zk0XxetRiw270KOainV6o5jnHGyW4zQav54acbO8silh/tLEs1FewiiR01E
RhKsLj1yw5LrGSlbIaL2QKAgDrybYswtKriMbEjXahzBqTWrpFqHfj/dr6jvNd2C
+vAxsYNiw2QTB9mPCguLJ5kNAOB2OPCqBx+kjpRp6p5gxOrBfNIzEnrBe/aSRHMu
Y04IbBs3HIFgPW9TUQe+sbjY6uFcdIp6QloUSkRezDMM3OpUBtydaz84wotqSVwE
Du+dPnGys64QPIkX0jwHn+HeyiX//G7wzck4AdJ7d3qc+shmoxaYwOLiDNFMNZn7
qW4vd9aq37jB8f6HQXURbglOtjudco0wZADI4kzfYsBit4UqZMTTxOfZ1xMPmL+d
c68ooVKPYuhUA7ROwcInmOuDgKyr3vnhRQqwS0QK/68i+4QGJrvXwtYU264K0Jgo
vxzALBaweQKqIH2IrUD67XXUez5RiNabYkLKOTFLDqTkWz+GNcBc3fLYqOBma+Ml
1Eff67Q3P0aY9wzNKMdjwTBeCCmVLXKB4u1TUoQ6+iWflJQyk2zgrpkaUHOh2tgd
L1M0wOQKcid2hjKrQvP+Txbzb1lW2MCqygkvPl+u1Fd+Fu8i6geTZ6um92V9wrI4
kF8SrCgU8By/jldx3Hw0CvCzD2nWMjWTs4NJlk2vcUZLys5dXHt733nTgyXOqSQ3
D7+NwLmo2T4SINcgtUfa2515pp+864CHLM/AsLbCqdOMcG8kyT02P/Zs+pdcC6zh
Lg1g/Hjb5iHa7EGrGtUKcQ0cjdXeXy9YMQ+arKYL9KgFGLnzGqqdEvuLbPSr99t2
WNN6sd+wIS82osXpnhluG1deU1D3tZ0SsNUWkWJVz+ChYmn4SZ5NZTPQ4MR4cxKu
ovn8IXPGlSRdu4fxDyPDvntb3l2haZkeTV5oCmTJ1lsAqUS4iy+verzZTYVZxziQ
O7jVm2iHK+pInWULTOC8jbD/lzhr5wCuXHU3I/MK35NgK7/3+Q6SKxx2VNtPfLt6
mWNwcGLKihAlki7c8QOHnRl1VOPEJlc8IHh5Q39XfAdm1WakLnI3q7dbd2zj5+VZ
fKjGNTo3pQEilIaR47hxac1VIHNW7xPqBpKoNdeYZ84YwvjHY5vu7AcDRHjgYBcW
m5ZcJl/hcCFsTkMNLhd9p6JnyUFctOYsXqvhbQXX+InUkK64CxON0YgX5KfrRT8F
Oy3HXm7DmnBP8bIKWjcoI49BHz3Bvbq8OcjhZWjs+e9IYgvF18mERDex4g+uRlYt
pf849DTYoRkK8k4Ct7gw6GEpzcb/h0/yftVjVD2RGRH03lbZN4ZlFNfNKF/HTbtr
xlB7PdH3bbPX+cWI7+1ZWRP6f1FvIPCNFOyC21J1W+by7T38P1mVxaJ02Wrw3dDc
VdplEaIp7O7J7TYdpyTSVLVNZmN9XzzdWYt29wfrqZM3LqdF8GuZ47rGRd6A9wPS
Wr98Ju6GityxGjwg2deMgFNfpT/Y/OaEj5qoakNjSp2do0BhdfGpWkEtYOZS6eki
OKXT4AGeHQoMyvW2dZzY6BhIxp2XcZ+I4wTJXbtIANv3LmhiK83mFgKeaKy0Q4N8
8NgkdmZhb7aMI3Dqln8LQ9es3X9W5iPldBXfOMv7bgxHEISUinhxbkNJfUzSKjTj
f50byEnYJWdc0VRrRPdeWel8wVQBUXbHYA4sQ6VJeBUlWrQt4iE84+44aba+x6/m
sLZB2KaMDDr2bRzmC1WAK6pZF9qF2Xs+dCmFTPd0hdmxgIYnNyPqzzIUqLrZz4H5
8Dh9xVhIP6V1XLWTs8XuNs0u6a7GFZ3y5RrNlPSl+ef3pVpFRUfmpthfel1i53uH
qAjgRL/QSx6jlymindnSPeFlDFsr0W7xO2Z23zhugnEZaJI+9tLE2sUbNhHc8BBv
VwW00NhI4vjJmkij/v2Sj2tZ5MrdYY9wpWtwY8gh/xFFqrDK3AvghmDJcbS7r9Z9
YBmp3lftBLCJXfBMoH+VU5nXr1bC7I4tt0cHhLyfZnAG+JucYon5EhYQv090FTeK
gZKXcOgtfpsiVrMqPuc6khZc/F8j4S05nFkaBN2nQfroSHzoyCj8QuIdcB5gkyDk
WKfu9wZKxC27tojjV/tjISYg2m0084jkzx3Z3yrW+dLfQwVbAboSWJ/4uUyEMXCl
to20rTt5CKElx3L6HzVzqDe4zm5Gu3NlwQf16LquGssM7lvVY1sdz/oiQHdrHX3O
Gjxsaee75CSpJ5H/a5o9QjtKHtJ5qRx/d/kuwhlLXW83bjCaFtEqKRk0FZcoASZ/
7Lozsg0YsbM8bdEtwQ7uRq8PiWQLnpTSskyp4+Amj32QN6QTJpOYzkeGaPfER7Xx
ddL8W7a6Lw9B7v7YhHmDV0oycMD/WH+gpO675rwPxzl5B7yDbvWKIYYV/g4w2vPe
9fLc/QevfmdyMLPnO0w9/3LlwOVQkm96OHW/q4qcK9VRTFmeONPOTG4BVLXL8JPo
Z4+sjGadsNzcUJBdPjTRzXRXy8lw03JJMg/GG5rJPvgLfV0rGcshrEvL5jbaW5HD
708NqvelYiZgtWFU36SU/rBetIDefmz+Y026Yxi4JFH5egkw3eHWUMpCBIm7oWRY
7Dx+0AiG8bH1srxJFcZr7BP0oBcSx5zDDh+y5xqJwMm0WLUCvvRt8hOxGhETQNaW
DabsNj3CrYDeFzQ3csDhQxZ5X4aslRToFbBl0orSSJAsJyojr8CkoOmwIQnh7xpV
RBNTTs6LVfHR0FEfFw0gwOQH74we92ChFZOw7b/5Q2Uge3oH0jGCSY4a8SVIDmPi
zEbwkR/4MWUo36UybDi4Wk2B2X3itDxsEtjOg5t80kNgN1jKxGRDaMheN7KgKh6t
siYh5LzczD+2QKHNWiKvTGrya0Ssa2yiDXmat74n2Z89Z85rpDD8SBtzJ7CKnIOQ
mRe9b7xxCUG5nalnkEszuHNXdFTZuDS8NyEfem7NeJ+m//neo9bbO/7kkS1S/uMz
L4Al/dZ7o2qrbgsz4XQSApz/W+MUa5KrkRbjZ3gNvN+H4U9di7q3KF0Dqc5QvTyn
bTfGwkUtLsxI124+WqMB8QTbVY1UR7n3Q1aSa9K2+ZkSL5mTJqvimWBFZ/Kx5OlU
vqWsy9fKmi062LPa4UaUDtGIsz3OJGlZxR+yqjRS+V9xV6At/pkPStwxuk/DDJUP
NE9PSh5aCPZ/O11ifjp5d1/Qtsv1uu7X0J59SePlrs/+aMKj3WWg46KtZgeyt3X3
63XINURdn8Kb9OTy9xQq4+4OjZHtNDNKdYY9FM6sFN5wi5x1T4j3PebWE7s0xxYm
hXfb7EPzapf+fMgfnLR9rZT9iGY9aZHVHbqac0v+g+VOV/8l9u7FwQ480y4U1anW
CAoD23Ra/hORIpJKL6YUxD8mtby0rsvX1QLJ1BNnm5+he1o4uHNp6iyjOAoIEsyD
CNRep3qAu2lN9/zhFMSBT6Qx24GVeu9ewYQN/P1yfcQLNS3zro0ZO0Ch3M4sptup
gP3nW8Sf6GTkE97Kuuyjoy/3w6J7gPrqk/vIau8eLh/305IHf6+/iU7CO/M6X2j5
MOmyRBCk5iTalzLtNsHREqyQufs3L/o7Ff8wz+mAJTFvVUND0GBNBhhH8vB5Panl
pgh+WY6Uui1ncHT46b/xMcDhOvrWPaw3O0Goy3XnNSmw1WvbnNTkBHsgAgy3tJM2
ID0EWzPQWfMarL3ziy0VnPJgV0/moCiEv4mZ8TPSHBxV4YaKPrMcDQb922eF9Nyb
4UBSRkU9UCdbUu8PjPAdwjkEBFAEFlaTFZ/DvWkOkm5E2x7/zVvWwTxlcfVoZ0Vg
RfSC1Mf4bSZnOJ8LrflEj9OUueIhkxAnkovtFCRrSw/7zYstcXTAapZbK1yPi9/y
6pJbPUvRHIiShIjvhYNikklhjJXBO4ebzVuqa/gIrQeL1QqQ/usphskiSMoxb+pp
FMzfmaxHa8wYU02ZlgiGqhYISNEDKEG/68hBbpWXQWkN9MokCOw92VyLM4eImn7Y
Ym29jasBdfFvzrUO/5rQWNciXj71PiQIA3wTTKccpPUjXL+hIkdACG16VyRRVjHY
l4qywfdjPiqa2LhuRX0ArKYAoO/7mhmRr5zND80+H57uqSXvfxP4vyMZAljqjuMY
n9nRIcbiOar1U8+xHuhLZ5wkgUdEQeR5epjYsumHbcq94pPx3Nbbyv5EUey1bVvF
f48mKQ7fHpL5GPT/rP5u0xA0qSTdHbtBBlNf3KINfB/k0S+CW/6LvXi3PSOR+5pE
D5ExMhzhQ1NK8jNdMtviHmSQV/OoMPNoLUZLUJEe7ejb7/m55MA42i1rMRysB2So
ZoxQF/naZfgc4ml9zGASbLnqH6BUEPwpCfarmUH2/4ZP0VdCouRWeXkZQ7tdCw09
sbws1tolBZxpI3R+/9ya60+ZWt+1AhogMiDtbGLerIYOVE5p4jd2Q5iW6/lKRpCk
xg1gByi0nTKh0cjhFp6bVg1DqJG+JdNKvluamvjRk74d7yjfn8sD0R4CEn3oXnnG
KrrWA1fXTrf6mW7f8tJJoapkYX24sa5dp/eylzNSw6YNqjR+ZGl/a6RR6wzc6bdE
gw7X7jjp8YUFe5KCFeN26MO8J5nyO2CFQFgZ/C8TqS7HPcDdS1VlRjB6gJLbL8x8
H3nE4ZzYU+G66dG5riQwyud77mEeQzVEaVP3zb/JFB+Xfz6/hbBI7pj9RTrhjkYJ
XH1Su8Eh8OQw6ld7E9CdcMVDTA8FXRCqZKuQcf4ZY3ZybwUiD7YAINl5YpIM/b+u
0TTNJ/Qr4dyjOYoAZGjfRv5Dj+Q3qYhd6WsIT6AURTOsgBiGzugnLiye4qbLv/pz
aYjobTNQ0vfgjXh2Cf+wrcvkcCjISeTXSVEcNFSQvKhd/vCCAhhHrs1ZeHAwDDPa
gPTKIgqHxg5cTSsJ4TnTlx9Hta2dwdfcLfnlEJEzn8jG/m7PE7vjDDYJivCCzY06
KDouUZNuyqxfWuiMfYL7yxB3t9ULVPBySNQ4kNOF3WxONAeo++ihQcj7G+PqWBw7
TTtOHKIG30JJnx2TANy9i4UBIUTqprrXAHeyfUzK9wf7X0cUmQViqsIIpusRIL6D
L1p04q3iMYxpmRkHGBvADOaFkvB6q/QS4R6jU2yRGXw1MK7bVbGRBpdV5PtPHcgu
AdOH+RUjuBnZgu+9Tzv95DUY/F319rbkfmx6NmySjkn2UXbqfMGb1javUGD7ZhSy
Djv2TfhFKBT0pPO8kk8r3dzrOSmhhdAI7DtcwTQQgrLpJY8IfDVqZhklTOWm2JLM
0UIddgeHr3JBiMI1kplgziLT7De2lTGKypsu4tLZk30GbqPUWs99KbPqzNSUQsPh
Oc0BUofvtUpFC/buXSqjPUXrKhR5sEKO64gNSY3mle8/ZyMbAMON0iReEBOPHioc
3TOUpdn2ym4qDawvsXrtjB9j+qfZfOh5QZ8MnyfP0KLqONnNTkeCG3rr+FH5i0vR
mfEbbDZvJnPCux7xvP2o/Ld14/uMswZQM7FFJE0NPKifMAzbuLjnOGFf3CxaOGQs
reuqEe4sviSZ5bo7h23nl7JvDnLreeLFAZ7rK2FDsIQXRDXSUIpdtsvNv9yg7AWq
9WKmU10mAjOBnE6iUXDzBWaEsAxZjcQ4BIBB6VPvCrEruyAA9pZbol/LJ0NPz5Y1
AhriLctkt5/QFM+NQaAFGbKhISc0vqDDQ3dkLzv8AddOF/qggRO/0rrh9NvfQ0cG
D983BwNBRxfYzBXx1JAP++r4voZGtqh1vGvL6mk0KM+/RAKLxrqrYHg4FXqvZ5fo
PKUx3oLGhy7AFFGReh+m+Rh3WD8sRx2LWukk4qH16RneV0pD97I6566bxXJkapM2
XsDp0R2WSKdW66qSGHN0QZ/d+wr0PZD9a09gXZ0DJYbH75qjvqlI7u2IKbWlv+Hc
0UZ1VAT8rWMwPcIifsftPkQ/L1F2A2Sd/Jh65g5EHF2ZTgsCr3Dtc+eQL6KTC3s7
Wsct+w8gsFuRUZYUThDrATLQkjWlE/KBtn3RlEnx5IaHqmoLXZJJUX6DKoX8Rt2C
oH2kyl146LjuIMP6Aff2c9NbxNDmcUNODgbgMR5Oj4jPTDXLeIyR7ZgSs5wKHCcA
MJG24nCQYh2KT7Z4i99nW6N7viRGPGGsXze8UFizTbykar09RiN3ewl00cXQ5+Q+
GUOzJAlxp1H5d2nNoIY8v7wSycxBidBjCyuFNqYmTVoihdOulnRw2aCsLP9UFVJ9
FzNOAau8b3vRfhwQG51zmRQTt2M+DnBbbP6CZGBCCUbsPibMq0fOReOehWtMFP2J
1UxZVo6L+qcLjUiTAtvff6t5B3S/ViBt/daQVS7bzXFq4O1zFz2EZSjm6mFWBX8d
hfuF6D79eyrmRd9mfr2Y21e06ThXaAsqEUrSLKdhtgEY//ft+Vm2CUgspw6cmaq/
ioKCYQd63DTNCO8b4x2Yrz5PO8zVJiXtNAn70cqRe4HGqzoy7VWbODBsSLS/LIfJ
6ExkfctQt+4FSo+Z0WgSQGhotjW06Tq7ic+9yeKn971za/ohDyEastHCq9GCNMSx
XfXnqruUNv/hHTo2Z1T3cCb4qgApH+TGp7jTSanEmtuI1KnXUk9cAe3w735rrhcf
ROtal2iM/WblcbXuqwDKG3P5hvmK7m/vMKgFttBwBd0eszMg6j5HuMGB5oRAKplu
Ko4Qm3xLi39JrUpO7o5Rov5H5dIIMKkOd3Q3ZxDzpduizxmCLhviWFhg6/0Bj84o
L2EWTpqbhn/WNbFDrEL1t4LR+xPMckKR6WQFVAyoiKcYKBUhhlYbQuNY/YANr5K7
QpDunhVBqHn0qUVa/LLv+vvg4V9DV3eZkca+ukTPgHIWzHqL1W0UsZBD7Kb7A6+a
vlDgcHPgO+bDXeKbOcBcspgzzAvKgaTZjl5lhAgHVIH1zZWq3jNh2RfLqeau+mEn
hfBvFmQ4k0VL21qwLU4bg6LCMMHcA9914AXWdqZGcpTaakN1A7H7DoThXnaCDVC4
kAtNktlA1dMY/oKMMbl6PWjSgjWDEstaxVeXDeyvwaeYD70roV9MMvWa2F2B608N
xiOOjH6tbbNMrH7e1okzRtKt67HKW/misU3iuva8mB76lXziKeO+wv68v3TMweIy
x6sTVNH4nRMYbx5xNercV0qHqH8bQR7emHCLIrJSDN3xUQImZgHPl8DeZrbeU9Ua
KY23etIpm7V6u3jNLWgfL2fdEFe+23LZY9PYXdlPgwt0zvvbQrGaaCWmVF2lMzhO
qE8chuC/iD/0Gll7fMcPWKV97tnVLvKE1vtesyJBB1blAv5V9SRj/skjWFTnNMyv
2uTSVYxAKW2yxPbJTq7+AHP0iYkM7vj8iyZ0hLmDFTCRVbrqkIowYIrYjbJmBqQ/
TbTSzAVZZfKvTMi9AtwNekfNh5ngtp26lZpWYHuB7y4pBF/AZcG1optjyEmhBN78
PnceIGuVh2u7EAQhwXUvQFlMKKVb60ko6dfW+vD8IqaHR0GEr3PFHi62DzBL3quK
vekKc0Heos1W37dDNH0EuCEv1lMPym0ZA5ocPJXqy0xW9jmjujwDP71Rs6k9/Kuk
n6xZ/GezYKoy7zYcWczYWqc33uYRPSA3W8aEkplR6uwE7tyUypTeAFYKIYWmaCnR
qf6WyDSg4KEoop+/LxOqKFrNlsDc8br09KDB2OrJaupgVkPQaM4BfhUtBFdQqY0t
54cBalIc5fHshYlE6rtsKnVRyL8RvdafObhDpVbobMH0hvvj7HaFOeDRLR+87hD4
YdaYZt7NG6UjKk8xtGl/tQ42Ernp17FHYffOjxeSVoQuXQ8ePsCkDIKQ7f/tNUuI
mAH5jC3uRTsNYNNKRlPBOmG1oHuIBAz+fmQ2zQLhlSyIWmBIz+DhAra/fh6UXorH
ELwkLbXtJhDnacYEpRMKPPwWeH6XcJ+mXeSiZtl3biMlnDb83yXTV1wjJ/ECKjPj
FZijBPbztr1Ehv5dnMlElqJ1XxeHFNkDSo5PdfTq0lACI+sbKymCEZP3gWR/B1xr
XMFjVTGG2O9M4SHfTVLZ65wdL3yXrGt5Jn7gQbjLDpZ4+43rEuS3NGC7616gklTo
kdk+KL8Uj+r6FV010OVbT5gXgujjopuCWkID0cTUMCD+iiQu4ExpiZRNLnav4CeU
nSdS/K8cLoaMOcTZWSSqmggd/oYHzfvv82sfRdBZbZ8NW70YAGm63TzF7RUEobxu
MGeEf/09aufG/opVQRlDORTqVKTaAgwUWyvvt629xH6t2vL+2fuuFzMeQXv0U8mC
MXZTIu8wnzBeMEqgxSDrud5nKc+dr9UxF+JQYXc8+O1rkktbSxS7yiCPw4TLslfg
DaFtO2sPsTxdJ5P5RFGteEjYPyc8UytOzbebu0KJUyATH9D2sRR14fwQkXGT4R47
Vxz2YSdA/ebeohHphl9TmDaVyTysLIBt9aJDPzs4vIITv49iB2+2oPtmHGLjtHwT
R47oTPfSoYwVVRp5t20lAT+gOtoGifgOykXlF47ObRqNYgp3k3d2JHHNQfMsspM0
jLEb2e8bNI9l9enjm37gZ3wswDPRQW4JONVi8/rRrtOHH4tzfawT0zP7oW/i9OKF
RYKnWBs62uW/hvVwRL2K4+D08dHIYg4tu9qh1JQmkWx4gpW05KmP6U3ejpo7bJes
a5jc56SYH4qiF0eWghPSl9wxFXf94ZApm3XP1D1S2xMESZLC0l8+2b96BQ2Vuj1J
M4QgVDMtTFpyHPxLimWUvoz3gqoc8+BYHgaPFuPIBrd26cxNLhFAvqvwBMeHiekn
8KXURwk8REKK3akr48tXbHT++Z1BB1vlG3jEgsvC5h4dkzVdqJEC/wBFvgpnpkPr
ZKOuvThP7PddJs4J3oxr8N7rtl6/lPZwxvnL0UfDBId3SQTYeL0iqXEE0yWGWqQd
dfqWtnhKbxM61UxZ907mfHS2XKXlixP+VqLiG/1j6nSm6s06l0FmepUZIG+0Bwub
ekMVoM4c+95jDi5QxBCX49jhoj/bgiL7Go3i5VGUGfUbyEdCIAM80lS7lTZ/dR8Y
wCBK/c7KO2Jt/w1qOUDYJPFy5TgSbxNqvZSTg2JtU3463jcevIcpPyfqQjlk2+ax
UV3LpaZGLMAmAH3cP0Oi9+Bo+JiLrdwmVkBMW3B5ybFJqgi59yEES1n1IiYXlksX
0NzSkCilcyRNuL+9ZwvzZNw2+cJQC8vI9nNxe/rP2d9eil4QE8wbulyhbug3Gm3Z
QKK+8LCUXgjgW1jJ6KJPwXYaC8Uh1Q2VzXSOPAmrT8Sf9Lt1IF6Q1lERd4Oranyf
D4TcFiWCqqu2atbwplUEoB3mLiUzSsd8Zjkqr3gJuqXXvAOJ21S1+0k3xnQGvHhI
oe/eGKcaqHj2JiwnJMIz31lV3dWxsJQtQAdMdMh8dg8hQPyyDcuMybw/LRhyNUdX
JyArdfIlbbQ23nkNRAPWTTcGB4tFHPkVz7kF/LzOGoT58i38Et3cKzz+ZkxFW1Dn
X75PH/ODn8u87SfWJZaxZSoYwfQHg3/SxT/hWKrNUnzgcBQScBK/SkvNmYve84Sh
MNJZFesVZSpcIcM8tTg+n/i2hJPzpSvls3yKOt1K0MRMgTt1vgHW1k+T2u97bRRl
JpAFUXq6OFkMsPpzHWyhJYlLjmGHqsEPajy1SC4aqba+65ULDCL1Hux9Fz7v8vPT
z2j7QP4m/481FAhFkr/dJAiVHMR0aPwvYasiHEByuXGvzFKx2CaYFyh4RnB64Cku
yCjRAtoDGH7+AsJKbxPznTB+cbMuaJPS0MuKHI3+WFHVbYOztYUH/a7nalyDL6mh
QsXyH09vPR/k4hL3RA9ehsAoaBBvMM0GfDSeec0BjjjC5XCXc67H/Rgi4Pv+tV17
/uKxoP8vthnt7OvA7jAP7iZ6PF31+jBSi1KnK5AnqhNN57SKNRQy4ul7aKuhSXro
sIJ2OvyTkPYDchFNt2Jy00YbnI5Wtx7VKuYUFrLHHh2Ga030Vefhjgdm97S7TtxM
KOHsnpriAtdqbz828EG44uvg2Py/TTL/LtA3greuuute0SsBrHnnTZ+6DQWVlVCH
Nt34tWfnjFkqWdMC5oIFlwPadXnv63B43E55Tef4O1EHk11E9hy50m05RyNp4QNm
ZA7ZqIC98SX/v885PrmnxDdP/OLQikwa+Ms3ZKX/LgX4OqPhaa8LJdz53U/QE5RW
4X0zNCXSE7fRYZQwFVlYHbY4BvP+l9rfTx9HVUrQStdubhkbB5Y+GjTBWi3PKGvh
MXwLKCh1W+tcFcSG/dJ+FeF7feXUcEyIP6J5gDFftIh9SkEYIdIP4q7KF8GQPS1K
5qLIdQYzOH7CiBlHM91dPY2fxSs5bf66SfC5FYh62L68Y+BYflw0EitCV5s4H0ou
ABul7oj2HOB96R/1Om6g5OJSJayUbocEyuwEAEFIRP7YzP690Dluzkb3To2s69pC
oe40/d0RiUIYww26LTrRUfJOEcq2q5drR7hcRJOBg1CT+kNOfGnzPN5Vx5fWcdx2
+MgDJRC8XwAiJ3Kd6pAZizbcBB9JXqyH6OgTv58Cz/UYna2HIX1uxCVgY/wxRs9i
lRrrtaA5SU5H+tiqbqqv/aJ759KBUU9MMNYz1Xj8x3YGe2dAmrxiig38tQ29DBis
r4m/P0LP7NT7xjfqfG/vRSJVAu6tdC+jY43TXqUEKIRoe2GAiWCfUpGT4+ZoYYNI
I4ffWCbiGzPLzXHLpi9QpbDS6PtaBtkBzQs+b5UPgqFwavpqGsnoFaqEvlDOh0En
PX3Bv/HdXgH1vDmRRxqrjYaHXPuUa5DF/19h8d6fkL9Iz/yQmBjTbHoqWTat8Vq8
Vs7iO3/JpJL6oNB+xWAuIAbLfK5aase1DAcCc6FizhyRG0mskl4C+i/HtEtvWdSq
yuR4XKTC0AZB88VkIvsJuu/50zliQKRZSeUDUUxMYd0N7Ha7Y5uBM2D76AVPdqZo
xRY1F3/yFwC+bTkIpbi7RRh6FE824OOQg4RlR080qDsuTdCyIiwt1Qcg8eY1XAjN
22b7NlzK+IMcW1ipMX6pPXdnC1/oQHICGhlH4YAhK2qLtnD6cjUWuwVH77eqXGuk
Vw80cr9godSjoBiPN21K0NJISMtlt9mUlkLtjjgr10KTVO6el8Rwa+Cim0vkPU9I
pZguh9a/PYbrw+A5fctZ6pGO6uLR0RsTx2gmAvM/OChR48qczAmHQAkRzJWMhzIl
TPMd5WsrkqgibWmbhWxrjVND+Iai/8byr/ktRf5gPeJvZhTWNIZnUnQZm9b0oZfW
8+0wagIk8Pi027mhFdoR3dP+XDSHMFQArEGQ4yvjtIQxVrZvRgHhvzD8ZRqg1Sat
Rs8c0hxmNdkodr7ms6Ju8GwrLFeXPccvgisugHNlcnV6P9QyXiLr5g1ZWGLuW3KV
5JkptisIriJRjCS4tAIPn9NatiA0jRK2EswcCURrBn5cXJKleCRyg3pD2y/vi9wT
q0W3DhN+vX6OQuXOGL3LuIS0Zp5OdTJ402u+NP1R3Kr2o9RK1zHrnElgWpyAIC6y
riV/bvsgmCfkIR+r68TK/qUtdwoDFMXRKK7pMz6VKcMMLI5O52PSst27EaVSD11q
pCeD4amFT7oxorsW67VE6C5lXogS7v6oR/Xgx6MddKzAsUXDJ7jK2G3YAYH2KZnU
PbIF4fK1qhev2h6FTHvUygEfvHvUsHcTuTVTre92rXurFDZuhU4uICsn9p9av+Mi
EwkPzCeSc68weYToLc6wN/rsVK6Sjm8dHkVaNXO1Uhrs7dr9tAmdgupCCeLlb7H7
IWj5/f3hHDOg1I9SNyNVF+Uol5aqNQM/rHflN1BxEePG3ynV2ldzkFXZ/b5ls9p8
BcWpwMxrc6ApME8UaYuZqYmRTsQpP5mQ1I2my61vE5jnCXoURNte0DWvpQd76/zd
CtEs9OqeupvTkr//71BDMMTVBqXX+rTnydkJd/ugcM5f6X9oamNS3tpgpH6Ri+xd
+x5YFR18r2fXM7NZgdWVt8TJbjTDR4FcAbyhHLd0GHRg2Vqefm/42WB+xyu5FkIL
HR5n3cJzdIIEsYLhl7g4aIp1mF7IwUPDNW8zL53OIMV9/WUaOscoXrkw/wOSAXN2
MZ9bT3w/cBZetEbuGKaGGM9M2Sjep8YiNE6HD6BpNNC1wK61A+61fc8pZd0v9sK2
d11RLm4S+c8O8RHCyUxGN9JloIENb8fcKNZDlTZcJc6flgvKu0Qk1ExE8VkgYGKS
hV8Kx85vQSBKNF3wvG9Oz+ha1uR6DOFebjEhRhNHQz5dlikb5lLrcs/79pbZqn94
tP/5xTAmhMkclD9WMhJmD3qhl8M9yqkV9Q1dHrqhzsDkj4k6AdyWL+4H/WA7mTlG
EQffKwP3zIKH7T3iT4WsXQVAvmCUjbKmo/XV7JUoXiyaEm5hJhrvcs4FLnbALziH
ITDzIacNt0sZXO+cO9IqhNECuQQ4rB7Ql0MdlfAZbGK0aN7n4cofs5bWkYCtdaMc
EqrNaPV9j2QYtuMkSpC2OXRBlAY00IWyhs92N5EYl9C4oyuIoEUT+Np8N07MYHS9
XOIweKLCWVQK2g4cEuNyuH8ui960GDnZ08oFqlD+bOOQxtJOU1ws7pK5GJcbA7XD
scBUruBbdBvSt18ERE37OtndCo+m6/CFZ1OtXSeJlZWOj/l/ygBvx075ovihh8/C
wdiLCG5W5bFwqED2jJT0/4VOUR1TxMpsOOpN3T2Tc9ZOpWl+oKhgbs8nvV1VW0lW
kmAph92/DDjCYTy27wdSJyPcta/nZdxHaKC+UKg4Dl7AGAe2Boovu1V9SwyhJt5o
oK02i16kMVRdtzJGi5hkHA0FhGl+1YwqubOTvrnOVoy5BnA/4W3D3fPrdHdsDq1a
bEhDOsA0CfYPNRqA1PWlvAcPizBijeSqUf5h2MgeDfh+wSoo7FfvgnT07xZgi14+
dKS6DLG/S4UMai4r144C1rr8jM8E9zPQRTvj/3d2qy7MpWVSACdkXKFi8Wk14Q8X
mbdMic3FnlziorqzVRyUKuLMfJ1K8eR9LPmzSCc1oVMMpguIeCgpi3x6EgA4lgFS
LW0yFKAzcBxj4hi+N39HmXGVpbeMLpFCLamP/U2KFk4hiNQNqq7+GBhjte0UdIIK
XqkL6ZaIV+AsppGDaloci6X3KON3WMzB0psKcK1k8uRW0TxZ2AkC5x52yeINMBwu
sDSUKI9gKaEEpvMFTVi69LiRPBAbi9Rl70GsSqK+4DnEpdxLP7+qAP9yKU6M8EY1
EJyFEMoKo3S54KMbijDBpzO8vLbsE4Gndb2HTuv/LS8vuWnOJlq9/YZXljaIgxHr
I9IeLH/z/CypvG8GL3yk6BEEoY6QB9ofemraSPCjILjKmFDe216JdyFsP9CuUK3v
8wbYWDVPq17lDwlFqe0+gzWDkX7tI+3PHYhqyMXVKm+eP+7rkTvvLeIzc3xT7ShZ
DW+4rp01wf/R78qhKLM1I034YtoxB1amCBRM+fxrULPX+PSOJW/78KV3zEbAjh/u
HhAr3OCrGY/xplm8IA4VP7TPQIT1v48E1FBOcN5994yPr/jNVxgxnVlvld/X9MJI
yzkMV/z2SHWbzMqI2V+exP9QvsCAm+oXz2KHCP9OpQpEbT2QND6XVuv6rS/jvV86
FsUyS7R7riXcxQlwRtACnzTEAji30CddTaAdaf5175eGlLHrUq5n2Tg8INGiGgkT
aZY1soZP5W6tmNvHDu7QTl8rmy5kWuVq+PlNqs88ls2gPFJyMa3Mmj5dnY0K4Bj0
TUILQ5Qh+BxGeBC3eqqTBVeXgWp7Z+um86VPGedLNInvP6djgp+esXwPp4T8Lxc4
6w/aBWH4Q7KSAZGbJUOFxt98fHiNWlYPKHT6GXjoR1AdLAAMMQ1dXgMDnXD+LaWt
I1PAUKCUTir7mHHKbnqbAfEQuVkL4Hmfac83u/tg+reatkGbFFvT9IWK0wEieo5Z
hpZrm1w4EUQM4I70UHpXb9gjckck3HtHuHLV3YRL5wnEsUk74NQLc8V+JteW7ZUk
SKhdI3AP11LO0JHOHl17ud+etOKBtRSuZ/gQk751Nhibi2cPXEW7XS4PLOskqKVb
nN0NtCdpaASt5Yf/UX4+gaNOY/Nt5PYpgbBLqJnDOYBRLnqZJc45BNOyOzdrGCAs
t8qTMJVCVQYgE1C5kMWR/33QHdVpQytDhOZR0qwL5SDTJFubs23yen1dIguOIrx9
JSZAs5GfMYiTEdDXvFuNNuS8GH9yOOCb3VJoxPNnSIVtfBIqanfTEOaFZ+w43544
6mA+hauuegSlze+8c1CIRSWEaEGKA2I+cpoloYI89Sh5tnLf9mYDqOoqzS/QW0RV
SAs91zgPbdiJoTn8hsPQPCqoKrSV9Dej0Q538YLBEXY3QMGoJcz2wy42pWS7+dTF
QfWrtt0E8/gqeNVP4oGJlYXjRz+aGdpono+kdTmvUtNk9WXwBMc2IsHFY0sWD/pb
GFfbff3ZnlgDnp6u3TPytHrKVSpKlVJ/lJf7qfBbGx4MNxmaZwf+eMwTKadlF9yI
mwMyIvUC/EKFqlhCU6VzEIlMSolbiQnn5krU2ejliOiXFkgKDQhY9zX6JMKr+la+
hsfXFRVPOXBCyPgSKLXfWc8GxHIYlbTwfMZtgpnYjxPlRyAHj6IFjTAj1+jO02V5
jSYpkj2TXwpKIgQ6nYVj83+Y4v3WQN1TUwVBAJhmAKISgu/npXGKX59oQmJ5p5dU
tHgjwOgo64Nl4230nm6ieP3W4nS7m/cUNMXHesHjIhn0wymUp089msKpi7CfkQML
jAlbT5WALdRVi4luo6znhTDR45DAIAV/oHE44fAIK9cZDdlpfAQ5vTAaXsI3vJ94
X9Ml9YvtS4y98OzpMNuyq34gFT6CsgHqFzTQyROwYM3wnmwfSC3jMZQfyHA/PaOL
sR595kA/VG+t2mnwE4PeEuT5S3iiyMvoStpMtBuMxQ853kI3Q5EvQU8c6uoi+GPb
R8W5dycR1E3A8pBQGDT0ovl+8qnv0MNd6FW9R28eSngdcdpAUosZ0PMkz04ISVc1
w/AjYh6KxM0H46pOpVPLtT5TsafUSsH6oj+W8wV9bqNagaQVvvOhO9uvQFxR51nX
uBnNA/M0jJKPPZuUjaF+b8+mWYDy5nCQQODwNCYH+/acr5Wa3Hx9Iftr869GRfrk
XZKO1YvPtDoZL5VN0ajHefNE/Up4V7RzNBZzj6EjvH4NErExsIlDUNFik3ftyi4R
8Jpd2+x4/WnnZ1IrFp5NwKgbgbw90/4yd+l4qBNWJu8AEadXEq+aO7JrXr/uMUi5
LFafPvIc6gZrGDttRi//RLjpv3Ia4lPb9diWPLKNYBvNMAJfhXgYNzgOIEX+w+0i
jjcHDGRYseAA4X3NyudjgWKGnutJt5/ibqpjZcf6sAW3K9QwzO5bViy3/7L5jy18
OPdHZhVJ4IaLg/fwqS3tmPAcL4Yvmq03FUdQ9f7FyNA6KivST5FqQ3H/d6CGYtBC
9HDi6LSeeonTqsiBWcbJ0iZvSjenKZEGaxyZY7Td2CqGnIAWMGjjrfv/ictYQmKk
7s6no178KSeDE/5Czt0B3k6W+1zXs5DY8nqujHoMoon7bEIyvdZpXL8lZO7cdCsY
z2ApRW29Hxz5DYAj5JWQ9WAq49VPxwSVU9MNbFv4ywoO+NirhxiOxZiraqdM9oYX
GNK2qylB1gJ4h/BAqJNEClHkY+v+Be2Hj8v1rzSrDHE4Jfqq26Zo3Ljkzt4Je4on
kHZ484CAndsY0MkFYUrEo3vc0ni0sLIZzGNvzKYHRPthZ2mXs/xxaIy+aT7FvrQm
cm/uZHtm2JwHf9zy+XLBxY8v9DcLteiioZZq4F/Q+zQF9E2gunAUD3YWuWDYrSam
s6mBtlxXgs0HOJ+i3FKlVlPrYZonXN/Q/5g0ccvNNc/2c6ZcN/fGIhDWLMDIvsn4
2mTYx/J6Bms/pWYDOOF5Bc/qzV9eIH6ewlWUnMZ0km2k6wk6YiW1h9QBDCcR11F9
2CPdGEntdi2/yj9MQQFesl/i68anLF8wYCgqlrcJyIyGse+zh0MxBtkG8uCjVTmd
dc5l1Emi1+bBg8FzxPyYtBD3yvqWATy9Pw1NBeAf8Lm/Yk7RS7e9bA+w9cBjksFx
ZfzbVmaGfXPC6g7zHII6V+Sjnz1cFDPWVMNRI89zYQ+rgN0Qod7Z9FpqQSAwuAHF
biSTZBpln9/3RinpEeisjhmEk/g1tVo7tvOu5t1oA4tKWaIKt+3XmU81kRn4MvzE
VNr45HeAi8pFNcNinjZntL80ZaBQw9+shqGF4P9WgJewnslO8ZsoWjPhZHLi1ZXM
XoQf956xaR3IBirwfc8OHFZUFpEWMIKxYPjk9Vnl2yfKgR+pD2shsxuA2TqVaXYW
K8Th2cRaMA/3JyRpJEDHPpbl9KbiOwOwCXbHlNc2niaENcdKWtVM1FK2sroxrw5U
yQJgJxJJLRFy+DePSnLQq2G4bh67hYg1UnbtMGb7OuKShr8Dt1BarkbmMDRBwuMs
PCYo8x1KB19H7lrn+00ujMvrPY1EPFp4W9cXLRxqeHfcXNOTLsELz8D+F5mgrvKe
+vwIH/NUF+maRNBciPa4SrnLf1tRtRTiUxomrlKZAe7D6O0Cm6AlmqN6Imlmn/xj
VQJZwh61xsh8EqmY97fNCkwEgFCOzeBsC7O/Vd2pVVa2kcVlXNdZmHgSSBz+Hl3J
omzJcvu3vE3sGO4Ur0OE0Mq6PANj+qVSH62w2VuwGIl+xqvreY0jD0/LmnNmjK07
iMCzRAibWou/m0PMmBoK0Ru38+xChgRgDxvJ6j/6TRZs3U29B4IHmsFVIVPvB1VY
+d+hsrRG4ZK/D3e7WiI7hJ0KfUVr0Tw9S7Y5rA/esi8TXXL2zzY0Qn/RRbs04Y7F
aUhyqcEspIUTlkwCKvZLg5xbIL/Ss/ndmyTXuaJOl+5scdsCHDYoIdzysnXHjl2I
FKYISR95/L8p/Ha49WPCOGYHuEZ0O1rsWxZ3ILD4ja306QQOSpNigfV8aBQzpxZ1
0y7qUU+Y58yf9S72Al0Swr4DxMnPyClGSKTxZuMXGdQeoe8tjgXoDisKNs9Me7uJ
2IYxrc1b55Hkd1cPjOdtf72oLnFNVUJ8KzPaAVIQn9OUg4SvJuuwaFBP0HjKjPhO
klcBkKZx7bbVDZ+sHgZdQypsyl+HA+at+sloevT9H9pkEzwmWe8DlWZlNDHBlK+K
bnkI9F6UBZm2AWH7uVk6zaYQAd1RA9cnrRGmT2i/0UvtV6qO0GHTny14wCZs9LiH
HIc7MqpAQQX5y7iuXQhLo8omwDTPUn5GnP1bfYMxxnznJ/PawzI5sGKzz3aLnlpQ
9mV0szSZBWYcxdgmfuWVYaoR9Sa4n8UWR1rPZggRyOWhInafGBfusVPS13B+0YrE
sZKTzYeK6obxkd0dIFqve0mj6Pb+iTVQbcTpK9A2QDaFhWy2B7QdeSVW/+1jTIr8
/vCvgvDq43YZK0ZYBY0atb6mA1ZSDb2xKBYVMwAZM8hT8WVR/AU2XU1MXx0kiwhG
92xBLJtsCJgT7mWY4Spb1CW6DNc5pr5mw7FenI7B1f4b4d7Ik6l7RQ+ZlCFJNCRc
BWAYE9C60FVoRqFDvgL5yfFcULo3DKit9j9RNNbyJfAzVJ61Kkdi2U4obA8aEbKb
v1HnElYtlMpScOykU+PjGhyYN7XZDWGYbz6301NgZfSUJLPX2Lf4KteGkmI1goYt
uXJyQIYih6llbSI632sA37BhOi3UBTgOyU+z+TBZFbm3qQ0qej6Xjgn+Lkh6leuq
F+yxC0+lW5CjwWYN05iU5K/3y6mgwLVjLipG/RSxcxB5tSnAb6O2NMnw/3JzHSPS
2Ol+lUBmgWr1aqYbUzWrLgVA5Vp/3fT3+exo1R2O6SR24EklQ94PRINdUIWARkGe
f6pWSaL9Dlq70vo40vn/vNrs8e9uSBv3SBdcA2WdFGAX8MHPXfdLpDN473cASZrI
NiRLOPg61tdVwa27uejQ8v5/i3neGXZ2jZLxR5d1A5wbR/K3KdiOzGgG/cl9lfDS
NcvZHYTR+L6Sy2fvrBX2eWEryCk8J1fLsdAp1paBo+iLz7acjE+Y2OyAX92hUwxu
x2Kw4huP8vKQDkE77RKMt+/3Fsk5uNIa7yIWj1ofNrMZ+RaKpkKkWcfgZV5cDzJ6
Wm5TYsG0YRgq7BjiRuH4yQSS8DXkY+IYp5ePrQEqJIpGYdR9BCc/6qGFBRTYEFbv
9yLbG+6TRcDK8kGXRm1guUR4PmX4+YlK2ujmFi/7mozjFTpRGRZ04yA/P+fmSsY4
6iwEihxBe0q/LG/4GJoIQGkHR8tjTLiulnKOEVB3A04v3Z0twNyaX13yHQe01Ekx
ljZwVf+VY7m27l/2WlOmtOb/kUqwPcCWNE38SsthS9fPXRsWQBEogJtksJubkpBU
g64x9+p3W90zQYovz2tYt6FpOK7NoX0gbBf7mVonbv0IwzQWmMGDC9A4guicdH1h
3+6g2Cyo9O8Hhf+uUak82FD1ciRjCuqt/Ihn3k0cqzulq4Bw+xzzSJ+3xCPguf0u
/41jhwJ6aWY49AFT7OdUWvNu4K3IW8pu6hyZ5ef2eUXt5eH166nYqQouLsg4Xtz2
nUwl2AoCqM0ExVs6RBt+B+nNhxHz9YdbhZotkZCzNDveFfse5k+Km3o327LJlg3Z
5c2czIvS4zST0awADR5PZ3/z0sVziBKzNvlrBf4p1Fdh9aMODbCzkxhutgtewVO0
6p5ih6yaBtQOsYsXuqvgoDpke60Gvhx6lamPr5twD7haLDCRM4bINYNeecPMoAxy
zoXhTEUswZPSc+IaXLygHuQ8wOWW3P7/4htSjHE6GnYqii//RI5g/VYfM3Qyxm9N
ZoSg6D88i+Mk35UI9aMYsJrykuVBEC94tQ/Bi9USUHJHbbPODN3wQYPHlFHZpEXy
QsYC1P3v3GIyOfQpnCKepuNg9KIIAc886N05O8ONwUCIhnS796BAdFLU5s14HGTB
uxQ7FiCBqO0kmKd0VZTI5FJg6INH0H82CD1NE95MB+syyWH+jFC3wqyZEGxJSzGk
0cGcWZ2PLCNVXe1V174pGE5UNS0LyfIPwRTP8dtr1BTS05eqgjLSukROkt8PfWer
Ojd1x6+qny/sy/tWW7WHdFhBjGMWgipXQUfX+fOiqdtzEFLld7xvDqWk4W2j+SBn
8SyPUQA/Vbad5SyyZxIkg1v7A9ViOJ5/TqXklizwwPnfidhw6/xfYlh3IPlRq4bx
cRQsvpruSkoqM2SU9PHFy3DWmXLFiiH14teIskeSOUPMUtNlrz7oMytkvAWlwZuS
oymZbDzwpBSXBy+yrpvednMaxaJMpAnP5O/4Kw37p49reoSkg3YpySlUyxZ8NiTN
zI9BGfd8PcNCPVTOuYin9CASbRdQagbUtfwBFIPy1ej9jx6hvQhQweYz24LE/nL5
/Qy7EqAoecGTypH0SvMJqAJvfKgs1LTs0C7F2+n/6ldx/TSZlvRHPWjgHlpeQfUQ
Uy5cvFLLY/17/2sFXOYTORPmnh2NcPOzIMx14dknNpQB4bHtbplSFqOJzqCeZo6e
F/NMZ5BavF20NHBbM29R4iGJ0xVOiUdGyNBzxoCF4mzrnkLWKC32KWDC0hEVZFyk
H4+V/52Zq71X44NSuAAjsfsJxiRgqGBk/HA3qQsI0DZtu3bn/XAgfq/bTEdwWIVK
CDAg0/oIEIJljs6zeLlXPbd2PZ9/sLDQwLCvJvUNu+bYpkJJI5z/PcgYGBSwQxjC
qQFDD4QauDIdFR+UKdpxCFmasjgMMPwlM1Uz2RZcnms0P9jdxdkOBo0RkHuaDoJx
t572/bpg5Q2TfLvJ++SEHBIbqyDPwYEsP2kBc+CzYV/x1RMDcgxojd3AItv4QoIZ
o7j3ZGLkic/p2lg5GsCjtscIa5mpj5BQLM/SeKp97nuVGNF3juMFSysoVQyD678q
6lb8LPoWLmhVd7vMVGbMPyNpOw7qsLKEwDA8JRkY56hUiCnehzZYz8wiD7yq9Tvp
CfsvK4KClOLJhXCIiWxsbpd2T60XN5u6zr4EWz8Kq/wUyhpBXeUw+6cZecmTBPyc
xq7j545NgQpr375U1R9sfCBrUUPeqxBP6FrTwG6Oo+FO+XVqGdEEgaLYKGd2QEZq
MEBXRBN7XxSHJ+gauKP1U6/6P2cElbQhAJQD6m4NytcIXARxKdCoyKkNGisiA8Ph
ciK9b+AhFMeVjYuNs8DdISZL3nrvxrwkHxEjtmlM3mjLiHuH+kRRZzH5AjNFtkWF
m11F7ab47WG4rkbsZMNXnXZrC1b59DqLjPpOjE6EkxtOOtg4HcDZPKyI/YgMsr1S
WR4pm/Cy3R5IBePgobJY2N5dEDFeQqfNcqoDx3rVQdgmPlA17eoVqI83JWvv0t1Q
mJKRgLjsiea4IpW70hdINBR2raL6wVQsa2AMIA5sx7TrbBNlx7279uz/EsKvqY7l
nRsxz/u7pj2VaZAPum6KVndCppon6vl8gIWjf2+/j2rTXquFzR4XxugeAd5g26oW
Tm0PIu0LGSn4dk26GEZzq+9TAFAWaLQrPCzdW6CRwxGpyNimCGnOp3RJqKMo1spi
78A0KY2UDNwUgu5Vp6SVnAqZt7XEikAuk6FEL3758Tqp262kza3sgp34P4HO3Tnl
sPcA1D53kQFO3SEfyO5EJCh+X0FqD5T0I5BDPowensjUJVis3+J7fLW3XpkC5fAr
X7ttwnZHNzK1nnboRRr2Wv0WtqOf4Orv0WQhcX6Fq7pmnjUk/r3Cmc3sVOz33SZ1
fBzl/NoDP1CHnCpXlx/i5gn1dZL/TZR14ETv+VC3UNQWo0ISuO61o6mgnuAuEpPj
8gkgcnIaFZ804o9Ubw18UhO4nMiuOpMCpKz/udkbyOnohX9QmTOJ6Gh2i6Yij+QB
etiEPV2fNMc2B/nSkFK3N9WRsNcLzz4BBmqXn4kMK3/ILaXkLFdYiOAkYGerAaVz
LIsud3/qDEmJekGtzjltnG1CwPDsbeTGh84XyJnW/QJqjjs5V4+BBFnMNnQWR7ki
PLu0LWqoWtF1N5rSQe1b3HvzgQsclFiDkkar8n2NRkHrZZSs2RD3zCh3vrAtV7iO
LQbvoFghXsLItaGuB63kh3wi3lfGPMTWYfA2FxTMCvu31yk+afJMmrOkkS5OBRFo
pgvHPhY5VINaci1TinKCKwfidOzL32SwNjgpsV0tSM+W26UGr5UTuNuD4KGSo7zJ
uEpDFsvuVFhsEVY5LQwmZ8ZlUEem/xOUniXq1e59x1NezKXQYYfYiExSNk2iWsEs
MwwPfNyIA7UD+s6mu7KHPHoVNuxrdcVXZFq6opmneAZIr+vdtQQ2lLsAI4VcHhXe
sOVYErVWJzxdLImFmfScagkGoXGaHu4CmVe+6jztPKax2N7ld4kpOc0xoL8XzRmq
XIJcI7EixcMBw9h28aPOn2CsaVzncfEhYTPiV9lMOBIvRBvxNvYjUqidcgp5/jRF
wmk2Z3sN6Ia+ZFU7ToGdYaX7QpftcpS4zrN07Y+MGW05SDUjgrWsTmWpoULzkT6C
ZVMpUoFJ4jkVTVO6+hRAU060d6Sh7LXAH1ENNx4HMaTBKqvgJpCo6UGGXuxNPWy8
3D2tD6niO1SVeE2V9FUP1/cFZviUbkfMt2/J/yHJjFAtZqOakHBKWkNHbkjd22nN
b8vNRxCBW8VZmjEeV31SPKeUQLIuccWpPiK01nCCMSF+t9fo+uaqU2lRFShmMzIU
dJ27T4/kEGqsg+wL/QR++1KEWampso2El6SkmUBHjAOLSzz/nbyNWOfLzxeeqQpx
vC3XXnnQfZr7eiUTcdU9M1o1n3eofXglVOWqhCjzioB1rr120m2druvqRXHCqsil
5Yj8BIKEpG43AVGE2YKxTl/Xk1ayFsaF7a4Sx5qWmxkSXw7Pa4hNo0zuTMaH6e8q
z3lkB2dTE9YVDyXLgpRvwXdw5IRjG4MwvwoDucBsiqzahD4WwANIY5+KUMSd0TKl
YESDrtvdkFwOBqclMCeH79OdRM+NLGO8pGsQ6eWBUgYZ82e3e2nQ71CCgi1eLhjC
rJdFtif/Wsq5VvlvGSxrj5dYFqhYHJ+O5GESA/Q5vjchZbLqD9JLCtZ6DJV2IPC6
5YySOaAxe1UFwUmxLHD6P19zsFXxtwdQ+KK0dbw30zg8X6cl0J92TcCkvPeTmceH
6glFR6IHmjrzDLzm6G3rebf4eDOEJwPqewARbvyJhIM/N/dID2WDiNDu58uoIGHG
gdfR9IpSXtFOgF3snqKD0XD9LEft1Yc4sso0zbUQ+acILKjN7tLmfW09D5v/q1w+
hYvB19c08LUXReGgspgVO9aZp2yYamYeNhOjpGkkwUHwU+qqUazd+cycB8D6of14
rGh6yhsIC2geYc5LkJj0LG3iMN+Rzc6xW6vmK6SAL4MzZmKICMyGgV/8EgxCQp2D
YbNp5sEEnjMya2JO26Ry4g/QNlvLPEeuANolNsCnGlLg19giKlMhRAqfJqL5+QWn
FqfnBOTlPSEv91IwE6CqWGf7sE8zRUjjRAXcVO2FWjtqu9wnItVL9uWz4WIPfyxv
iOMIh9RMHWzXuKGbeqNlCsuosUj4KsVcsjhpa2EcL/nL6TLrfuXENrbp8OebJBgo
oEtUOcX1x2FkFQWW0/ekCTOfzqNWXg3FmwUmXTezonc+ssNC5iqOTJQZk0VMEbDB
/4V6RTa0122+XmTS5ftj0o/jJjH+PsA/jOBPrCk4IbbRPPx0DubuxEKQRxRMjaVF
wWXSwMEjaF8ynRf9P9GLtv6SmYaIQ6DBsoHZ4mnNlI/yJRANgQANRah/UyHH3KnL
Qvkb/AIWmqnJCWmkAnDk9GVVEXVkATpNLmo2/pX0Wkyt5zWKDkqwJTzP6Ox3PHdT
ymOumdcLHPGz32lwfY0+/oaP9tqcBoXa70/SW1JV8N16K/YdRS/fRZ09YieuL3Mb
HtsVyQXP4CkGHsIw8sKozJDuUsHzjj/vKlVS+RiF6QPeoxvEPHqv3ynMjgsSBqQs
dCBX9FA9ajNCbiUIaG6NYzpY7TqZ1cXrlRW9AMQLeUyUbdRfmhsC6SO98FSrrSXa
2eL0d4eOXU3Wfn5WU6L+OEsxx1OxDaiMq0jdp9qeeX0Ib/BPgl34TC9TDkxYvC/v
rcBpBtKsPlWpukgu521IB6IGTVLquSgUkdzejDJGc2YbA4N1QByr+LvaZaANrTgs
ApL20r9Nyk9WaknZiYAWotBNaq+jOKpn74ZjQC7d3ZZMcDswkA1CxoLqxY0avgXa
Zzmbex43pUtbPpN9sfBJzcXfYS8OdoRfwN0WEZ7vPcV9BHoCyJCOrVlUYa9kiXBL
PFVcRPfjb36AULBTkYREqLav54V9dbM4Rsg0gUVK5pvZL9vQ7UOinsnqTtwV7yqR
0i56Az9gs2oULP0NFjF5KEFnVWYoIAuKFTqTUHNMmchE5peYFlxEfSgtxaZkXYWV
0DVgvIC697uXf71i9NLLecfdng0UQycuDekubkOMZOxc+Wn4FC7pLqbn83/L6CqI
PkYjmrj+FeI6+CdUuPmi7IfFYYBipg+OWBExPX4NN4/INNFyk1LGGZ8ii2+3EyTb
Z2FewUfbdqfF4ddKWSSjJc8fz19pENQqjVQkiKupitrCm2qFn/B1hKb2cYeDjF/Z
4YGXdGy/UqjAS6mmYTlNHZu4OHCfaWDK36Uo9VKX6IBkXX4cZaBNlFLJFLDkmzzh
reqVo3CaRTjWu0mGrMn0HYKA4D6ym45WUZ5+qSEKKzo7H354ax5YMaVcy4FXd+WT
GE3iMYKYn92e5MewI1nxoQX1y+wy8mVp9lawcBwuCm+bUjIIlTo1T7jzzKnUSxWV
e3WeAjfOENBsHMZwgOCLDx5RDsJdDeUXi5o2MQcSwb5ts5xCKHQwMXh94Z2Afvs2
+BlWBMiv9Jv4rGdw8zNcpN9qTCI3WCE5h0JfLSvv+hKAQsxjuXGCSk5mFKMsfORc
fxugMpfNfRaXL77YzSL5ZE8aCBt05exr//Pczj82lR+jVbHTqit88iQWV71+PHEf
e//eIiJz1QACjkm0/QPEa3IXTGsP8HdXBWDOmfbRoXowtpEqQkZ/M+5srrrApdem
tIjPXjYbKdPv5/twF/hYkG0ZHQ8CjnkZqIZpXLXeM/Dws35pkuzT1bJSBtH9DqO8
xCQ/xKabeHcKe/k6MJ0xL8jhzm5sHD6qjZc7/z+LZ7nPdxS+riw62Yxh989u3v9P
JsIvYO9tdOWXjAusuobXmgR3XLDPfLN58xMUJBMtLjW3aK1RfHwf1e/HLLzGeXdQ
uH01CtcfXyag9hIwjaoRX4pemG1hPG1iVRNsMDD9qPW7zKmIG4GQFAX5Y5r5LcgM
GTSEWu4NbjY85GaCnkK50U5C0zhnnSDUuh94n6rOPenELP3dIClHaLmcH+Auf8mm
GDnn/LbUhz7OQrHhW4EyIKmm+4gykdvtbSD87rxxc4z7+F64MpKZP1h3vyaikVx7
qzg6wGLilJNPnxoHRt+iA7gSwPuKSXvrJbslFMmbDJQKcE7rVIq4WiiqrQrbztmQ
6XNndeObtzh6bi6Myd/IHQgZPwMgggJCncMbCOou9BbCw8DLvW9yJNUwaBWIhWjm
ejLDPlib+Hhp0iFuDwkWW90b6F3NXI4SyLrchv1LkIvusqu2hZ5+LXzhJV/tifq5
GSMccQbs4VxWrJMSK20uoxMY89PjUk7eKRL4ljj2HJWtvYWaHIFIKaWIX+ah5ypK
nd+si25U0Z+BDsRG/MJespCI4NSFdPRol7Graj4+PenK39evtH7bQaMkCeYrBZfr
0+6Ls5V9esL0M6TBTnjtXqWTIbZNZn6VrewiM6aIIDsBoCUdPe8AmuDdZQNLExjk
CWsSpqwnhmvacsjrHZR+J8BANL7OZKHW4zqgOSxF4RCz7Q/IJ7VtXdZ3XuSljCpZ
PV2M4QY8Y/9Wp8t0UBUHpszca3CMR/5uOnPluMxTs+unKgSBqbFc32R2eDLzmEbD
zVcZXsYDANvSVG6ruz5zmaW6jcR3iG20sRJfJGp5g+UEM526DxR8dl51fmuC3Z6O
VpVuVyb5lUaqc1ofIhuHBcnwE7S/V0OQ5kayEHl7VaKN5dBkuADztcn0taZ1RIH+
kahP16jxjWXfJO5UreJ1+SIAyaY+RLFaUtK3STMJT95oGh+9YBkZAyo5N/73D8oJ
upKMweCltkPkAfYAwfE7W8ECdqUx6FRAIBq2uqW4nWc4/itLnYVw+PdCbin33npH
AvmhrR2QVSnT4XZ/YCq7dGVpmNCxUyL6IM35Elm+Tre+xG2ITl0ChYWw0DII35eo
pVlW8SM+SR8rZ/PoKKuk/DIHoivIS2nR2V4I2UxyRjq5YkgDbfhPdrNUYS4oEH/F
FvOSlF87k02VjQFjpXk4ek2S3oLhJizlvYhXc0hmn9J1zOytia+lTRIi2NR52F5O
8lCtBHFI+AAdTy0Cd7s6pno1Q5GbIO2yyK1uELZ+HZPEl1jZ3O8+eiRxUGZOr38q
dPfCbCumzowvQqLVzhqo1l86bQrZrfKQhAx+3OxFFUkJ3QhcR2S29DFaciTHCczL
vy+SrSfe5kjOyAaZsrJ7eiOOZnYdKwbuyFHjB8/LHAJBk/bvEId3yo/Y9UGCmiCL
DzVK837HwQV8cB/i45xpRwfBJJloEqIxi/3BMDZmEfMl7cEWHO1Poo2fpj+G+5r1
NpnCvrDXSq/wqLq1gZFwGxq0gCvnxKmVdnqQEqxE/TcVBj6xR94LED1wDun4HwLt
uJ6W6TrfHe5T6MSCQduT3YtgrnQzW2TEYzGat2M8bEiAIre6L0K9TUP2buZ5f4j8
HFWVzkKMHvYdE8oqxu+tlNweqquXm4D7V3/E74gEtW3kYpx6wIO4uaXAqM/D7caY
pxbMO7dBDr+bvSX1oR/bMnoRI54PXivOqDNC0+MATc+P7sIXu2wRefjhPPI8qAtj
LGtxlTw9RbZllmAlhmITwfPlijNZ5iUzc6/EKqYuesDWMSLsynMNo4ZSv6xlp+7k
0P5jpWboJKpX85esCzn+xFMgdVvn5g1JYgc3m5Fc5BpIszSREoSeRrWSrOM1j4Iz
9X/lOLpavaMq3jMFL5J+7OmOAQGATMpYFa4BHhPXq8p8Cg0tJKI06yL7rj6RYIo7
DDi3fdNfuEBbQLwlvguv8TbMPGZ4nKFps8y8C4X2aRns4Cry7Qu84Q0BoNAmR74W
eVNvFVOFR5mDWna76EHOrrzugl87gLTs9wE5f+PMedLCxDPtQztbtFhMIeKZrMR2
6Cxaokze92C+hMozNIA99Pe8Sqg7qkArr6iMfXzeFNQWJXO6iG4bhKz3STh9WJIF
te4P/uX1wzlcCgpjekmwzpgMfYToakBbrTF1+Nd/tYC8/l3vDy/2vW1bR/j2JH8v
SLhWdH4mLRGFj/lFDTjZIASLKpLaYFQMXBa/94re5RDL5v51QX6I0zjqy3VWhkdW
bs0km2aZWQdpHeREC9qx/T4roPlfpu/oeIskMrtX3y4g0e2aexpWKGz4rp6cmOwo
9YdPeeFy3q66c8zLdoXGorvBtcLL2rw876PQLsGrsVR718/e+9teSet/kgtuqMxz
OuDIixo1X8ioYt6Wo9pm8GzWlpORRcGrYpElW6mrQpiNwAtW9nVRAZlnLpp4xu6l
/dKtNARcOP4SeHd1gOV227fR6Jyxd/UR7kBc5k+ofw4bGv1I1HUJs3fPSTjoko3y
Gxkw+RQKRR6VzhO0s+4eqXUhxzyUROThqJnu9jrRHWPaNmN5WSnUtFcpWaffAQMH
wcI27+uaMfJapHMh3qjQU9VCxGVja5kEgaowIRSL35ZQBTnm431vGnNWAbF+d93O
mwpg9XJg+f9KKHCwqpG5/xwXJkBmGMfqhhdprIaWinGATi6HrcUlDyl4PFBBILY0
9o5YnQctBBq1tNo/2ReHDoUbFHpCHSfufBPEG+BaBIHmmBq4eALSUlKR5CGmMcgZ
QC0XSI/Glc/YtipRz59qNmo7vrUGmoyyQG2VAHthJN2b3ml8+x3tNjNEDpzBWBVQ
bPqgxMspzTtK4KJqCNlZOZYguqN1ALbiN/6bj8HQ6aAc+TThYfwbu5buNnuRsAzv
Md4KwaE0y3NVCDCjSaz9m0kGYqXLd02XL+z15h5XLejYPfvpgjW0fAlMqfU6IYnU
W5x+Kgj5DkVc0vXNocpanIILNkzjR8dZVkoSToauzPqmKb4JIU+iTsRhJIL2W+8A
9sUZNxYg53eN5ZOOvaQYlGFs+WITb+YmCjrii+qiwE6Cwqzwwe54acJRkLbpei4T
Jwgsj7TPEmMlLBh2REpGpcE6IvkXVbocJa9m6XcQIaqiq3rLE/TgR20wcdRK2CXS
tKosL5upxKZ9Yk2ESqZWgf0AA1HeilFW8FJuzSbJpP3StGaIgby8XJrNntjeuPSE
8BOjBYr9OJg5H+mPFCXGBA7hx3PX/mbGzSx+hvYdT5yNJ+ERlxPd3CMX3W9L7k8W
07XclxlZQNf//mpPT1K6OEtsuJEPHxR/BBBfMc5WzYXepBM1zvkOH2uSF0l2Kv1C
YoXwuN5ItYasRiWPRXhNlCodpw6QAM+DjKr+KvBirbYhzvidkDPJEksQlLwHb7j0
Efz7NME/KYbi0fcwVapGV867G5teT683pv0n8zTD0VmMdoUqdNUjq7Q4/m0Wz1JK
xDS5tEwo777MFerHRxY4pdL26ISFJXT4oYwJLWek5K5u9HqQsffG3aWwzqaSp8Vs
U+kRvtLW0kCzyk5JhE8L8K7LNiZFNbckaLB5ije/UQUXLEOHqMyNgujM1yWqi3BE
kvCd1SHLYqCbP5twtFw9p1D3ONhmb6qe57b1QKEC6EE0JBgBPDzvvG1zLZ0xv7pW
Q6haf1dXasYOlIP7eX0kcDAJjPc0+5L33H/283aVYfoBetcERA7zoi2LsHf71iTr
m24trfCl1aI0Zk7fspitW9s8LXGSFafZoY9FZ7QR2DVqetSpU5habu55FZDyVF0i
0w90MECg8S4fMlb/I23cXOZi7uK3qEBR4rBhE9PZoDRKpb2iqc2Hg937HdZafhvW
DuVUlCSMG3mFaWsyriCyFnmrUGtl5tc5ZP+wCSVdrludLMxvd0kqHfES+FMxDKwx
hpzZefyW5MbiWCytFfc5j6ZSuLG3oaHtjKt3zKcgtURk7yeVVsDPsyUEP1tr833m
v5KNpN+RZiqfpI+rk+tdBjcwZtTMpOb/GNzE8qv3RXUGLEtTERJfxo955TeDetiU
j+mdxrwFfufsXF01D75GqgWB9KS+ZLcbL4AdW40pLUt/f7rqdafzMWQkHHGTK4RE
KRPiESw9eSS5DfAYRvj3N6BOxvDbjL26PHDA36DXi3Iaa4rKg4GomfHrm5Ld9lOk
cjIVWLxbTODyGpoLGXCnrx2eqN/eyEVWVX66B7AvoLjwwwl1jbYSa6yU9KEmIMZG
UpzVKqC/7fUMToQkM/wwnVeHcWnR4korn/6wzVYKJy63YtTBcFuAJggTGaeg1PMz
S32nXl2uyP9VeRnh2Zs2T7lno9pgKTdEKqHmDIxM0cDRBWk4d3EX8cq5/hYSVDaD
3PJsgZwV8y7qeOq2FhXlhjdbL7Va2VgLHomFwhIweffWHnbg7SKnaOc+7b3sOKN6
VTNINVSDw8tFrZXwk3pd2rwKbcgQ4Tw8dy1yAfQjYDgkxJDGUUbcdtKGu93uRu48
1SfjTiBHhbdK1WGv7OLiWrGO6ZWtLMoLwiH/7fl9b73xpCoOilkl5s/V5kGUJCgt
3gQ6OBTkavSIO94YLKM3U3GKRXstWOWQMEwCKin52D+jagKDlF7KyBSP0x7C0u+T
NqdWxDA78BXzxg2V0m9nAtsvG8j+N2zxdAe11N5P98gzaPoMNCiaQbOWaAXJ0vM7
/Gas2DU0+e7sschTLANWGvAdBxwslpQ2KNXwg4f4Z6Pz5KMvOJm7rwZfx3qybLXy
b6obdCK3Nr2wmdNQmsbwUk4RptynnnpipJrOkysjCkYo1guQ63ePRoLMUclx6OEq
AkL2jRv9W7YTyi7FjphDs0fL3CODYY9tq9LX38AZKeNmi3NxDXHleNqkc25u47Cz
RfpQ4DmLnu3rnheMQx3oGK+4htFG51BBXLOkKpqTXxms0chSi8D6/7jWEBFBE+dz
tG/ZM6BLToZw+9dSHWd1hWo/lDAr5y48izKKYP9FBVDvMu3dXZEWlumW3BmPZ9j9
a2F+0LHvz4bp+UP6gAJ6fuGBAYtvrFUmkgBAg5y0F89OJAT93oq9EqLQD5pGgw72
94gr5wwfYn9zwz8Q/j4FMbfmWNjaB6P+4noK7n2UlLp1RteQtd4ikkGdyueDmdWz
N8BHspp1/M8d6EQrCKkF3U2zPaY6sH5D+gDWhwG1e4BxHn2IzlaeKKzgxw18F1Bx
Rbi5aKTitNc0Iyj4rlCYG+gm90+pcQxCDxD0M9id4NwUu1rbA8RzFznsITHqaOv2
xzg2V0TQYE4AnSeNAcxUHIxPRqkFq41uDSCevWp7y4M0Ugu7hfoHwvZAbGoEkwSs
a7oU5+8BApa911u80MM9Zrote+5OQwBLd4CJEOw1tfGjlfRGVM/VRLXKp6ht+iMj
aHn62kEnJ2ab3bacR4gpzZupznAoaOTb4lSQYLcK2Dhz6Rh/MjFyziLwKnB63ozX
CE7bcNQLVQVUPKtayFpLfqw0XBRbct8kPq/JQHTZ7KAt+uO1cssVV6PG+LWAI2ti
PunY6GMv/9x4uBZE7tzODM9hQmBsV7pam+ptsEZA4Xo8ul9Rj8fsQpn7cvpxIL0B
8WfuM3t2kI569XEyEYI+7iASbQL6t4RD5XPopsmCT7JrdgGn1i2w2Qm45YYh07AM
xloVMa3WTsbZ5mKnHiYRMo3/UYRsBh+ivRUCko5/0AkMshJm5XEWLxRH6hq/S+/Q
jk/R2/uthbX2DYVPmZ2SXX00JIhKn35F8jeDK+aDxACEsMxV4B6/CFm1eqlOjNXU
6F0Mb3B18K8oztWIv4hdX7GqOYZsd3Sq3ZOZQHkhoRsXTDet2m+8ORvRruPuoJOi
It+1KXKr8Oz0wvFGCm045hfygwOIS30X7LwXnj5G6yUJuhlfqYqJDlFzo9KECVrY
SOTjvR9f/xnG+D57MbCIAmsBbrFEN+juj60avyVIrL40CYLd3nZjvNM/TwEtf/T5
DVCLUrHaTY98opgUFN9NvLxe418op1gXlnuZnVnw96aaN86GXzKxCQ14nGLzKyRg
BN0W26qGtkdp1ozBI2jC8ILW8Wdh9X5ymBLsHl/Azcrw5TdLfvbnOd+Ss8/MvqPj
MXjCvmgsAHqJMMO0zfZ1GFd2VXgF8vLxEvzp5243rpryzxFQy4S6GgCs7UJY4Vh4
dpXm/l6Chw7kTC9gVENDsEyQjTop2ADZdzEpBokAzvJdd8emX1TZXDiJYGcEm078
3F7ezlR2ugKDSTwESxKdfU0iSXCWpqUvHkBchZBz3SO4t/9ueiy7VaI6q9w6OAZE
nhG4Ig5SOVtG8UX1qJC7yhb2r+QSMhElPx4KcPqE4G9xG01lB8z2LyFcy7zO+R7c
kTXWvMaSkuBJjx7kJWDhRYw+f8/svXljKb9X1xd0Bt2rgxAFN7F5VM6hoZ1ZKve4
sFUPzBsQ6g1uB3+N9D2fbHXPvu32rPGuUiAwNmp5sxP7BkmuIacD1rCv+LcsqEaw
YMS7u6dydTmtHqZDBew2wwOJeaOoBhBymqQ6wKUBgjdmk+Z9YDhVtuQDl1UMEIfY
C4K7zXTj/mSJAK1qsO7UdEHbAbe6Z+nqHqgljLG7FwO6OccLM4qbweFZOzpCFMQa
XA2zUd3TS8P9E8DPhMwP8Mgoj++zAlY/EJ1WgWbIZ+Wao2QA8FzPgMxJSNPKJvIl
3Zp4a9zi4DivY6EbkoPETrIZEzY2WyLEky3/sg0e8rKkAcSjSH39lFAl3c0wWMNa
TqtsayrJ6z9QR6Y44YC8seCMx8NmJO0Tpv29zSnj0osoKsFol+WwYh1VFBxmKwTk
eOZhho3UgpU+NoQpu+zK4qdDhtNTCrGuS4E6JHG2ghW5LHQc09hOTnvdy3AYW+YW
CFPWFVAZboUZXJBG8oDz5g5Hn7tfp3Pt4jYB/bPZskq92gSChinz3lrg9slmhBuX
s7fgWuyCao31br2jhofLhiOiyX3FyMC/Fh3HP2YEL8TmiuhRrlopLHhlXOIXBRz0
9CLck/vo7Rv0k+WsZ0Z6RgFDM+gzDcLzHmMNZFvwpcJJGa7lUYDJZSIJbnUWl8FB
BMAK6VwWYlGPFJJDcYluLS7LfXfEaEz4BwtV1zge48JhokzQC9Pl+Bn9rsZAhTnw
4IlhYyIuRQ+32EHBe99BrxVwp+3/LXXFNOVOOcSRJu+yi4kTUArzo2QR6/s/uhzt
ZdmDgXjC4p1ScUqhSptKG6E6rhc5OkyhnMCWLOLzSZE8X8VjGAxwqSEajVlflKNh
uGe9fTP4FtZN/OrlMwdmVPrqAPHZkCE9+eJr2nmX+UoYwvyxJ4EtIYFRZjfsYTkW
mQrFEf2aTa8ffutonzsGHtvn5tteAWE3J0/ZtOSIK8aoSCFnZA2Zckr5+HeNc5op
DxIuOblEXtXACPFAljHrcDQ7gmlZM+rAG/m9E9veO0UV/EnU6EZmQp8kWCpWEntO
LJqozhLQLsFAMxrL2p9hwErr6IGh88j2Boy089VZViy1YWu0RHxu9yV0fYB5RY6l
Hpq4EcrnJeru8YM4NBZWkDgv20TehG/6NP106bSXc9FtrichTo2QDqoFgMVCi0rn
vtrK3cecMURT2iFqYpogEcJcxIt5HAAbxnrLcX3WgxukN0hjcJpDQFiDUmyJ3YC+
8Xzfbl6vnusdmhPiD2BPA96igN/Xj3QX82ZYc7t7ZZuOJMPMleptzzF53Pk9RzfD
tOUqmYPq9F/NbykLrK5xVwzQ21AYSz+K0XsXaQTTxkqVZ8PmvesUBXq79iQ//5Kh
uKkaidLZhwnJUfzrVM1H+CmWnKlYHA/fiw+1d73ykjG70PZ9FgSug7mieCmpL8TD
xisPwKiHZVeLCs0fOB7z4jCawEGMuAxhX5hdBfkZ+Vkuia68CXB3vOEAxU8BBvHW
WwwTXdhijeTQoqjxl10YkhfI/4QJC3saxy+SZSvoldgWF4ES0ZCJQVxFnLo/7gad
58EY7bAe+RcyOKAAcSM6ZdaASshldiLWzsbXlkazZgfsEwfg3ZhUdT6Itw5Ywnmk
lTRNe4d2oLXwmN48c6Rl63kOtxgosGJlr5nuCElcdPnzDDdnQkxXQUqPomEehnjX
V+fEd3E8GOzADvfaoGmZ2DKvlk54Q8gNIbeezACzEz+Q+vj+QzdCXB1VDXAcxSK1
G2D1SnY1kOgR6XvN3DBzKm7zikA72/McPJsnkTOeKozRW0oQzSNDKWSTxAzYxRrh
Ht/vbrId5YgNtbWw2zaX4cDdPEcOPbh2pJ3/GA0CL+bvzhC6vBmZJ9gZDYt3molr
PPtWjjvGVZqKL+TIOz/wq4qoJ/YvjdU7C+waDjLZoQATgcQwzjrVIADw5bn9Ph8P
sKb1y2XnYwJ6+i2NxsYaKSQyam/sBhiacb2igxialXSWnU4PJO/JONCGPn5UROG9
iGYvIsfUKAv/QAaNJS9nV10UZ03LhI33R0s6H8IoEcaqzw7M2XUyUHqxJBqiPTUc
jhN+KKOyMitfJtN5fjcczjT5dIhIvKE4jheJMF8pKU9pXLfubn1I2fXxxVY7sJaO
aFbZk0RJ/74xMq0ZyegIVWrTD6zoL1ttXtWfXCwFPfIjSPm87NWKErMC+6U6Ni6u
IlUXWe9vFZE6Bfp+XhORc6bHVmcam8ZRnXxD3ofeTG9s1O2ExZfXr2tBsX7DvC9k
1fxNlhGznTOAggEPn05ZRTpIn0yQfdmPA3bmmIf4yEpQc0Y1rGhnu9hcmYO+KeKG
R+/hFxJmCO3Uswe42VBvDAW26zBuXxWQooHAz0ScPorYvK3bf4r3K2rLADMsWE/y
tIEJLQBMIer5LETuDcLnte5y7FvOBodhgc/x3liH+4P+ba0S45aNsDayc1zKprre
YfL2qe6eDeHcB7U4CZtfV4apr/kKfNmpqqxE8Shyz0qPnsg36/8o/Pv3UkrJrEf4
n/RhuSk1vP/XLPjv957+KmY+ccFJAIhJ0FvYrEf5dd7ovTCPCU84uFE8yCmDaF6k
s0jx9ui7Qcli1GYTvvEg9Mvbd9UJf9Mw9ii6kqdxuPOgcNympQ8Uvz/vRjh4pXWA
G6uA1MAnmRN+VFhh0gRh9CaO8nbBHCp7tca3SUtTMaJvdVf75JRvhKaUhQKIkwEQ
hWUn0WJAvrBs5eqgZIjGamooOF5OWIBl+Cfm68CZ5K1KqZxRMYgVoPl7B8fx+kYS
Ch7WQakUxSy40QajEqVWdYDtANkw47+I/GJpHQAqddTz0TeUMJLC7pT4fdHv3GrT
2EkE2QXuBV5RyqwcDUYqZiW5ybEzcLzrbCcLOXKsRtXftbugrjufrMguyruBc2oH
VemTDWZ4A/4qewTCvVGlzkHi2kGgv9sOWHsFrcX+fKt04y2RTNikCyHwsgItnA9I
gW1esZqx9X9ly0/FjlMx/DDHd+9kT+THClWRUYItFDWNPymuyFwfaPSn+0TQ2NF4
kliIkzO73ASY6hLwsaYFbcqaPxhTO8HiYme65I5qcKtHM9pHMgcPyL1Hi2AYZ3N9
Xs1H047WO8WH3Z2oeOaD7b4p5RW4a+alE/5q1pxJriuhqgG3ynwClLMe+0X/weHe
fop1iaStFE9QQGUH/osgog3Iuil2oz5TxxClfXchIlXk9djaWB4pUoMgR9AlbEQK
KaqYDHgkrAze+TLZVtByA9T/LCjMoWYYUXxyu3fSbtNgdbNE7fbu8dy6zvlm5fgu
fuAEqa0lvwu2ol8tPw9H9X657ddojZmYjeDKI6DlTp8C5ZfU+w6ExEfT9bKbrKpQ
+cE/RyO3WGObA9nbLg15bapdGchUEBAsBdTYKIdm4twsj8VKCDI25cjtEClwvfbS
od9w+r5aBCDOXwWYGrRFlceVCRmAZ+A4l1e9y8+gUW7BRTRiXgcXh5Z5qW3nJNyk
PfNYM4giz38Zwed+kaIB8lJf9l0EVG9hP74r6EJUOShhlig2jI3O5zxj4kFjbkJG
rX4Ssu/Oef0VR2u6chxP3QUfBJF+S6/JoVgNzQCqWzCZh3fHc5fvj0c+Qztr1V1K
Su+oHqbzXk4w3djCYcOKwCOurMLkKhpnxcXB/Q1ju1l+z2TQAqCgqFL8O7FUUg04
/fdVqsRRd6yQc4MxiPwLBSZtGSpsrl2UHZ4KC7Rar6ZCn0ygtvB1FF070kNm5rYG
fsO/zFvVxiHx4ysL6gyMRPDlBns4pRU9M4GGnX46CaClhO3U9bMmgvPobn0bfkrK
uhIkOmBl00FxKHI0uWE+56MxaT4iWcKa2PhNTqM7OjT2fdsgIxsfcb6+Fy1Hjk2A
XfLIofhqLwI4LD7K1PM4JwK+QKYxQXakUW5AZ9/0B2IDQW+h6MSbSBn4R5xNgsXQ
2TV76SRvdhgtTl2XlsXf/vMzMxugCxU8HBigS5SgmMlzwHheFk5ArD+NZauzkKz9
sHSZVdDosPbvkMdcAM9TBzFm92gtFrz58i5ujt/A/5MwJvuifJZ9tcgDsMJQVnhL
i80hxUVpajOIQu22U9ICOfQQTG6DokLAIfmzIgcXvRGcEv3c36blYhmLDhIgQOcv
rbom+1QNrfGs/1TY7qkUw0MiRcV2nFL1sw0raLHztYAv9fTrnXwCsfC8klttYgkp
2S/KXwxJWt3A07aYHrd8TaprlxAFj/yCoiJGu/lN/YK0mA1FB/BCa2lkxifNAGIe
nzcjxR2pcEMFC8norwYS70fdLEJHSxfHtTkn0yjAZkoZhtuCaFfS6TBwQMECOqg1
ZFvvc6SzdyFE9jQTqhabdI8iaIYcTZN5wDfkzafjLrSlanSxsA5rnmaA4kcBr9nx
XbS0RMAs3XoEN7EOHNm9hiS36mny0laJGdjWMjNdLcrtdO+B3w3/QOyA+Le4lnaq
qZH5ryNNg7pOyQRMOyHECsibW/t2x9J5pkrmcBfZ7UR6h88dsCz3F+2aWjR2wxmD
89N7olGxyeY/q4v94aydEV1sojrXx3qi7jzNjk9w+Sa1spZnJ7s4S5PU3cle0SXo
oXMTjh/fHDdzzIU6YxzsI4pybHcrLEDPM02OLZ0DC6vNkdc9AksTzc4ErpQmLXKU
+7bRpAJSigcC7boKhLZV3HotBs37YmBRxyVNYDHQIj3AHYLujUXDZfLmO47W0NNJ
hm3R7X1/xONYTXeVf0o38zYYF4FODMqywOnqlWhMGQa4p4P8dIIJfuaOC5r/h9sq
a2ZqbuBMXuHML1Ztd80sXfHyg2VGrzZGWjuom4aw9KDO/0vf16F2ARfDOZYPrEgz
Sm0nkoRlcP4CmxAySPjatFwyTxJINXg1MJABpZdsarMOWlWJoTp2i3rXGEUIn3A7
SEhQa45K1lT6Zsff3H9EUG/I6fWvP3cYDQwH/tyuo59Z3ClTwAoRJNYCeZOb3OJw
ugxqcs//U6jRo2e1TMeDMxzVca6TQNFxU+qqFD0bFnQm9VM3fR5W+hrmRAAwnv4j
aOLm9IgaZdxuCHrax+FAmQ0cCIKEOeUxMaMT9/gtBhR+srjP2c/3Zeb7Aso82VMY
3vowOtUV3XX8z8NRuOUFu0a4FrO/Kc6omK3+P6GxVbqJczxgzYCDB+Swj9pd1HOH
4s0VpJ98Qv0io147r5yxo/IDUFqxnqhxeTeSqDiWwUvCD27WtWS6kBP52KOi29p6
q6pfedjBROJtzxOc4cqMW+cXz/2rJXiPNpviUHLbLPslG+po/eDp1NrjDLYRedfp
8+fBc6oqlbavygZO/9W8RKl9CBRK/rPfZAlxvRbNe+YBZ43xSMA7clNoVBk/2GWC
Usuaa1VxWi5EiTmIwl8M6PFfjKSYbsmFLoG7BYkpso3CT67K6PcNrxUOmMWwrZIn
x2ncNXt+m9JmL/aAf8PJEym/nANn+NFSlu6UyVuHT1uh2TaxWX5l3/SqPq1vEE8H
ksODMWXvEobtqVE6R4/xp72kpdyATgKxlRre4ChS3rVS/jAtdombh7cDpRQafvB+
HmDqeUySadW/OFxRRfecHWFUsHbcoTlE5IxlVhTXv4o+iu38GBHsnD2X8toz1i05
ryLHfaJCNW//zSxQs8I3bYbfHxlFQEu/mfuOWtSD9YokQb0dV4ZPm7/X5tNXN69j
BHNgz4rlwHXdseL0xPCaa/TkU2680yr3IOWQu0Uf8lL1lsCK/NIN4/Im4S9TioKK
KPSJr3lxDAGg8UluwouW9Bp6YjWRuv05m6U8e5ghWlyzgRNpd7AL4S6Vs9Y9qZdV
c884r1Vs1YH0GI3E0FNVZy0exTSRoLDoVLyNNP+iLByBCjoxawa4T5eQlUGROJuC
R5qnWtHKV+s1ZWQsLR30EzazePoEd8CKslWY/CJtU7dr1yKd5D/hYxbOg9+rI1BD
Y+Rt1/Qgtu+Tc0BDNE3QVRS1YLed2lQpztdEWDiC1kCkZbVkxJZJXYU7TC1WIYpb
jBkZ5VjtGACUI+Du1foyrjW8dDp62pUTAvFT9Lor2hkGYyajs9xjut3a5q1PfT6Y
sCiWlCqW2DBOblLAHp51GE70duvusx3K4TxWwK9TGK8MYH2SOPkUyE7PPWoXYDp7
t4sEb9Jhqj//EAWZDEPIa0zdX4H4HtzInNleG/6o4CPRQ890YYDglBzphkiMrY08
nLtwfmZ1hz97/VbQxW+hV3LURHqEDv9NqyLkKg5jqQr7gH6McWADpQMXbG3IHKT7
VPhrN/LbAnd7sBAw6P90CCi/SQMGX11uVAhXLe1zMKxOc1NuU95i1gDKHTw2CgsT
Q7l68ISL0IJ/XWa0Ls5WJrrHLIqQBefmSBIIfG0IsMEQu+0yxcDmjjAy48MfyHWX
md90RzwWjQO4s/wusqiPn+DEEikx0g69yPl/vNCH2s1vg8/bDdMAeHGWCTBUayR+
gFiVHHLt0xL4Kk6tdPs88p6UikVvYC/+u0Qix3bX2AHxwXNv5SX5GnNfzefJSblf
lt+SMlEbP35DyL4b5qQabvlly+Mr7KQtiAJ4Y0RbHNxqRUaj9Lr8RpcYJWvJ1w1E
z4oCBWoLRz1RpHXaWovt5U3j4KVWEWk6p2CvUnkyhuhVNweNMtRafnI3Je1vpx4H
ke/z/TE4o126urgvnJliyr8bPKR5L8hLHHIcrd0sb6Qa3g+clq+xe6NFcj1s8jP8
yNeS8/6fmuqtiha2WT6EZV+Lx/FJpiRO+ABHkgSdBENjYnYdTLHxdLt9Xk2od74G
fhPbZ6M3MZCzDGB1L46xInX0NFG7/rjoy7rV5bWrHUJ5PTZIX8KUn77qR2vPyGWG
c681fyNjxE0gPWpptT5goPYiVEtKlkQFUyfVD8djXdJ/lvle97QRdh2lVGmyWL6l
/z8OBcbyWXyWwAVMSZ9txHzrxj//1tYLH8YrMpojEMSPZwPJx62+rtn5jA1YYaS0
yImnCuEas3kh9/1xvzBBJYrFE9gX+iZbRyGdrCONLQ/XvGxiavFIAlKWSyLqEno9
Js2Q8vX398SzLcJDvyQmfew5PV4nDyvR+7wJHrNUEsX/Y8PqXqi6T/oMSaTsjz+r
ICjevxqvyq3RatIObV7B4KWnX6g74VcBZ2W9kUGvIYRm8jKlr+z55dTCkrJC+/pg
SdPgSKFw/vYnA6SXyWxz5W789EPuabVjVEVCvj/uBU40lYZqdkgRj+SuQolHLbaV
US968OgBclYj4dT8ZVxu7gvzodFoxEo6TdwE0ZoTeTTvaMN9uBjPsiFPWI0nS++n
Vcfv+NA/NVPb1hk8rEuYIztlYwAHDixPBuM9tDlimBBWNJRGhpLe+6NHb6/nqOCQ
3KevH6TJJrU2Mq0v0NE2e+ngLH9F0rqP2oisi4A2WgMvDAsfUcAvValUp0a+SAXT
6lfNB+AY5RxP0G9OEFBIKfmCCJkZwzj/DvGL3funz3zxiTucjr8gMO8a+rXSZGmd
xOxQnazbAc9ZMBb8SuE/Cs7GTBkbSkk9xTFx2WxY5DZNfBCwu49ARJgBbBnxXsUr
0imwuSEnXirl2xtZHvJUOFjE/c5y0zn5xlPeRywScqTMhlEU/RqmVGv1g4HRk6Uk
iwUvum7Sf4CVUMB7S+growN7i4aJ2JaZLFEHWM3gBT9JCGOyVO9wBDssGIAzH/6l
qYRdtfAuVsJjJQTlySotg37usHoEtEYGqQHpKJFurpq8Jq6z6NL2jz0+BgdzBmyh
yHxiwYmleuOLXEPlxTbGJpqAWJuHMDKTbd3BziPVYOpcPkVQNZfOV6pTraC2WA3t
Bf9qulOMc5HBUUYusFsUc8z1oBVdUgz1FMTFp+TalMknBjIRV73LwclKe4541gXt
KW4kNT/dC7pJwySC8h0F8NBYn/AzPQuApjYHHS2WfAvNBKTfickEiJVUIn77EcKz
1aZRaf37nPzfkeKkzBf75If+jIIwW6aNOXOfFygF8lLH22H9MeJH1Vgx2dOw1SmX
/c2J1M8bncMUxKO0CEJABFv4lzyXMQECPaKlGrTqWP56U7zmkRVoF134eSxQOwlK
MTCPEPLvjAqi3ZpMbVLXJHCepA0t5wCuSZO2TVN/rmSjWoLreZvZbzdAzfFF3sdz
TeCFco7o0RP+cD0CKSNgwzihZxsNm2UdXeECb8trYCDTcUdPogLYJKaDm6l9Tpc3
HvBi4yIlIRkNZeynOKwddRCK2Ugz78GI6RL1YBeAc216j4THNKizOslnJZTTET/e
FAM8cJZ/T81g7LxgmspW5G/bkYXZjzTB1FsLYBnnR1WBl7ktXKS27W77rVzdi5tV
BwuyAfzUhByK3gGl8Ia5GIasyLq8fJ/yOQzZHj86T6aodqtLCRrZ+wHgFrDuW267
W/oYfG8Z9ENudZfks+YSz90bjcIuR7tI/ip0ydvw/cYa7XfkurgVzC67aVXODj/H
4BhIleGA5A3tSbSHXLv1lutWR0xmJoBHRJFsNhpYlquEEGqDESTPixLF6D5MBv5f
o4VvBgV4SlZTiPFzLIhHutdzbhcqSBESUft8x3jUzorWWQCmCN8BoeWrkvkCH9/Y
zfKBjVNKMp7IPYsciRMMMlhbQXhkosyN5HlzrBUQ5+GUhrl9ipNnLNlVIQKeonzC
7QFujx58xd/pni6UCICqfabYSphFegvaiMA+EekrYcy9ULRSB5PLQ+q18kNQnH3A
xivsdmVvLFFlLkLQqJoyRVD2Tm2f16+BWAVAz/We8918IMKO+j6VHEFatdzSrw5d
q0G9+cmaz8/8TevBEmsTaE7l0H3TzTmn8noocjDXEGZIVsu+Tm+FaScwT4IztbOs
iRybZsvO9GvgrVDXYykcVgppVkcNZcRLBgSe+FzpYcBCz8jcshW8CDE0rrqeuXgS
1wvkG8zn7PAL8/hTxMlEF3VRaTZChmQz3DMtOnMc/LVqOw1l+werSFCZODe2uVVD
+GSZJnfPZDowVKG5qP+4aA8hJhQ3PBgMAR6VwLoUQyObPbN+uUC3Kw7cyw6Y69Mz
7ULKQfLhzgqaTv8sX3ZZxHOLuDX6YJRME3Nij2Dvw8UQ30qs4BuFRJWYif5HNXul
+coY5teNJ7Lpt8Vl3dH0Z6MKUYejo7Hgugz1Q0plO6Lf6JBbdxeoAeSN1tpA7h5B
WpF0lmliQvk8VqP/fWw4FMCh+SepSR4K/wsqSMJyuXkPMoDkwYzYF8TrYU0xrDnt
fserKSmxRM3ocnaMdXiDXFQlpOthz1D+866gQRSsCp90e3Hk0s+k0lD2LiIIWmII
bkfWtINTrXZfX2ZGBertcrGwpGEJEDDvpQqaoiP5ILc72bUicLXnTWFdIk6Rs/N4
bd9XNJz8gKTnVEAyXuGE5QxeYqYcGvfkF09mo0CB7ImRG59RjvWERr9zVSAoa/13
O+QOJseD5Hdx1UUPNJ4V2exFvP4dY3rzsFIHVZR6QgxnB1MQpSVqLFUG0iAjkXc0
ylUEuB03soLNezmnIhso2f1aq3/RlUuIYX0oL62lCaTUTm8xLDOfQQsDv4DgBBzy
aZVn2UuAwBdkOGj3tU+lG6OhOHXDMye4u6pFFfqCnK5M9G6xxqSx1yjHZCotzPjn
vXgMJ4f6jv7KK6ptTYu+hlQSaTT9psYdbqHEr1vDFpsMFKXh8xfwZLPU278eSB8q
rRhIqwJI8ome94UTzJZPViU/uk8z6IuyUF/bPGGUSYUzwaLQqFoI60qVIffr8qVa
/GwX4t+EPSa69j/luIQSvy7dbMtwGpaCtAI8hM1L3JclPQB8pp9hyLR4X6TZTMJv
kejyQC0aP9PGiXJ2zBfXy013WRvK9zFleDkYkaoXjozZrZgeEjzPWPGsBcH5byzs
5GolnG59YQmUfP9pV9GQl3SIQtCvfnzyKIN0aNa2osIQ8P92CFm0/fzNCLeVKMmc
UfFvvI1I8o/sfSC7/sTYC8tjljX8AVYXSvruQ7HTvnmlLiizS7Gq07ZcuVLXKHPv
ds4Pa3imKhV8yoecDSaYDWzQsOeOppIcmYQnoaAjkSmlL3iizmwYweiCJIrvSQFX
JS50NjsxDVfD+9D7511BCRw0J/lkjNAHVIxBouqd2Bh3MlS3UYzqzZDNsyJDcPlx
2vIxFaWI0Gyu7H/gFsCKsd2ffcipXzJvn6c60aXUveL8k5+kAQz6v+rJmfkrRrI+
dhGyeQOfCPcGaaz6x29XL9weTIBmwv1P36EeQDI68NaJaR68CvCNVmWpWx63B9gk
I4N0C9Pofe5Y9moKtWHVcQNt+Boc3x52do6Lf7G/+Cp1s3GpyTEOscsWS55PS5O3
H9vA7uvgxVfOm+qKgea5XgMG6R+SeEh5GmBk/4tqfDkA7GOeJf8hJZ9Pk5ciB/L4
uSIzidJcs7hH+hZw0rrZdrh0DQ/Ta86CKDySSf2b5dclJWJb2A0yDWsw8sPsX6Jo
O+KQU1+NycVMqBXMZQnDW3TkrU9XfDPgm08z49Np+d/zPj6wnMzkW6NEz1ZVJ2ri
CJaRwkcV7ckaTunZrcjdknJLj5NbhlXARDS1e8FfNmMvJKQCAokDwgSDiSjmIiNg
l8D+9Un6pWnT9eQasAmeC7VkVgC2BInHN7O7BOpgeB/6IWJ1WkW0lrLbgWzIPlwj
mifeNk9I0I7tJS88wdRoFY6pTF9kzCM4m7WVZKH9sPKvReuIGF4uzpKsj3+PY666
UcmcR68C6+JMdXxZAZ9pMkdtOBD70yW5C3GTrfMOK7bxOjSlPueOWje+TB9Wydod
/3Dw6HId1mnJNO1mulO57oOkQxpMei4sXAC+hs+RaXihH23lyfYkr5anempztrEM
l8WwcUKBItPq3gRJV27BObaY+vpQ30kuH/GHszOTQWqrM8UlxC7uM1RdzeJojT1U
UrvPGJUnZLzg1tbyh+gyc6/G4A4LBl+xlboe7RLpS646Gx2UVDSbw6Xf6IVPNtFQ
zvMJuT5PPE09jeWbVD0S1kATJvA4nBO0iJJTi+Y5YbfMbsBLEDP7eXR6I+3uFjaN
Rv3KT3Rw/Sq42Acf6Gv7qn9vDhaleu4jaJ83s75VIKbZehZ0W/ug81YM30vqnrWq
c02Y9QpV7GXviFDYhUuyU1EwMWf8fw3N3zAnDOJ6hvCD1YQCaPbIuxvVea7HAR75
T9aQd9sjA9GdESnb6riuC2d1Yf6g3+6Tx41OgpAf0XHynGmbtCQCu098AupS1+RG
uD74o7paCs/OMj4qjH3VI5uHEQXg42BFUbHBoyP0Hhz12wpX3vWKXU9kzmVyugRs
iYPploxvyEJ9VPsgl/K4GjCgu2R4Ddz03Q9FxpzHknEKNtPBnR1CpjNBdPttiGqu
QodRvB6GUjglshxh2vPki6nW+HtQRGrHRwcEg6uw2InvhTZYi/L5GuQkAUqVKH5a
xzYsJhwCLWIQtYMj8k27tErODeLoDwZXj2sUh9hgs++wxZ+FJA0aGN7Jx2+2aQNZ
WKCgsycd8pHvsxEE9rfg9G/ogen5XeaHyW3iSinjwMDCYBMtNLGcC2adgJRiYNld
GlwSbqw3bDY1NoXZNqyKLEz+ufLZYKRGJNO8leSUcn5so+t9u/6OCc64aagngW1J
Jwzhxhd4BpmrOxbI7U09zds/xobMMEjLd+w7/LO2UmByR8sYFN/u2EGmJ6JlhucC
cz2q71VrtBjLMfccGe82BBAaEgW+n7UPAyverJADqfohnpCHGcbSXPLz0Rg7jdh4
gT2o9vFULJlV0jeVJ6KWWt+sgB6Fm41KxB0ALGBsbibFpPCbu2UmBHfdXGhhVeVq
j563XUTo1TZqYiA/gWhCcxosOT//8AQZlVUzC4u66mP4PY8DekhBCu3kZ6xbazUU
sKHSetoRMWD+/FcLYYvD2ta9XYDXT1o1e3BDDWVumLfNKCGdm3Gh6tjaZO6xD+1C
IVdskCIlHhPXpV008EkLVB174OiM0TDgiXeClslsIqOnfmzdLTDTYUCSYTnmeSBF
f+s53Xsfeh0zzXd9DTw4MDh868mjktkVY1BaaNs18+QjkGeBqH+Eq7pBWSH7czGh
jgJKLHN0OX4P6z/FIoaZb5JoIOn/55QnLtd/AEevixuw3OkJZ2vzEyZJZSatkw/p
TAWek8Ooca+0Wnb3I9AoDIHIiGUdDnkcN3i8GeyjbErbCDpQaXdxrvRO1KRd2xOM
c//s5ZhAdlqC7je9+p00eg+Z0q6yFI7ZRYY4rHE/AFqSJR9K6eVhRMct4v/QjECp
CfLAKnb4Gnkko36JA0TCpHY6d2XyfeT48CJv6jSsYYMjOziH7nk4gFMnftcwErVS
bTdnhFfP5rb+LjV52ULxRZZyRKmd6mXzX4wkx5bhpm0f7CBYVOa0acZdj3IymAFC
GWL7sIY77XUiW95CfNUeBxYn+f8k1ZjSZXyvvQnpqa3RDDEds49vqZZlHVHnSkYK
X1kudCtU3MH2NXmUb/YsVnQOQjYc/jShxMyUchfr5v8ZahC6dgacoykG1iQjST1o
ZV+NE5GW7irNWcsvpitootc6jnCud2N6MJ+UOajrCEJImmy/2NjQLR/HBjv0NfwG
L/CjvzXP5HNJIZp9QgH3sM1YS85DgptYaJVYjOr+skV8DWSCAWOKoAUgbikBk08w
ugoxXq8UgENAymvBXDXn3KXSFc4twrogAVg7lajOg+DL2Bxm7UDTYcvSeGcsTiZI
aKtO6le+IEPb8ier2cdc6FgTM+GHu27UN93+y7Z7ybpl3iU5+aaf8KEwoHLf1JQ/
TK1UPkSxQmFA29L74/2igO5cqZbawckkO+SUbKRxV3m7vFgxsZx5XGhz5Y+2m14n
P0IpEZMfALRWJuvITotU0DjnyoZ8MyGeMsZVpYLhCF2tar8CIF7/n2MAAMUWoRpv
fdm8mRMrmMuRbuDOmA+pX97cxUgUury8oFS+d7UnDPrkwwGvIfH4vAaqvE+TJXVz
jfyusYjUnLmzbNJfDVsYVsmDJ69Yz3H4fm4NA+N+rhXJ4FElbcoj9iMuYGQSOv5u
dkrx8mX8NQwkH/FMIL2LYI+W38G15wLeX5kzkpsEIuNNQ3Tepw0HECT/6ulstEyE
wl9Jzi3oBJdhUoHQiZAvW5vGBBpi3TEiE7ZYnOaJ2GXdUCjEI032LdcJlahFfEUD
2Yy5E2isdBDzAmUG5oTV0e31Fa06CUNvawwAXS0jqPth0Aomlgv474K2MImfAMgo
qIkYXPWkpYYP4VyhWDAMNvzZWNPhTWGW9JTRQMFwLLYXTFEXocZa8bQJ/QMyGesP
imr9tjxVz8e+byyp+ZO+aiBW+/Xvz/p/r2hoTz17ra15HWRapef+2NKxPs5h5LBx
DBU8TLKh8OUGAP5iqUj85mEHDFNAYevj0rg2KMyRupfxW6tY7f1Mv/cW9P2UIy9o
/kAI8MqdX+LwJHE3jQcycq+cDEvUoUNFHSamrObrSLTvLb3XxdtOKI6XLc84Msx8
lWXn/okrDTenrxtBE826hQUAV0B1iW2x3sKtDG6gRfiQ8lcrzBuNqJC8epM3FfiY
uh60mR92Hanz6rkFVYUfZZgSx74oooUYC7KQqOCsomev3nhZf4bmhcUT9IBfXqiL
oBfkSeDs4Um2mM83lStl9AJS6227Fm7uKjaRuD2rY3NrYAHSBEwNuyQMQEe9A9fG
r85IDCnOLhnbcUCsKDEeRjMxjCQZf4kdm8Mj7/b42iaQ4oduy2RcQaVJ1rsYw5b4
dv9cnzMUMeC9+49z+647AWAj7LT8pTOFFlCDiHfLbIxQ1OtxtLjyor2AAY7Y/znG
IB0tj7HIWL97CifweB5qhuQBV6VG6U3TX22AN6vHFOXtTT8UOlUXgyrQJANC4HVl
aL0a4Xf5PfvmWGS9rAfF2AMiIMKzN7aKd4I4p8jTkqkOox47x1HONEyZZYYo5ezI
izSSOs0YheNsrpYid53+stsZsgIoA8FLYpcwlqs3xnsR4ZNMvbrQzLwWoP9WPeo5
RLzVACijSl6RsRvjkFarYn2jJp3LlspKINDWV+ntPPUXwuEjO6zFkJjPXWsztZOz
3ESV/ix6MTPsH+9B17mVDC1XBfR9+zx2NHrjCeTzTYstN4kmkrwl5z0xVSS0tQDe
LFTS8OFd2zJL+SyHCEktTilMZJoffnelsgXkgW1OzQJ/MWhaQN/ZQlb0yHKW0e+r
DDGUWqfMxufbEXvrYfxn0heh1z2XaW7CVnZsEKTSt0OrtUiiOHnv2bWXEBegaamq
o8fYVQ56L3wcO0UoMyztS6OXyaDdmrmNiB/DdWP9uo6EErtNme14W0widy8zII9L
L0OXqQSzCKEHMi9Vh4/pSscgg3Or5qIE5iETEefkC/sj2SjkEtMqHg2/fa4/B9P3
kbuBFLQ8NLz3z8wy6uCHOgGIdI1gWpVuAnMECbRDFakv8hddl645zCduHRLO/ROA
TZ3+nggW+Toy0MmXqcbH7gpZ6Af2hDLTK0DqB8j61qITYOy0sincbqagEyhYQHA2
AKiLxE80dhIL8JlDT1mpA/fkWY2qnigfb52mIc2ciKBrrlg/BtLWJWVh9aWQjk8z
ZTiF2SAHQqBwVhGl0YUckPe4aHAmhIitXNB13LSGxr5Ct+xzYLlRSNMZ4Hb80p8Q
Mq0pqLTaWmCXZoSL5Qs96kvcvOL0NN7WRUGUpFofqtxu0iLAZs4emt9wPbaOuZ55
ShjWCJ3/z/0t9dk57t+t6Vvlpio4aJenncblQTVjFtdkmWomjT7QuIFprux8gCOJ
Ag/A4imKdGb/aRu1tXtExP/ObzQ2HOWIh9pHSGiNY9jGDWxof0sZFBjb7NJ1XuvV
frcIBZh89sMp+t9kOwx+vlfmX8CuJ2XS3Ju8rcARfMifRTqjAHanMEDZue67FYYu
tOcl+nVb20YcQKPPaxSd7LhgJwD9f7FkllRdGQ6ixgJKyFtInymVMx2TlZXgwR3I
3JgH0+TVRAsrp1TEZ7Xzus2O0Lt+1ZWzqMU7E4F9v6qYYhTe8p+QOv4hxSO/ndRP
GFHXeSstaKNKxM58V/xq8l4EMO95RHPZCm9DhuR7hm+zhARHvZZWJiHoPcW5cxNk
2CoNKPzIPh+2NCV+a/KYf9vigy36mTcgcWQY9jnYz4M4T9XC9bZPyR5tBQDzTJl9
F/lVATWILF8b3YzzQ8XerBELWJ9kBLGQuEbJZ4A/T1pZLgOtGornbRdB4OsJ/+sb
O9S0ckgH8s2wMm07lV1WAKvMbsbOrw8IBHPGHFNaXD0UdzN4IaviCEnvBiMFFiRy
qz3ZXLkFu4wHNrDTU269rofvKF6ns2gWaYpqY41LDS8KuSFUVa1FEjW9zTXEJSG9
kUvpoKcDQZaj0F5DyFnnr1oVHlUSWpNPf71Fl2o/50cN6iCEoCbMW79BZKPwh4Q1
8EGvI5prqKObBw0ZRC8SzDBoIlxO9jo0TMG3+bwyFbQh8kCThOOAvvIaRQC7iYR5
ahuLCnYv0xqM62kdE9sWzKBWoWrOr2EqRss8Op+GA6SbkUorQRV0s4e0HkuO7Tlo
BYJgADc81Sg8HGg6JTZnV4bzuX6xRR2TxolPE4EcH5boTdE8G8Is9yekcxs+Glzx
fC+UgU26UH+ELfb1pSkwazgwsm/kf8s3/VRUbScFwctr88YlbfCT+BdpxbyaKd/S
IyokQ7Dm9ZkOkjgA4+ztPzmoFCVSZwWtwd0Cwcl4t3D+Vl0k84BuGHTh5D5uwCUd
2jNK116v2857BbgjV9M0hsz34Vqj49qQRk5kWBuvsT+TAo1uG/AaaB+hRQR8B74H
3/Jt35q3a5t3tKtmxO4PsTbFHq2jpqUCgPvqGUHbWL7x+yCMJY4o7G+p3vd70xLV
I4GLTgBA5dXJ3iSpoD0tMFhr9ye+IpJcFcmUfEinl6ygW/NOHf+KfYKue32OM80G
MgK9pGeyOFIt1k8fu4fUxmID3/sd8PXoe7TH0YgS/Gv81lIp5YQqmB/mAD/CWs0O
h4PVCbXZIlTjnDRVf6H3/QOUsHB6MHT0BZGzu+h0Mc3H1n1jAscNEeJOX+VgHF3w
oLRc2cN51/fo6lQb+n0q8NY3fPT/RTqGYfCx+gr4tavgnLcvf+BNxDYeFKrbcgZo
MHt62gSIyofgVCQ38jcZzzch/Owbpc11m7wYa3nCabkqkEBP339kbGnq/vdEO9jx
cdDjqmFnsfdoK75gsZ76stHNenD50RXiuFdne+mJz6p6Nbirz7+EWAjc4VENN+O/
wJl8PXkEtLOsYgXXbTkwNfKlUTVV/BrzofbclDkEBSa5dDaG/6XhyB9ynSfvzv30
5x13txTTxco8vDkLjcpbDoh8qCQi6uUCIoXAZwzeReU4C4mc45zLFbWBJctjwwH+
MDrtc91SbETkvBD2KPy6okRLU5htH0IKQ+W19WNrfgcDZ2BCLODlJcqLYwHZ+LP4
+wlU38KcW60XevHQLlspQOvjHiasv8CEOLddNewLMeLzoui9a+suUT6XRviheRin
+HDcNJN6IkafT+NgIoJPxO5x4F8MWG28tDsEAZDmV/3CObw3oZMCI5gPuJJP378/
pW6G+NK8xJUYpOIjuawNoJzaSk2EpF8lNNHRlpoaRFS2YiLwenM2YecUCVmi94Lm
iLtQFnv5ZiRzpot9wvnHgkLNpD7ShEeqa4720Jx2lRQFeZf3u9ePAQylYAb2x57u
kFlKSzdVj42Rnw1NooPUBO4T7r8ZJM+LBJwZXSIRZT84Ka9i9dE/qonXdninDx55
XEkTCaVIefKXuJnd513G3p1FH5wBvdbqpVyX0YfG2JbJveryqrm+spGpGDIDe522
fcL7L1MELLheyy8OkJYNCSiQuBYXNCmps+CnK5Fg/8nAnQgRtSmTp0TGNcHeSXvu
nrzjyFt0P6X9KFuiRVPyoAAapnh+XRP//MrYo8SW+1HJfbDuzWUQjsck2mVoq91b
iTR3fQGFdReSEFG9IWqZIYBHn4SDee5wj1JYc2AhgxkDqBGxKGeXjQkQUkVOPjHe
RHh9rblsY48kHZSYR/haeyrCIWNUfF8luJq09KlAMsk4R0cZv5BiSGO8KllL0jhe
G13xs+PpyJaHBHZxv8yfmqRoCRYx+WRxQTE+g+d2lv/8RL3a50FhLwfzcAeVVXDa
rIChkYiTfJrQ2uZX8RQyar2gZ1lqHb4ZKXCnxw4tq+xi5w25O8dGTj3dc53/9pgW
69TRselycpm9J001wAMcMCzp7Eho9f6qTAUdxT9Rw75fMw3a/gKYCb8dIrP9MFJh
8B1kDurcRt6T1dTFcdH3gBeLbtlKulIfVojpT8qY5cLT2SebR7v6SUGtlL+7Xzln
ixjU+ZERonR8tpYNfrltKkIh9poTeMgEDTiTIoeVirpA/QATA6ZofsHvEjQFR8Kx
9hBwGtSl0QzGMXWb0uruyay/qodEIZ4TmS8Fn44GA7rzIUewqh9p6nJyUWsZxYh2
xeXcMN/qizdAAYEf2VxVvR7rKPKUQRy+zXPydRQZJrtcA2mRk9EqRo/4mdm3xg8w
BUKhPVI7zq085z5Vn0Sh9PnonIkvEhzRM9VYJQxfuO8OXU0QNvyhTa5Cxax2/gRr
2QcP8+0azr8395NN157salYM+nKi5Kv8no4SBMScUSLCDF/1kAWRAXlGTtw0iORb
UvjxeIyx6PtWvXuzgdxlfKObx79W9YiXkqqC9dzoTAuYsaLGRpVDLsvyiOqM9jZT
DyRhh73Os25ZyvECbxT3SDsk8InKTwZZLyoKdEcNsUa9vI7zyR554GJajaWbxo3Q
Cwp+WpEjjX6sZsB3MG+OTJ8q+AvtrR83lfPjNc+WSyaU2OAItVo4FTDf/HP7ihsS
cI5M9HccWb3vNNZ0kMua+dQlso/fYawJTzI27VuFV+K3wAQNSSxDFeo98QHRNNja
YFo8JojtxJp7tQhgwEfo9CaLkxN59+zT3NTymZC95Pan/W/Kj96nkHCzwJ5qvX8p
vs5gFoG+u/NVpgws+dYAG+Rrne3ss9cwiEAhmSM55zARCeW5XSsqKJ95VH+2LGcc
O6S0dCNJoE5xXwkz849uHC4AeE5uRQ4rAktBQPhOMKKV8KTyRgTAXhe15+ISc0yV
cv4rGRW8qynHqy4ALGW+IPzt4J4RPjivC+J062TmqQ/AUcSPIMEbKguG43piwsH0
fFRHlHRFS6rUBoiABsc5vxL2gNIDOlf7ULImrHu+NJb5R9w00vX0p2X8DCL9eRuR
BndCB6t8SDf75ubZSZXeV2rpf6pacFGa56wkzqw4WWIRyUZyBHqvyaOIf804hYzr
A/ZPF7FkUXMJuPrW9W02G9QrkpevJ2dsra9HJMgRzos6s+DEkicFq/+9RNUKE12u
MYq84v3EkQvgFh4rNZyzfCZsMHFCnCsLUc54lB7rPNKFj1mhrWnJGFarSLsvCNWD
gzI5IBnMJFeJU5yuf56KHzenLwcHBvlH5h29oAIJHRsWrZ6Buu83AbzGk5J+zmC6
FA+zHGv0+zgX/Q9ILtepSJeatbKh58U0br9vQKvjtzO/+ja3pQzb39v1I0YHzsph
46rvkSWfL8iZhoDdL2wG9kgyHCneTEc/8aedC9nNvRgOXCZCUmGEPjfgX2BHNAKq
reNFS3xVkU1zORr46WpUhrjK8xui6GSZTwf9c3ENdNTDEUhhTqtttyhThkupYm9l
RXSG73Lp6NxUkQ1PX1+CLaDdHSZz2Jb4f2p0JZ41Nw2WONIraBbc54VrCcsBL0HA
d1iYeCEhzgTHreCytbVcRGvOnFLAcJ3wTV7wEwpz/50KrH0RrID0WOTXbaZqdDsG
df3YKam6zABrVYB4JeMaReJG/mqbERddNUnvphQ5EViRepOxCP7bpHFoPovxn2ij
CQtIwoz2wcY83T/OOKxG+hx5Qo59JtemfaGFiQo44E0BVHbz1Fmk9m6x/8LyiHlT
U0DxCYXLnJ6h+WWCmyrRlh0a3o5AuqIvpzaRyz6MGe0yzyphgzjhuV6HfUxf1+7x
xBPLglCTY0Z4Pb7SYB5sDQajG4urx7OXfZro37k2E7sNYZQUpjOSZqStlGCMapaf
ilmHgpE8BsGKN8fMRnkKV5guN6uymL6vq7l9QaPG0ZwLCHUiFpttuUcdlSW8ZtxW
Mbqc0ONOUPpzireu5HeX7RrNGquz9OoK3FwPLPuabYXahqanY+YZmM40+7zq5NlZ
ZMj9XLa8/bb0Dn6If8uI0/7oi+X7SixJ+VFLHiZ4l2xSvasEHiWSsj9V0nJ8I3gT
5sSl4Iyye/w2zZ7/7C33j2XOjZn83/bINV+ivrqeOLnSjuKDSC3ycNbrYjaYXIkH
Njb4uz55jNEntNKam+7mLty/75P8dJOqDE6C0MSS751E3NFLk5yDduUv8YCzWdmZ
OES4YXChDMFlimnS7A4u1FelB62HWLB6npIgpwJaEH65nHvwWdT6puhF/Px0Tf8v
YFGu6zMzPRZs3aHz5RJnutAfQ2eoB9LD1mO8af8lRy3xJdyfVWQgCDbcuaibtIFH
DQeOx229i1k3jJC4z5HLwshBqL5ECQgjMfU9iR7eygTWq2GVaTTFnC9LaNvqY8in
EmqLU7X1V+7tlkSu+W/jKuIkXDNgu6ynJNWvxIw4v5FRrQ8pgOVP/e48CCCSBTr0
XVbmxtnC7+04f0WzCgDZ0LFEgJ/swvA3+IKPLQ2uDMoTVTVDI++26dILmjm8n5YM
iJVGHRRYAHtAesuSslVt4N+pMCyO9MFrOeXaovofiszWdcE2xfj2DxX/FYmL4xJf
z3R5lNQunrrNfgEtwv5r96HE04QHyfIMxP4N3/Pa8FidNbbgs63d5UBsp8GPA4Oq
2x90OjpsOL1vXiiC+/S9eTYh7QhQmC7zEIwmsVoTDU5I5oqqE3Jk0SNy1UYyoLaS
kuKuQtohN6D95uMObAvhR9zOZw0xmPfzGso2rXW2D7+/AsbxH+q9qoqhEehtspOq
cHY7/feHvrIKyCndI+rmk0mRG8S6tZJo5sipRDK/ON6KSH75qPZ2ZAhf0DHUQfPr
480glBKZ7HKH6/aJ5ebArXNxa0yQ+muKTlHDdzKyZOz4fienFxMZq955OpZ/BdmM
Bz8eOfVpR5tFPi0PPujLK2bh/drN7Jwm1+3WqGYFIrlL2KqSEBLzxosfHATtVCcr
gxmDfMgiVUfrlThXuUg5cfNdELU23/+yPnpB03ikWp/W22aECTdzQ8Cj1VqUdN2r
ppHvH0mV88DOxlBdo3GRlzlyaAQpS7Stp9ZW2hQuubqEwXN9ePDcDAUNOq+nJo3Q
167IP0TQipEWZanz44xeIJ0LXwcRTzkilv2iLZBHvmo8/+9GpwvxJSp1SubBmS73
rEsq3RRHOc7PvhtXKoeG0KdjK+1znkbqTQZSk0l0g1CxfI6X2zLcYZ84a0A23COc
T8A5lenftqugbuKM1usf0W6BpR3Em5C3ZrSNiLlqwc74GfJE6WNky+1cr1kOnkhH
YzOr2o9MDwL7Az5tbkyj2JzNmBX+1Lmc9sQ+6lH43vTZotgxOHnr63hksH4+cSbD
JAQlrTbDhewrxieURXbNbD0WY2/vyO8XcghdbmBENp2Rblx0hEmCc/tMio7RA3aC
JTkvLPXYTWfSCI9veN3ToWgD65bhY4fYMf66DvB84VW80yPG0sC1W5BnUYPgDxS2
I2VjSaW65H2kSZY70dV3y1uLnyvVC7GEZH3le2dWXZ81q45HIFLemWGtbp/FBnOd
9xi/1qZEfIqA4bPx/vfgnTMQ5V0WF7mStNcn6qat4smauMjKWMKWfp5uSPhczNeb
6QuH6v9JKuHsB7Pxf3euyPdNt0ToFqyTZbALfBd5kjNIZxeLh5uARPiogLOwEEJW
Ry29BNIsBXPJCps25NPRW4GVYpubNjh6M9GKAduPFAPPvTwrkGwTz9mQ8MBtXd+t
7P4KMMbZlmuPWVkNcQLXnAL1Uf0mAoOeW4Ty7O+uN5/HevaXhP/ZPIsyK66HCXl8
x2hWhqZ5/MmOAfrQz3Ym6BrIoATJIrWbRNXMAYgpPBjBIr6M3IitUxcvUplOx1+a
v+KivOkVYp1PpOi+YMYHz+K2znavad55WEuVsjeB+JgaeCjTbFCf/HinQ9rzDGRj
UUxJ0N3sloroupk1YruOSh4sfjOuxN8dGzp5nSonryQokug+/3TYDb676wf7E5oW
l+gESkIkDuCm3dxcw+PJSDozcP5C5LfjhQvzEzxOtySa59a2ZalIgj10j6rn9bHD
YOH59MSkEWPbG/jHpe2koYB6zaIp99vObFKm+lcYsqbIVQm9GGNJvu55UnQOOdz0
RSSahoQwjur/wRs1muyHazsm58ykFG8N/5e9iN2zVo47gZpuzRRxQ3Eg4pUNwEDJ
cIX/jihvZCDN3kwqqp5IBlnzBgA1/MzFP0Pwt+Ia8R/OttkZ62O3v0axbrv0mOoK
ROd/DOsQZwh+/wrklTiqBCUu6nkX81Ox9Ct9ssCj4Tv9MP6xVrpOuAF6BSZxMrsZ
n8eK4mGmWFVT36BZB+gG9u2ypD2jrzU8s8f+0oUEvtzGOMovEFBBO9TCgFAjT+zS
kthNdpo2LF7gK+0DecDaU+R1nYN2gyOhUjxYpZQuBhjjckB8JhfN5oWLYdtttltK
bvjsmf8ppuEKD/8La/18skrUddg3KLmZfCU6UnQKzHIBr5JL09oZE7UbUd2nuhHn
EOZhStQgR5BZ0f2Ffn2DOJhC80ySB6i7luwfYRbMjfH9hdjjxOjKlcGj/KyW//Oq
WVrFGE2j7zProkDrUENI0skoD3sPcAoAQLTR1Yt+WwPcYjsn9BCdGxYOizbVu2TW
4gR08+S+9jC1JMQiW3ZHJ5YAQ1fz24kzeIrDpc6r+IorF998+BoGDP/am1SWXPME
gISbtATbrW72bv4jyq+JLgTZhLwYzwRWtO+2ykZ1SzUAwGo6WTiYvEFwNfs9RSif
LhghWxkP33Ivujw3VZ4dFbexOimqRQyxaEULszX5Xxx+tFikvpSWVT21lTu+TmSL
WwBwfaxSspvg7fJXyasCAQV9lKz8S6FMpRingvts/Nu3lcuYGW4G3ymTdjmN2ryc
IniuO9T2K3QqHYyR0YuqxSATob6qvSiToYFkVkrkBGqZ/jGusFb41K6DZVHUfSzS
Bhheteq7XSFUUxtuI9iVJyuh7MZ4flYwel+qXRUq0LTTj55eaSUposp0uKNPZ1MN
Lby8NrZhSXk6yDPW3vBJdLRDhLiuPyddkZW9uZLR83Q/+8O5rAfH4zANmYbYUAIU
js8DKOoBqbgxy2ZVAGHlb+oG8MEfNzK4RRHu4QNgGLSDwjZ0g1nufuJrOEaYNjI+
VB7mCp5BzKx0gRPDish0+RndbmcvZaoXBkZMM9tA8+cT8RspTksQa4/3+Dgjg0gV
kvK5l1PCb5nICP4+fWI2kmsjwrLA195K/QREg15CpILZ2aANJZD0WCwBrxiHTTY/
PoGRL2DSLG/hmyFotyXXfoKTme8pGcDxdGjPmbHPN6ytfHaEaIaz9HAzQa5zCT2S
l66/5glOIL5zEeBnW0haIAq3FCHuBkuW7Dr9s4G8r+QbDZ/Whh9ZDIiKtDNPWnk1
YjYyMqV3ftCgIfy2d51PNAMW+oJvYDkKNmgESjQ+ToJG/1DEg2MGMWygqQ5q2gK2
O6ASDb5Jj3QeJwBiVPzJo8lYhaRu7lTJR9lw9pkFHjIIVRe5s2Zqk5/MaN328l4i
w6XYx39wHWSfPqfDpYrjYPz4GG5IN3Y+2P8ObHiRILozwsGopHOMvNKu++IaIHjX
gGCQl+EyCU8tYHowN2rQlQIALjkDgo1MV++wiAR87STs5hxm2kYzaO5cTq97l8vd
jEaiePMLp3zyBOmYFS77qwbQK8pIHDpnn5gk2tDzBVFt39adMsSpXiSguJwd92RW
ox5xN5SXV8CZT2K4OlEr1oxG6lsmoVd16vc0O0cj6QNX9HDYVYBxjKzx7IIyUFQn
RYpxszpwzI2WfnNJJZZeF6BSvPVLFu10iQtUzQAWEKan8KpH+67jEu71QUYJPDpX
M4JOWTne/H5nZqjMecmxPx24VoxKFrMEnI29b2Opat1ccof7xya3UYvTfIu0TFaP
C+VtmUR+3xWgpngEtni1CK1gubJ/juIh5X4A2QRyWgWRznh3i3zTSnpLl11oKlSb
XmnWPofLt7npjtZuas736ZI9esH2yB9WoDLN2rtjs3m11QHY6ixYxwUgArENBDXe
4Hgg0tM7C3zYD3+XGIEX0s7Xhh07Y56PHPkM5n+NZlSszTESDHNI6fdjV1xX0MeX
9lZt3lvzZLa8yeYHrPmb4Cm71Mh0wyqySgYXc5OaJBP/YdXSl5AqqhlyKoDc2msX
cU6MC5brSMKOpg32aN8M+HGHJ1hlYO97RMxVOfraiWvUUP5Keq990NVnCpS3zmwp
fzs8h9YuYYm84vO/4JKxO7QMVkEpnxCv9XTbwIVOChU6PEa/VXkfsz55sODR8Drq
V1ozJYlnv+injljHELSbTbh9qJSimlNuGoDZUqNjF5Df5TaAXLiHTM3777NYTGM4
xcbJ4Q3YrhCnwME4vOC7CUkxVKBiUxbhyhbaqW5ddtNVVTxW1y86mbJ4Spanx719
gY9HrIh6/GAD3aMrCvX+oV4Cve8jYcnWBzVDAzAPP6zmElb3PDHXc8iCsMxerKia
BzIJnUXeEqyHmcrWOOrixlExAgOz2RPe5e51QxM6y8SqEde0VMZMkM9rhN9/kYHY
1OydKAVRB7nOnjnw6SyaW/7BYhS1cYbeGoRlc5nM8s+izfnhFj4ylqGmNX34YRPl
v1MOaojPn1b0id3Z3RLRTACwicfiQqnJ0DSzt+GWkV2s8bx9yHlnyNbTBbMVv1ix
zoUuVVvFZQRfRHtvjc9tj/bDpN+lOC2oxMATCBfkALDASXVOYn95vtgPsEwYnvG0
PBClut+2ZNdm6zfxQApUgXR84JWT5xC5zGLo3Gr6I+MXx1v77d9pQ9HqGjV11qIv
nPVIzcKz3jcnvGRRyWL28Ojfiicq3Qx4zXg53ze5gKV4pJ21BZt0LMOc9BBY5GwI
xRmjcfcqpz2Q85h2XhzxeXfG6LOAkHH1lvZsKWWnsN6guU0c872b7siPLbdaQtL+
ayJieV7jFNsgZlrSeKgNe/0eidNhDjz2TE94rmfSJhUuxk4fKS6DhEc3xTLaf6Us
nJk7qZCaCn1BWdZoYIvQfUXH97DVN48Pa570OFztaI8pzIvq13MZTGlEDgrtbaBw
Z7v40D45aDK/LttzAj5rWBIKjnvc17hkzz3vQcfxmfIfF0XXpmeruLRtUxCg7qVG
FH3eHiuO52ofeWfgZIbeAl767sGn2s/jLZ6rWWw18qhSNUpxi65mOAMOpPu8tk4V
9EpSn8ifRg0E33SvXuCO+QWy0Mw0buMw0cgRyn5HxAgEPqaPkuuoQV6RNtQgEKID
4tDvO1TYOaoz4lWgVBcNJdn/Oc525SVgwOnGSEagG1KBJQdkW3eDoac1HN9hT0dQ
vDlnVqVonoNqU79pIcM90VFRAH1u1jMmdln+IT4W86UUAS2S4E4dyZGBMpy62hVf
0+bW+5+TVaDGM5H6m9RFEimLl8KiY1s026cni/Bc0ITOy7Q6foxhLBmRYg447f1F
6HoNLkGswmEtYI/QpSB+dk40E+mQtu8Gjc/2qlOLwXTLjjOdfm36kKATXibcVfeK
93x4MNZNJPT4CyNO4jjFtREtOFAzNAgnUA9ORJTiw4F7CX+GxgBtsQGHUlvBzpqW
0KYmDQ2EQqsq/luVIjUvXpyi9xm3nhl1/9ATtBC4jt+edtT+f1kgTDdScuQjoNSS
QG041y1M+AJwI3UCjlYgUUFWGcrBZqfW4N9hCvnwKASQ0bM9GqYbSpGuM7Tv6ZgI
uZ1Uksg3wDAz/kp50Q5DLG2tOYV23zrLmWByQEvxQZ5mthQExevRTFCJoFcwb7fs
madY51JLljubCyztR3zX1EwvHTqUbVB2dygXC1NP0Twvge0kim2TwTRzu8YiCAVB
AepYWS9Zs58s1cHjNjMxgGDcd0ftiBiJXh2yWTt+pmG0zuo9dwkcBrdhFDX5E4gW
Kd8Yz6GNVmXXhEbLdZxVvTxZeCaYoC13ZjH5140ejL1TOlfURICSZgi2d++6pa6/
8u+7/mAPwjb8/0M3+d7jIT7R7LPksJuIxTeekyRN9r15h9IoKBT6MNhm/hrXicdd
2L6WdYwUH6LQUYt6BwjsRvA8iOvqKldYp6S4WCTmUnPZIA1P7miEn7UcgZw3G5y0
1Kj+IprSWISfpmYo6RbtNPe30MivyEYRKCec2yYUhapr1ZFtsDLXaVoU32rqvrtx
+MqLRUmeWGo0zX05hJoV3l/FMSgY6LAK58NHK3dydEO+p6O6MF+N7/y1P4Ez9qvT
rDcbWypPaf+CbriM4ZmC1Xg2E6piNjtR+T/voR9LZAhCuy0Vu0ZWhrQKayI19CDf
qlTvBh8uASxTbZrxbDaGZhcf+aNTmLO5CWmqcN/IP0Q9ybvnIcPSFtc7x6nnJTdM
dbim9lrUHWuRDctKdImnbEtW8ZQYIpyk4IuvXc/mjtsdhhbvxZwZtA1EPvpaH5Ut
3HrDs4uBWf0xh19wQfvlGFxZsdY6LGY/wnEnASg3Qfib63Bla6tKLOyrd6Fo7Jyx
F7Pk64INjnmC7HXq12NN8bAEjnEMBNFV3OpW4aSmrsGvq9gsBTEdzPDClaWGYpL4
mFl2nG8ZdLhuvIfNxszGWyqE8mTm66pICRVOQo2lcJ43pgFAxPW5oGB4wUsqBsUx
eeZUV+e8B0yjhN+qHob2FBKX+vZWsGpHlGs9xRJxHRjgobC+L89vXmdXdIYUzWne
ETv+wSdAawUR0kYbiC6fPIff8fGuA1HjGQmAwqimAuis4w1te4ysQze5jf+bfZRu
Cfxuf/DePljEBbZdpGOl6GjLiyqUPApEubX1Ck0C4c0nS8cOIDhlj/8cwQoJ5hbF
AgdJ8NHhSFV25t+qEdTmVRtv7TSr8GS/ZUWFVciErzNVcJJDVUPOZ7L+FOkotkJb
DVEvYM49pQOFAGE3+prugJeiOkQBFwbar6mPKuINBtY3XdSvCaSv6JuMEGQ81LeI
Fj99JHGRrZEMKTxva99Km7Y1WSSNfv5g9dls0QK9Y52vbWxGkBUnN233fkWKGXL3
yuxPM3SCbDq8XAltAd40SqACYvjKnQwA1LEnClcE6DGjGy+nw123xn0epivZpQan
Yt6dTYKhtLvvcmZGBTEVaGoarEqaSky9z8V18CK2qQsoARBoO62e+/uHPKkT2uST
RuFgjw6lpIb4hXBYNrNORNE3kCJtnPtBkxP2nB7sZHZrergpDB9JA/UwpxXQcz83
AU1pWshLAmRCK4WFwovWRAxoofROdW+aLoLnymevex4OiMcAlar1l6qtRFdxAx58
DJ6aOIS/uO+3iXnP1CzOm08BabT7EmIFJrgyUMVJulapt4S0DK9xC3UOLpxcrIq4
b1xMn64VyLZCI0ifRtvdRyEGlmR+gFRfuiR833COVzrvFRZDC4XBD5dU9B2PONaA
ufnrHMipMq2fhBoRl6ijfes89HVQzh5aFSbGZFlwJniSi2vOeP5fDQYXCi+4GrJN
pQS4IU9iQCcL6c4Y0v0JfrB5gd4v8Cg1DEoLUgmVm/PDqmkVoA8DmCoGgaLKHdlx
LjbzBI3ZkHgBF7cRH0fG0Q97ykdvj98vjE55EVAg+2LzK6qIwwd60fnODaaQ76d6
peBvgE2RobMquc7PBQkRs32Ddu/9085pI6qNDiylVAX6Qndyf0W9p/xLXTARPhkS
Tar1ykWeXofSQjQB2vpE1WRD13O2X9IEhhsJROeAFgnp2UsHlPIYl1cjmUbgzNre
hcTO0uoPy4qyEzWqfDifX1m1zR7an2+XgxpK1zWf/oyAbjl9Pk0MZcvHrwZ8zRyn
OvTNauEEn4E5ygYq28ypHARqFyYE/gMG4jVicikzIO9xFcpdzbaOT3ji01LwP1pD
HfIMaD74GPOCqFfkhYluBm0Rgii1uH7Z1Aigplt7gzd/v68ZT/+9J9bCMOyR0kRT
xu6ru5WBhmSb8O24aodE/qrluH7tVNvarhLoyy07BGTMyJb2JaFQOrSpDkhTzx9y
/Z/8mGp3D+aEzWPpBpAeS1icLs1eIryPdMSHU6viM4nDur96UZ0PRygOIGLnuwVT
/gF4lrcpvhsxxB229ZrDvwCPcjDEoMReyqI0XtXY2wkyTuoQPdokloIjDbVjpRKJ
olu5gc+crXWy8DVeQF9amdtwuktU6C/XvoYE5XalygLFegOTUek+pjs5mNNbI69J
bsxOgms/ASWPydfXFRhaJJuYeQuef+oKwC/PjMpR0ZHNl7ADkXSkCiNOrap0Dnak
j9b0o5mgjohE6+unroV5j2UYq/TXlGjQfojwbBq0oYcL60lw+a9ZiMBoFGlclnEq
QGf0pLkTp93qQbIHtGY4LSfhovGBDjpRcTvQUZGHhyTVgcPJgrEuU7aiCkrQ99an
8lZFluMt5WrSGeLbLrK/sSXYkQikH3WWu1Mny340meJgxy5SVaz/kY/ZE0E0eagN
86y0lh//mL6MlyQ0+ye27xs3ZRynpJOL0+SQjZLb9QJzFp4pt/zA93EUJknE+N7d
82LaTR9oIChJABsn4r3DDW1+bLuJMtU/H/l3RtW8E609PL/W7oDzg2iOzhPy0FEV
9IhRO0/KJMFfqB8YZ5UenRR4HeLGoUf1wVEKghZsupRcENsIUtxQkxDXoV8DHwM9
GTNEharDiOiAXwkC3S/oImbsGb8xh1pIFh3prKej7POEy4bSl+ufK6EVuWFDtxSM
Bb0QTvEAHnFAPrlBxeHCV3Vk1UrPvQ3S3u4EXESdcXCjJyiVP1UfkM7jFIxHvrMm
s3NEzj9qE6yxYIOj6P2i3K1bcqKAiehNuAB+LpxgAtSRKyDQfd/ERPcn7qZoR8gP
a8lFuHNiH+FKoFibmLL5XNiQ/E9zvT/JiZSzFzK2mywd922Ybyird+d2J4ZoXCh4
xz/12Y9HlFjrfeQCg6NMEPR93KaWad1QeZtLFheiMFtZiFMBeZjCLEPdXREJqQZa
t6htSoVkUxZMuTiR8hBa4nhsYF1xZXbehrmymbF0WqZhohW2bhoqwKxT+2n6Og0I
g/liT/MynrXEC3HoPhfr0MVJ9ywCcRuHl7f/7eZNYa1lqi0B/CifZg6GUj7HjCq1
iEP0LyBvDRM042whycP/daKHwQxTBTNQ+LCHW6ImbD5IYrYMo2AsFW9bpsZbot8l
hn2/fizpoJJgv8hM802hAyWMKkwdOF4QvQ7ob5Gz93f33EqxlPiejk3nfExWRs5f
w3cyfqcvSvfJS7iqKMKcxAs9zSRsvDVjjRF2BLoFBtlbvHRn+6UJFBwZyK0g7OdA
aISHhPiPKH7z82I9E9ZdkX23TwvBaXxthaKjlkS2SR/PKMs+SDYlZF4uw4dEmZ7E
Z8P7ljHZk856P8vUS8IwcVhXpgZbRvLGn4t1hO9uV/6pjjHO+vWMFDBpwtrQuA+i
khVe4vRQxhBBLWE6dUhBAZCRDuNIDUm2jzLvRdyaI9xsSF13kE3ziAgTCdoJH9Jz
+M9Becy3G7QsIGxDmZQPXa5jwz6jXqL7kGUWEnbzgGl4FblRvFGnW82kgBIZ6XiX
H0pwOjNiwBpg5P5+HE/7CmXFNBSq1TLfDvZ3GzJvzFCzY+BNWJM7ARxFmwxDgaQJ
gg33XcL4aIaAMpVFc8CiAJHu3u01BmYkUhUk+gwsApLwt+bzD9s+nWNfT9rI1E3h
KE62+tMuM2a0vMBqlslHIW79T6+fgHJJu0m3dYXOjkmpwTStWxBGUcewca9TXJrX
EKnaP8h7uulA19voxwzL8WDreGq4L+pmcEGdgETXgePJYGRYsh5eg2sY6HYKUt7b
guvBSJmHYAf2TIo1ns9MOYCjs51ZtNRpeL+FM83s6/frixxXmhYMyYZGNP6wgtCX
9mu2TOsB7ZuI4rtfpK5Uxu0Oy0FHXq+8jSCi0iY3IIGqG1NP2L4rz+qlxfQepMft
7/M6QNR6HXD4Jwmuu6SP1fy/TmHmrKNCkyawC/1BzBJwvs3Y/snLy8P7ZyUuf9Yz
mXS8bJDRe62FUt/VsWFFIx5BSVk/nh//iIYdrOlvLE9+C9Lp0Qmqn7uDtOV1ldNO
EmaScDZTU+aEnpuSPDawIiModFWe48/38/WL5Auk/ueehiREEo1gLuwrjL9ymBzp
/lzeVmKqUXWn9QJP5I5O08bc5W8sfalvlvIi0dmbViXM+a7TM6clIr0amEBjC6M3
1WVVBE/RwRGRJjfZHuGXYwDRPOOSpcueG0bRn1aePFcq8oIW8YaW4QhHG5CdNJvB
zkcACsTv9IvDAoOidJSR+67hOyVUDd8POCsqX4oXAM+BsYIZAvKJ52Nz2EWAdKYU
CzyC8d654UPsHcJszUuDNHOnAN2KsKDxplIx1HL20FlUhkt1dmPH/YS2CzSknbmv
cSqCzEPk99orHl4x0ODpT8yaEGEbdLEeMbVEPsPfTjG/adsowZEvCgYNMVHu0eSu
v1aLjW1EAgDI/RU/7KGQFnJ5s1GGXe2skabi4gizhVfhBCzRCRB0noy96bfIJcAb
91Fn5KQ/qSkAUX5UDz0Jz5Y/o4GfJLtqduuVpAMH3EQfrM+4OqzbpBq2ZPxWRe+u
WUEXesAFMi6GPPaOPOZd6WLOL/TyUx0PQaXHXzacUzE3YeUKZlaecKWcnMuYjWbf
Zcw+HkKWmFnRsZY6YE7io5OchSfAlAs2ee7TQGS0czJgDNd13tiqT2QTR+J6cIzh
V0qjSZSf6hwld4fkAx76Y4zpIZxPwYLLiq8kAly23ZAgMmND+jex5z7Bc2snCORW
ElDaepyFNXuBCz6EWP6YQAxRt2+ppXGKIm2xHStvPDGCoeYKb0kvEZJR3clB8kd5
DroHdLuYFe5UybpfcxMuBa+91iEWjdKc3+kQ+qcBLhBKinaURzKbl3a2D7/M7qoe
9Fv3aeSamy4E6Qeo13TzkBMJT50vaWmNDGQY0iQCRXG09xe+yiE8Kb8bItcranCA
iClENvgqJsvQKDeXKsaAm30Wr/OWscbCqHUaYgomuiAZAd7eQy41UKmbBOBEi3/s
jToKk9fWgV4pWazCexXzYd71jTj/ezMmXxxeuCq5NOVkUeSF9L/qG3fVvByZ5OnT
4n/xTvO1whqPoZzpuQUHYlbXyXXpYgJISvHVgC6EkPz4T6ZmTHhLcCoJ1rnbY+UT
HjHKxYhp+YzV7kS++Mp0/OotwHb+CnNCcSKMt35ZiyD1YGO+urneEFLx//u0V8xK
VCkbIp3m+Ie3QMnIsz7h53xkhwtMc1SdipJTiSQkmKIy24whmiQetYq4pDqzZAnB
fWd0dc7tzyTvkEf1r4P1t68prpqWvrpQsovhDq+wpZ5sRNyxbhmFX3RLsgg25W7G
Bf7dcKWYP7fn/bDrtZiA1Jl0kfuCrQQ2cOsRLc8EYo4wbMg8i6KYXUNOVhCvtPob
LDEeMBx47y8CTKieRr65X9eBGRYUBi56hLIgkHe9Pgzeqpk02SxG7qJ5xYsgL+U2
ZedToAWEVUwrsplxDU5y7izOKhYdkK4xmzlinLiAa1i3UD85mYdfTx2+NMiURgi8
aET6Iru9DnytDKcCGoTz2Eqf0gcWsxqVArar2+xzikey62lGip0jV8yQYPXmDRrE
vWIy/o5Z4x1inOuFItEBGORle+nVjTiMrYmBtXLcoV+kJRDhen6n7qJiQk/FuEWi
fYee4o7l84sw58OE7IaaIXlBTjKxlKCHW73FKDYpl7DJJ2RIpNEvPLSNUxBPHdtM
ga1n3cUw+nPPeLlgibIq2tr3Hr+NvOxqjCprWxGxtOLks7ZM+D9XrCdW4hxbgltz
wAuGvO+dQMGZ94nB+NnD0udPE3qsAhxQuF9vKJ98JX2mhkXzs5E5C5IkR+hAhxfe
S6lj4u2EUUYVr0EmaeMp2IjRa8T90Umfhv35xvGlsHUYblR+MOIQ+/mXcgF5mT+k
1hU+jICS5MQsC5De7UiJfvWkUtOq9E5qreEqlIaMiYNq9SpzNTtnVjJsNHeIm136
Kc3wkjCoE9evchfN9W/pcuhQKniTzk5Ggwx78q72eLmgLoP4kMtye6pgTjKCCTxS
qiE2JeTzZBkLJiZuy2ilNnlCqDHideBWPLoiZ6HuOdh1Iam8mr7YSEp37/df3Bf1
o5g/4PgXlibCv+lXaOmv8Fj02gcbYws+8RYqXheLT5O4KxV/0qMZl4W/tjgOulDQ
JqJvLCqW1ihO1l8wi9exOw==
`protect end_protected