`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
ddtXksX2+yylW5zu6QL2Lhnb2d1sD00763mmSITNX595NcHTEkwn0zB1Dry37fOW
FufOhVzEJp80NC5qZ/+F0Vk7Ik02dIR0elf3clrjeJRK85K4e3Hoo4xn7YbFUIms
l/8VZSb14+JVGURjfswrIyCUotIzlzVYZ6gzoZwDXIi5gQIBf/gI+KxNXPaKV+PQ
Ufys/12rjO6aI/pPlqSm0hCvftmBcnezN2hk1UeXgOIuKZnogjOsf0iJVX2aOOWE
6pD/psybjbnsNB6kH5uFTA5frkzIzkzl5d9+YDm9OyC+k84E83I/7/j+rk4L2dah
QJOvksSIzN867/4Qt8qYTQ==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="MvBXkzurAa5VTw+1JJ70nePUfoQXBvZOku/SMmg4TwQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
oRtzZL4VJ4iwysPsC8SXYCzXS8Fw2gtZTOskLcDV+1B9Nzn1zTyNtlo6lNICRmmK
ZRVu2BmCc2G+fmzynYlNTnSa7C0Cuel6FYpxCBlOuk3OF2tzAmLAuDyOH3Z1Yjzk
a0aHuoCdIRKv7BrZCdALt03JeUmXKPdOmIlkVGFl8yw=
`protect rights_digest_method = "sha256"
`protect end_toolblock="Jn9CQpRhJt4rnzZPRk+dOpzAubz7omckX1MrFd4p81o="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 29712 )
`protect data_block
gD6l00tciPUa6pDNTk/+tzLxvdHE2s3DQL3/JqqujQBC/Ei+vcAB8wM3doqg5vTg
mdfn9XB1bLOis2CVSfu295W2DNwHfMSTc/8BhCDRnTlLIX0UCJs9Za0+LoM0rMrV
T7EjVWppbP+Em6PkVKCwlmIQ7JKaifJ+Y+kjw9HCGboYo5074hY+K/CBbfsBQY86
AyoN0MKhsIx+eViNgnWjA5lZYArvsznMlXydPA+fMKVzkZk7bflfsqunZcYo7vUX
Z9iA2vWXoAnxIELRc3VUSFAaTQ7ipZNE3yaZPVhIfC7vr/UjVCYaQxi3E6GLhCc4
SB32mRmKehqiUGBhMxry4liDfkovyH5ksgLIxsoqbl6aT8R/zh4R4A2zrZ3QNQWr
DUD44BcVOnXeQZ704j6D95Ux+KRXqt6mfgeMlkDcpQC3vHO2bKGyzzEGTEJ0qt4+
qF8Cz7NinXCuO3ZzJ5w1oMVklsMl5FSWHd5ShmvxMLUKfJUjZaKu31cTUywTu7n9
rSRZcC/JejjFvrE6qlihJjggCU149em3E/kcJzO9Vf96hxVBnTf5h4uZPfb3hDja
rEKYk8kUCtaSYYSKiggRH5Jcc9fF/zXp/QEPcY5L8P1IFls13qI+wd2cmJC9l3jL
ttHiwESW6/xUgu9I+LaUNk0+rUqhWzhDf5EQp1VcR7mPfpmBPvehqRx/co6agyII
GJeevtGzxAnmX9HkWKKgOwlfUsqlTJDAfJT5Dv7i9jecnr8+thrNtZ6gkebut0jK
8+ZBKUS2MW6fVW3R2iqV6Xc3m4n6UfR1XFztuToiJiiZsFnkJxiBziyas/RtHBP5
6CLs8Luc9CGszRUO8ggDuXTjSfgWOqphpUF9L8cIx55Qi/DL7PecNR0GwbusqV0e
xzM9IH+LcGNE9makr7uj9X2vWcxo2ME6eNhhqmbi6q1m2ZZELkzPOSqaeG8Jc18H
lsBmRvHDdL0L7ODK2Igxbq2OakZ1Sp2PkYu4XiZua+GcEjN4cGrbyAGCiB8jl9L4
pCeP0a+shg2QZeBgSYiNfqUP7G8sFowZ4iglcq6UiqwnX4MvwxXueGLPLM7Bium4
4dMECvMSEbEK3wTjoiInRLqVt7iidTzldFebc7p14a2t/Sp8TgOrJEkiWwAmMfHp
XDpNbId07xWfudHQr3KOiMfw/zEflywJyaL/JhpFy4VBzas9XfEybsJ3APCcTrLM
pP3KCH8F0MPsK5KNzkU4ztvERuuh5QBDqxWyIozfddLGdLPTfGNAPuXxcmoYPhk8
GaVEr2UPEeQ7Ofy91dlGdF0uanjD0xhXVGXC86w0cAgqsALwBwCNHeIHpB+i5maa
wHBKdWN8AxVE7kFq+ZZ41UHKhyQj54uroIq0PCU3JZqGvloQz9K6qcHE3AvDiF0d
TXjYFNW1mFwF3czX+6aG2w3IoAHBEJm5y0S1OWptNcG9z7+5EEXBe/np+Diz7Gqr
7VWZiA559qwfe3VmoOBRL/ahNhrIBYczsv58WmxGk5txONAwWhbvhYOYUiLfcudz
md/+5uzfUJT2q1fHBgH3EraMgA8acOpfPh/2Hao9oIgFyOEbgebdx/4rEGc9FW5W
wizsOGpd8Knseo4yXAfvu92DqhvnmJoS5cReBma81M6NUyiTYh/0dGlmd+CrCbez
iUxZPo7S3qZH1awTEONV9gX4SHIJU4+zvwLE+cYZD1+Cu2D5Dp/raACF3E20j+6N
Q9ATI7MCLef6evTmzywOtBmpHd2vNEaWjtHTKv10restlR8t/lP8pGFTyxguQfWW
aC9PxYs6Kxu0mV+EkG4RURsbxs5hKTrvaR2E7sA5J2KZbqcdq9JEsQNZJ1N4ekli
Bs07lzpltS7tk65t4E4zlmVrnLRjaszaZ51PffIw0Yp0RXeDI23xpzadhd0hNJl8
j8NQAa35/VHzKKuMIFH2kL6IfIuAl7lOIkHAI60Bey68Zh0j5SIMhm7xN2mZMhpw
tYvYUsCI8LPv6gXRXKdf0m4IETdRpyDY8/di1EmTFMoEXMgnpZolJwp3Bq34rqcu
PjI/pTS9Yh+RbCFoMpJeQASB23I69wcMgeuvyFsgW9yIx8rYtqXdyQedeV69mi6y
bzGpKQzUOxjO30ID/hTrmrfZLviEVHC96v7bkWrnNPuemFE+jz+/GOfhKbbDpe3Y
UWtf4dI2obPgyak9Ncl2a6Xfpp3HMyNYuUumOfrfKQpx6kS1defDYFqKGew40PgX
HUD/VDgZ1/cFHjPSVjqmuL3cfrnEDWS4KnWm6urXUqCACW4IFEmnwf0D3xXl890Z
NIxsOTl3cI0oYPMuomgFk2zSRl7Lt/a47reAM7OcoQ/fqxmUpnz4gRzx4qTD1cVm
Re7LgHV03rCBkIIch2uUwuMZjBqOCm+ziBZCE1+3CTQ2th0zl/rLHhQMdaeVU1Pf
RgJREldijty+4dpwN3h/6G/UcPNpM9kBaHw8T9ChI7160WSP9sFffIHiTlqgpLQ8
cIiR8O+uXoOtcjIn+orZxxTitpYyrl9oFxv4JiqerRdBHMyF8DEJ5xVaseSPdenY
CwwUATrMz/SaQrlrRHYoZzrw87XoRqO9hCmPvyWAFYF6Gd9QK3D7X0h+cDl6WiVE
T5Uv41wZPYd0I9jdNF9epaWONjZRUmQx6LL2rQrbOntWj4MEssJJXq+sT9XtnCA4
eYRUQXvHxMKY8SHzRFXzY0951i4vC1dkQMnc11URJKfSniyE3050e8s1q27ziyJX
DnI6K3DwjOHs04ubYiaCHhgNKUZouc4ZbghwojkToeDg2OXD38ahzVIk9d33vklS
bpkaasFKE07SeqXalFt9JNKoZ51HMy8n5ExOoKvCIdtij62VG9903MY6gHgwWYxo
Zy/cFPlml5O4TYi7eI9lYpvCN8BUx6RbDBe5OiLKhk43bVDmCr6arOBai1ky+eB2
myioDm6Hdd144BU5oq2vd0YBApkRCFlcKznEpONPTs9CayoV9CTcoDHnSmZCq43H
rYkjpFp7MFZJ51yLVM/lDXbJR4+mlZLjyCyKbizN+P1VF1JdU2cFrKdYr3MdYlLG
2kJR8N2vcVbOF9+7ltbhTmPh4B0g4YDzHyiVTcGAoi5b1LITXeQTulpFQHcGyG+k
GX7Jh7Thfg5ll9zDAjjyjXhG8wBwP/Hs4b74VCuIlNMTWk1luYPxJz9YsHi0NaF6
jzIITqBQXpOtuDOi0HNn/YLIUdN0pMqmfRqoB72dqZovN6jDvQfd9Yj+Ot5o8Gj5
ga1PwGtD4ceCuCva9P849v+1gB7rPTflzm/6CwGNjDIUyYyEg7bZKByHx3+Z1qBX
ZM3LOCbr1PjCXEaNwAvuYHlpkTMOfoONTsiDii05YsODYNAyIRmEYwpQ0bLGTq+O
ddlU25A4229VxUfdMnEJKoZiXrx6LyuZ05SNi96HKDTi4Q1N043vt6MOBRaEP5dU
4gsJUiJLWDzpoqOTB0kU+pnQbSlbB03SBCNlioZGIDAXnML/EmtDekwRhYZVmzNY
TIGKPR2kM7soPfm66Kazpx0QWIPPm/FqIm+ZYTR+3+sErSavTnE/SRla+Mt7fAzj
Efy/RsYV0xpLMJ2FwxMuUeVLwnoJKWr5SmjFf6hYZwMRhylm5ZF/ucFLv2hhlCJg
Shf9WdWxmn6I1MAoHBhys1CgNYRKc+448L0MA9On8d021DEKBcCcBZCDFtby8LUK
UZcdwJ3Mqhz1W+fxyCOefFY6w95dVnznaFUL8gWR7ikGiHaaC55fVEPfjUrNZHEc
n/xVUYeMK0cJALgn/qHBirRUr1CRMxLw2tvv+GszNSmR0V2ndqebr6XexOvd6LZe
CSSDAsXH9NdXKKtAIewbxvjOgjaUpRi6i/kEkPOeBCyK68kEXW11P9oWDodhCP6q
ekFsgyL05FZUp78lb/o9eb8tK4DSx0vkv7hs4RHbFCRm6AFhjKEAnbkvyWltaQUQ
CbWW2a02xtsilWqyBjOk8UasEWohIu3nVSEPflUBbfaAGbkEcNXyQYhGAZUfvK0n
SwxExFerO47HN2wCj6PwUHLHwuGBKE4iKRTWALermW7kKAGW74wGx+DlWb0ZCD+f
ffggQWhQ7CZCJDu7jfMuhq5cdm/aBqbyOEzOcVDoL0dpfHz3RAB72P7yv+HpIxJ2
NpBW5FEXh8m5aXwy1y/GTieRyayIx5rc+0RB5jJy55DxqjR8dIGeXDbfOoDEJJ/Z
tJS12bbMJHG9fG1Ou1kqxSGcopBVBrrV0ovxFh9nSa2JRNHacfXUScHE31qK5Osz
r7R/cPi4Sjem+v/c1srjIl3LYbsDvhgDuCC7YmkjdyXBcVwXKhPEJcBwXns/WMlv
FffDnMKaER/6pe1B/Vrgbq5+h1uO1S6ui3kxMjDFJJ4kwcZ7jTKKJc/DhHOQkBcZ
Duuo3R2Mj2EGogWZqrTZhEClKCoPmIprwff7I3pe2s28ivwWHRNn6iMpX9llxchw
3TgaEP2of0IhYCgEB31uTIy/EIlWMj3jDIC8iS/hK/Xxwg3RRf+8jel6oJ6kJ8S3
DjjZs2rJkOtXvIKQNkOJ+nP6MoZkWuLs6hdCoF6GekcBZBPWiWFrfpUsGGUZqghA
nGFe8lhySk/1doX33qiW4wwv1718kOoSqmQmbmhMsQ7TohIuBgpM35atSIxMs2Fa
ym7sBam5OraoMKemiPdrJLRvMRAYQI2LZTEho3d8XpvcEsK4TMFPKum+QhNz4V6w
zAqoiXZMugXmRmSce1YZv9l5b77XQpyDVTyKbKVJVcORHbaDw7Bqai+yxg4tR41j
xAO1HH0eVv/jrboQYUlEaDrvYZP6lVPby/DkgLNbUVOO48WV6TZGwT+zrZPJL9Wd
T5POFt3ixrq7Ukl81QytlICPY9w7MIEUj1AoNzhXAwdvuf+yo2HGhvZavbj04iAu
X2T2aFS4AZGz8MENtt48g6X5qfMNXyRe1l5E+ok+PjZ1E9qV/Fc8PggtX2CeivUV
STV6WRI1AmAACVbWyXe/6GXHtgZORGHSCVetWxXweX4khfR8X3KqxbuVVGkhHmq/
bWTbhV/BKY1TtgJIiAlEWXeuKyqUjvxL731/Hm5NDmxHMg63u+0RVCwjEALhepUp
FYmjbZzocNi/D58rSDAm7pxdGRdgDBdPibneDCzSQwK/HcQJBsBwqEBDc2cP2Eg6
aNKiQJ413hb3zfSgfu09xKN6eSCSgJ8P+3jiiM0wi5pac4C7heRMNMMwcwg0m0fS
iHB+Msf3/dghtoJ5RBRDdbitAKiB65+mN1dOOqTLusP7QnXHq4N0GrsJWtHgSshk
CE/k1ahklGotTBRl54Fbzo8mPvXSJj0SzD4oy2/H5ALbGDsJ4zijwsAwwjEtoaF5
17h/3jtrwtkdzuuslgDzpNwBKn1Lu9RA5/s0CJQeNbQrR7VHtARVeatCGyJmGvKh
Bn4QnaDyPJwF0zHO1XAVBoem0TdnTWcZNcya/NpKTMeXL4Ql/0gz1zjlKTSU6ZzP
KbicbG/F9J2P0Q5Bz4gksQedFft8LJ64ZS/UcsPvXrtN3BTiXKaPRaQrTgmEVp2Z
xpm9qqHjW+iGVygDw7rg3EFGHb+mxN17MZCjWGzbBCVFtCdIdEAM72giALyWkTdK
6zoA80xp43VIAv4qZAynVQZTKRR0dFYT20UBozdfEbchrO5T+siDZ761aBjL3jpm
cqSjw8/QEZF89XK3sQo2yutWIIVwpvQ+RqXFS5K3A4Ri7haAOcTo499bhGSjQhJx
XYWqj0XEcoCXK8JKLpBQEtJDKnoeOt+tXW8RFrt+llFzgs5KaHixlPSLXwd3w45I
oLn9AogfnjHIRa/1Gs56h0DtgbW2Wkiq+NXTUxPKm8iY03xPH1vNI/pCpyZ2ZHtU
TS3RfgR7bej3oYlSe8B/MwzbKdZaIT9ZqXprQu3bNEevfn62NxYYFu/P0s/FJ+Nm
rz+GWBHQgSelWO2yCw8oeOMloif90/Fu0yUllp5pLweKRRnuvlcHwlgI6TBZDYqh
S/u2UnXoe0BOeQ/QrPntLdgW302NmsNvcXtFIID6SZqyNx3KexVJqCaa3dg5IDRY
KZFaXpWq3APu5v+naq1gEJGSsjL50uTrUL0d2uWXGsELVtt3a7DD6X1/+k71Zbmg
1qWbdwND0llNHUpjLaPchQzj8cM69p+w5RvzjotRSYL1KejpQ0n7rbC4YsqgnabR
tphiQHsp91z6iqUbrSQyD6wAb4NVvyp6CBdhZgXV8Ws4T/RWLD9UoPfjAFqqyHt4
d6sVPga5KVSCb4iY+A6dMlZckVUaiTj+S+FDrod+uAY1RLBdIaVQgm+4L2zVY3QG
I0zFfvvfVZ1EBBDhVrIuocfQwwJUkni6XfSjUZaNrrniLBS+jjnMME7MVyO0c0+O
JM8Iv1PN/I8nHUqstFcP0/+IYzDp2vYJofw8I4hd1I51hdEosx17I8P9VhGWTOLA
wWq47q9O72OsWPHB2voJ9/sFAV6+7XjWzr0mYek1/dscuWccTgTKd4w0F98okvMe
fji90p7Zr8rp1Fi+v7uBrcg8aFh6A2vy20TG/aDWTIS88i7vo7p/jqcDxMckD6O2
ruLW1kW5PKvIh18VYTtjS16IFDF7yQvhTkiFEzwpZTtaxvNuiO8IEb3/n0vQaQ+t
RuVGb74is1Ns0p6pBEYBgJX7ZelrheRZmpbvUvQQKNsXnR/I5oNdbtK3gagtMDbM
euToa1aoeTfpPlexpDcN1a+pJka88Xv+MErKWWrC4l3t/gOAvBCWRtAeMPct4vyk
9QLuJ7RRfUltzCnpxgqycm34OrU1O7nE9g6YDwZD//MvTVLrKQUrNALV/YXfYFqK
Q4fgI0vW6BjuYa/OY2wSCm84ZGMXZEVAJbY9wHpKdcg426tNNs70m9zhirf8FNwk
58Hx3Wo0sV5GzlY+YNy0Zb8oYoNaLrA5h49mPl/8Tq+9PLsEohMAap+Q4vvuVJnH
koto1HlYAu3/YTzXS6atC6DLG8Bcis4PAHL/1YyQg5wftr0wnPzY4mlokEjcGZmN
6bxK1M2zrgaiR2SKpatQs81BejjQW2JnOSJPhauYsOQAquxP2GudwHirETgV04QV
kY+rYujh4WS8IzvSIzeqibaTkU5GKFLY9zPaChJ7ZNKGu1Yp9ldKH/AgGy34GebR
PBNnE4VvRDbvHmLrDCgKXKKHDTOBBxgDmsPgf1x1B/efKpqPp0cvnYmg4MqxWpBL
WfMSOD0xJ35h8GYdDLNMGILVn/QOcDei8WVhFp/qhTOgTfIXPZRUc+mBumYvpJuP
4/1VHm7q9bkbMnfKQh8zeZycoq90RHIlN9mMlLJIfLAy5klcwbUG90v8QisJgWbz
WGA5CNzD0r/itz8TeVXyJ3mzaRSLHOlpbrMVaF71JOFxtBQOehTn8Rv99DQusNsJ
J6Vt2wEmgPyH4cMRJuOLHba9BlldaTymvoIZQydscsdFlZ8JNv7TudSFk8frQn/D
b11s66H7fuFme7wNkYeR4csryjOUTJ/OxqCgiigqO2lraNBtAEXTRjHoWY1gV8ld
R41dEQaCDcJXc6atmxMzBFk78fBhRKwFIDucejkQtQDN7bXeQIZtui04BBmwgR9a
yRM1JBLWNwMAyV0k3uzRFD01bA/YZfABpAA71DsECo10fxDlWLj80iNxa+G4Of1A
fth/zy0ksKN0Q9eERF9i6Tx3xh2eMoEno4GqQOwewI2EQPs7NV1LEOgObpSVWXZR
iSlZOYJrNbE/nvn4Qi+kMAGa6CNYhvkm3Klk8jxMLasbf7kxCGhaiQ96VFzybkYG
qfXN3GPRliJC/6L7xBYuUS+4JNOZBnSYtctcb+o//DOKXP3u7o+vi5zHbMB1KhbI
yggiO6s092N94R60ZLXXuvyvOBJ3PvmjbdoW3boTzSYADJpulWml5Gbp4E/D/ClP
H+kfz13CDYOOGpK1jxzvATCfSm4qaKlfWnzjW1xSMYqd3XQurmbHphK9OPIrEdfP
HSObWJwDh39g2sU8r/HX2wkM1Fi4YfWSc3biix9ei9SAHRo/zagsNX7/z4EFDRJL
jYySZx7Etu407BE46OHS065hiBrH28HMN+l3NOcwj9M2TxE7IZTDTi0OgUWowmHB
zBe9JZU/f8Esrqlu8mMi20Buiu8bfColJzlGTVp8kgF35OXSqELkkDaCQ5014TFu
HdzpP9kW2U5qGuN4Ss628EcePtYYfx7XHEMpryKqtn+nZzX07ShXnwLfXY+YWxO8
Iq147n+N7XX7lZEmTuHAymvBhGTUH51WizE01PDmP85dlPQ20h4U8ODuDxSI3OdQ
doh6aRlptOjC82BofVfcopL8ZLlxHZ7sKB4abMiERVracg/fYDzx6DWuJoAp9C+F
ra2rw3Cdx/uhu8eJh3UpDBYrZJPiXPAdL4n0t6pgW7YHkVOaI/4vb0sqXBL5SAG2
r6rvk9vC316I7wRI2Jx6Ewh2QDDbYX3WRJXeeQ89XQvRIDXJHDtPY7MnxvTsBtPe
db6JNFU0GO8awJmXKRjeqhN40NT1JbfzhGuhmRvOj44AWyp+wfF/kjPWJD32n05y
KP/SecHu3muXHeGD9t+gx84+P2AziX7Pkm6r+WdHrJg/0M6rCcfVPoerJ8vcZ/62
K9spVgBZwSSyPs/NpD4t1gieB/DWjljXMCDKhCmsFJafR3qELPmn89WtNvQyBz5l
okz7Mfe50ycZ94Uj9jh6ap3qytDh2gmOHYrPSUOF9TGfBMipCVCXGoQ9SJ+agqON
+UXylQHdr0F1auKRJ0ERr5IPboxRlBRGmcfopxepsKzOq8GAJranaba32qVUxOJ7
GeuuV1P/UC1ZfoYsa5B/2frIF1SnByQ+pJdeVQ7Kyxzhd6l2e1cOVL8MR2VvyWhl
58r/LK2l0Nr5DsWIUnNBN7HB0wBnh4onKjGTaWG3uIvx+o8bOSano9bXyvdrNjfh
wqVts62nubpH8UFRM+PAS0CYDlBPencM+NWzd/Kb/zkKuD1Oq2qLEpyNi2jdlYFD
s9dHC76XDiNkWf5KYzRe4WK1IcJ6sftp0X/TBhmKN2kVQQpBPbsva8zhRS0DyOl5
TH9Djfd4M0B+CWYEMkMNd2j5BzutdRuD9SI42fiPZCSzQW1K+WdycKqVDhB3EeIi
Gr1g3dkCiSG/Ay8ZKniD3jipTavvAy+Q/JTylVly7cyJ/7KLVZGFZDMK7bVAVx0k
FHBDVoRS5MYqr7AFvVPaLu32ERofXMtE1pqclygVSyFpUcaZ+/Uha/uREbJ7i9b/
8w1g70BzJ6x+koaJO8jhCVNIXElsKG2jy/Tv/FcoZYtHN9RUpuUqK0BbjVWj73v0
DZPiJfZd9aiMfgCzug1/4num3+ErSql5WMesK//ozXl9P/AaU0X9HMfCZC4cNG4b
goKBmkjoOfHA93lxuzTkMixa8WNYLDTVVbfYbe3q99PCtmgGiWWk6gtpAfNyWAIp
lp9HcNC6cSg2ze0ZTCodP8CyiBbWvLipsuCBsOGZA0kWkYVAmD0VCBtAwF88F/U9
WI6KosfSE156YqGIsiSbSBEOC0eKJwf6vEQKHnsfuUSSATqwq/apQy7eUMBISlGm
eUNwXRtWRTnNlshIlGltFDghgqXGAJHTrI9xVIASBLRTXdcamQFdqUjVKCFKNKxO
IE4Y3POC6+oKueDeE1P/cW2KYruvkl63yFOb+H4Pb9EhZEuPI9HnAti8ovE/r2Qh
Ymehpb+H5c0R8A872mpH5IhPof4XQQlgXfM75OkHSPVu2qK10PpaWAE0lg/dpiM3
L4i+sTKEj9VVjUMma8GNxedYGPNQxGZ+X2u/JGR7SNplTl7qFyOOVaDFxhiS5Z+A
uy+HPlndRPPnyjr509ZGpqw79UCkkzhoTIAN8DH8TYoeizWjQBsU8F1C0I2dGVt/
WHE2gkeqATqFvBT4FJitbowXbdLnEI9gvdl45kbs9Na4Npcm2L2DWsb/9kSKlLSl
FYwEXeARWXlCgQk2ar/3I5ejKESb+rYHk7Wrv3qrOBx9LT6N2Q3RMz3sU1i3JBoi
1ny/NNtSrS2H9OnZVVpIMEEJALBFClFPgGInrihNoSPDgIGSwtkxE0NcofHvG2jg
9c9zUBloM56Xi783+LxGvmQvcDCKF1rFYnj0P1EbdCaMz0BHkxPJdjqRVQySrx4C
CNzqq6cMphi7fwlaBIkKJBvE51PmCB0y5TEJH6mnhbJjQ9PSXLbhTrb16wgu1wkC
E3dDq/5LxKXhtR2eyQPWHQiaNOVBto9Q11uNHUaSaTj/JTfhuk50oXBIjGbDMqTI
Ifb9iSOGqeab3agOFVW48nPbV2jUVWG27HOVaJFpBGkrnJhSxuf4JKzOz7NKcQ1K
YYcYRcX72qvcvUPZm3dZVSsZlI/rzbEG/0T+kpbECryYNXH+F1tCz6eXaIq4V5mY
P8uX0Vo8hquOiy0u/Va87zbEQeQ17/l2st2H1UwBAUEIwGyA0veju9s6TuWGAPib
NyL5ZDrrAjvo+15bisBgtTK6GYRO2iN2n78PlmI4Nu/ZfTSeE1pkVN3g5//NeTQy
B80348ivbsWdXDa53D/ULt1WH8mRALJA6QP/5quGDV0BCugkRQ58KeQE7NUV3mPz
/TFTKTpcoQQejHELtyfHqdOYGDEtLXVxUeRCaYkOqt47og2k04s0kmop+8372WNB
inS6zVVZ0VlKycdwAlext8JvIbmfrDZPaX58VKHldgPiqW5H5lCDwhuvY3rW98gu
CNPEfNNjJHU3inmd82Ts8J5z/IwNfH7q5FBtPA0X8Lc858FliqsYSp/btZTihpLz
3NkWQGNJ5UJxWkMCtR57Vt9MHZ0tpi80frB48kzwTqVwJ6F1LntIQ1ofNPFaMKfs
QY2oLvf/4sHksjmwF4lVYNsc5AidbBDVX1UyYKx4Z+k8CO0ErLPYNAF7GCxiGSqT
1POeyiooq6iz1RNbGoRwV7pdkheq3OKu0FGpf40uLXAUuPKnv7/bDFVY8f35Usvn
hKYf7f9hprAlzpor1r/4SGi905X5uGyb2z6Jd4RbUa/rGLeWDnfoq3YUayuEYhb7
GpdPotJLbl69/1DaYbxmhGm5xVv9Pb19F0hW+zO4VqfDGn8/ig8ifZ9Ko+5oWOO0
4dD1fuJATTo5H+4SmTc6rCDAcTdt3Ja9HBb6SNWFIH28EF+m8nPQafifzKClSzGf
aPuq/sQ2YjBGMdFc5O/5+/MeoTy+liVN4TFuGbLKl6ydRu+lXraG8VlcEmhi5etH
2dEH1auOsnLVz854IBlC28jPQCLbTvpBr3Y88g9aK5pyq8QeOEfR3IQNaGDYK2Ce
EpGRkE5ZSilJSLaBicg78s1CxTXecG0FCKeKg6ZE5xIQGPMOPvwJX1S0/zvAULz6
2D41Su4qVufrUicm70zLkZ93mpm1c4seQ7AkGcfgWf9/CqdR91WbiNb46sfmCG+I
LlcdXsmGHe+PsyALRqWSb7q+jYaUmitfX3WjfXPw47KfqLgmDHHPDSW7BtkeVKcS
UVntsuH8kjPWn4Zv0V2hnjpIdS3DVjLiqzyBuHiQnweVPcDIDHhE2cHQvsotzb5Q
+VIQfHCdGn52CUMGvV0V8X6wQ3r00YBywrqGP6Zo4mOnz2IKiY8OuF7NaSXOeANI
yawu03XtSu+y62xT97mSH/WKJZiojuOgiBIk6zbYtOh2nDHjuhVGoKyhHlFO+P0M
fXg0SbWPJiylET5RmfJ7esI/cv8hNx+JzYV5dW5rYN4kXTxyE1RoQUloQds2IdCF
gQUHbBHMuSHjeMnYJOIgbYBY+R5f9Wxg490OcfFmwVHp93AhRsE3+5i2agX7xE4d
Q7uua+kBhP98KljGZPwAIv4pWTe7CmOG+shl3Ec/yxpAgi+cKrSlDqjveSslZyEP
qarenW7CDS44CaWdYFtzSBB1IAjnmk+XY2eN0UkNGWplMvBJKd0OG/9hLEyh0uhO
O4T56UUBJuuHFGH4NlWMsYBsBiiutQwzIeZT9jpFeLe3dqe5qx8UMk/quALKzpxr
I2uOJEIlDUuCqPelbNgUZhdmMkyWK+QacVcm0XSfpBgOHv3NNEoOM9eF+vL6FiiT
XH15IunJ31sCy7USfE1t+1zB6Tdy7t8PXRQ2FdIWTzIOVompPwhG+rQEAxgM0Rck
oR6PTRjHbHuPZTNlNhcBbY/o3DPhoKfDfeyDidT7/7ULgNFZ4BCo6FkOb6mjNx0D
+iUnub2wiYljlUu5EDA+QBZMz1nHUUCQuHD2Uzp0jxpN/kai47KtRa/v6FFPAfMY
DbOFpmrFCgNCXNq6t4Q0xeDf8sUZRBJr/JNTKF0phm+iJK9vUY7UFIZj+zdD8qpM
Cc+44jvC7iBsGLosthdaFmZpDa3+afAFwszWMaRZ4AnuPsr2YQQ1sEeS7OTCBi18
P/oW8lcrcaH7yLJ0AX/V3EqaZH0skoodzY1mVYV3RfvbF9CHOB60YpojPUh1uSEp
oSjpMfUxiQfRojmSue48soHRPODWokKiZraAwpAnzP62MT9pWpZ/OpqLeoXxjXry
2vRxoMGat2InSBmhDSpWudFyucMp9yHKjaw38cEQ1hnZtCPWqEaiB1lj/oD1bhcv
2IXfwAcxy1gIy7v/urumqP0hTZmEOwko/M/EkdAJtV74ZPPQVxdpmiUQ+eejKgF9
HwEIs4eWJswcFxMrw2EXZo7BTfRh5fXSHeiZOkm0keLTrQibC7QR4oNWGnCKenrt
Q1EMpHOMxny5tCLg03xjBYZ/vR1+x0r472YFgvHBhvFkxwKaY4Hv3YyVfAXMH4lT
fJu4TS+Zr5+/ZaGN3muBno6s3MiTNOZhCnBtuIGdjFBtz/erhw0BphSpaQ0LWaek
fTdK47SfVhQuvesGhq50+K8qCReYDuIjGSkumZyaG7pfTNa8uhWhB3qQvHQhnJpp
CXko22aNL7qAx5svHgrcwqScB/tIMGbaENLUnRToesljWPuieRAEy8BoFZdCzqGQ
hPiU/GKYkbSCsdLBsWP+ZJRsl+wWNZLKOYRVhYNFa7cpMKongjV9NjtHuozpWzqc
hig/+ELtPRcvDDKgyitDuOzvxep9SWrObJ/vGaDhLAKvyXILYAEGpF7VON/hwXPU
1degjqTCz0WqVi88TecNxfg/14lplSCIcod1gT1xTfbBDf4UJItDhcZQ3J+OWqur
yI4oKIzwH+lk8H7erphNdvPzuX5Bc96sdLS1gbK+euAC8EQ97iKKxX1jC0Sta/yG
z0o4Ok2hAohqHUXO4McxUB2k393/xdI1Se3DzS5eCLfeLpt8Ae3RxwvYUK9V6jAA
ZrfU00D0NZrh2L2hSACKJ2OWnL53t8lteslBgV+CwbZm0qzp8Ao2gVsCE5mec+tx
uHiDC4rV6x0epwfNtfOYBGp6StjO9Z4XToIDGtXWx17k7xOPnpl/LYrIF9xDfoPD
Q3IyHTmpc/gyPR0JK7HKDVWxGZwiOwO96/2dDAuRYBBA8ZBU9olA2DvnGneTZFQ3
ETory9LlIfgVCoLk4BPJNeb1n+8gJkrF01DE+Dt5qtS1E5RcaJgQ6K+a6WyPfw9m
cJYisL+vbulz90mnKUlP+mvLFkJITvIxOTu3h3pE9ptfWNWbyLooX6Bl+NC7zg+3
V1AJcfmgZ5pNWgXPaAL8JFm0sPFNzMRXkDhIa+1nZw05nq7cGke7tfmmqwhKbu6N
9tBQEtnlyodAVU1spZnnJwldm+cqRFJVKvT1Pee5F2hG1xps2V99dANvZBNuglln
ilszuZO6hu5aJ2hn6QlA7HBdEqGbr1oQF0Y0YmJAOz7tiNb0UkXBiDE9yAvCVduK
hikvtme0JilkaGC3j/UkbRcEiDL1SGDYpqvtmFzfQ6FGR+v7dLkd2W9cdWSnmGqW
/PV/oQNLROt0dTDUkuWVkJWisRrYTQbugzjuc0ce0ntXqm12k8HS4iyMGF5PP9bt
EUzqtglhLXedXRXWVLoP7MMRTkbTTBBXPcHFkYWhmHxYIb5dxeRgsMX2NmkWLIWZ
L2SO9n8QGFIH0LpxWwnNIvTx47ZDYVPd5cn/X7+DsDuc5aTgcyt60bM/Lvx0Jsyo
4nttBHKGjTjgtAnVGKvKbOxBBhqHjpG0X2cWuV5NseMAfXnmcaZg7OYrdZT7BZOp
4nsMy3Add4SnIg7J+5e8t1r7hDgFf1kbmZ8Foynd5+27v9k+YDzdYjokrD49DZxo
yne4OxFDFS3T4GMPighcVvZkepmWYMjn5Rb0SibLNJ3VF2YRgcwyABehIqlBM+tP
BV66Lp4S1j/cC41d6uiJG9M5kAfR6yM2eP8IRDXqTNeGP3AuvIJDeSqRE14IiBNy
ldKihV6T7V/I9WpuLYoL5+OXOAKYZ8WccOgIcd71KBf1Z4lqWB2BFn+K6mrwc9lm
e1FPGj+e4sXeU1TfY4RGt2KgL7oo+Cy+E6vUL4ej5yTcJlvJ20ALFFZSeRq+w7qW
YtKVNpuaOkmES5LvIDxnRQH17FDYUD1x1/J5PqsUnas95jR4iZ6yj/UH5fb4s0Px
plMPYoVnJTX39b4C2ZKlUX4VFpsDa+Ply3B87GOVr3wXAzmiXr5z7l1K6OYAlHAE
hcSV184A6Q+Piu4bJY68C2yDJvDgd9DjVJsHYfzfazuP9jXRz8q2SY0xvJsfXUT3
HawJF28I7sNS6XIHGVrvOKdC9MpEmvC4S2ASnPJ7oqCzzKM231g4ctCZFws7ctY/
HSR+eCi6AyRVbnoUFkrLPjdZmxV04GNjRXbv2ZDJsyaS2AtNA7cGopBcadhbJsWB
UczgEZ2ZRKTuoHiPN4/x77L3MhdF0gisSPdNQ690ROBpG/2Bdt4Awm8dzpf1B7dW
wNBDpQYQrCzuJ3VpRetTJXsvmnACtaC2kS87Y7/V7x4wp7G3owZqNUKoPhIM/pZu
ZdXmTHEckJKfQpli6FkCcTeR+4WJorvDFgerE422K5s19Lhz2x3vJDvEV/HtWwYZ
XONWsQba+OQhD8a6klDcO63UXgX6UIpYLIMI1JAuR/02jjstYfovxY96Ibo1URep
e2oehlGcIgCbX95OcBMdh3TqxBPt3daRpnYYbqJdrpE+QWnkeuK7JJqBWZ4K29Ak
G1ROIXYogf/zwkU8Ofvv/t3baz32ZoflbtpUnCbLjb1LiiGdQqKP8iL+DgIZ1xC5
cstXvnEdSbqMBzha1NBsnZCuPNuHFP7uodx2DaWmXi97HxUAtNNTwnwit6BHSEB1
ydKYoX6hNxoCheAMUmzywJnM0zriEvYUPetUIUEAaqDVRFGUemxy5+ZFmBK5SgpN
0p4utJsxMisn+QOyBtDN9XG6tLmxCCgSVMMZ09dlTU/kQPXUfTUkX4bsojP4Dr+y
LPfnNDaaAQSuKff+I/C3palKmkL+xjUln/wTOWL5qaK/gMB6XF9CGr6gW9yPi559
NeV3l9a03ElTjYlBAaiOfE07Z1A3dYSmMYn8GCl5djmScR97UMevmBXpx1cfESOs
UECGoaZ9Yw62GjxuezfkCZlN+hTiMvUIkNE6xc1I6zm+OgWVNqoe6oF3ZcxsH55x
qhN7+ejVb4pzpOVKcoIFHcaMXb9lJ4KURt82pP7UJLkGoUM0OLgGs49CgmfiS5AC
TeK/CPujytoJzdrIGL5XV39EHS/9juCY2fKYAcLkLH8YZURf3hSH/i0u8BHmfgKN
MpAtcU9xjl3cb8dWDTtTUZaImR/IxNSTrHiugwCb0LAHaSVbWiiGvD6N/0FgRG8I
k6BcZPYKPcsdC/Xvh/Gsf3ZdyNivwQ2eLHx/RuUzdl0wSXXYOKFPai/sniWYevTe
XzIl8y6x0A8WnxR5xNI+i9TEJekPCw3BHdtNI9RcpnFvMBkxcByJ3B/22RaQj1oW
0YDzXlUg1PzYcikuEzm9kijiC0wOkla8bNOHHHFv1h142PnPhD7gR+7TzgUWcpO6
lY1IPp2VdSalHYsq5WFc73VK91xWUudSp+MefFjVdOe6i03R1A9pQp8LrLPJ1+gQ
1vHAQIxkscDkZX1SdXB0ipqqlpg2CvlEmLysRi8Nt/+6azDeaf0FcvSMpuGtTM6I
zssNGj4YRpZtMCuQqqkM6xixfQhfBN52xlltejQ4DF0WGiyjYy+b4HRMpvg2l13l
pUWfARXUDP/sigEvrme81ZdG3FpArrAhyPVRGkFKOoAidzJYEyEjINds8VkbR3EC
tD7nRFzWm/VRU1Jq/ymkNhdWeXVtG/EhljRH/ghzy0j6mfAUSSFX64wtfoK3yq/p
reIPS0JZko0Gi9QN9HzDlaj7eGjwI6Yk4kCzGpq3anBrfA1KYH4TLL3p7Br3M9NA
71dA/ZrrjHhMgi5vALMXIqeygqBNmr4RFiBb2DSz2jQE1x20pY7eBSA4iskxp2J6
uef1oiWip4zzzN0XgNAiiwoLMUNSjWvzg9JqVwOm5nqTwNKjhGZzliTVYBa8zqu7
Ocpi4kuOBwsT5JCzpHqeMJcjtO/ac9zD3uU5/mvnku0UADxQu8zkXW8BFKGOSA+v
mILd/2kb6JvnM7VrYRdoR1VhYWm+D7TfegNYgQOJ05eqatx9rIjG88NpTLJoWfek
t0e6ESZGfFzzQ43kjXK/ncszRQu8/UsGrR0K6qBSpdPcx0si0A/c9elW2BdE/bxY
CYmNrmbzwithDSVZv3RszqDxrAeEXsdZiByirTj/tikSDwk68S2FbKWN6Y8Yrq1V
GFLuVbxU7GGfT+NdRJv2pabkwel5bwTDmOk3kbfT/A/Z/uvJude2VRNmW8WKl/us
X8U+zx/nYCQQXjffLq54vRoMJxK8rJghamrMH7inh9jELTA9vfdAa3+FiRyA4Isl
+2dNetaJDljmB28+xeNyUxk3ip8COXmbEGurvd9P6Op7m4UslTXCLXqtF9NoiCQ+
Vkh5/atOPgbXWyQLSi8+bUbCLSOxbpLtpMeqC6uljiw7qTB0fRVmxIzLWITWMWU1
soOJSuVKk56kB/7t+IIIdTty2aWZAUg/dmEt7eRaoBT8dfUHb6oSfr5iGZQWMl1d
uVd0WIZn6qD5sh++7IqjklUptrkO84qw/ayC+B2GI2uBsilpxo7f0D/HjtZaLdOu
5TMPM7IHVwbD4AeIRnJ2RLLwbI9CVr1vn/+5AbSJ+iVj3wMuoZ7ZWWuv96HQLQk8
RE1knEV/erQApGKExoJzQDnhRVOZrbWGnWsjXSzo6njQ+x0PHBUyGxsjZI6rBZJr
uWKkXHFx0lq8Nn01E8qzNULaVBtCSqG4hTvx92RzRLYnn8lq6c7klZmX7SZHOUfw
7otfLE3jqCH5WOYQCt2pqb3+1oVMw/LJWPQtYrlzArVjDNH1PxhkxvLmQqOtrSRn
MEuhizgPPKI+SGigVdvTOicvPFDWQaW6KPhNC+qIpEI80IQgDhOhu7jscB1yArck
Jti8Y393RcW+oB+aHZgzh+ax8vmK83BZ3eoorPgbarKWnfeDRzcs2ChVhrU0P7Ra
Q0UwyV4b3OyTOHRGGpPQucsnE+X73WGk+QiQLtviLNNK0RRxE+uxbZC/lIYVTyIF
6brRyE29+roDS/CGk7sutf/RW9euic8HU77FaQvMtYTNn1/1jbwCwxq6gwCHMotp
ZhYA2ggaHpQeXIL9TC+f9QxBS9dc1DB135hjfNV1mj9e3jwyFeXuMP49KlcU/ODC
NMRNHuubL6n1iggw8dtGsndDCQu4WX2sluRMF2UozjKrN+ro59q26XZceCaoJ04R
gzQDNQh9IvuKMEw/ZgyDHPBpVXO6vSgDGFtw4hCJ/Z2jhZsx1VkLr6KivQTDg0yL
7JDY1rdZUxsUFXE3VFtkVhOsGOAxLatZBTjiKvQSjmHZg1zER9WPiQG6sztoc57K
fEuGFzLsxK8cwyJ8laj/zJFleF4WKVqRMfGWeixI5ghEqn2HLOFEgZhyiv4wuJjE
JkT6qRZhXQ+yOE1fFWlb6/Rx7PQaRmJi5WR3GsRM5wHA4ysNf2q7VzH29z49fgnA
4aHLJWD3V38xLjA17SEPcwZwZteYfgdiFH2Vi77tgYbaQ2R//As56h22Ey6utnlP
LbN/f4GB+tTQMsyzwjmghUNADAQWmakYdipAy2ciCdTryNFMoGAS//HSIZJoMmTn
vyjXzeIQDyzx6BTB/RYKz4UbUAB7cJyzVrDKaC3HnFWGyEo3BU0PejzuTQ12H7Rb
kkxu0XVLeihMumYmHW3Lr0YzUVAJKTvAHbSde7qes/ClZgtL5nGCiIQr9cScxmE3
sq3oBYcoJiro99X0WuGExwHIQroEqsu+x0Rv+SAJJoxhM8E/NTqrj1Wk8IaucItX
eex6xNtKWxAfEpC+rm/41LNKvb9fD4+HYjJgCEsM/+GiwzcWeGpnSI+VXNLIPTlu
spXJ59nazLFTm5NntKe64+UQ3gxgg4Hh8yHXMIU6m+uQFgzHTe7EBycp3Tdba+nm
2NoFuJiBJDOs4CM8a4Pu+x3CXBnICS2iZ3fvoN3CYofCVOYt9WbP2w9RtMfH3t9S
GdSOpTU6YcuqVAuccv8RiNij2dY1fw/ZwyjBZw+mUXk8O7zz1S16KvHMSoS+Gyo2
j7GgymYIWOMS/j2OwUolQ9d7rBdpcHWlbIg8X5OJg/DJO6BNpsT9M4cpSKiqV44U
k+Zu9Nr7AB/WfFyoLIRCY1VZgki0efTxaWqNluF4Yn/Q5WCNQYKdmxecntDb1lV5
/X/2UZOTGfVgMVbOwCqE28oFD+yifF4mNmYXnFC6ChwKgTYvYAA23JPbRAGNE/zC
B2E5Mlg6dFFCEjCd4ovNceywk5HKsmOaN6X1JSBCnVlu56oiNa8kPxPt/+sZ+5YR
xzKzIt18im08mX3pBV3OGMmUlQj3AlVmaYad8IkEZOR39uYoaC842fZM7RtdKwTM
NF6Pc+Yo3j/0Vrdtk9pHExMnejQUKaxCEjZWZQidxeoyh8HtKlaxAz7pD7whifig
ayJh+D6MerrsjLe7IKwWZvn+VKpr1c85Erq0kyHRO95mKnckc4sgeTos0rucHRXL
mhhVkQwOhxDld87DgRjI0RRxxJZQMRKE1eyxNMbuaL3J5urlNV8tuHkicZuMuSfe
/do5RMSxlTP/mqzrIFQcpklAETkc0to3aC2Q75OC67wsY02yWGZ2fRxJp1phRa9+
cxZQBWl/JGjXMuW369PT5Zrk+bOo6WX57WlGE8R7pmjSHSvfDJbo2dC6SkfNP/59
/e8MZZvppBONJkTD2ME/8KudgB25yoxb9LRi22+tgAjCMIse0qo9mRRwvMKRPsw4
JkAbFT6yr6946Kj8Zj9Taw1bE51tOjppujXoM0X9gnvT107ov9vejMG7UcocZvws
3RDFqEsTFCQciREDnmQTwV0NEj0rFV1KTkwMWiAirFWSLu3OBzJoPeWLW7rdbsx4
4JTikU2PerFeHDYLc+Xr/pBth96dKtZJv1S2W3cD5Whucz2pX4bqwJ5nBdJHWbF8
mqsyFyUNgJPLuJXpIDsEc0vmXHi3sVFZoF8jcjnlTpk/8AECc9huLVByO1lt+3MD
ZyUaHMisYi8LgBCELxDIZaxfvYoK6zwkWT12dsJ/eroamKR4YTHT/eciwEWd63Lj
5qBa9UZ8ZkUJqwzJDcL9Mw/q6l0JMAAoRP9ne/klZ2e5mhVbbDSRJ1cyIXP4j+pe
K2qlvSmcZwefJPKjxaMKtj4VvREhh0Oro5WsSKd6g79pwcS1Z3gF7ClhUQ8976h9
+ZgWW2ei1OYiIgrlgK0iuhKjaDCWTQupXsR+GCryqCitfi38pcG0jTVn+85j2ZZf
JLWfSpR1x5JXH9o1iduxWlwNR9bFEOqSOdZZQIbGytU1IL5NF75nzTKVY6HTR9IO
tIEPj9kk3IlYUUO7awNtRvtJ13RFDb3KvsNWMUde/HrYIznRpoZHjk6Kc5YW1C06
gGr7lBTPlCvCgXrdJF7aFsE88bDoqm7sg20rqkIU3a+yDKT4wcYHF/UGteZJwplp
9FSfG+S+d60lMMKoxJhUcdhlJ57OlQ78bASMQFo/eCObXOrBOMwnsR34uqs0xVA3
Nn3PrgbWEpHm4odysOq18rlUavK3bEVIEhYy/zYfbuOemFUZcGf2Nvi6QEXy2Mq1
CFWTucrrl0+vBCOS8IHQ45NWN8AUrdQLxQSQoFEkkB1MkwrETS4MhVg5hAyjDjEr
gti2YrXDrWuf/CcUSELfxtwr1nx8pBRnsxrOMLROljrGTbyC1bAGyoLomYmP9sQQ
nAKUnjo7xApUxOkOH4OK7/nAjnpL82SfWxr0Azccia4B0mygXFVsqb4zysz3f8cM
aYbqfJha2mkcnp0iMkKl+NCqJK/93k2mmtGIsFgScUYf4t6diJPkaTCPW4eIOLYZ
s5eVd1F1NRV4ekSmRnO7AYAa81TbIveOKCP8HYI7RszxeMJPmcxtKV4ERE+lrM6i
qpVyRGtIuxc3gTpTK2NkeKt63/PGp/TDfdZiJstddtpPttHPM0hoKknGJEWH4AGc
rPaPZsHkro1u6yXOyWI9uh9xfkoDCRop0miLL1HKXz25fs+zN+cNThVcAmH7V2OV
J+fbnY1M53VzGnFDuz0396MsuUA1b42Ji9aXroQSn1dnyCj1I03CBy9XFDFFw8rb
iPOUvqp1/+uMMomB+bnDoeSissNIAcoUTZv6PrKF1+9bYt6bJjC+o3jR/k7f4azs
a0sVBPLteAu+OJEtyJejV5gmOxINJRfzNvuFf0RDOEVmjX5BRF4l5wACHVQn+8oz
N+5xgpvcUYf9966EDGHExTUKmrrOdvUjy21wOFfirAlK0Rv7qr3ho0yyvMjfCxcn
69zxG8Hbc4a6Gav+gKYF5D/7i3zn8I9vDWVGuSNYVMEzSdci0sMINdifxu1/+cku
vcosV7Wf232+4J/aCEyK8WKMSuT2PWpJ2A3gTIG/DzSl8P7r6DcDVF5913UfKjUJ
og0/8/ECyLWq3qG087gEAud7CXdtkIDVfkThxO4DFGDBLqs2FW/7W9cYVkTyU9/j
lmkLn0OJ6BvIfts1iUQRLfTc8G+0WA3zs86Tfbcvsi3FwNKJXEqAtOYmRO4SbrYV
stUTxMi/f43fEtCU1jAaCpPeu9ErQkLkg1i/+xeCSuYEdKF86XlGw9wYYlDC7qz1
x4TJJrJMGxNukoZbBHW6zoYC1HvaBs8jPeqyvdv2FfNvrXSA/iE5Yfq9mgBilzoB
ylSlUfWF5eQzWYbVxqfuF6Pfrz9OllaRj3bQmCFfxvpJcS1WWLkfqmUFdFtcbprM
+c2GJCl+1VM8PGtrSDjTrSNsKr50jrndNpYmzC6KfOMQ5FpsGA+uuUjUxa0NgMPh
4xdj926gEl+vNYDI7QE00VJUicc9gID4BWScW0VJXUFDw7Wj6SsA4dJa5jufd4yy
N3DKSjGyVOm8AeFl1whP8fxkrZRutNbMW5D0miPirNq5reBwS3xowXAeWtmmEQGt
l9DGUjcZ/ZpGYwxPyXm53fDvjw9QxUG0fAQu5kl2bxL+S33ptCZqPn76ZE6wxmAG
VqXxpfkTScvLHfS/bHlMXJm8YHlN2elHvFAV04eIDYRffa5MINBSiXoUqx9SHvBE
rLMypBrHCEPIGASdYSeQm06JWqbHy2S4EgMNBGw6vGzdgNaEDbizlX+lNQ/mPoNW
nlUSQudBSLtphClCTtugF89jkx2CymvTtN9xZA76f3zeNvS9voaKRCI0WGM5kHEU
+HlluFdfUHhMbpcuPLhZ/AqeEs/m6l1eoDP16TNP64d3o/D6mwXVuvM1tcTPzHHx
3ghTOtASLE8J66GyGNV8Ih/siM430JVMc+ZCT5JaEZ437wnyvH1hoKd/jMZ8cxnZ
UxD6+FoSf5hR7YJ+04qbMM4XJqqb1pTBnanpzh8QAAxuXrr4Wp2kI7u/MD2NcLmv
EAOKdwP7E6o1LeeT2uAnmyikqRxKuDDcgisW2zY9GCV5Z7CesQL3bUWEDPDbof4i
dphBx2Z4pR+xm22Yz7gfh0+MOFXyJLWCjDGUKXBvd5VFOEKFW8N6ZmVPnjv8WaSi
yE9SQdqk1VAAezFWzZ1O1+me1ZCX4R8R1Lq/6FtDmEnv8xv0rjsfb03KTdCBNVDO
G3AFH+AXod4kzEU78Zvn6PI37kchbkrtkm7vNMY07ZhE1zULnZMlDrZpajy+5Yu7
XXaFELEajfoDUVvOQ7ads+SK/kOLc90/e8GS1uJgV2Wkvz6oEtTN59NLwumubGcF
+7UhGPUMgPqMOQ89gbAV3HTodOzoQ/0pXBMKX/NPfA7ubtWuSGnMy7DOQFEZ+Gs/
H7UFsrykJlxnRGAcZPiPeeeapHPtorJ99PH38O5dcpMc6yTqCYUi2bHPK7k6Hbtm
QqNRjqNMUw8XtmOFIDncxfjQ4nkP8U6SR9tzI1u449e+4e7c+RR3frlmdhwW8oEJ
/FW0Ij7WfydCQyq9aQGcy0mlW5BLJ3AgC4VqWrhAzhZeC595Ncnq6KWI5XrAQgdL
5rmH03Ipmqd4WgrCqj73RIEbsyBdi/YCKq63ego/0iNcwgP01J9e74w0WCGTj+7q
A8JtpsJyMBcwgTsTKfBMGm/NBQx/d5o0s2OpXgRtKul4JwE8KoTiDWDQYhPflbht
clleog96z/r7ZPl+Czfwo0NLJSA1OLzfohiu0NsEIQK/PkCXdAaPasyCAdNDcGwi
/RgqjYhGMsb/OySwpk4rHNKwPcN+jpIQhmOaQvaZIeMwnlAVLwOi/N3Oe1zQ6EY9
kL2+Q6e/37mG53U8OVR6VptJcpG3FeFPj2p1sF0fuDZ7Z0OGEh45CPvtmfNYdXXV
IL7VyTQnjA3iGtJSrjPqSQ+Vdaov3zgeAwOdrRdj64Cbkq4oIsTaa6l4q3K9UyhJ
G56lF0tHURMz0qxH4QqvLPPNXBbel9XZEmMJfv9ZKZBsAQCnYH1Q47PMwMcvJPCy
Yil1aO5vTB2o8c1qzjKsfjXdrAYpgDremNAWU9POuB0DU2WUd+g6pNN9R5eyIzc4
phvEq802lxhsTcTOlO8LL/bhhqoWzFUc+HfauN4XwOo6wv2qV3EsxKKbPkI37cTI
Ykmrou07bARSljERWQB/yZGsf8LXekYAvaxQyjNFO0qT92V6Fkv0mEi0evuyB4/y
vXld/iJkATL/S4+EemjesVnyHnS0GA0heqXN0F0CDNEdV0R5gUZmHGdTmXlfcFmy
iFX9jpvERo/VRkLIRTCRtnGPZdCBWZSpFmWHxz960fO4oZdXweLZbOy3orI9ng91
61R4oT3QkY8RPZKYoYf8hg85jHcyE7xN4ukEaug1qXFm7WHo1rZxbH7c6kkiryjW
NWWTqUIO+3SGmRcv6GsD5ksTXqX/KIeYq3f8haeNe2g7bc+r40OAUIBS8txI4lhc
zGi0rMaEMAca0ZXzOFcMt+mBdmLQD3Xj6xD+Q67GevxfjorYsdDxfHm28v1MHOKU
niqJHkHV/wiahR8LYBV92l9UauSgu73350zyueSOdmvy4OS19wk3eDmef6BbooYq
75p0rfshdvzyYoTJhCkNVk2igs8Cjh8FUQ864XNdPJZKx4DuDh7K/PX/vAPYYtVV
qlyczD3M66/d2N+VQCj+9oBa6YRYAUMOKFYgOomjIoitZ6F2uXmGau8nYEbU6cQO
j0jvBEsbIM/LA/J0mn5v7x7bII7QXHQjXjeRAnxqgdd7Q6dUYrJr1emuSAa3+OQh
lvIEqjAjvFQ1RKifzcB2prk0GQrO4RjsLMKhpputYbwlwV+PA99goEwXqizfBuCF
HTyOVsMQgF8h/Tyh8CmAYRbW9A8jwcY303HgKzwYq5oP0Tm+ZSsaKl+oD0mg8ioP
2QvMC3sgp1VXPiJd3Fx87Pw4B6mcWSBuHwVou8HUsjF2Fc+CkKvkSZTpolY+XX6d
9ptF9wYiv2ohZ5BeeV1nAuoaFaLKyY9xP3tyrtl9a1HgmB3x74oswrWG1VvOZ58E
3/zo08OMkZQa3F2zJTse/igeo5qEucpG0OsQeeSHTZbFH5xC7YPp7d+suDo+fyP5
9ekPVwUYpnfjEMiRiHJLEG8W1DgZ8iwI3hUbzOyK/G5TBzZ6uf9sZ0tcMgb/4Sqf
VMu7deQPBzQ0YB3Zn7elE8GWf4xcOP0/DwwdZ+O7PipDncRkuCjgajh9CKHgzRys
w8DzQ6vYKoQLoH339UyS7HsGZY393WgtbDUFub7pvQO6cvxoVXsk+E0CiLbKacod
DxZHSu3/vV9gszSQvqnpfXX9RD7+yq2sbO3fe2YTYM+jiA1aK/65o39mHbJolsJV
fY1IDAW5m7cdre+qfkDcBRQdIw/yuHBiJuNDO+7DcbDLE1N2YKf/Mj/aYclxF7NG
EzzrhTl16hROscTMdKYFMRRDxXiug9dTw3X5VurIpC85LeodgZxQT56eiT14anFD
tnjGgyRquj6VKrbbPWMf7E7rdHCLoBceaGn+BvvY2tMzVZ0a2EKy0znk91+uLkmE
8Ab4r9MekS71KDprHVQqKiM/dgMYtWkn65erUKCGbA+RlzU47TR0Znj56cfyMnG2
5AXhvh8PkTkG75EJxfREkwI05soLC5t3dLsI20IHwLdz8u1p/db3as/kJ4yKqEGI
M60Vr30tLmRNu41dbIZLWFMgZBgioGZ6MqfBOEuKSRSW9sFtqAxba0H4rBSPTczN
jyuxH6rnJ0EZbxuqxCE0bQisxTxdMuYeasR2KIljubIWarm/N3Bu5yfyhewE7Vyt
hGNFbkNyKv3hzE1rID78VNN+yG4N+LYDsB0Q5/zRs40GjoBbqrfF5N+MBrfFsTva
l3HsG6+U81lbxSxLwyt5u4UG/uIfoih3+g0Z3ul1z5yIqzhp1aQ7J7Kio8i/KwQq
0AAAV/GEffijR6BwLWzCPLmGagh8DOlHZA3VSGSaaryFqRHc/YQA0LdXLEEAFYXd
d3CrVvjQ1bJCA+xtxkXymvfM38kZkoV+22b3wBKuomR/Ybe7850ehbcsnePhoHKu
U5N7u+seFLNWJB8goncp4dSL6gCaDbRPB1BnZlfQWULS1kT/FChXVm9xaMzBqC7b
GMstkLEnOGrdDbrW9YjqiI7jWAbdwccKtvV/xgPwE/llY/hOVhRBC8cAIfFJpkOw
sPz2v3G7qdoKot7GtWT9bozrlL+GX7BEOEhUYXUO5Ywmg9fGGBp7Kg9muvYopPQ0
SIA0DHQkxTkLmVoxvF0A8ehJhMRzBDPhxPYygnJChYZOLGC3k2hZQ/X3RAJ9EaS7
kA4aQNFq1W/vOQOJJS/MMbVpzktY8kyzXHqHS81pDHbIAtNuda/I14MKiRlTk075
tU4GW1tg5CFnWSUzQ+0P3SAQzivzNcY08KHlfIKrm5GVjfnY90PKn3T/SSm/14LO
D0WSsVEYOfZ5RMNE2TIMlvGHvEim1Pxx2mqbocg3jPU1J8WXRkxIKc69ZfLFEmPE
F7d5MHY3+7JsFjn6bmk4dkxhNqbRoh5Jdf4131R8c5aj4cdnAzdvwhw8x06LmIKy
4rg5/JNRFEa9h9Qerhy8wgisX/cvXW1jvgVYpJnI64fZ7jOlr6dzkMLBZIxmrlgw
AFqfm+sFRyl3N0ITn/M0gU6lBa+ARW+edkQTfixVG5Xb1ChzXgxwGmBz5n8wuX5Y
bJpXsEpP6kO1PI1WIzAtBsgWFICDBmoFlOr8KxT9HgnnhjaVNw+JpztRFyedzCrA
XoBIRLNzc9xLw2z0RqbLq+eM+xEB4zHgV0PweqgPy7SWlI5lyDaxOXHNeGnRO4X1
YgUxFWeLhOomwxDhVDe7J7keZz7OPomRef1le9AYSj1hcnZ2lnN7LsxM9pBCykUn
8G5hD8UjfS+6md/3PePlBi5ysVksn6MZd3jHZc1IlWWa9+AvzyX+ZLSZFFcE08Mu
YYCJm6SagScEOZeBZaIVjjIzsCLqidNF5Vxmmkxco6npk98JcLBRPA78VLAls7o9
8Qmgy1ys7k7/BPykDUng36tLnCc43ZY/v5yk3pMrsEYpRXJyzMUVO0l8GtuHvKYN
lI+ovN/kx0qEa5AWQAVMXYIpKk5rN/QY/C2kQKNpLnm28JM5SKB5gK+G3i+xUTcj
tnQ5UmpfMZgyQAxGqG75MJL0k4M8maiZYPYsSziWJd3HSrg6L5Te8z6h7q04gDVj
SCaXhV2P1qfYEoHknc8eF1zloO9lCjb3lpYxYv+DnQ74b4kj93suLVvJThQVBhV2
TX4rjuyYiMVf94uPzADqwnKgGOkih2wcBHD5F0V7W3d7RWMEMS9m55UOxGsfxMEw
CyQnphvdhUqzqmhYbWgZIdnE7gwxmgO7mXqlMja0A50KBPd6TvfWKTugVRESY6GO
q4mNwYjw9SqzN8AO9yOOXgUf5qk0rB/0BILTlGDxBkbsNGbi7OWStAYXgrwuAcXW
gGmY1mMk7el2Ki3MfGjTksLENHyIVj694njo3nLieVomsE1n3CtBF7G3bpS/55h7
J5CNvWTspRzkuv+maBr4qdNEQnRX3o44Kha/tUOt+3eEA2/ypLlv+WvSCUa9/wBs
fSfZSjH/zdJ2ZhMF8TiqCj3NxCbEsHbFZ1UQxj9zm+AsiBMClt55P0Mt8D9+TskB
XcmZeTVOfQP09pQnsGnp3fiMl/z7I8U4aX5v6W9+dThSNhiDQLcaTOTADce7HSiI
ul+fFdUTKvsaa5STYof84Ep0RD5+VybcYahCTLGG7hffAojGTHK2jNUPFtEA4aQi
Q3nesuKt4htgTl84YEU21DK+IdzuK5SOkdjF17m+g2RgRmynaFk0iUJ2v5Y/o508
YfKE8+NyBc9lLl6ahEc/AozmaWSDebn8c9O1tjQC1XkqDJPv0Lnz0I4Q8nCVZe6b
xBPCSk75eaxOHEgg3Mvnpo9/ZshaT29jtfcJPu6T+lgfWSYKYuwvQA/NRu1+MIkc
m0svl5G9ggArEu6hYjvYeCgFHeh93cA+146RfOUtvGUYICx8yZePtzxezp/nCNug
U7uPnDyLSBgjT9l5FgT7Tp76ac99FE/QmaZHW4yan0VJu5KbbbadW1d4zWOLx+yN
Hp9OMGT1E1sjecIovZOm0QYkaIjm086d6SKrpysv0QUlPk6WC+xO7akUeaqVO4Aq
JwT/+R1N3mQvKBwNh+eFiBZvyllvlTPzxNK+bI0eie+hETmOkbsbSK7Tkmbetcn+
7Pu8/DHGQ8E5qJGO1BYvQFw+wQaMRAM9c7/jQAWKV8ofzIxdtXTHxPhUJ5sZH2vJ
TTeAJ4+nwOWtJt9s6nNK2jF8iwQm+pH8dPMpjPKVMm8IVGJSPjJ7nT1yr4d993iA
DM9oIRy7FOEJQf3ctWD6t7qJTL9Re1ZNH/aI70CvOJjN5Ja1jolLjk1EDAxK4ns1
X34YADvqijAj57zdQU6S2rm75y35/QTjaDfsURgPstZHS7D31lNHeB41gXMZTz5g
2hTTgXHcKLm/1byKHOIlc6vXiqYkxubgA959OrPnGVynF5Tk05apt+5mVFpwnzGU
Q8Tuc1adaRDLsalsQ+9mEzH//3VQjqquN7TuKfRA06W6zUzlqer3KqE5T482/G0F
SOXheHDPGvf5jo01x2HFKmsOZQE+J+9nQ+XEyn2G8wksvzaewD+uJXesvXnwLjKG
vyh80N9PPPi6ZxzbtznnLxszcwJqEhDreC5obILGUKp7xkss7xh3V/kcszHBClYt
iYjlR8l5N2Ytd/8cbu1R1kf9EqlKDsNLXa1IflSKIo4jiOUXbM12/8cFBWrttjhM
Wrc/703cjImeNMaTQs2Qpn+Z4QAecLaDBLbwFnpncD/9UrZzUGkaQTlvg0V2DQ6w
tcqKuux45MLsemeAVSLiWTNWbfmWvt5g5OYBzCUO7pkyLi089rcyYiz+uuDcMCPK
zT897c9msVkyaMy34xOQpRZpq6XihC6sg7oBoM4ASUuw7b7W1SWGP7HbOhBrI8oJ
AnZfmwA03lFtbEQqNFNdZopk6Fc//+ZvGXfX8/LdJ7Lbm02//jME+gYAwsvwZ8bg
ybir4XQr+uHqfWjblOCMaz1crVsOCP5wVEH6MsufE2KVMOF1I0mnwrmlgVRNRkgU
qIWFK+batpSv0uXRfbW96iZSCwPxwqZ1lltFwJ02lx+oJ/KJYdbjfbvZ1DGvpRSD
0h7LKrZy6o9ZnbTxDc+TD+dn/YKC99Rj14cEMkYc3Uk3EwrWhhXsv+4gaHVPQ6Is
JaJdzpRxpItUvRHsS7VjxFtJCmPjB9/GS0yCXNEhrKDzfI4UzwIBijCCzYw9WqAn
dPc+0Sid0+peUhsDjyUZq2BG553l9wD2wA46+TqOl9xTyefrBJ6Jhl0sV2CQrmgz
of9paR+GZJqIragjrLFdD/aAmprirwet8FWHHMZcqhZWd0GQ91QJFrsTLrnfpMHz
Ugek5RB92/Y4dbuXsma9F0Q+2oiKYZ4LfLjOcVpkUq8jMVRKfP2n+pEj8g4J+IZt
L1JUu8R1Zhr8m8qwPopPZfgjWS4wZjGi/exRXeQDhj4rVYFHt370mctF0EPAFcXL
RpwJ0M3Xnbl9z+iF+eY0l9Du65QjK4xsep2oFVAthngfaT56dV+YBAihYEflvgCv
uhpwChmvFqYOKnFxcVceCzE+V5eCrZUhlkj2F7v3T7lIdgwV5ma2+Q1JE3K+IsG2
ov+ORf0JErs0ZgSUOuPhDQtdEMAZLMMTcqh188b4p2By1iHjlPBxmEMSYd2wvi8Z
oePvDK6O8zL8QuVpo//Fb+SXnpRzD3ESE/Y/mBXewkpXdIljs/QTjsJgdIIlZwxK
3dmwthB8mtEgntag4IFBFoDG8FmsCbHJPW0CzZKSEv3y9EWBz5mSrblI4xSBGfQf
BDdW16kkdNW469BfIR4v8zv1bTjvPsP1Xke7ng07EOJgP0Y5kVmhtF5kDKxxYTQm
nfWe7Jq9RQRN83hDLBTZpYTfZ9RVV7BmdTbzGguUC2nQ4n7JOLgWANQqD6ToBLRV
oqnoF+yx2n9cMehU/QqtHdcY83CERINuyFCoJ5WzSGwaUO/PWwHWTZR6RU0aaPEt
yMO18RPZDq1q8En5jmxXb1S6qNr1+VaRf87Bn8PV2/JqJx3H3Y4k2C3Zk33+GdLj
9zdEkfn8KdfD/pRCiWTrWoR16L0q6RZA3/sLgL2eAXx5/PfZjIDXLsGoEOhl5bIx
tXvPswSMsl6cx0NfdbUmgVXLifV+qZzP2tEgioG1m4deqSCo9YG9Hr7Yhpvp+2KA
obKRZ8ZbFoUjiBZMfb7GyQkgzdkGuHdteUP8feaKejpqN7cD0k0xQY8/Q5OwtnZ2
VoTsEKRMn5bRMvxhzBoaLEfRP8e/bjEWKuSsdfVEw0fPY+zCr3eG3fsNR7po9w3h
62BHNhNXiUtCchm+GEin7CT+lTxmfOMizZvCqO9Sk4XOujTsrm69byfsyoAnlz8a
Zj/rKj8ru93NzHurHxZnmLhVPjcZncqYxsybvg8TNxNCMw0fOsCG2PWYUW5fSH/Z
3RZ/kS4ui2hXQEfvWIwPRYeYkrqUPJOmuyz9vLkltw/8igJ7zTFwPnIpIewL4Zn1
Y5+YB17zFAL2cHq1ky7+tEhwT/hVTpeOKU1YRlT5ScvHN4rsgdh10jvgLXVd8HqZ
MnJO6uug5zys2Hs7T2KMbfgQC/pvucznlqaoTWpw6qmyZyHV0ZrEhNob/seLDN9H
ze/FYJ0FvKN8x49dKQrC2Dis6ONswOgOom1R3Epu6tIjI8V+H2JyTyyjDKb/bTEK
oSZs2sY1nPd02ovR676DlKRIwQYdD1jG3jYkgYww25TcVyKNctIsG7AGUgrhnqfV
nETtabGz4qb+YyH0bjSA+v4kcuvLBcUCoaX7JG9NFd+mV0DeGKnTzzxVHhKcRqmp
OXEHgLEPJ9jIxKIYX8Ja8UkUKN3S8g/b5QGJDfkZHJY3uEgYccehbeh0zZH2c+xj
w956h+4UHPMoKhGPGvDrN/h/dm2vYr7dVWhmj/Ia8r5/N2dFWpoJladP6+ZlR+sw
chD808fpJRnHaJXxx5R2Ii3JYQxHIthgx5MEPakUsTv5KQ/5ZWOdAL6b5UVQktP2
6xNx0dzamfaLufXGe3A2x10je5VlMaasjk+KjOAINxBKQH6wr6art2g3YlADwAk9
77jJ2/PaR1zxAT9npszpD/RztTtFw4n/MWRd1O1BDl9I6xOdh6Tlws2JZZJWTLJ5
IA85/BMxCID27MuG+3jGT7RXB5forL8Ko9CPeF3/+ffBEKpD5fGj+MATrGUVMw7D
T/HdMIz3tYLtdWjjVyjy9cgdsHpZZ1JHbo8EojXy3AlXwEylY5j6VwvnTednI4c1
Ed/LvD56rser8av9okF6p/sBH+mGXu0cuTAhwVYoaUOBj9gEE6y77FCzUhvxVOGZ
oIh0Njb/3f9iWtECm0mPYcDRLz3/1eWUnGqv9jF285+XrnNCWS50IqO9IMOsop7y
pc+TlH1dWIuZ0Fk3LnUKIetKfoMk7XeiTvSXEw9gq+9MCYSYW6DaLcjgLkW8bxD2
UY+CDTMsoiRmmpxOjbq8kUZ9FY/bUomxEwOQyPYc60MYRsyYVcHNcKZllacj7uZJ
A+SiPinqmKuwPN3P3QHWwwSKIec/pTSWq+6j6Hag0KwqsBiovtv9Y0ZPfosfv89c
B/GVqReI0TnruANAA/Repz+veTW8sqXJc6qZGEImy6ytRa9pPytkenEQqUIh9tZO
6nDyDNg4WL9rerSE8JDzOh/AbhK9VbdYNHK1Ktzg0VUI25ubDjQ4rDpkqlwsWLn+
U958mdyPJm0WOXpZyAbuqWdywEh3UB+wowiQ0ChLoFgIukLJiGGHfUoF8RNu9v5f
6wfbXrTZkzwpHkYGI9+N6HrawsClIys/QmKKLzw/A1j6U5WY98WXklLWH7tszdJX
WtvHX33eb6Z6SmrugUSFSnVy6ldnp5u5vJ0lo50fxZ+/CqLtDJtkKfOwTCgc9GdR
AeNA5dq8bRvVFhsSVXifk41bfMbzKpaUPd+/9P7uqQlS4xYsZwAZGGYIM2KFA74v
RfVGDnLWoMkBnTXHZa5cKrklaxBfIKgRFNk6Z2CPVv0VyMFiEzkG4jmFzawjt4RS
LBek1onc+bkO/B1WF9pPvwRnWURAt1gqNhUnwAwO9hrzy/TTRDoj6txM8ruPed2z
L0D/PdXxycOCkvWQm+vK5mGnaZpNMfQIHq9ZQ6vzjQqdYvNMk+89MLpcGBCeroXc
kJJQm4ShwBuIgr+1s2TmGBFB8DWsJAJgW8wtL6JxIgm0gLZjYncjcS7d2NzIqiWE
4GAzOumLvLDY0zOvOLnvyjYZGReBxxQjm5At6PzmnJ0bupOfOOk7zausEBls5EyF
OizZR9/aqqAxzQ/7D97M/4ZxUrZfxevKSnTEV0Z5OgOPiMY/VgraJkuHiHKj1biN
VuuDMx4tk8fRPtkxzIYD4fGRetQpCNyP/g21+JfFvPt4PPjaBp5AH9LFhy5WTC38
aSb8niJXVzLJu7mzynw9w/Q6pRfniGJ2hekwUEvzsRnYGKzwqSfA7ZSdceUab7Eu
qDt3bSdX8l9bIN4yBseJ47lIPVAlycYH2wES1FDwAh8xIS/NFk2JRKSvGBAGCkYZ
QLBNq3yyWD7SybxzhVjpgHphRyhVJD7kcQ8mIcFFJn63VOEcxB/bhLV4R8IMF94J
IDJuJ4qmrX8cnrgNUmklFi6eINGRwBHBAfVmiEbyiTXGYGta5BnXlwX4XLS7oMUE
5ou95c9nQiLmVm2Ej5uAO528rSDm+UkhhGIW6MBOJVVGYUTuR8zFFU70Ach9y0zQ
X1Y9+KlKXpphsF1qZg0dOpbRBnjaZcG2fC4b+fTjWsh2dLmKCjJ9oz8moM4EqfoF
lWCofpCc3Wssg4/vvH4bQQR+BrWwJxQS7anKYjWxUPJfJr8RE71e7MKZ/MxIOeeK
vUoN8ui0JMei9RHzKa7NwjDujUHw/Mkz8G5EkuPcqPdbLlCiJbMxyTqyjDnPt0cz
LaMka2VWO66EaKf7Iaih1xjEIhr1DK5kGaktBVbG6q7TGt+YeskhaCd5dL18Orzj
Vf5O7Ei7iix58CdQJGl+LXeIniJsS2KZM2n5BOphFESjGC45KPUF4PRnk+08lkiG
8zKELjZCXEfmsArB9xMZrKEIJ+IMVG/m878ld5dgE+sc8BLyROJKqemWHxqGSBCc
R9PE6075l79muwszXGXGig3xyIlvSIVIW3ZotD2wwbNIG/KYdUOX1U01Ac+L4LV2
oLFfUfoeV20w5vXc3cPdjDV3fZwblORX9MhT+2xSn/olIRpGmaf1/Am2Y3HKQDv8
+wEGTSfjgFnVT4p7m1jZyxv5haZSPdj0ImYUgGf20dlgb1zJUQDNAquYEjBtdlWs
a0CO6czJ06UGskEIbBGryzVj1qlnitsePwwVa2xEEgG82xQu9SI/5Bjq5THHmLTx
Gu2dullKlfOkFWbIVO25EPsahpWwu/SLKUZWe6aOQBZtfQg3rkuSh/YSV+jaKfmm
6JMm1DdmHGqVhVrzMQYAP4XiU57MH5g/5RgTvqB0lfD+zDGkAbPO4kYZcqVmZko5
3R5OB1EyccucpKfG6CEPYGL5wm27JFPCJgNEpoSCI8Nztf+Bked1BnfQXA4W4c4+
114rkDV7khgTblhK/L4SDbtONV6IFPNNQwav2lPoNxOQ/oGOezdq6t4Eu0JMA61y
jTtO5PS+Gko6gI1T+EOQ53eRFcqSOvMLSQfb8ATtDqyXDzg6CGsHy1fl7lrTjRu7
E+IctkRncPQDHryMHgicuG4OyJTCFv7P+BgbCAz1Ey5yNjCxot0kt6PFX/TTzWLR
YjodGARhPd5h/H55mGTexrA2UXCDHV9BbWGfrVx1p/VSc/gKxWhfkrIk+WEa+Opf
s9ZOxYMnTCtLP/Q8LJD+w6QiwwB/Rx70e187phqi/TD/wSCSBdp3LBL4sfUI0Gdd
6c/Q9A2KA2r3zLi/cFQHWNOK/zRMFHOIMt0jtaF4JUm3s/dhR+uQzM1+e2QWVO1m
Xm7PSomjGQj6gj3v1e1h+SvGkNermoyy+NRpFwQrTH8mRWf4fuTnTYhol//C0SLo
nNA6sEuzqTl+zIY0inHG7XpS3SAsVxl+8W8mvEgyYB9AQaF2Vk5P3/xMs78PJwtW
xEqGvIdeD5cre4v584rmGAKUlOdeXlMf3sC5TLABZYmc3jUYSxhrtjwWSTDcd658
d28447899ej10wcss8MSB1iI+HztFfSiiN6i4WBBQW44eEm5s4qcDVg3gpDLs8pa
krSgNG64Sm1EsOu2//OXVfzGwpp2Dww23XFmHxcT+9kFq1bsrbeWJB40ScIJnO2+
JKR6plMNDbnjKAeS3bI5npGkfVQw94asFScnOIjHMPHE/gzMhaoOLO32lZXktT7H
ytwn261m9mtPjmYMxS4gzheQ/cZrpUcdmeDlR2kWuVYw+bNLJG1F8DYvNbT0Xuo4
Qx2yMxbMHA+kf0ZKHKRCnwtJJOJ83BngZdVRLK1a0W2kpyIRV032sXPl4VBMbkj4
SbeBvzpTwah3m+XE0Ob3LD/xCDXhgKfSPPGpmrSNnSCAsjN8Z6uUFgFHD7IGVE9p
5vCCn4z5W7yBFN8pnNyCRK2G1if4mOBSmhuCAZg4nsTnQW+FEb5PiYzr7wQ5tZ+c
F7gXcE74lnY+f0arFl5j5RTI1XrZkuGwqjyvnGUOgRzm8eQxaOOSBOGsx0KRdq4O
/ZJqwDr4IpZ+9dgoGgRBXracxJvTYhhK2jVl9+WePFJVS3jEISTePXhzndLlfoU+
T90vUcdYaOa9O2LTpVrm/Na50QOq/irxzjsD9sAWfu50/gf+ABrtGWxizB5qBKIb
g+Ha7qY1D0AS9qOuKBLbqL5HZF36/HWezMDaIHCtGAec5GB7ayD710oO/UYjpWXp
oFXzIg6+JpSw783pLjRQH0l8KTdKHMAGfI1DPS9ugtgu3Lp3NPA8cg/GgIljBWD1
pDCnf6/9lHkqO2bALJjNbnfzV4sDf6daC9xPtLFAzU0/skVUA4A7SAC1zTFcvzjN
JOb9rDINiMeLve1VSN9FT+qdo/8UciCB5vT+56cWpHeMutJMEfvaEMIS8zo30kO5
EvtzrU/iHBSOUk+YnecQlG7Eg4JOlyYXwwcQsxEAkUJX6utAHEVbzhTNEnu7Uvzy
Ogs2IeK9Qcc49w98vkMWo544kDpjraCd+dGpkDS8hS5hPO0UktknJIDqheMqYtX1
uwL2DUOaEyi+rCX2dFeWRZoMiwojJQcb8xj6wgbQ2JLmlwGZCOOxFGnb96Du/462
f00IHJJajciQqA8WH64uJX8i8ZTUY+clJ4qLZbihpS2Qc4LvHx7j2DydaU8+nLVL
RdORhLYqa4OgecQ70KrtTr7iZ/LJ71swAA0mDIbrDkbhLCuunrm4Hoa5leAVo+o6
rpmrvO9uWLa1lxddMJFSwSaOKWiHLMPIYikKEWONH1aEylRXc1Z8WnA3Va8zPsaK
YsfWBA4wHvJBI+WH0D8TuxmruAo+w2jaG8xQv0JonG2h5fw98rdY63LEc356Or8e
EbkSd8l9y1U1d2DNJwpbOX2eujcFKtT7+hJYTqni2Q+0Ofl8TbOjle4gNue50BWb
r3vbr8GLbA8GIY5B6I9X84gU7FkWtoLgn2enT5vny9lGpTe88r8uOMGITfBT1wqn
0y9+KyLIIXKzBloKIFgM1ob49RE8SgKq/RsGMKEh/br2HbufTmWjvD4RDTTPhfCd
WXa7oNzF+T6yd9vE7n6OarXniT1K9YTmNhgcTZeNN+U9/PnbKIuk8hcO9rIcGBzB
u/olpjBdWggyubZVyZrqDrv+VcngI/PyYy3XkavmlBhCCyzMdvutK8cnvWP/TfIp
KEmBiouObp8LOE0lre5c/m7hXWjeGCElrGMn5Ipx/sLOpgLn6gTBhTPuBMFUI97Q
dwXNoRt7O/5kQb7rh/sp4B15c9MY+1XwDaZLj714oLRxyWbQ7ktGFu+aFh5/QIsa
3kkAsEpoVzuOeODF1nEc7VWF4lQXSYkGUeKyDDjmTRKPDDeD80Qcn9rJ6kJoCdoy
+4CDX+ukBRIyUOHslI+0a+XLtpBKzXFoVs+OZnmnWEnmo0RmSUql5pPkEThEFV8t
uHkvFQdANweSEZiCn+9cqRMu/rX+bOC6hVIwgKLR2u98lglazFDNwv6Pg1mNYWnH
yhPaSTWnEDgs6cWDl8NsDT22sf5/pF4zoR9lgeTiJ1xqAsMZJn0ttwltb0Fo0N/R
UulKjKKtluROVYNNhlqVAxxQWCvvQrPsVxdUAiHOESJb+XdyEXdlXdQwQjAclMgE
j6/J07x+RyZQ6dIrJvMuQwmrmJkOWjrTWi7Bxi0RSnPdi64wktp8freKM5bGTu7Q
erp3tRVPM/XDyoQ9OPgfrmXZP6HgTqep9cDcwkgzApTwBacllEvEuo4oVhglccat
qkH4tWqPUxWD3I4rm2gGe48D0l8pufX53fLBQBqXOKFKIn9Nq17SQ2RltkP5nhgN
1lFCHAAvQg26t0t/JNFtf7PlInVHRCdZMAFLuanR58vIs35cM/AdrFIleBcIXKML
pL9drnWl71FAypxIqAEc7K1UvvmFAadHUJ5Wc3A7GxFvc1bUc4Pw4Fgcd/xyT9VV
nGBLTgduXB3JYpOGcd3khzxRJDkMbX1sv+dC4NnY0AkIObPXsb22Ujoy+4isshq5
e2b8U7zSQ47goKE4woGyHNzajcEoXRSBaflQZoriG1+ZgyYPW+StDQmhtjekOEaD
jxaT62UQj+xya0FDaUjxJjAjnkThaGGzjkcvkTeWBMxds9dZmxlsYbn6GLm6XJ5x
mpRii9+/Ruj70KlHiVPgPQt8PGvc5rGq+i0U3MxgB3PvW2SVuTrdGxlhQ/5CDRsn
zK3B3ha2/T1L6CjjK/fgfbtRKTOiSG79aKXHvuOQDyunb9Lc5iygEQvUVMc3nsO3
cFtUHSo2aX5bG6LMjZKSOHQbdFM6In/ddn53wpPnTOc8Czou+k5FJtfdUmRMPpcO
54N0MM4s+mgPNEmAB5qEIBMMdA5VMZ6qAdwx3U4eEA+5s7YzlXkPBRSLipl5GXSJ
5FtBkg4F1BJDat5u/YHEkhQOHzcCjET8draqiqNuoGsSHuFLWeT71LUyiMqK0fDX
7sqFEEjT6KHWJeJXOcACW/kF+Pgv1xpPjKjxK1O6BBNE/+kKJcJWv3RwBwNEG/hq
5HyQlwrqA/86Amkd5eApVx3VChMWM8vZceTbZHNRtF8Ue13BT2qJiiet42w298qE
gnC3GsxSXnDkFwGBEnFs1B7C0rytYFOyzdlO8KA3m3PmyEJXgcoX2rm/cGJaO8XR
Do1FPvcUXIqPvHaxE0fQnI0mOk/koLVwc6MZag2H0h9v0FSTes/Y92B1jK0aFLLI
jgWvb6Z9THeIaxkP/Mr8RMJEAT7LFP8JT7SVcxz0BcmCmM1dOypj3jQS9fXRPXao
CH0KA4r5XURS2Y0myjHtod+XslKGnGrTH0Jvci+8eLDQPR9Sz8R2T8zZsdcOixy3
ZrXYDAZuXXAF7ZEYy/OfgQC/CFYTdJWQGWYhDp6xBVsRZMcjS0CHtOBKJe3LL+N6
6zf85+IdYFiHWugVZUud0L5sud7Lfo4GrA9K95PVQ9kusps9ed2LuzdTfW+xTkQg
3hzXb1DFKFVqQD5ANxxR2GBGkyNJy3OXk83MWvpziHSRxuD8MU0WshRzoMQKDYU3
H0Fheg9iUxyMDPU/Gee4oo6XOTF3oFBFtR9aw/fuEpGqCrVwxV8foPbz+tNNbjcT
o/tpTLuBGCYPZOGVA4xP7gxpMW8rZcY305poKoMWy1znX792SEs2FCnNC+Hy47Zn
adb/h8hlKkxJrki+0StkOWVC3BgInBQdcB6B/Wka5Km2K7x/QMx1aOrgbvWRFPNN
TDiEq+fPvVjETSBtJDml7exOp43nvNIEcgGcsEK7FjMtBys9ulA+IVSZkJyYtiPj
TW9VNnG08wd0Z0/nlvVX3O3gKL4pEtoD4lW9OUPUYvOPW25aKbUslh6kRnMs7irp
GbFJkV5VvFlwXxkfG9qvxHTW5xdVLznyDMBVxybFF2e9jyiY9+ldWQKGaMpsemRU
r+6hJZ+9yFb6BQK5yTY3DnmJ6rUjaB0xPd8F4pdEFsNFmilGqRmUW64hP0x2Kfy3
ngXRdRp6ap1rUfxN4zUuJ/PWGZKhuTfGCPG0EY2AtBQcrExG8Sm6gWP2KgxQXwOr
wh8u2vxrUAQowk5sVYb72qubVtQKX0nakaTrsTA2dRdWLzQ6ZVLJ5mx4E27DJQeO
hod8xximhG/px8lYxWIgYs9p8U22T7NZgiPNuGfEu6Ds8jY9S5gisDTjL/MHocgq
9/+rdaXNyPHesqen43M7x6s0qdMmk16NdXfLWXjghLLgy2uWmiYNy7xcKDnZRx9l
t4ae4tVIzKvs4jC5bo33CaDjlhYgdYTYTMxAI9RQrN8Mkkrmz3VUpsn1nZwJkIa9
ANkAgTEJknZqnnxNWe27DYX+iXV9tsEH/F5I94dv8/A5+8oUlfgmochRLMT3YC8z
3VNpw6S4msNsdwdP1JNluxqCcvnOAMrPHPPd0deW0fsDYIsra1EVnp8dW4UgG8TI
jNvz2QosQLMirVK5S5aqyz65nibc9PtCxVcfaTokR7KF6pEP5QSWJxAURW5asb4F
G02UJqzSwllnYUs3gMu7nWUaXq2sD/wpHdcLYqQ90guOl8UTaGmmC3KLUmiYXsql
p7RaOZCRG0XCb/A08IAUKKwWb2bwCZiiNiIvCyA6VidXIQsQQIW9tu/DgyRlsUdn
TQr1c6NZhmsbafujVuXRIqeRmDbq6f0hpveeVj4zCw9Fr5M3mmygezqVZRQDFOF8
m+Qqm+gWdT7vErlfohIEM3KxFK0kFcKK4+QbIhhbwkN2HqcHVrYPgIm0t+NSTqng
KBfauYInXpoXmDL38fnJtnftrqdMBq+v20SKWK2yufuskilDXzZVkuJDwjKgxYJK
XIyF1lEXiZB/rVPu4lu++hxLGewO3KNzihC2wqGDhqvnQpkSuMn04SlhGNytKk0C
kSyhoW/mvctSixjknG5k4QXUb3D+woDofyndlQjSe6J7K2cMRMupJcVJz0092w/Q
QYwjVaG3PoCK8i64rWeDUXaQYdwq2jn9KGvaaYYp5pImACEfGuuHLtLJ8h8vIPp7
WnuYxdd/oZ5g+MFRqXEOPPQq0SAq+l3984+NjwpCQZYrzX6DcqFBIvene7NH7wwn
sSXuq3zivc7CsMKqHfNU+bE1t6uU76yDeAvrNFZAnSshpnQMqXFhm4fPj9w077M+
tOhIxA1bIOG7JtoE/jw0JYqmSsV0a1vgHJtzxZ0VxAywnsefqtQaXCkX8a+PNhhi
9IFMPIcZK/UDUMt8Vtr8iqNho6AMOgsw30ga6rjr5nO2QrSlJvSeNS5tkWfXQvAm
1mJVXt3ZHw2EwwHPvGtNXIKEipM7BpTPmSo+Ou3dufOuJfFNku/JA75b2GrxuGPN
bPWnKKn4TDtI6F+ubp74uW406T4p7p8PMRJH6BmNtOMBGMG+zjd85MKSU+ehxAzw
dUAoDHm7PL+wqjXIjF2NNVXc0jlti3V2IoIxbjknv/9Hd1IZR+9R7fs8D+W5R9Ru
PxPhkHoO7XLpZgtRzsuBesEixN4QoIMTLVGLajLhdrH/59Pd4nHej6kshE4ccyhM
MZ7ksdch563HAYB000/N4BweLcKVsRPocXThl1heWcsJCT1HnxbLCRj72CDdcpT+
2Yg+St/rHN4dbg9Ge/RJN0I728SYI6wOrrk+mU9CiT/hUh0OVt3BKPiJ5fYUzyUZ
YXtaKOW7K9IjE0erkWQaFjqlb3qYHlM7VLGKQBHWK67v5FDay6nk5OtXEzLXYM7p
Fz+GNhOL3Vwrxkn4Rh6s0faG4o/pdXRPcEF1PYs5sOfckYXHZfNClCLuWyw0UsU5
vTddcIfL5YK4ZqXb7MhF+eMxxVGzmbabst4wtVa1XvJBF4nkFmGA8g1u0F+1uW0Y
3D/hCvI6zBInyx4UitfY8G51iRA7blE6WwINmWGOpdw8nPV+3i8hqm3bPFKitqMC
df2Voezjcj+TiGGdoNyLFb7B0lVhxLP1mLJU23334Wd7x2J1L4vFtzDVnDzkx6zk
vhkG/qq/z5WFP/VhKAkZg/a22bDaC2j7+iAjDMR9MH/D2cmhx/luD6t6vSDq0ZjD
arHr2UVJqAFBlOWBnapog3UAq/073nkPvyozedUhTdGTbN1CeiN2igqexuojOcH4
ICFPQHytk2SqZf0+yGODkjcD8Vyy1rcIjv8P9UeQSY70pdMVN/tK811LtlsKeitr
KeGgO5av8iIRlcDNrnYuXnyRq0KQQcDxPuiaA4/6VXdo96jSNqo8Y17UjMsCwIwg
ogKEa5Tcqm1p/Fzg+p1HI876hpIpqXuLeaEujjY1ajbPP45Ge8+foCBGa8Yn12gg
iOl7BGon3LPP1+ZfAlfKILid2zlF5RB3GmXwffg88tuNpem/twBZ6CLOt2ZUktxq
fZJVOdXGp3VZVrY0s0G95qBO98C6Old6HzODIUpKdxfBP7UYAiIfYbysNOzE8Dc9
Xtb01TFMv9Aego9glX+4K4UTaC0VHJW/MKluPLjZyN0DNyaceofmpKja2UpCWtu6
`protect end_protected