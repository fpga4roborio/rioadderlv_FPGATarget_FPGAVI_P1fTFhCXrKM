`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
ddtXksX2+yylW5zu6QL2Lhnb2d1sD00763mmSITNX595NcHTEkwn0zB1Dry37fOW
FufOhVzEJp80NC5qZ/+F0Vk7Ik02dIR0elf3clrjeJRK85K4e3Hoo4xn7YbFUIms
l/8VZSb14+JVGURjfswrIyCUotIzlzVYZ6gzoZwDXIi5gQIBf/gI+KxNXPaKV+PQ
Ufys/12rjO6aI/pPlqSm0hCvftmBcnezN2hk1UeXgOIuKZnogjOsf0iJVX2aOOWE
6pD/psybjbnsNB6kH5uFTA5frkzIzkzl5d9+YDm9OyC+k84E83I/7/j+rk4L2dah
QJOvksSIzN867/4Qt8qYTQ==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="MvBXkzurAa5VTw+1JJ70nePUfoQXBvZOku/SMmg4TwQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
oRtzZL4VJ4iwysPsC8SXYCzXS8Fw2gtZTOskLcDV+1B9Nzn1zTyNtlo6lNICRmmK
ZRVu2BmCc2G+fmzynYlNTnSa7C0Cuel6FYpxCBlOuk3OF2tzAmLAuDyOH3Z1Yjzk
a0aHuoCdIRKv7BrZCdALt03JeUmXKPdOmIlkVGFl8yw=
`protect rights_digest_method = "sha256"
`protect end_toolblock="Jn9CQpRhJt4rnzZPRk+dOpzAubz7omckX1MrFd4p81o="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 10624 )
`protect data_block
gD6l00tciPUa6pDNTk/+t0OO0nC/UTtBwLB41d4inuAUA3i/ALrNyoJVcBnAmEQW
ptbcNp5fxEUJjnOxnedyZEuEBxWRieZFQnkRdF269oMxMHE11IsrzpyXuT30fDhw
cHhQ/sDAhZgXBwaN/sj31bFfWBuV/oMPixMdValhebRVGq/R+sEYof1FkgsNHtNI
vPHq4HBc7EwhWwq46Kthv82O7KoLY1W2p+y/KYldm9pw1u3P6ghLb2r2kbQ1tuLZ
fUUI2Ajd2hny0b38tQJB5gQ+dQmwcIVt+oPGaW0sWJVHef3epO5RbkZpEEvGOEs4
cpsAP0wCiggaj8eq7nEt1qLgZM9nu/6i+qFJvdZxok+lNAgJFhOYwMbhG4jAZ20f
GjJRq2+gRNpADflhyzDNY1F+qnyJ9wm0UnpGVMjPgVupqyN6Z4KZt9dxVSBeZ7lZ
vXxxmaCESM8Zlfzfgi/fIj72z6xOjZsr8x06j312wHRSfWjb91DkaQ5vgZVQJvCQ
X5xAH+bc2O88hSIYsIaMupZBdYzgwcBrh4CTAGA6r3DvNLBP0HrU8XkDz0GRSdbG
7jBhLiBZJl42dPlmLmOuJ8jMQY/tlaioMaLQmtfvv1hmi8vOziKgVhLnnCE7wLPM
ZhFGPDxyP4RQquia1GD68OUEW6dOcO21W2wNIcVCbFXPyrGLMP9nIM42Hsc9jvWq
GkNdsOMCmudg1W4SrVLB0cAjaSFGIE+Wzym8/pEbSjKUjnCT6No1QBxPvKHDwHi/
hDWWZC+DB5VS+DPdRZXs21bGgEDAoS2aSVNCuDiyzYVN9lrH2OVIeSZuUoI+Isna
NQ789U71sM5Lf0wb7JNLjprNwogiWdWR2fj3VXtdpugwjKW2I6JniGDv23tFVRn+
iCKAz5sKFRFrTdDF35f4mOW6DbwbNw02LmBhgLY7lg+Kp1TAAzZSwB9yBWnLTL8b
w+gzCkLWiXzaNalUFQc7mp8iCZTbSUrUDEwn+jfgGVHOFQAbG/Xde+OqXOINkGic
cOdefCKioZAmgpIxouONJW5FPJX5BSVCluuHUQm5up95rdV4lV7s0Xhw/pboJj1K
WTzKPKQWmrQw6NQxNHeV6/SRmFxv2gyexb2PeLvpoqwl9NkCiTZnlyJb7V1qOdRu
7tjHcGJBX0eGVdU3zbzx90kFhjiclRcikX5meg9g2uVODhOQC8JKz2bqgjesUFX2
el4mQ7p6Avq6T1MzkzugtA0XPSBq3PMBUaSOV/aXx+gDh9ksnqFkJQH9c8Qy2NCV
plqKjKn4Y7OBO+hQ1JH4YQfM9QxaOwLTEK1LDFCN7MPUCbH50lOIkSbDbmsTj7tJ
FaXtStHRzCpUFTjtTJ+ybkF6df7tEUulnDadMm0QC+N0TczcvQJjr7xYAEDRQmVN
ZFG1Pv2Px9PmMZTnQ//K46Oe5p/QySa1UFJsqwsRr72dlCbCrT8lFSDEN6mK6wc/
cAiCol+rWY8DsNZsRP7jMqd8fKKVIeTa4qts6eqJmtf7Je43U+KkVcb7egCxv6x6
gZmphflE3YGUvub45amWjV/Ss+3euphNIDSWf8s/mBPuSF/SCxKAtsAKbccJYq5b
F0GUTzEfUvB2wElEzX1JaNiGpz+JtLkYiHC8/pxkqgYjjVis9sOYRkXFEDwCReyV
iYAbyw6VyQ1lvRE8xjXx9Loi8GVneEFNLIuixaAd99wcm0LJKphdYgj6Y9m6cnSJ
19jLdUcVqODMEXwhJdgvFIxJaSSq7KKc+P+nbg93B7VHbEWuOZZBcyjR/yerAIDF
U7K6heA+Ce+JDjDcI2mlj9XNfVihnZz5Bcc/D63ciEWw+VvWLWLjImYEm8Wtzoi2
O4gO9xLPwXN9v4FBkxseN0OM3RdDeXNIQhpB/H5VSWF/VQMimQYNWvxy+/V2yIez
qdv1M3PphwrYc9iDSqdGh+Q2Jcu+DZOTwNzoWJiVaPidBtYVUwHCDFtaCok++zKU
A4yDxa7OqXcBLt0KSWja6X1TqGArH5Zqhe+s/c1IRrU2iTWMK6BXEvtLtnobBlVO
07aRwGI9HTPN3hkKYmRO+IRAfBhTLJdqPC4kM9QNDqrEAWpmJe+lj65DlOUGSJMb
2UT4TmawKmjhWaPECoH4Syp8fL1S9Tf6958vJ1dw3HDfV8M+vl1FOb6mOq1T86J9
VA0mvViLnlgQQ5+8FV8F+Js61rTqzA2iQhe4if5Azhk1OLR69oIKKAHO15M+9VCi
Xs8ppKTDd16lDW6FMhRVmwf3RKc8fnmH7SMQGT5OA1JlrXEpde2+QW98i9n99q+M
5ffsCWCdtAspfTRR/8Sknk+AMuyBqp8EHD/A3P8jcd0mDcb2/qaw+4N/zJ7L342B
HN70WTpyABu+HUlI2+repNgc7eSKTMDgEAZ4MCcSrUN3y10hIzLdzKFBgtgfEfXg
jHCxUeD69cjbDIjnaOhMOO9Y8jTd/WkcdV/wlEhYQowVMxl0hrhAW7So9lSAOppK
78nnyVqDLNvaHw6n+E9RGvHrCBpQsirDJ+ENW8M/+8ybgWHtdU4b4dfiWbyaCg1E
yQS4dZRN0JmeXRrCAPPLnOAGO0p7sslBvKfReoZAqxYwTrA30VqkdihYmcOvISs3
vUUvOlhQLvM2egqsqblAGnTGFmHowRYRJL8GiLq5+KBbndu1a/axN7jUiWmE05Oo
TR+UWVE/0aNHRRSgrqY+QGPHemSVaVNrg2g8+06VEEOOdGdKVj0LTf+paqwbduJV
U6174RZZ26SiIhYnzWHAeBBv7AQzfXl+YPKui9IIDEgQl4yLMPQ+SV9uiLwPbd90
tmU+KOGPxGB1a/CfZGRE4IgDbrwBWpXdQmQRX6q4C8O7IDhxx0jIMJxTzW/tbNwj
xWlRgFC6hRnNQX3mKfnxbxa9AFIs2u9NBxroRJ+e5DXgJzoFfkgeK1rlddJYN1W7
Sq6xNMn3b6Mp+u2WO4fexbObd3JqzD219A97pZiRFvImW9Up0yKF17E26qloOgQF
w2f6giqGK4Tneeq1n3BDgKHGbCf2CiETOaZ+0CV3Aesv//Qd83gNgt2709R671V3
9zCnXOZf+G0ND9w+CfNN6q7x7nCuiMOWvu41IaFKpnwBtfl+YcjXnpe34+Pc/5bf
2XWDNpr4ZlULe4dFEqjLcLAGisZPBxIRDGg5JO//wqKQjLkajKMC16FWCy/s44I7
CFeNSYmpIDu4z+w/vu4lSsQjY5mNYizDZLuNM64q0Ms1MGPDwMsf9neVoK7xaXSp
oCvo71ytwlXnBt4RkL6aaISPMiW7eIaTSARYcEvtwXZj4I0jEleclnJqcmrgjON/
1iHTh5eaQE2CRS+CLPil41gWiR+J0xGpDMqc6TZCY1CZjWtXmfpycsWjyZZL7QKP
CnXUSbGQnnZl4vBYhXu3JDtThy5SreWU1wBwlQ5PFS6G4Mu7o59I/+p78KiycuID
xd8IHvNlquJSgPw6QzJO3bm4Bq37MOU/gWt7zJA6UxP8zsxur4D2+ianeASERSjb
v+3A2BQACPrlT8eU4TJ0C0dTVqBpCmrY3kp3hC4ucwa4n344Z2hZGFv2URYQ+ty0
yGB6u/lNOI7IJf0+jf9LB9wt5aTzTm0nnknNb9xdYJ2NUzDJMAFQknSvyloQ6TY3
YVmmtr43A5DwGOF7I6R87MU7ZDCikVm6iVVwSOPH+8qyJ/bXZxQXAve49fJ2SoL1
G1LeRLsb/RtEJ32XhMAPmsdP4vcHXll6Bsvvi49Q/7pkYJl/7JTkiTeADv3Qea77
d/i3n13d51P4K54mVAIn73Bjv+vOPcWhwYN6+P+gtrDHnG9L/ZHr8Eg+c5SX4VsH
a9ErsFKowxzubulnIYKaYhLxM7RwjqiBU6Y9HbMcAJSRz/YZJHjRPc6bkASob7dJ
knMl2wElaG3yvozMlYqU5gZo2vgTXVBr60YBeqF7c+eHPkBUpFB9JQ1eWdylfpcQ
QetYDFLOIOR7o8nxbF+6h9Iw/dJ4cxyP4a9xCDJzANIUP3GDeKW05fMk8VO/2Lqd
SSeJfFxdH3MhfGKuaCkEYfqBET4i7m4J4AcVi8yMIhYwCOHdQhmSyPP36zqxhDPN
ZvCuNnwFADrXm/qVfruFO6tg9QaitB+gYAaoiJeB0dG3QIZF43w4DqLg3oi5aB13
Um54iRoCMY2py1MOnO7W9S1AGmAFnnYoRNe0BQ7Jnhy5INP3FRrp0n99zZUifq9w
SM094c4Scl6AFx7EXn6VGTDB6h24I40cpNrk/6I7atlIiB4K6a3q/DI0BZtPlfUf
/4QKCQG1dXnfwuZqdKB0gov6BlWhcBlw89vQ9BDaEUuB2lDLAJ4VAR4TXGACRV9O
OGIyrfmss5twLEWtGbpp/zrzrqEod/No3UJh/l/31QPCjPfyIrLnGMZ+JbsDF7bx
vJ9X+u61kS3mwFTQhe0zcfhgOnFUfZ+0+b//XoOQwnTi2IBQEd130WP4nx0Dn75Y
pfkz3SOPkZnhie0dX7yojTqnaMtnmoBjUoCz+J8DrJHwUaBYoKLg2E1+rOvBCjPE
u/XHmDDV1+lt06Cmv5ovk3zr+Ix/zXdM4pvzfxmX0bMBqb02vngfijaIdY0fXRhu
GLUQ2VNpcNlOsBKE1cMAkznrYJM98L7L0vb2apRinBY3dMMlVusy7IrEpkhf5C4r
2nxDLTcLcVp7ZRN2hX/u/5tSqaI2RX181HkdVQ5a2tuV+MOZ7eEZtFno3iTLSoeb
jXri+N3dmiVNIguzmBSUER/3hMjCGsKL3yMWqi8VLoot/7/VUXMSouBuyFRh3KLR
AnEVEAX2Ek5WJuGjKJ9/0+jIDJa221IcNbZJ37k/rDzNfvx2nLhlUr45gwFn5KLk
YbTYVTvvMTI5u7Qn0mkJzIO1cY3WSPWBf70E+X2q6RsHoFHqq5lQb6xvqNCcbEZ9
mfFYKjcEy1JjO8fE4ceOSVZ6hL6ggqJyBPOb8id7TMxtP1f9RPqq9ERcO/o8MLU8
PJrKTzjsDu63Byg247joKRYyWgFUCo9ZadBcrmE+IylwEIrmwujimOmt2JIS3Elz
Wyh8YwCK9ck83Ri+fu9tJE89lTGyiAiAzrPckHkRwHFKuhw0GiTFmgcyqX3Lt2YN
3POr+b1S1yq5hxRBI5dVUgPzLLFbrjrgSKDbfd3zlRiIdA12wCV6waoj5JnkL6Vs
C8d49V5QmHYROuQnduyxKBcP5bzcO6ktrudTHaZN9jUGhVg0mU+rxW8/a4b+D9eU
iqySD/61oVp9eEH/PX7xE6C5Q9wXLMLlmNGz/KgFR5iQVAYpEo1+b99Kv0fY24Ha
u0rySG2Ds92bbsi0yv4kietW8zTSu9xAsx4Jtf7a+TthRxkCuSZTpPoq+Dh384T/
45hIJiDP702E0RWsdsfSZoVuJSpZQWLDmibqR4IJU9IgrYPVKQOUgbuCL39TB7rN
XnZRemyFTWoyV/Z9PM6cvzbg47f11IoZJHWBZUSvHKImsSfgSs1aPc2GMwuwrtfK
wlwYqX0kEJvr7v5kVQdO6m7gQMi4FYUi6nnIRxHlGWatKBGoUFlGoOOQtQLPTH2M
BNQgc9ciFJds6+XXc+36b8maRSg+/2Ykt5CanZAzuhgk6Hkkagld1ZdU/arJqnDd
5tLifez03RX/bmS4EK6IP+wNWAy5Fa9Hg6FX842BDWMDNLmnBpFzBKy6JZxQ90b0
/INxPKTwNRu7Qz0gQB3Z5X2TNRFosOQIGBDa6HQSIiqMURiTiEd54JuLM+IIP8cy
+ukKcycUEiMBix/iNbQXzbgJgb/SMHC/0cWiYiZS2E8V3lMcM3Rw/Yinsc0c9nmZ
fKp9mPSSMosaSGc4hdRkwo9J1MxFCVKYKb8y7VnBrXo5eh+Z3HmUQQpaqpczLN0V
x5RW0d+t38Fwfauo0wIkLdIjT6iYk2Suo6dw2xW7WPipE3WWml3HniE9tm22sS4J
GkXHfUxNgV9EsBAZgh2n5zLvU4OfyrOD2HrlmZQIKqKMl+lm1SccrQoJsGpk6eWj
U7Mcw+Qyhx6v9oNpfdQOXSktqREdcHCNR+sgLEUQzc81FZL2cUrAKAfXCAJ0An+F
XzX164o0E51oSsp1yjBfzdoz7dCvd9q5bcCeIVG0rxmcg13UB9n10Wix6NA9ukcF
VW1XiKOMdPwyT0Yb9msJpXIVihegO9ggWzRhZD/YVC2wZY5XJBQlubXPYwxWksia
I9isgGzqaIShabmfc0xvMsCycAfGX+/INzAp1Vpj3dOjNFzpm36edv1IlfedG/oh
xKbWhRymXTOMJXyqqVzjKDRvhxIg7Dj25hpPJ5svm7U+ZgtbNrVcNbc8WAlrqajM
JUa8w4Rmk78QtzhxQeueciulBfX9LOn/isqA59XkIP5CgIlrkw7C8+iw+ng7wa3t
sv6ezrg4TOAsfqyLbB4rmh6xVzA1HA3vGvVEvCU4YvrGYofEUWbVHheeSxarzEjt
DW+4klUM3hpUg6VBHTXHZYX/JCdF5iiJo87gM62NOESTjBEXX07CzlkCc6ZIdcoG
CxqI148yDyYIq7euSJZPzBQLiq8cr4s7SEZPsv56VMAVJivIdsYC7p0llq2J4lEO
VQULkkySpn2YVoCUQ8OeuMsNM7QWRxLgXLjbMQJ70xopNQINKizbjEEgh+fRGEOJ
oMht8qGKbJus5NSDsRR6k2ebJuFvvy+aWEhnr5cz60PU04n2yqhXHYqBIESTNga9
Qu/Ylv8aQzdXFk4OXnpIwG+/s7pRfnNhT6RSSFO01PwlfiGfJbgUt4rPdrQhkGrv
rb8sHqmh4z25B0MauDG13DzR95gO1z7vLBMuXtZ6ZoiiW3s81N0zz57U5VIac8FH
3nmgWlBclAwA0MzmumyVhuhSHvXvTwQDMrwRToJY0a/OmYXmo4ZeoQW9pXvwEX7g
kizdYD/fONLprU2DzQ3qLV1nFYG23On7FNihCSmmhBh60GYj3g7+3kQ3ElUd/ZLW
Uo29mbxIIB1epsmkJmBf98vzbCyDSGjqEI9Pzjl6euhOs4hNGaPawIQD4bHYbgQQ
JaoIRdPpTn9iLc5bOcY542XRgs0ixli3pcJiddTAZKHgz02+T3drStnsDzrZThNU
/zPJUHjQFVeShAeS/ZgWyz8eoF6fmV/2eovPfNXau4x9cfrddTXxjexvQ6nGQ0+n
+YQSBTYqTzLQFXlwAtc2KKCm/R76mmAr/diu7wRLmgALyG/ULS2ndAnYXZGlpaXg
M0OVSn4gxeT5eYpNi5Ao2KAgV0t+OfWDssnRTK/7dGTfp9egWjJFiEb13KoHu6h/
yU55dvj9Ff5DehrBYSGfd+0AcbHoAm/QxFQy402yc51wiYRptvFPZyrI4rCk1yyN
kLi6ISHgfJgEsn1GtwYli9eFvQ4awhqVUDORDmu5mTLb3PfrwB+7tQLACwP3n8EG
yILR/2uu03AXVNdn4E1Zd+lJecH8O6GIwQDVHe7cLZUCWvCjpdqXZ9gMwhEhXnI+
l7WL98jWDbt0t3FLtpbfF0IYh6miNzSb0vjfcepkHW/HReSzjxyKOpjLVppJShs4
9anVw0NBZD1IQ5Lh+W6PsZpDbosksiG0wFeK1UhH2ioeRzBkZzlOgWoeBIHnY1Eu
tZs/7BKSgeuMBp+/67ipb26EJQdoNFnkkkdVRJStvGT3Xw08gRR+d2XtwWcNVj2p
Z1r+TpYH4h2/wGS7TR2uW1UN3WQdCBiMJr/+hcYrU3xoeuigZ9C3d0BR9bqdRKwW
O88hK/fG3D89JPOYjjfnQOl8T7RycvZwDG2YAZcLadkr9LtdCuqp/EtHbhq3nVWG
dcS4O/a6WJZgJCZNCmfsoemJKOZNZFBpU4HTSqGqkrYLZNzQdlCfz1FB5uK0jcB7
HXdrxA4JswaT5JPtxrEC+uBX9HYooJQwTYjnVcMImiEMx7x3/0QXAlUmMltJn3Nt
Z/orqRFbzAiOiNq66hePX8vYrHhAeBdjkPQVU8UA29JZCLIjdQpLjppjwK5nqE9F
lvotrACAf3jwQYIlTh4N+9MhRA7XTKGAZdaX0I15km+sQ2thIRO5jLrDWFE3YPue
63uZcBfi501MNKmvMJUSAqfrIR8Cbv92WgSVgiYDLZ5LUuHanOY4bFCrl4lnrPoB
wl4Zc9/ZNgqZIL/7JIQ1a0wQRo+JNOKRpG4djJcJwwOcHQ3J/wC7N5IHsSd8ofdI
PwguyYwGnwfR/+aRHD0lW5ULXac8Y2FgsNZBJ27dEZBE+lmO7QwxPV4MDJrBczRC
wVRrY7CDD8aWLzWk6ts2aAs8aCz9mvaHdnK/3hZpDUxksA+py8XXngMIvTqnVUA/
vrfhoQ9WUIWAs/IQCSrKEY0tp7Ll6zxGcmUt6mJUbsD0sC6T580ZqzLL71vQEoVf
7qkt7kVOuILrYyBHu9AKvoB6s6/tZragX3V1HXe848kYFWAiS5vW7A0GMBOuR4+L
LTySfJ/GIV9rg7Ia3LJ0MRNfZLLYySAgvYK0yrOOTme6jVPw2EOKAPny6OTZpl4e
wt3jZuhEp/DjUgQSKMgatD982j2l7G6FDe4znlZROrCs9SBadgN5qwZjLMD4XN6d
gP0vGVfR8fI26AdXO+b0E4rIqAaNJwROwejTRqiP6/YEP+3adGjuNEVx2kM67RPA
M2fnIazdJe+TrSeREP4bFpU3m7xKPRxsSZjULLpR/8enm5gdKHgPk3W3HqGYGH+w
zBvAcRIrN0D7NQdnS5xyJ7m5m4lkWg7cS3Z5KLhPv9Q8hDxiH5ZavjoWZcWnf6xk
yK5p2JllhYXtJ7OlDFHK/ZWwZpa9Hv5LfqlrXAJuL/Uksy8201LcU9C+YZXu+CPh
9l5bV0ZNVJvcLxj7aMD0v8g25eKuOyIGE9oky29b5Op6UezwmAo7vdlfgmAZu7JA
GqvKnk9xbO5phu/JlwN/FzoqUQNlnFJQdmfQvW1AAjLo8qBVskwFO7TRwwHI7l07
5cGyCdnoAe+Zn9pPrEIvPpPKj7bWI1qsFtdn7oodFWRFjoj6Kl0XyJSl0oh9G2i0
l3Ok5cedqQ9Y/hjRWUrTBVnHezZ0Bx+ZDMryWD8WO7oSigsfvGINfoMCXFW5V0RH
wvkMWYYFjtAZn3Mi+RYRe7f9mxasxB40QaAa37Sz8jUyp4n6jYuI6MFSVbs0/kVA
W+ZtDV1ZfVZh7pj16NPvL5TJ8mQNSKc7rA7I7NMa/OdstNalt5fdvulXini5sL4+
oW5OOAuoRguZ/x3KK1/ireAMDugdjJH5cJKVzuhj5l4FOUm+wYrJOhO+PlJQrQap
t+w9LbvZxO4PTRxDA3zBrfa0S7ubuAuBsJJ5zJfe3uN+OT/HaGv3obfog7uACFiH
9STlVKCS68cOMALH8JbKhBjfPMlsi1rdTip6ZOh+yN2xOGsDEYG7sbyI+CihpT1h
uEfW1nUExgNFQk4biB/SXSVm/NYTnqWQvndxkGDKHjjqEP8vQ2RYy9i7NRnvWmkd
gvFms1WpYB+rKiDiT91NuO62EVX4MBLyz3Si/gc32tfMSQKpROjDDcoWVIOaocjt
y2EmFLIFNcP9Bh5rUgx0qvuARWMWyrSioN8t42DJTyxxLJc5HlUEFgQRN0cVH5mK
QYbVBYjIBXArUAnJyoecfO2OK9WZpRfIhY8ifeeVRWgWw9bcE2UOy9BPPfaOG3Vu
apW8sNtnmgpsIQWn4W222zlpdFqEsf9AAasIgDCbaKpkAux9OvQqeKEAdBL8Fu7j
bQjceZNyghsvO1EJzA40nmWa/2eEx9c4ZZ9xWK6AGoIiyvuTk/pdMtMPj4SbOghO
naOlXEqZmOGZpRB1RCWLcWzKZ3JEaU3QzIKamptdSDMnf0WH3tScACP8Xy00UkhK
mr9VMMdq08kALXZ5kYsEirlxw3KyrRSN3+/UzjjJx+9/kkp3DyLoBx3Zht92zNOK
ZA9wzaqE5zqi9fJhw3k0d9YAV7reEiiTgeOyrDZvklcd+srbKJRz0saHe1DjZuGB
6kLDK5nvfsUJOaZdOkTKcrJLzN9uWT9F+kznh3OD0sitqR5bbi81cfhrRC0DOxC7
Nmpgc4WD29HDfKbmzHACU32OGrrENBSyTI8sIILRnlTqzJZL1qT+d3aaAupGAcQ5
8IByyt6wo0EZFfTgIeVVql81D4FA5u6+1umyqtFpc67Z/xVy7XuIPi+gQVd5aP6b
OZmxS24llabX28gJG6AlhWMtBav322CHy2YGWNYBc+pJfSokAPvBvE690B520nHc
Xu62zP2cKiuV1SkGuiwXxba5zYC+PYAv0C1JRuhiUZmtcoKx5/FvRJGuv2UcItQ8
tQaQr58pjtMyNIiLQHg0BHM6RMi35yyzusgAiKqZ248G8/cV+tOVChStzR9w79Lm
RUADA2L3Zvl9nmEjwKm1+CJnOhVWQd47wlwiItZypMjIaHZDgxFSZDt8kgNP1cyi
L10bB2XpulkFHGnDX1MWnEcRrNc1SNimYp/IQ0FPnrVszSvM0lEQVPLHlPbwCXl0
XgcO3/YVcpKamu7nyjCRDsi+8mXQnFjazB9hqBAAkGfU46FYBNBKoNhw78iiFX4F
+maZTk4fJLTP2xi+Pa2V73sBK7i6tsb+twn/t4spez5GHU8LBizsocb9uPUkn8oa
bcFNxkP6eEcKWEgl2NNociqogtOm4PFPqs4ZjlaehEEVPp6MgW4fuFKgS2Aj3fN3
2saOoKK7ILlDizmlWK/YiIyPhNWa4kldBk+2fC7E0lsYwVjoiZdUPenju6KibQRJ
zOPU3JmHRDUyOM2E58IblGMkBWZIBen2WQcS9wOozMoswD4Rh4PDoH2uYy74YBe/
0YseNcdQQheozZkIvlIyaWo4mrdzB2YTa1i7G+EtXw90vGMdmIjzR92kfnIqJ6CH
P/jbQ3vESv2eyyhmtPaR+MnF3BbCD4kOU0SUsZBOWcIpYNjJAcjSvrc4wcR0ZzAi
PXkclQ2RFJ2SERBaTYiVsssHvJxX6VvqSLMyYiWNmQqSgtQA0u0ahwCpfY83xcWm
ng3709AAErBWqQUClp0leyUU99e0JDrOaO98iRKYkJt35AXJKyiAzr1v87B8WMlF
8Aq4w3hoPtmZbKK8kCpBulvqK0Uc/jw328m/YPD2DYj9qkGuFHXagkkVk5Svlvwh
/dAPUF0q2BwyGlIGoxRUjHASbTOLQFEEkodppZMpY1jtE5m4Klw9skOV223pX10/
bd/vgotUB6bGWWTQZjysj/VKk6f++VlDJl8mfZnjPNoxhdQYHm4vMKCMO7aFOvFl
ApDGdo5zcDO9WLr7mivDI1HsFggAvVk6G9EjQ36VEiw95fG7I09Qeu7hCowJ7VaJ
feX7R3FL3PiCImvVfKqKPlFccO2YFwIjYMr0khR+26VaTbwaCsiQhLsfpCYNERdz
9UFPWZ1+R7wGOqjg/m2K/Ad6TmqfT8JOVp70acYx+3xPOZvXVBZFMIydwqe27GCU
wWCFQDUFDe9/kEFuvTKCUQ23xEnC42HVsAQTJeLraqudMXLWZaUxiSAQiEPbRKMZ
vClpO5mKb8Uqhkg8oKuIBwm//dTSzrOZhA6wTDMywKZt5eK946at//AnFqsSTBqn
gPsIyw0ooxMFEY6uYZAx3XdyvFI8Lg6hiNbc5DQEGO3x4wD68d6LwVGDplO4EHvY
0zUKbLVZPXEoiAm1MwiM4SDJ6tyNMvlTFiS/ZRvDlNY1uwAZD7ugHkep6qdtjzKH
/haQv1O9aNMvUtXHlDj84VVhjkskjyazC8zc7b8YfIwmVZ1ot7y8PhWWhNCHzqm7
+FYQEWFdM2vAv/Nv2NvsAnXvZiRTLDfb1oQxThruBlVzVPKJRAfjocbVwiOa/Da0
FMoCIlfW5Pmi4pxCCGY8DP0E/APVIdThWtrUlTPE2dWcWzde24gIKrNjTp2ZKhYJ
du5MqsB3PmleFgY83/eqNYZeXZuVjbxwnbG05uYevwa456i+dMEhgGyFwoKgRDNa
jk+IWT/kzb33WTyIlAwbRFNUSiIiwnNF2sna5SeAeEEumCVyArhUMXhrLSbyoy62
Rt11DqbHUt0ZWMt5RTgRSY/xxVaTwZj5c56waPs9ufSh3dmrMx3bmZuUTOyK3cGT
thZBHopmZcSNPCpumczZd/SKPBirBS2zRkl4pK7ryZwVCAkEDsP+vzMD2AjPdnEX
E2Zqi/ryLzRbYuwXN2FQ4zyA2p6ZJERXLpqDckQ2E7gjNR1u0r7Lk51vaEu21Vp7
jN4yBqB1DtKlVoeqhZjgKpYTWQVxvK17OgDw7VJRl8wIQ7AkDiqO/o6Ixwd4P3y/
Aim/gsDWSbs26jtCUcLFETof7hdbfmwDGhZQkcg6g7bsbgXMf2gF9HzmYVUQWgWu
OZHyUeug9qn+KDiitQcI0ZMiFISWCzeV4lQa0+z5sVaY1JqjhM5wMz+3ZDyBLlIk
h/Xh+3JdRUTPN6z2oworK/vohT6Xn1sJH2u6VLxkCDmd++HMcLqW1EgC7o7FL9pM
kqYfC5czD5+AzTyzNdyYW0YNRDxAAte6j/VE2aj2rYfBFaL5QpaOJPpQAIo3qcjX
rfAtqnNrAnNHfn3mi6k1vHo6CZNdHHi3BxuHGOo45i9rO6rOvBP480t5PSuXZpN7
Fy4w5YzsVlvrioP+ZmHuZZg8gztdHKXszxBoAhJBrr66s1mD+wClGKDo//avXwT2
ZKjBuhy3PFhRBW/2zjl1p/442q0fYA8waZJPmcaG/EYb1Zh657sub01AVTb7I70/
iGEH/G7XOj58S0lXoD5Qo2SJ8oePLTsGRFqWVqtP/7q6EEjD1qRlj+ydIX8lstle
WrRxjFUUjzpj8iDEsb6FHBYlIgQ5butbUXWfvdfRWLxWfqHt4Dwo6wqu+NV1CE0B
qWfLiOxe5RTPCp7G/kxIp+ghlYRGtSZq5hA5JrnGgeN3dAdrDTdCOzzJ/HGDOYGg
9wxSq202Xew/R+lxm+194w6Mf0pEtSiw5uOIszxOCOUxV7SOOm80/i5Rg8lLCtQP
P8PRX5Oc/2jVYySX4OEXNFwqX/90xATCZ2Ju/5H8ju9aIPJwdIGIYX4jX/Z+xuem
pjKhzFv1XB2/mnaQtlFCHFzZclYR+xkUY4NKCe3nkswgaz14RCZ9YAnlp6za1RAF
uSYRFA6DUaKwixCU7VSVAm1izfUH1Wm747pQ9FGnc7K8WxHYRpVCqY2k1b+j22Hi
OJs/Jld9b9R7Au2EicHzxRFMto4iK3ckzM7UdxqtME8DqGXTDRzJSQlBlwrI3UvZ
V75RSGHj9B1InILBZXlxGXaFtm9//u5/1uGZgxJKM/ajDPEQQ3kGwlS1w2vhISvr
kZ1ZX9YC6cltBPEhSsicaoRhWsLTsGrkpoWp47A7uuYKFLEkoJ2htGlnkr6eocrK
Us56rkcjtHpcm19vn/66l9/sFFeZS/3Wm3Aw48TOWxzFd06wpTK+s1Xu+DW6cz8i
xtvDn1KfGOpMn+MOH1nvasAgqTBww4FiOiE+7fGSBoJwMCoI9gTQauAv7hjvrnwB
tKoWFx1ztc/YdlrRMnJF+p6IHW6d3hK4GF3hn4jf6XSEg4RMY4i1hI4STF1WT5nl
tZbmESjEjRM4p6e02qz1sPMMSjtIoIP1tDnSx6t6mC5vWvaHM7D7R9txsERrV4oe
+tEAcvLu3us6eUsd+9d+/W/ABquey4heg0ZHH7gn7CiV0x9dcrJOfyTv3o9c6xcc
7SR/YoiaUddURMvnB8yz0Roz9bp+ad8HDpDHzO+zi/yB4nt8KP2vl1uMSpEr5ppb
H+ffwFajZwlwDFcevtVFwClhTK9FpDHWlZmZOIyTDkturpINcTWwhFL6ExZ/7ds2
9n09undSsKWd+AqCjNWA8Y2EBq9P38cD6jIN3eo+hMQag/SYjTtHhe+uI22lVaz6
T5hW9apNMsed/VBAof/DBolFCFA4nqnDf35g8jSG1inn6hJpYbZ3zrUymndCJvx9
90j/1jjG/GdI7QuyGkIkSb06w7n7qQEVIW0u60QEVenIlCbpaH/lf+VKYXGaB7Rv
VeD/5HIenQkSPy+eos8WuFRylA3qfWof7dWD8D4xNTvofurG+ubyaL9cBxjMGEq1
+M9cAlQHo8ICGULbl254MBab5IQkgmftx/RoBCfR71/9+sCoSi/hfXBpJlxz/7NX
7vgCrTYjjZrtWSZ2lkHSrQ==
`protect end_protected