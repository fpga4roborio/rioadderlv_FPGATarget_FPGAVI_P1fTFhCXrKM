`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
ddtXksX2+yylW5zu6QL2Lhnb2d1sD00763mmSITNX595NcHTEkwn0zB1Dry37fOW
FufOhVzEJp80NC5qZ/+F0Vk7Ik02dIR0elf3clrjeJRK85K4e3Hoo4xn7YbFUIms
l/8VZSb14+JVGURjfswrIyCUotIzlzVYZ6gzoZwDXIi5gQIBf/gI+KxNXPaKV+PQ
Ufys/12rjO6aI/pPlqSm0hCvftmBcnezN2hk1UeXgOIuKZnogjOsf0iJVX2aOOWE
6pD/psybjbnsNB6kH5uFTA5frkzIzkzl5d9+YDm9OyC+k84E83I/7/j+rk4L2dah
QJOvksSIzN867/4Qt8qYTQ==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="MvBXkzurAa5VTw+1JJ70nePUfoQXBvZOku/SMmg4TwQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
oRtzZL4VJ4iwysPsC8SXYCzXS8Fw2gtZTOskLcDV+1B9Nzn1zTyNtlo6lNICRmmK
ZRVu2BmCc2G+fmzynYlNTnSa7C0Cuel6FYpxCBlOuk3OF2tzAmLAuDyOH3Z1Yjzk
a0aHuoCdIRKv7BrZCdALt03JeUmXKPdOmIlkVGFl8yw=
`protect rights_digest_method = "sha256"
`protect end_toolblock="Jn9CQpRhJt4rnzZPRk+dOpzAubz7omckX1MrFd4p81o="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 21328 )
`protect data_block
gD6l00tciPUa6pDNTk/+t0OO0nC/UTtBwLB41d4inuAUA3i/ALrNyoJVcBnAmEQW
ptbcNp5fxEUJjnOxnedyZEuEBxWRieZFQnkRdF269oMYqYwLJir45fcqmSmqk1hc
qS8WdiKnh+Pmxn+/y3vRCaKNLMPyF0nSnSgg8djFaRh6ZelAoQCZJ9ZRIJK52cGH
hCkYlc3OXPj4aF4ul0U/QuA7BDMiCgUyCp8Li5657XiVDi7A9eVpxVtWvR/q89py
zPY+juVEH+SVFGr/UC4cMP7Dn6g5Hdgxl29kUHBQNna6IprKuV8sCAIseSroPG/W
Mgu7RF5XeMWPlSAl10Y2Oorq6pE1vZ9XPtaesRBRQ3GBh0NCLPkCv7qiAtb94oLR
lDYiJ+Bm8hmF0nhuhQU5uLVPC7du8Df3eb9hfTNE4028GH2ik2oVpzQCGnBx4twD
8WANa8sjyWg0uc8KEerQxyTofbK/T0aTJxXHF55PsypjNHpHO+ULD6uhXxXhexp6
g6CHwQ/CJ/GqJ+jmj98vXSIAt8n04JhRNoMswuf0dyOc1dqEHaM7bNRTEF0OCuvl
rg70xctHfLPBXSentW7L9E2/0RS2lvX2KbR97o2aober4QDVm7YXBhrJh25IrWCE
vMrqGFCK2ahXFmM7lHEhwoMbYQ+rxedH0l5S+t54gSoUnREgO5w5R/8O86ijsq51
508IaSIQEmnNyfmtWqS6aw+i+MuQJw3L5SPbpu8KbV3j0WdaZYQj761eeqgDp2nv
mmH36Yyil0L4Pi3nUTgnItkNV33FkiN7lsz0mqIh2NnHv1ztDHj1HAqqRr5L2bSf
5rXn/qnaPf1X7DjRAQZv/uLgPEpgq8r7V+Lwn7Sas8ooybirUpDmC5t0LD1m1m7O
bdw4g4MD8RnjtWDxABtgpSN9AyNzATAfz48Q10Qi0oM4oewmOmTFg+ZrOMuAscRj
OYXXaXa2hOt5d7ITnrMaJ4w3d0LJ4CVOYe2pb8AsF1Ium8JrbcAIUYCTyvD9FRT2
gYfWczpAq4x8Hnb4tEF1OO1/wI2n4Y0wafEY5i6Sd5OCdYGmEv96S2E7xvPXuVL/
oG9KDn33bN8OaB1DikLA+7buu1VViq8pxNk3QVmFVvNP8D4gBCHHiWGOp4pswP14
nk7uByG0lruwZJerLXpNVTnKMyFeN4m93UfBx1wEWjMu2D4TvC4vQ0AkoGXmZ9vq
5cbytbOa0R1dO4lAbvgkDD8EwCeEeNxtNYOQVJRe+NlnZs0e6Xs+Obl8lhe7Vl+y
BEHjR8UIk5zUxhql54N5MgwJj8f4Unw6dcQQyWF19GBLQ9eRqw6mbO3+f95kX/ux
ja8mmererTH8fkCZmbAtAq7doOaxtkUHPaCHFkavayZRogCP9Oiy+OdqVmpS+fzR
+l0GVgsXNc9lAeNTTQX49WGmmBlxtIA1nbmzsBv/XRZM4dzg/0D+mkoErZJwm80u
5sV0ukaFHYta+8gSnUhRHCVKROSaDuUNCWmtN3BOYlHINTwspUAUpCDZmTwlyTiA
O/hndUz1jK+KOp1j69oY1xBRXCbkj1T83DOnJExnw0Ykwb5Zp2dnxsaG1nNKGJI/
6kYPiWN7FHlfPVuYb7wZAcpx6vQJArJlQpt1YM+J+SEPhFbHAzH3N35NfTaILsE7
A788sZK+s+N0fBIRKx+ErvTMwJoAyF9B23zOrGodplDjt8YLQl52pj2dIl1Pn+5v
cC92/apnH2ocbL3dFcuOu3La7uJA3MTGPit48aXkuLKEkaof1qJucYGc3tqHj9TY
+VpXzPBz5mYbCcnTrV/5Im2q6o+z/GHX5QUX6f7+yXsidI8KJqZfywLnmWyK2MtU
2mY74a28WYOefgTN5PkkaivAhGU1Ujl/BktT7VALYrCHgWlGhs3R4nFRGoePlcPE
O67OW/JIXU0JXCZXhLCsa0lnDD8suiZ0RrFQzyFC3b8kSVnX3rBZzq3mV12isytZ
pZ5PKCpAc4pHLp4Ce4vf7tHDWe7ZYYX4NMnnEnaoO6r+BRosKfszsLsDK/VkjN3M
G9hOhnAhQ11k5CDPovZVzwvSs3FvshgplR+AsCmIJV/3HUa5KHZTeoNJtiJJJRSA
n5iFmxwrsDb1/9FEaaBjp+3+OyZDdJEsLzAuXx9yWitoSDaZLePdsG5aPXFaN9x1
if2JBlSGCRyS2WBV1u8hUT0DAYF3SRrjy2kiH/AbeNaNxSamSLTVk/FI5YlP+xuE
EvARooNHufoXnQ5/GypVXCPORnTNesUKSNkvMJjde89D8Jt/41GUi8Mqs/0cKdlz
upAvHX9hu6oxzoRGYkDpqA92M3AZAW6sZgw9QLgQS5wDbBXMJvw3Khsd0So0phXB
i95lYjulfzWCwbRFwiN8j0RSlJWNG0397VYezGBZUURWcgehY0ShyofE+Uei3BQB
IXVx610asQOqd5tYRswDgRkFoD5JrzGHN9TqTfP27ZGRIo/t4YZmfUXQwSKH9odN
fju20YZrugPzMuEa6rHym9Qc6TyM4vLF0f2McQE0F4Xh14Zv9tnHdqUf2lqvUm3G
xJ+r2NPjgxmecLQC8tWoQoB1lOZqz1PYyBVMHbORxU1fMtnjHz2hFtP51kqsV8bk
ZuPAxfqJDcljyvACIDOsK6U/WAEjb1UI264zizHsPn80BM4g5gh34XfZ9vLigDlA
j4mAhEWpn4NCNL1EWKoRW0bZdqd3gv1xUek5y/cMGkdhRpz4dLcJsUFD10YfdLi/
+ID/5Al3YB/+bbrNBR0bDl34Syg+xe8dqQTQTf1owVMIBWDbqvoLrzkAvLNceVSR
nIhStb/9DGYDVeUqRV4InHSLTXgffpi/HMJRtJdtsyoM0/c5mtgSZcKfyuQSYMWd
QDEE5iFG8UPMxLm4EGxaw2QOsIyFhC67kM4gb1aJTd5bFkBs95wLI8+FixC64UZz
auElJiiV/uvaRoGsDhffTsG2qbkSg3NzokzEp3lzmOxgb12n8e4ctN37U89nX4a9
1aLcf1++bYkcfxCstuvPrOLX1wpX6EnNruZNmPzVxpzpHZevD1OwyNVrI8PzYzu0
oUfbrIqeiTUkYUng5QpyAFC9VZLY6Y29TK+/vhhwbv+rm6s4NHPpzfC3dEPbfKGx
nf47BVHuzr3vKD8YaIOegWv+YdYW7JTurjHT2Y4hPGX7cumd2KyItFOIDkuo2/pO
vxToWrAfneWrxGt2a0FsV67aAZmt19sLTJT6zs30evtVU/Y8sCS4b9VboDDlnWQ3
uIJP/JegEntI05SrGLKWaY0WXwr8dlBj3CU56Q2xj3+lsw4TGd9Lup3qD6+0Hw/Q
1zvsq4T1LOJn4wfkEabJK7DNW8DwKaDzuAGabVxN/HGm+zx6bJma343KwMsQI83N
DU17AfzxMG9RWattIqSnBwIhaBh+mA3OzyqF4O5Qkad/lkAWBqnpbFD+7J913FYA
Ythd0p353YdemzHnsXXAk18ot/KsTIHkN7221nMillzTk1VrKtNowQGFBJUqxTWf
kbC+zZT5fo3mVoEXG7D7k9C0QVuFTsGrrJECAsBsUUUhIB4YGVS/Jq9R7QVyxFVH
ke3GnryDeJOWx9f5dM2QqBxO4SquGXkT/t6YU6rmDjoh64H6vOG8g3p73amHXLhg
O8YGTxGOF5vnox703tsOvWQsuLuHEDcPVhqVppXt9I/s+YULjqMXVSykoj1sw9yS
G4TBxN0CdpchfmP7/AA/ySsYd2o7bXHsVgV59bI020618PhUe+fPUIOOeJzxjI/w
Ew6ZUZAAuzF0XGUFRIQOL9mK+912YsFva7DDOpI7bK+c9ATY8LY0NgHy99jkZwds
75XjrypWZTfg3SxvJ25oj/XF4VVL6Y6Sp62XiibDSe1G8FN1wMBsdKMLiN5mSSJc
j5ATDN3WvXf2bGwYcpggXH6Neupxp6Zan/B5G/6YAyzreC8TBQrdwkCm5A0gYJoF
NOfOyZtEX7cPgGrP614h+yLeSFnXu+/auekGX1JyrR6yxhMYib8VnzcZfu9M0VTG
A75D4TvShJrgT18DNY3m7hzw0eXXFdEFl8WBGpKwlFPrtDayNoKMrI/cyh28UWFY
SfPNyyeY6/nI95qscmiASw8w3uCFoMGDAV9r3DZx5r+Omxr/yUkU0/UI02r9cbD3
cdoe13ojR0StqL7UCA6CdIpJif3Hc0JHLV5ByfY/TfNLIpXW5nIgPcfkyhma5y7T
pD5xgFDrEz251M1TZtdjiD4Za4yoxjpg5oiCz5lgzE2qP1UURwCLNZom/cEoAVBU
rZARGkvFkoMZeR2mH2GwcY8WYz2i/rwk9MeUnQX4s0MfzfNUvNwFDSax3tBlQNU7
4HstzjOTQkaCJro55/ARQov/dFwZ8xSswRyzrXGf6Gj/YGwdPuWfZw6I5/9OOPtD
qwqJn/GIfwEQ6vb9A/DLQGc6UEGqM2kf2rmn7X++e6jhRwkN3VmEQdgTPGBf/Ldi
QStByOQcUI/4x4dH0pHuTO+k7ILM3zQSds8s60a4SbWU4E64MRISSFSd3UQAzwx3
MrZITfTr1fTto4lFnkan8vWfm/uZ1G0BspGAVfscIlcir9wzgqT8gxqeXcJ1ylTH
0OR2aEcBCHKUenATXOm2LyqhXdcDZ8DUabhsWpso5Yf6GR6krtQPIbq1mqwIchZw
UbnsEdp1hUzuEvjldGVEL/XV7gr5KJonhXPfJzJes6IrOh3Fnr/KWeTwcVzhkvVg
jvQfIeyKW80uPH2bXW5aIwoBWgGSrBnyyx6mzNZm4lCcikVAmtEFFtEJa0xuihFh
ubm56ixHK11VJreE+5uZO6pmdgwLiMKNBthYHUQJox93wHkLunq/KTUREGMzwhr+
cOISGU6JAE1Gh02jmgzsS+vL7vKyjQQcSDIL2tOeCaWkf+DOkh6RRrMdKm7sgXnJ
80eQf3FZJ2Tsv8VmGQnXGNhZox4skmf6A491Cl47k/9DmKdpqTmhUffQX21Kz9Rh
HcWxHh3jJhBHZ7x/JKTho7plYUX6yXWqXcWaXFfQ+1Vxn65AJiTfk6X3rrxDkvxH
LOMxjt5WTwHpCPe9UlBZhC7F1OGg4tItmAtVJBPY8lDEq9wRUqTo2DByZITYdiWz
DmetTW2+LFroEk3LbU7ltxZBNty9gFHJYELGwtEFLf/Rz6ffD/RXVC8JGKHPxhvX
E/iSB3Gh7jt+mOrfG+P7eSIFu+oAzvRjDPWpZVVPxOHseO9zFgtRQI/XijDPWDy3
ocbFHm9/tZyXhHw4ytOJRTCSyp8W8qw95ZfOHKlQwDbto8IwX0dfYsaS+pBHq6ci
6aw3niH5aT1RbtuH4mOPe4O9PVcxv+6kz9y+Q/CwcW6/6LZtFFgUf66T4bjcaRwe
Z9tCe4OZ03FAas8tBqcsiF2uyD31AilJQN9hWcL6SB6kt2AJ2j8GCNUzXgdFeI7x
Iz0hnJcRHw0clZHqOf8IoeriiCjOjHaHExfzdAD44uBvtpws/l7I24nNWrDQpUqi
dOfN5ijdqQDHiR0ND98eTM15W897J517TvzsPqvRl1eK4xMxkhwcZBALD5c0t3sT
/3zBgG7QSQ7ttTLyZ+sEY6TeWq3jvplUZ5rOsJsPJws2lKPXoXkfCU9FyFAD6eIM
Gf9K9imisf1RcwHYS7sn/fvPA43Cmed95NMD+NHs1LR0NpBdo2CElcjeZqSetW6X
CSk2ZF9MwWmy5X0jbzeUpXkwO3eWWqDiLq1Ooo4pTCcmRxZOTmWDGB8hMeyJ5YQg
JmBX6fHw+G3eqio2ZYKWXmo1zhadbzHaCnlseNaHnfTMV797JIfVkkBetom7Rk81
dvffB/AHx0SDPEtCL7aRzVij3DvvJvH+4cIUlVYDGVNqSCtiEHPel+HpsNZf+BCr
I3mVhHM0/50rRyuz+AXIpCd+zdbWImgU/I7GWuW/rHJdOIaurnJBnnO6L8tsYfH6
YSlupkfOrGmvpey1DIm+SKrsCCwXqenNpy8G8DSmVRXR8iGZcstpg8Lt80QwP6iM
17EnPbf6uEzwo9pDQeP3q6/F1e0fNfgHFSctUrMcET0kMjKdCewKDlBSyyByo/ag
qM3hxw40k9l/kawRdv7W50n3a/BMhcD6RsoSdRBq/HC5paPXerCqte6GYYcO9/Uz
3itmMSWLRoKiVptXeSS9iqb/JmWXUyaOxBOAow7we3nHJqWElReww9+1IdLU5yqK
uWhF6f3DXe0psCGgGaAk/hqfTe9v4/40KkiR0vz/uFzXn42Dz+y6541BBST6esN3
Qs45YoXyz5kA+7xUO+Ui6jPHsSGDBF9XLsrAtpokSkO5MnkteYfR6EB9kW1o+aUf
UdUuBL5o2ej0Ai2+hclgX0eiKWjY+Dq4hg4rSrO2U4wqYWbxPgk5mVVBpzEdyPFw
AjolvVGJJTCrlx/0BARXv7OhoqK6B87Ms+4og7QbPAmZddbFfMZmZTlpzco9/Ige
TP/Vt/thkKr+aA+16GTodKmfocKdPCNEFVwEFqAYFcxNbcW8agE21p3R1IubMVx0
dqAPq7WuDoA230pIIFTBSsg+E0RsCFJ0FInl+dvOjK1+0SzlER2zfMRf9ZMCKRIh
xTfnEgN+Wr1hjfHuooW1D0hCQ9zucv7vmeP0cggriLOCrD1Nj119gBj0Zj1mCtDa
ZNFteDxzilZCCKsdrKNJC7vsHrTREJNu15LhMJL7MCooy3oP0It8B4zGDdEeSqGj
AT6sAgFujxgDnfZSTfBQ5v7sQr6o9u+83z73zOoKAmT0esUfsALXZKDHJdZhudse
9xPIyz2blWo/vFNPhxf5aI+3yItFIKYDrWiyZF51K8bVLLY3nB/LloH7RJk2HR69
gvJFs9H7FZ5nTwlFmAeWnZOJ5jyHXlUT1NXsaI9GhNlNPmF2hSgKqWVy/hr9D+l/
PuJeLtY5EVhssFVsc3ExyhYKuN14n98ZAB8XIfZyEW8rnk2D5w7i8N430Job0zJc
HT+oXncgqnidc5o+mkp+UfXrKZVdSrqZcCdxZBldD7IctnBhEEXcS3xNg5K1z+70
yllaBPd7AUQvcIDsJkISuUDZxd4grdc5ueUGXVOvge0nxouNV76uyXagbcPKjmfY
dzrYI/smiwNJPwa2qEtveH4VxNf8yamKHqtfWcWT+l0b9UjLJkNg/P8tHMxmpgMr
7AME50qBJEeKBXDd8+M5gbXf7F/OI5hIBLk4sHvqlerahBZVz14byy15pRLACsO9
yu4djFEBj9NwftEPjA0g1uuhI+ZyDh8WMLuFSHUD5fFnrrADzg7oY+bVwPX6A5hP
l/1gUgbAPPcGy976+94XeI5TmG9FLj4umeczTupy+3qcP9DgMqa6euzEZCADbf+C
JM/sxfkAcrtb2QfDPQ4jCxce/sVqW8mOAhGkWqPc4SwDKGNZtSFLaQ+OgzTup3Xd
XA9Pkq1GKdAobgZjoFqrVenxrDr4rHYZj5jGNCePIMaZqMtFH1Rf+ADquhZOF3an
8y+Sea0p8pmB65E3tDSuTYs56WJtJvUd/C/ChWEWw3am+VyXZpNBAx9iZyP6yczC
y3rJSVJeqiwIUQ4Oed5qMhGvq2nDpV+hGIH6PDshYx7K/JhOlB+HTnRVRqhVRLmz
Ip6s+GZy321zOPYZxdbnqFy9G3w41wZlzIIzt4zG9/dGXeKnaLQTbq8gsS05aRBP
VR4y4TmC4R2RldD+33mfLa+39jsHiIrnvLk3etkTZT3xYdI2oL26NEJLUIiIfBLO
rMXN17IkKENKvRSM0JjZBrK3MeyV/DB1G72hzVw0UWZs+9e5saIneQjtX5oaMsCG
uJslvnTxgYmvsRig6x8xI5ZXs4zN3xFxKSRosIP5fe8DYsDEb2JnxCvMmEZi72fW
kbjBG7VEsn/AQHRMTDCRIHvK1gHD1o8wBojhXdyFcJGSULks30R03ao+PCU8GSB4
lZ3LCFcqifRN8K4DhjwoTVZYBvueizAv142iadGhJTeC+nBBpQShMhC2DHGlogoe
OhHkRbUSwDACsJKp/FglhohJ8IysWOcIlqVoKiAHP0UBPbNQnb11Wvwv1BaTbbDh
PAH6+l3r+OSbnmmQRDUl0abKEP1/tQzGVZgP9keJuWS0jbpaXNadIgrYuLEkWq2Z
TDwUrD1Q+pyZK38r4IrPixRhGFvTMZ9g2JpG/cRw+lEXNQcKMpQ07npH1PdOlfL1
1+uZLJwZsJZPEjMoNYPsNmul/C8v2KY9qYPapDj/sCLgdZZacTvGN8632Y8IVkHq
hgz6AsNF+wWG/W/uW2YgJ4o4UmG4XhzhytwyJxB5yMqvWDZzSxt4S3sKT96flWh3
1r40URGDjj5CqZ7e7JcJROKh3xk3NgRAa1qmoFtNQX1E5moRRg+umhlofj6vhg84
KbF4T5kJH0aUSmZlvsDjmdmf/StvATjEvyoWa1bvu2CEkLRvIC9RN6K8fN4XRawq
/4bE0+vsCbgGeR6tl2wEx55hhUU1ixyLRqcOi0N3drxXL1NiU46RX9DwudF02aQz
jaJoRN7NkcflGLUgq5Ooikz7zUC8vv+DMR9F0HtllwjHoGSl8MCJSDFR6K/32/10
aQxT50Os4WJbMyREHxbu6Ed8f+dOEe5RitKFymG0EeLUbWc6X0YGpCP1BPrMI44r
44I8GmFb9pPQgIdZ6K6rYC9fckud8fsNPiK6oVKzeRrSy1LQ3n7y0PlY6Re5zX5E
LjW1Uqa8UvAWKQQZWvE1Ud6n71xHrC/P/ZlVVzD+xzuEWOr7FsMGb+7MU1BO5aRR
pMFpJR09l5t+UBbcCDpRnXvy1iN4W8OVuNN8BWtOfbc9Q+ZwHhPiiqfCQG8QuI2/
SQ9vNW7mk98RYz1FXjFQQ8a+Jq2gcnpzFw5xbDAQtKxIMSDOYV8e6/p0S0/PsJKP
KDilcmj5jnmsAVn/kXCwMlPCYUgwRjt3L9yorogEVP6Pgq5JmsJJyZ4RQmSfKxMG
OnMxjxIjwgZoyk9YEQm5KOo8c9yWtgCXbXEv14nbAeV0iO7yRs2dbr/jLFJbZLHy
Fjyvec3Lj5VMC+YNEJb5AI5K9uDP4pev6cVtJhvyFBcV3FvzoQ9/J65thcXtAr1k
wE5IgCYQsqd2pIYBm8aMrKXl1XaLJM2GsJ2nt6pEgxX0XJXjxjADj71bYJl5PrVc
t2Ss3P03a6B+JwSKU2an8HsluSyiAcjRWJh4NdX8x51dbNi70fZ4DGlc1UM4/ftd
/UrB/OqwXohzYu24mxYuNfn1FJYMizz/5dSvZ1dy+isO7G9/TaC1h+5cpiLp+VPX
lnHXkZnOgM8jDoopNmvj1BgrNkmYRyVAsxAkajjJ2wKK07yx9Zw6E29z/i+dEyiK
8iHKU0IKbVG+DqCmCYzHuxNhDPGODj8DqL4pN5hgJiH4XBWAbGCSToYqEMRZAoVs
FGjyy1sQa/hhAhSiExAc5XuZYR79G2fFWzbLo7mYM57S5LTWyGtj0bpm3Su4wBCc
y3TwntPY03YOdTUToYjgzmIRyqWjDMvKHBKLNI7n7DaHoFAG6AGP4uRLhazMucIu
t+oXxloW3giWudPhbbkFvv00ZKImdVadQleFfal5ZfQDXIkx0qzuR8gblIjbIgC9
s7WyUoFdTbPkUIkfl38fElJ65jUO/2FGi1fRwW04Y24HFCFsjsHWS1V/ew3NshlI
Z8Y1kbmbkruyghIh5fuQkO3JNO8PjqFnvs4bihzId1FQSe3s6LLWbyx3xLqT+Pem
0s0r3Y2AZ256pzPvC4Ex03O5GNLVAlOelHbfbmjznT/U8+BcJQJAYK98Pl1ZClp8
FzXXI0HcDbuEr1vGwnlb9taKTvTVXuvW5Y/iw7JHi10Rb69WlaDU6BMWeD5RfnMn
GZUttsHvua0SfZArEitb6IzeyM1ov/U3XLKem+6BL9PPreR+qSeKWSZTN9/HCaUg
8tscPJkBX1ctZ93fNaAtyqZ8rKkYugQGs5JC8wEsv+kJgRwi9Md88ATkRuetRoUr
YUdGflNOUHpSn626It0JG8qg0o5/QxM3KMnJsexuySc5g0kDeHN7Da5RQzrSYd3k
vMMIf+IZvBVZQiIv9yDsCv7Hvgm6S4x3ayEVmlSp4OxOCDFtvkqThaWozxk5iVwV
i74w9T+Hoz1HMfr0c+JNttJPKJnSbKIKzhIrMUMkqLWpKtO8Z8Fs6+aPhcv5udoj
SbC/wbye49pwBvohrXooJOLjh8ag96VApWcY/991N3DjyYl2/Chw1pGAAFOX0zGx
26YNWAXoXGkqtU3Vliy3eLRnMXSPkzuMSEW+4eprwNl/caWrnFfPNFOFOPAsqX5u
5xA185ybOp9K/BsBPqPF2frYCrzJmb+Oo1cJPlF+GDSRXWRgUj/mrhQ1GK9AkNs9
5zDenJSDzQJA5RCETKGoeLtoonVE6jf8kxLFRm+CYa63pT9Vw3DZ221j6hSmS1VZ
v7dRWvYjrhwQbCYAG03YcLmoXTHlT4mDSWKG2nVhGvBsjww63X4fGsryW5v3Q1Af
eW95VhARHq1oyoWDfrU0vwNuXJBCL7HUDNMWQHlcFCRV7ytfjShl1hw7X1iGltR1
7V5bX1jV2kIPflPoCPeqbT/EVnc3xGymmOo7He4ArR+y/QZdeLXH1vuhzNHkhPsi
v3BqySUw7Um91nwdG0zm9kSGcEtyJAQaQZ01BdLE4/Y4AypX70XN6J3n9HylAD+W
1dP8UV4bd+hOjtAWzpq13c/HJ0UBaYFf2oGsMOerwCh28Vwr/oeCNTwyfOtQeSFA
uJKl43pp+0NR5K+dTXvYdfhLBPjNhHSVVp+C1dAus+XtUkq70evNNFCemdtiBy/+
+dx5qtuKIMGlGDAn7vjb/8CXufBsQ2v98ouStwEAWe58yqCOE1ZW46ljmUZKXxjd
18Hen03XoFEDF1Lcl7Hp9aOsuHYIXE94Dl8aVBo44EsV7dZfd9jPQC/L0eYDpJeI
R5ytIoveWIrpt8SKegJcP0M4cxK8AZQKgt0cTfCcLS8wqp7PiBN/AZL9Z9bW8liM
reQC7I5TM9n/3Qq/uU0Ytsy10k9A5GhR4h/51kvXedruULhWJwYJgxDeNXBSZpPN
Dz4IH8KQkwaVDLjQczCmgyxrNNL0eNxUS0fSB/E9wCvzWBzwwy/AFikdQBcGHkxS
Aj2zB9xbWBKVekfHV0hClhEkd5rKOOuWGV+JI6xQccvQNilYbU44WmE+ZGdERl5C
U+ZNyf7IpLjTTNQ7an25KbBHOxJY0oKmgUN8riRkdRcESH6gjrz3JSIFl3fS5SK/
mzXuTjzoxUfTE3HCRRbrCPf2jyPnbZ97N4yZfNOrx+RBV4rzn2y2rxb6w3MezV6T
NBiTKZNqSnHCpw1XkGoJz1eiMm2qSWnxU3xbUVsguj6v9P7SxaINXNGdoF7QrikI
36IhzWNDQdQAPlYJX2lZmk5QrPGloDeDrpZk1fcO40fSQl+bipZmhy+rTE32SH6R
u7cpTM/MkCXVL0XmPQhIeislh9BV3ItS72STner2gfvjqysWGbl0mw8sFOlh8haX
8VFBdnLZE0vHOCpfoNufAPdQiBkv7OXHa65Z2slzdui8lxzHxEO3q7frrHILHUWC
0EtH81oFEa/YfHazngJI143Q5VdzqvrQzBNlV5mbgvYlNNvOmGwsB73HTlczKvb+
gSBPsEBbxSb/uNRVOdQq9HZKiE4DDrDTkJ6JzG3mVwF4h2zVUCcuU1LXJU8kwP6m
7aEwPBLIQMKSm2pOu0iX7Lgqw3//OXBTgh6ge8GArt7hHX32NB0640mZU76RKaoa
HsKMOk1em2UpLWE8ycBRbbDHhur8gnbyATC7b7iwm+05jg5AibJW6Yh1HVgT5nzP
+PQhAdd1Vet9A8e9raH56pZqB7QRqyvSN9dsSxC3tN/g9P9cs4kZHcJppBlSj6vK
fHN/gJo7UYgrH/PPyMQC0zQgvk/bK202RM6t9rRVn5Fl/8hSOAMoRoKeK4uvtaho
2nqBAUIhpmfQVll8IjwI25eLTCCSrczdu8m4r+ectzpGyCGDP6Mj67WANo7CF4L+
auzf+hYlfz/FxKJ0Np+J8OiQskp2ZWCq8rPlQ/LiRY7QhSbZu1AX8ikf7G7SBwGB
e+r2Gwjx7rwh49kpr8aaVLzZUL9tZmJl7K3TO8xKT8jzJ4UgJTMtK+kNFV+k8FZW
sgGWwLCnYrVzJBKDRh4PhsB5v5HILwybjefZP+uMYXanxxlIMraikJC4FQ7MJYx1
cLP7OD1ZFBYz+rmWa49jilQnbEkDz+HYXSNSrcfrwVxX7wYt7hvjI+Am1GFnv6AJ
n85C7Pui4WWabjo9j/gzBLVZucTce2V03NrQspTtNgK+SNw5MO+FxNeROZqmJIsi
Xqp1bfJaSV7Pf2BwvZsseqwNwDcpDJ8IVraY4TXe1//j0/NYxnK9wVHhB6b5nFPg
7VEZYXH2YWoD30gUFPT1MXRz4MbH5WNUehP38AfDiLz+vAeyk5xmo8Bl8H0aUglU
8LUEV1HzZCSQPwcIGGq8Gf7LhivE7Fn7iGBSf6vUg+VN/hKjkA07ICoeoCJHfV8B
nRhL8jF83JG1WzYkOORZ3vqH5NMGGckkAORgysmbzYmhf73buZLrelvI/Ku8ZgyF
FRBcSBAw9YaPih+5yFxIXRvqBoD6ILY2t/zAys92kdZ5gzZaDWw36CHSBlH3xKz2
lB/AHumMCFu7kOYXBKW1JPJOOfaWTeXVh52+GbhSg0TFH7XWymYynyR7BnA2B8c/
MHbs6zfsesfvGinzUid3/sI3vtx8NytwVNS12WyvgMpR6mwvjGz9n76z253f4kqr
jBVlDfT/LMWANybWxDz7Js58Vx+SLXI2nTOpnEroseeCLckZoQ6b0e7X6Z8dYM30
GTyeAQNUp4iRont+pYG01J1Pkdl4xj5UC5ZUyLUyZkGaXLkpeaas1ir1DUi1/eJE
etijA2deqJAr85WwKaEdNo3YREruYlv86qH2OZy8LKY3Sn2zYcWx3DnkhowC4IIG
qPkZxk46+IZZweMYFpBBJyv83ZbJAeNXNWkNOYqZ3ABU8b4fSK5vvIaIrxC9TiZw
ldwr245kG9bXhs3U98DnMGOHebLYEN/vqszCgH4JfOWt5azyFi4TKUas+q6RYKXb
vOcXpfhFVEA9ji5nUJgvZiil1u75im/V2e7ZAJFrKyBJprrWC2kWNZI4qpCDSSeT
hkML28Az3PTQwc5wvvoiBWJ7iTVP5ZywBtDxZHQlmToV4xGpHpzYaYtmhhT13UEK
R7TABgXoEYLVq/tKSRrtLXndntWQ81ZZ40vRONrUYO3Lt7SahymWcJFzuhfRQ2aD
pedBpQ0jIqMRH6nh5apDkGJEcKD9y9tJNm0LIk52BNun8nVUN1OtT1xF3BRylRk6
tBTwXD8hmD4a7+XcOtyew9ZiTbnTFgb1MbqqsqfB8NnGl51lco+tHpNlEwFptMYZ
pUMzHOuRwCyc7NmxEr2bpO8O1nqhCrSwxrsZZJRO8n5yNBJLPzI6IzNLszf+aSXm
3GR7czGi07DRtnmLW3/oS28tzVh7sjpoGR6tUCEdBb1DkP+Gf4jwxEZBLVASKoeM
zsxmL9YeylAybilL1MSEJ7mRlLR+GatXa5v3kVb2sdX+rbqLWey4ZJfjwbW1b8Tc
QaF03kem+UQ/QANl90F7x0IAxSImjgk5zr2FM3yE+2HE0d8byA6SkAG+kEq4ojAP
iFXosqxto+w98X9Ke6fJ4BgIAMMxbxG6Zu5iFOyJg3dgsNhNHbVWynPFMC9Kc0ey
4/UaDKul9QlGiZMNddyP4YGsGfrbND2n5G0I17pHM4n1BNowhIx+zasvYaFEwDJK
sGKIEMs5D7Y1F/gvLGby1xoGTwFGAcwiLrYIfXpTRrAuhuPCWD9cTYZKGTK4OI3E
yr6+O7NyG7l3p2xMC/WxNXRXf7itHmyDj53x70fVRbb7N59/N9NP/HWLX1yemQkD
aqPhRRL6M4C9rQDitcbW8k7UMA1wio0GvSt9vxwI9wm7QCmco4Ziz27BpY+fFnpp
p96dquPJesEUgvkNEYpzp/mr4CRq84nbQ5O9yyePLw97QuJDtoEVeX5tVEr0QYnX
TZr4L97Kw4cWz9R2LG5Ag16mMufjcXvWA4RSGZ6mbgCsSoi7UgpayY5BGWCUcNiI
pnQq+mkMR/s3/cKUYBNGa8ld71UkUvD5LGj9/2G4947UCs35aUUTd8lpyNvHm8Dp
oYnQje1v1hCny0dRFFmDpNUGboNbMVlLVu6rQbllz5odnoc1nvZ8/ZHsL7HfYTup
lKRIRD6R/CZSPesC2lZIR4FryfkwH4/h5K7AH6HG30BKDIiiboCA6xGbWcwKgrlx
8FpcLX00UZht2uZ7UXPocpRGgcrELp4dAJouO+LcIcfqgYzWZb52BMSi0rITrQg1
/vRAGXHg6YbtFcYsys7FrLUuJOR3gpH/7XLDtkB7LbhGUC3ZqP1415N3E2FwLWPp
Yd60tiQfgYj50Yv+UdTkC9Z3Aqi4eCZBeNbx06i4KmvM2wtLaK8OcTzkOnYFGkDu
iiFT7SfD2rjF+ZNXpoME+Fitc92CCGHfOcNpCh1dOLX/Ji+PMTxJgEiFFpCuYMFX
Nbbs0P6rWDaD/PFNTxWNi0oP8Mtwabj6FxRva0VFo8ONOIwocCDogMAwcfNQ+ijx
iI6XXTongYhnu4jp/pvrA6Bbn8dJWj+8ITFq7VmLz4MYl222UPLiqlWfB6LCi67Y
SaZNSzU2MbKymV/hO4VnAuwUF00gxEm2CnzEDv1PtIqZ06BY6bV4IgTPjDm0xrP+
Zc8A7YvVwOl+ewG6rrw+nXr+j3x+WoydvK9VrP4KjxHfccHulYhrxf+m2TIn6LZs
siEb9WzCYmQzPtXiKi7Eg80mrkbwurRSL5rTx8JBWX0an57dJSCZQE2IaVGIVqQ8
0g3LEDt4ZPc09xnURNlFPkWbh38JR6ikTI9C/BKjvX3lly2l9fUx/ghESGOF6VKo
i+FDkxFUukUZvMoe2DbptUHOlVlUpzm2lhpXgyk6K84B9uioVAe0XrUZelNUgUzC
YSYiBd5mbHSoukVqcZIQidTjVuZeoEHHFY/ZAd9/e299tfzjTJduOHuPWirC+kj2
iFcFFzeuQnbdIwdrIPRS7mg4oOlOXpfeQRtwKU2pjP53pMgQl2Xyqn7e3Rv3HdYx
qC4f7rEMcJY6jwH8YzteHCFrE5a+NDn4ogHjQ9CB5X+qRanyiNGKIuy3SVlpC8uS
CeliupZuCd0yXh/88O6J+flmuBkJUyzS3WHGp7fTvuQS0/exMcinPnr/ztYrPJVL
7cizR/roUXJ2TKvnjMuZxr3+512WDKzcuDENTzaYOWKH1HIFgI7Jk7wUM9qRZaJD
OKcwuqfUwRR5AQvXbj7oW+mCoiqpdkv/RzCIu98yJ2EyixnEGyMWrSbzxPq089uu
gnV2POQ/sYZoeIQfjZfAgt47MfiBXxYfeoeGx+YCf5uWoUHVtygfOgpwPGyFpMT/
cqW7B+vKfLp5jFXgJK6GWgtcwTW4MZQMkaq4lCpq1o4oKJdElqJ7UP6Gon2J2pdS
5TGikuiFF9LM/3JtVeTj7yVLt0+G58jhMasiDJ5rKJ6OVXKVETioJg5DuhXAaZsx
fzWEQjbe9SJbHIW3TkA3fCLmfnk9KOctCdBbRQeuXNlGdpLOmy3cDP9ZRfF9/5Z2
UUSY9oH5naW3CxRUX/Lsp7OeuV5ha/Jci6MqrBJcpI/6VatZSlc5+lRmMbMbrX6z
hN5hS4UkaWMgwGwOgPXUYYgRoZRO+hHdxVpoJFFxrI8UP+IyGAOwF0Nqr9nSFntt
eKDt6nvxxu3ANPkI8vq+4d+K0z94qtDuiCJzqclfINUqslborlerFyw/a3MFtjjg
0u4zFUNFafpNAn2LkPmhKbj7ZbjiLOcciDm3xw0Ee7ZYSAc9uEfEnXbarOyZL/2I
2QPn7Vad11wpSSKndXwwKgG8sozOtENDgrpuztZUsvQY4xjWDYCAGC+883uWfDlC
WidTrc+OhOKLZW1Z+p6AXit6D7cVsVx19xWv9wPJwNNqIBVtobAjB6qVzly8n5eS
HUKQlXdodmvOX1p0Z5dSejv9G79OoGT8dZ0UO1Kzz/d3w62rw5jePQEc/55s69uM
euD/m1DTil8FgBaKjoEv09utj/rv0MvRGW/8i7bK4cRDTHCE16HMT7lTCDgbowNH
W1H3RT3mQguJnFnNOMlRAD+EmrXZffDQIz0aASu9jHC6m0dTORomNu16uh52pgEl
uik9E06KQRAmXJbP3SJoA1Xve7Ka5LIdedJfkZvKnCj577SogM4YTfVVTxwqPC1U
RoAXmbhwSPOmq8xB6G64SzPYC7CY1Xe80dbyKXjWvaecBIbNqTrOMuP7zX0Vh5nz
qNmNo4prTCmh/n4eDeHa0h2g5M5pPFEshzMftNfgWP4moOzw9sl1hdQMfPD/LrPb
5B98Ciq2VRO0BmzKJ+a+TYh+CjVk3srY+RZRlqMPxHAl1SYbfoHMX0gw5V6EPsQZ
vDrWIs1NUBOdUW9AYVNanYhvSKm+st+wpzjMWIvKGqKHEuw3XXXz5DTgB3GnbFFw
xl83iKraIs3ZXgqkHi1uYraJ/T7tunQ5Y4w8mhwooJP7UYFS+qbWQhpNxX6ndv/v
v15Euo6n5HEiMACtpVHe91jNFKMPf1Eg+O18ICDYdCWmYC5IGNtrXfDrknXWzjaV
PYZ8FHtJ7TgkUmp5UZgdCcaMHBecrVjyP4fagaVS9DqTi37VhufVifz56qMrMAHW
mGDkoGhj018o2S3PKAzWbY6aDH4lO2xPOHbnq8bnKs9AJ/msOBCgOe6k0LUq+eax
a/W7t36WNnWUnCmmaw7v18/nRnaZjtVd2UoaJaa0yMBUltjekfPeZSxdkasSSz+o
Qgpl339MTNuAKLevjejE8d/LzQeJDZtlosA0lAP3Po8IBrnV4gQlOxqwAvoKXFek
IUWzlbPSIHMvR/mTeS/1soEu0lMussQdVipXby33h/Pmr0xEkAv7amfDN/wojqw4
6cU9c0HZusHLUn9dwgE1KSzHyPBj4wutr4CIuKyKMcUTSwz9tRetqieFEJYLs/qL
L9zPNByUfImMWDICzPM/N8F1lMCNwJEhwKvdrSgFr58nz1nHeEwzFHSq9sOxpSJD
zJaT9/P0Qkh1fc30PsA1A7qKLyGYJYFu8p6anXby6Fpqcqd6cRPna/YAHe6EvtJA
spdOqekXSVCffAc2oFcWUmCzIqVPCmWrfcqtcJ2u2UYrpjF5Fo4nyXaT85Bmvr2m
7ACBXt15hbFT2Re2+T8tVLy3c6UMVNVn/6Whc+iBzh6uvUqu8E2LefMy+9qqKHco
AlPxbHH9h7j4s2lrz1SW75AmsmeWMJQkO8mZiwEf770u7/3qZnKNE8LF0YC1FmkV
x4Vlgd4GLSyaTWSQujDaQK412yt0BSrWweGGAOO6raV3EkIWipQb5jTJjN7Pqp6v
mPQ94mylacX8E12SZcT5xgwmYCuOa+Y+yAyV0k5CrB7NQNgRqmY3loo2lmzgtWqS
Xs9JqgmMsVuqJiKKVOnoQIJ9DkOyveezuPpU4/D+xa8UtEnJuWW9n20BH0ujWKoz
3REygqo+HttzJFLlftlhhmTb/z5bKobnBzftNNJIquVw6i0dVDZ/4YyHDane1BQ4
PNYps9wnR7P5GsE/w7AvnymIUq4WgWjl4Va3i+4jYmkKNUYSyG0GqBqLltrG4ttP
rNjYbp5jKzk2q3d74oknjVNrxydLR9crxHW7gzrswWPApYtzEvEs/3FgIOJc4+pD
ula3D32UVcimN/JP/Vk2hFsO2+6gWac6I7QVnQyZXyh9eW59tvdhQa4lN5VeB+Wn
XuXCiTQsbNXnkf7NRgmqaR1zVmgEngYVgJWMAFIfZmQbZHerrvD1U6gnQE8FAdbp
8NClP3/wi7zc6okqBr9b2PVpoy+28TB7tXyql8eSbdPNZSexpCn8mACkiE5eFbEz
0+TmPMV8OXmgxwWiQ5nv2TrwRJqz92Bds99gFR48hSx3yutc77gyN4ineNKZqxJh
Jt5Hg3o1MSR5r0rPia1XkngkAig42Suy7RdihmXoHBmjqalEExYIwbIHLc4zIGiN
0NBpw8dkESF+DoML8qpALoJGHqq5pXJ5f5S0SuaBL2iGK1Xmm/OcWnH3qJFqKrLY
Q/91QD3Evg1o6exjSq/PG9/jNhsLr25y/UD7d4oghRxsBV9j1Zak3Y/Y2I5NlhJa
4HmhSubY8sQk9eCDVSpQSUCxHynOoY67CEQn5FWHYCvmSv74svEc4ZkpjnqtEU/k
bBDufhcJAicpUQsxSPR3uwcR/C0n7nc3TWRpC2hnJ+uj1hQjBMzPGvjC3qHQUgjY
jMoseAJEnVLa04zjK6CnDTTjnJmKXoWgifjtS2Q/WresdoDEMxMduiGOpraNjDz+
5kAGE66PJVR6DFiQTsYRgqsBOmvE6UVJsyzcCE/BprsxazdQSl8sEqVaMF4QVH2c
y7rm2KfXrJTg06XnJLZeKpQYJdzL+CkPpS4RL5k/jbWVZ5wmYrQXxwUFAoboUSHX
+SHl8foh4i1moUZBrQUEtqPho/nZ7XzvnUbLXKZFa2b3M6L1K69zHoYoMz+HPZIj
OytaQEf02IuEMCPGZDpC15832+kC9aC3QXsiNv7X9EHJBfe4wGvLv8SCkU2toW3c
PDBVQ+q2XqTjchOHYBpDmt7xPRWwyH8xMfK5lJRCaCkFwJILfGgbSrOko6gkz2Ip
Wwg3H1fafVZAuEWfw6ia3/vOLIsDJw2M7LmnfAvjWB63Qao8RhAx5sFM8lSxc5qa
PAAxtu3HQYSvp9GW7wOELuUvXb5dww2ri0tsBslKM1qxwBLG8n5TFlv+WeyfB5vz
tTXUjPQcZMTRVuGVEY6Yv9tPfB93M1jLStCbd6oCrlGqjsJObhsg6lxAt3ybCR6N
YuPXObFr8p5PBJn7YEP4cBwgVenF5tRVAKb20uoCi9VVd4xZ/e1uNq1uRm4rd6PG
mEtAwkd81nDIGMrd55d3cCFfzxcQPJaeD6OqVoewMnJ1O5OrU8ged9ilvmgD1wYZ
d+GGbUoRY5qM1VuS5b9acBRaTbw5isOWRsXQG2vJV/uDSFOUlXmxN2yrjk0qpE/3
iyTW1GbOXXNgaF47JiR6c+8XfCvZ1gEFrycAw7P/MiXyk4wX4Uy6zAQ/ZJuZFbgo
83ZJOZmMEx805J+KJ5Y6peiZXaH436HQCS2I+IHAx6O0J5Iyco0fJT+9idCS3VCY
a+ZJt7CtI1MBeGOrPbH+gVMtrK9urgWJYgAYp8SBP5gE3aNsmrim5xjZKgihNGoO
UQwCy/xHt8/F75SeqT9nXaY7z0VJ9WNqHNxTVKAeCO4yzEU+K+LI0hQjnT++Fy6M
Cnb1PHW9wPVxWbZXVqvRcgc4m62jwzT4cmpZBwGxrvLqHT3JXYg8TVpOvZgXl9Z3
RNYhVjIDnjV9x57SDhYrLZmLk2rzCVRwp1Spynnx96Z/b/vG2qRMlbMk6oh9VmQJ
O+SjuSYebjHmhx49oCheIszJFXVnm3NPRGe39CixWobve4+Yv5a3cFjTfAy3PC+Y
5lhRHKzR1+MNVFUb4VlkQUprTMmmuh1Xt+ocWKAjenYdhRM/SaaojEu1EqrfuZlK
NZ+AvN3CXUnH5EnSfSj3tPPq4dxZ1luaOFhs4BP5jsKFt04Nynjpd4MEezRIEWcy
pe/tI1UYnoXG9RUmxV9TOIBVM6usyOST8mHmBlZPvM0Surbka2ka9ccd+XvOkohP
EDiML5fxttUsSDjRLCLj3Rf6sUxpbxsVUYfgczHqfPmnNNEgQ20gDPsFDcbpbJ3j
jn08creZMVqU3IcoeR3IaYtnEsAA2haHBK4bx4gWhd156TddSDIZ6KRoeBng+cOg
6W+ulrEpXx9YD13ROtsGc5G7Az5UAy6FkfZxOkTYPaQziTLf+7sOJhWtsiHOgzX4
kkAF/ZkxweVMz7E4R9NxHGbXNxHalyCQyT6RtzQXV0/qwGNfB8GwKD5jCa8PiueG
wqVpcvNradIZNaK00HO4pJqVClTXcSTaEmWBTM9+VtZ9xCzN4mYOIcmi5Wou3aYM
o7bRaLdNGXJQI7G5kAphWqs/IwSe/Vn/Erk+gDuOGvmzWaqocV5LBReRPGaElZAK
iEnEbUMyrI+p6fhyyqdj1L2EPWH1i60LlCs3A3HSmOHl7NuaWPNJzj30ftHtL3zF
3j+WQviZ7DmN2tqaUfA1yvwkPIc5VhYP0Ne3qvy/eu/WA4AXJajTmjYhw//HnpbU
CH6mKtOJyJgcnmnT7rPmg9EH2tw6PFKIiF0TNmz5pIlSkAJVLEysrsbOjqFor8NP
6GdeuDNJexrP03qpLwqu74VpznzIsQJB5H6p0nOYQmhllwP/jOChEVL467ZLFvQo
595j+hxqhGmDV55Oh031GgsbySXkw0x4Lx8G7gVo2nP3OgjO/mVQlXdLnudcz/r/
E2S1bQkQznW/HoFXGDLf/yM0vvtaTEBJ0280MH+n5N4WA5Svx/mniqvsNPYKef2S
csj6ZcNw/Zs8N4HaVgx0bdku4RQTOpYsF81L4JhB870ULhum9mmzNtqPsULXqwqs
NG+OXBRWvw/R2LjGnKaH8Mk5Lj9O2vQ/1YbLJGndGMCSwGZo79EgF6eT++8X1CUH
lSyqW8/OEldIvqd7dol1jzG8uK7BSAZ5bNdxbUDsNycajzcSvD7PEY5qdPq7bp2A
uypkAt3USgjv5lbfGJ75yRLwRGRq71rWoPUNkMr4z9RE+cqugg7m7ioKUE47wJqw
O5hWmqiVyVGBfkQfoMyUWIBawWisGEQBrAdSq5encHDBBaJrHzgfBKZmEBPI533t
FMnS1qpQ+eXSOgWzRf8M9d1VnuPcHUYQw58+lywjlYcjGbGY0Xr/dKsxBwgQpwfu
cwYxlF5zdrzACWwGMzLsu37kPUeneSQB0mUOqdTwIPKg5EmCWcITEZqpP11I5W13
UMzUOMnX9x3u4oG+StS7rJLt+QLNl8FcadDFFC37btt6OKK32tfH2+8/Gv8ORrwN
ZaBaPZbxUSUJb3ZPofo87DDBJ5VxnKI+jKJZ/xuF+Uy3i/gZGacwd0UnSPKw9CJy
VUCNZP9ksDj53OqQuuIlVVPDpM3KKbuT7alBFuYBy85gvoKhuzRgXlqRpcjq5Cb8
92YqnsnBDQLTIe4iM60lmmlTNJ+HO4CDtegVwu10mNBivR9r2FQARlLAksccqQSe
DmTqB2VN3if7ATLiHUi3kNJc2nKetM2FSgt++Xqk4Ao3iNQk23Nh7g10oLEKH+Ik
SDeBMlqktbBtRRNKKJXQRn9sMX/McXpXMpu443CHv/eJh5xWYINZV8CpzWy1QLA7
cO97VpA2obI9K7d+o85/sWO7Genqc3bCpVn+tigXZ7CpigxnUNVyTYxj11tVWpFg
SGoHCGmqGdZKrkWTYrfkn3iqT6ZE9iSIZM2t3jx7r1thrDpV+8ima7RJdok/6vWw
Zf3umRhDjJrH8QRgAfoLCYYXzIsoV07CmeUDPnPfY5TOgGbJaZySbOBaQsru0xrl
KbRxHzuN0KqosO2GjE3nJh7XPBfGf4gKdbG0QozklBh1zJS1x3KEHz0uuqQMzarE
+LqaTJQCW/9ox6y1PYFz3W1QX+QDPM7+4CU1CQiaoKfFzo5yVW3Jb5Z8Uft5vDpl
YBgYvj+8f63qSyCeMIKnnuzVJ3T5ZrfauFMk3Yn+UdYCl7xn9o+6/RZoDPamPuM/
H6tlcwz2iZB97PZ8jYR6St9+jVJ/wFMekXzqFDr4q/hjZuBfBfPwYbGjgA//yEop
U1setjoP7WqMQTGip6AKgwWJ6DyJAPmEqQyaVUgyiUWJry/FEkK4/ugRsEG2xWWL
Tw47ea6FjzL3H0UuI5c5ljbe3yay1oY2w1Vp5133t+PwPte/UWhI3ecbOg3zVzDy
0OanfwGVSSSWCnrXgz7FZXG/DrkW01YqF+uXCa63I8j2TJdpmgG9pVDsGWHYyp6V
ieyBpiartFawS62QJJgD1BNePWJt/OYq/XwlQRRulSs3wNPPmrG0hrc9mZOLWaVd
W+HfWcbCPGLx50/7KKcGAEA612JBNn8Biw3YpvD2Jjwyk5khtYHxVbC6usBB6i59
Js7i7NXhJDXp0o9fKShVqgcBFMDUm/rYB2J5iT96SlTOtjRmu3YU1rXWLcFNMgsr
2eMqWAzhgO43+EuRhL3skXUgjRzOqIie9lKwuCLEBVGemsiupdEz1OLirdXttgG6
tMJ959BcPnXij/+DED1tafRidzDIUnbZhuE3O6exJUQcoyj2zIVB6XTOPm2Ve39N
E9Xw5sYZRIX37mb5tAdvuHg0h/TXG9UJ7rRps9xNRfnMo/09+6a89BXcKwWNIWfW
CplIznQaDNcoUaNjXkMIDw0B76JCMsRFNg0lxWybLHOdIvdHgwyyYFiaPOPaa7pQ
PG8nCK8AY0EzvPoUmOkaucUCl6UOktv7XnQDAQTIKPWt4ytm7q9lkRcvaUd+ILtn
LvRu8lSumFbLyNf0T12hlGxKxEN6cC84WXBRbI3dlehEFrq1Np+DaD7OOIiNo4qV
xjMqhkGCbjkQHPBmTt4oZN8DT2mHCWoYSPM3h4gYTkqxHbxVIwaYw5gDa2OZJq0Z
KTg1OtGay5cDscvoJNJgiTLaMWp9i6ePDaYRPsrbteeE/x1t2L7F12XOLtBRpYVM
lh6sViBDpauwEZzos5lHjLS6nVH54Z3vRqOsZoJpz4HM/6FTkzeFRCXkdRlfM7Dh
+WVP20jKgGGR2z4yx7tuOopYp0ei29jXx0/M61+mP+3TqHXJZ69T8xI3rUA0iAeR
BYbp4um0tjiRtSKiYOf/7dKZmaybfvbsLMw0GGPS83nCauyZiZmGRo9CgBGvYYpK
QII5SacPm4QSs0JaY+Fm5YPViZvCZQL+cE0Hca5pjZ+hBJuWoHSmLMc7wdQ65g78
H+1TC9KzzngL15ua1gKj+SUImlw6FV7lxWx7SxXlIAlWEBEJifbkhNn7CdcWY2rC
BVYItmQehZsERR8/W8a4DfDIIZ0qmKuSR7hXpfFkJmUE79AqaAEjeUedUrC4x2uX
4gHZmZew6FrdhqNvA0aClzr8geQOAGcGDGHeUZ2pcb/ra2maAZHtjmgAtH2OHApj
M8GDicnbgjZc+E3M8IsVlZHJe3gIpnfRWDLQpMm5s73xY7H9z7q7HWtZt/FCS9H5
b/CskMCfduOgdv06e3ygMUSd7FyR0JWqk5zDmmzo/5rIZIGRTrydmtXxKcz3tdUz
P4t0s9jiVuxa9Vr3YJWX78XSmQMWBZS8qOanMvRKkaQsW1k7UqxaHDbJTtXbbtfZ
K8gQB7hxBRfD9tSL9gP7tOmSm7IdJO4+mcUhVdcUmbr/1MaAcK+R+9hYEIuc6qCx
1qP16ZmN/LC/Jywzbqvz9FtvfIEesmVzR9FmLcc7DTCObrAkxs3MpObzjU0ucuyN
dLB+PCXpL6iBrr7NqeWyD5/KeR1sRuWvBUpBZZm4nMxlQ7gq/tYr/+KyGdH36qXX
71ekLxVtmeuWnQRhmwQdGehDeOAz9znWIDaPuZ/k5LEwDf8cpQ0rv1PYspuhIzYv
N/1RRqjyxyX9dSN9RTsOmSAyhrG6HNjqRmf/6+1GZMBhm6Xb6iT7oTqnEnld6mKo
sSMXCIRS5ma/z43WaZAnfkKTpsXLvcCRFPhVxVtKEZmsi/la923wxZrhr0Z+Gpyx
Ua30VM1Fyj/2w9FrQ1elfLA93FNOn3+dbY5nwGy0hZwgQZ1orNdKFuSJayHSol1i
l1Dum+3ceqMUE+yMJ7sh5d89Kv2bT8fYIAYuB5fXwABFGOboUO064iHGLpnn8nfq
KkULk5z1IIfcIIOBFooL/Up9SRPRw7Q64i8mZflrWw7V/bPTV7xkZNhiXxRd0TCh
Nk92sRhz1RJrDqBilWjI54CO+eFgPW4Wv5OcSBV6bmBoNAzojVlUjuuhhvdBeiqZ
5tmVDWTg/ZGbbk33pOpwBBvct8djLrk9UOfDfMJ1vhyqstwLoPZouk+silMysIdM
6hEhV7otB4cvhxFdl/3aAMH8gQ5r6kAat0WFfUm6mCoBggNIBW7rlpxfKlPlW8ka
p7UIdhESL06evTXuyZz1zDBRmLh/Grmp4YGTKtVgUbXwhuLpc2RNZnT9Vvm3Cx7U
ShciERjaPTpSlULarzRAFpwfj7Tsu3rnwmyNv1zU6nB55FlE+6BcIvi6pbhA3beM
CqnaSS9ypcX1pW6uzrDcCefYxMdK2D4loyVkaPgatUS1bspFX0/fHa1XlGH9zYjg
qs3PRljvJlwQEJeAYffPzIoTC2yhQaIxwNPEvk8j2Bl+q4QFHSy/RJQOzrmQQ5Up
27eQK2ZwtSvgXrPtZg9vdCn11+/nFTjUHckFQ9XfyFSxN5zQq6nP66DOU51rk0Mt
QFTYOEGCc63THWl+oHt5/HWo6Nm3WCH2OK8uA6vPeek6yUjrh8g1LHiqGALira4y
lGYRGzhC8UThZaFq1Yvc/5vvcrq4RgzJUnpYeGm555Me6ADZzB7Qtf+2YXXcKxhb
V+A6nvMa+f1MIvqnav9bJQC8w0IpsidmjqF0fS920RtQX+JgX5iD3teBkqzRne0E
lViQYPBeDFK3pbL36CylEHs1hWFuwGblulSvfa+kj6HR9JUXeTI7C9gFp3Mkdi8U
VjkGrANg/uNa/aSOjRjsIb0A3N8sIQF/A6O3gcCWESQ9ATJ7dJVy5awzjTxDeh+c
DG1Wgbn3/T65ls3rsDViXNGcnCU5iii1dTNaXG95n2qONIM2iygRqp93oO1eUC93
YLCUXVX64SqI/AQq1zPe7zcILLyr/kNv9KiSlWCeC6pp/ZtbJtQXU9MtVNDPZAwO
jrAax6WIVAyeCOJLumxnqShH+hJpKWNfF1Ia8k4ws5iY7vg9rnlholLe65P3Ltoc
EFU9Hc6vgyQ2kME/Tv54ETu4v+d5AC/Io836HnCnL8CIND3RmuCqm3pkRSDllcYZ
XZ4lqAwxk2d/gc3R3nueafjVXepla/MlDbyHOlH1T07y/Ix7dYehgyN/80UeVD7A
oJHh3SghNxczW4rpR+SMGjPUDyWztwMY2tN2dngTuEQwh4vEJjw69QdcZmW2ecRN
apF+TFfJtN5Imr96HRcH3n8ikMVGUuB8xo3e9uyf6pkPQeKrWAvRq+Stz1l8oOtd
Q9hI7GUznODmoCoCInjLxX4XlBLVOE++aF5bcjuEMol71IhVlDwd60xJDsJl+W/Y
eeoye4D3acrzLf3OzIylIRI5nHldbEUftvQ54jHaK38Fl4JyFUoHw6XWuKtTyp4X
CQQDK55Nhxrz/wu7niupmxp6NOwUHziXLzg1VdFHRQ19bZ0ZZZsh05vVsWkL4kLk
cIr5TtMqL6+qeKqDGfFJUJcd1f5TaoTqmPQz5JhaVj2lTeCzfmn1dJZdpAyWEZdK
kGp2GLaE6ihYlF/Di13KApdrLZ7WpBsKoKa/fRnLWveusD/OqdERbWSsjuKkPmbJ
S4ow8p6IcBYYkkt3RIPu7x1aTHr9s0r8YKMaP7ThxdnSxDwJYNaeUJLsxFDJbo+I
E3zNbaHmiwrxh+/1m30kcnpjDabHm4lQgLTKz0iCOpuXyrPf0vsStlXkb/WM/pAj
pKMWysDHpOVaQjcltOMBJrltc6S0hHwIzV+Xnw89ml5nvNOt3HdPG4NavZ+L3uFo
LtOdlt9H6YdVaAjcmPxJiyZOMqGigQKfiJKTVWNEuylu/63LB5lDysxQM7CKShZq
xn4fszGA11UuaGtN6owATpg1pXz21NDJFR4Xse/q30T74tqrPl7KR7FjkTEKxcJb
dxdAMWggODQKCejOJFIbajr3AeK6rl1FvisSMEFnYuSiC15dT/vz+crKZwMUW7n3
XNAx8RS0Je0th1WPPAhQiIVvlHGfyUYUdW0ZPysPu3Do9+810354SrKRHpThhS5V
+BUfgSLx5sB6rQnndRroUsNEik6hORY1PbnSAvx1oRFw26f1NdE+9aJH8T3MdgBj
CDVJjMWwS1cCvxFWakrcXq6K7u38Q0bd8nY/YE3W/qkvSU74rgP5U1RnKvCqrv6j
20sYBxMmDGoTZu3XKwyeCJItDOH+Ny/Jgm7QXwmirAe1TzjdADLUS9JJGNUXMxoO
POpjGjSp2CQI4yo9UMJc2TEhBeAUZa0sRyRrx8PUZu2IdHZstpJNKTz0RNLrcx4c
quwuuK+9c84iPLTTJfWwkVoSFndSqmzWnPK5FiPzHvtOk6EFQbgFK8SEJ538ComN
084xex6ALUjVHSamJEvby7DzDqpSRYMu0P5F2IVZguzBcn1GBo88qaPcjay4Aog6
lZQ9FuKYXzpN5eofWvQ+9BWVWMLdY+s6o+XRe9XZQrVhAmZSy3GZepb1737nxVol
X/K7ZaE+uYwQAhsD/Jw+IEBNp//NX96GrG3qsh5KkdCUq3Vc4lpxxII42+d3EXVo
EFnSSvIUsI2CVrLQ+k+AbUaaz35Mr+Kw1vg3QvU/j7L5Wsm4eOwDh3Its/hdGnQa
HxnRX42REgJ38GwKIOs2QGhGJaUatYMIsLHCoP3s5f1tvo+Ib+xOHZ9D1B6Gr7OA
ihTGgzG5FO07IjXMIMC82mrOPr9yCy8UYgY9hcZAePKH3CEk5e3vNyQk7Vory+mL
1nTwL0ceF7eELdZyhl7BKyLh2Op2lwEaBTipWsp/2t7NE4u+d8zcpF9evH/zYP4m
T7GNON9bg2UVTNJ2f08ADEmITjhPWmuSxhEozzTmL7Y9LVpOwvNB8DkU51K3eyAT
trl5mJbOHFfXPXNK+xSdq4kITth5e2ImowAZ4iVJ5+kdHuqyb9yOMF7yIMChn1vs
WrKJd3brpnyKvvDKw4O25aWGy7Nr/DtoftvEusPaQhNbYD7oOPlpuujVtAhaA2No
CwOjrU8EOV2cXXNMKTxzXMdwL3UB5/C9J7nbsPoAYdYwl9oFNAey4U4dLlH12izw
1G5XaWiDSfe71LN7PojdIvqp1IYhWOrFPajMp3ihI5hskpIAtLeuzB0U0bL9vW2O
z5xS8HQcrILUszfL77F22Bkwl2WYZlPEwT7G7XhFdUn+r+yFhPmi+jSrN4//M5IP
qo3r9LeHXhS9/018ox8bexQLkjPozsp9LZydx+I9uZ+TXXz0RksqDBtYoSNazMkz
xUubZ8NCDf3fTTxAD1wX3BDEE1ZLLfJ1tdxXax+5LfYhgAQN7XLYV6WoQowFZpQ9
syCcD93jGMnQJD477A6hXKESTIZ3pyg9pxdhYp8NSq7sLUULwJSq5ewrDfB8m2Vb
yBYAJYStYBNeZsIo9vKOl2TavWqiGaSmlYunBNuZ+VZW0502RbJk2/+46xZG4N7z
EhgdAftet2y4+s9vrX28F4Q5dqe8NbWVVJe20MFomvhHTj6QEUfdq4J3pI63BsQ1
hH6N2+og3jf8itcK31X669+zIN/FZpmQi+afB4HxV33omH7bJfcJkHbnCNhMS84n
cOjufbhfPtWuxXfaIFs6MDRahRFtcKPQIz/pEBdDWCmF9ZoPx7PPNXRnbqpqKQil
TAEcFiVKSaBC5ZK2ZBP1v5kcc1lF7PExBlcRwDJv9SbpRnhQLiSRvFNi8XeQyEe2
GK8Qt4xlnUDLX9HbxxZzZXG5YO06T+Hr1R8tASMnOz6RB2fX7lH0vJyQjTGQJwDE
JIz9q3TQjKPzYJjy2EVs1V8P9C+7uW9sJM+LfsJpCTOF6HIdFwpOltE7EhgGY0Cx
sENWOTUeiRiw/8s8MeLmcZt3dx6Awq8jvmRE14849wWGzgW77SU8cSVtmQfdhRr/
/T8OfIDet2QDffi8BsXwV1VYyk5ieD4AgyQlFKtLc7/iO1DXFXesrjZiJHjEZmSH
8QeHTNCH4VoIP4y3iyINtUHZVqr2iKNjf4QqZ7hXki2UDISAC4UZyizLQn+fkB+L
ScjsVNJCisUPtjliH2J8KMi7dhJr4OG3eWg84ILfE9jz6C6JiHfr3K9sadZtTleL
xITW4+EN4eklk85bBeEGGNku2X+cs4UBBGiRgzeG/+K73aL685rp8qhUuEvMA7Tt
SznMw2MVo1L3fsTIeJNvSNQpo4SK4tp5YzcFvLbZmpNUBKWHx5jp1kzgcqzhPZjz
jAbw07XtGfGNVn7KuiwThG8yQzZPzw78LjcDqBvpOTm6HcRImNoJY2yEhvKSdSbf
wMY4PlDUwyQXIKI08tc7lYKPH1oPfteYJ2lJFNpMqVdve9GD9a1L5Fa5SbkZBcM3
emR2ksw/vMYNTaovCGu5XWY22Ms7KoAuP103PWVYO6WVIVNC+msqyCK6fz+6BW/w
4l8q5sQ8A/x73gBT+gilz+/xX+DSrcb3DswzHbl91x5ahgTUIbQuWYlL/jIYOXSx
66Ce1SaNIZuu7nel/gapXw==
`protect end_protected