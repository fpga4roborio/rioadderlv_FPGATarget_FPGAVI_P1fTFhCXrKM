`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
ddtXksX2+yylW5zu6QL2Lhnb2d1sD00763mmSITNX595NcHTEkwn0zB1Dry37fOW
FufOhVzEJp80NC5qZ/+F0Vk7Ik02dIR0elf3clrjeJRK85K4e3Hoo4xn7YbFUIms
l/8VZSb14+JVGURjfswrIyCUotIzlzVYZ6gzoZwDXIi5gQIBf/gI+KxNXPaKV+PQ
Ufys/12rjO6aI/pPlqSm0hCvftmBcnezN2hk1UeXgOIuKZnogjOsf0iJVX2aOOWE
6pD/psybjbnsNB6kH5uFTA5frkzIzkzl5d9+YDm9OyC+k84E83I/7/j+rk4L2dah
QJOvksSIzN867/4Qt8qYTQ==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="MvBXkzurAa5VTw+1JJ70nePUfoQXBvZOku/SMmg4TwQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
oRtzZL4VJ4iwysPsC8SXYCzXS8Fw2gtZTOskLcDV+1B9Nzn1zTyNtlo6lNICRmmK
ZRVu2BmCc2G+fmzynYlNTnSa7C0Cuel6FYpxCBlOuk3OF2tzAmLAuDyOH3Z1Yjzk
a0aHuoCdIRKv7BrZCdALt03JeUmXKPdOmIlkVGFl8yw=
`protect rights_digest_method = "sha256"
`protect end_toolblock="Jn9CQpRhJt4rnzZPRk+dOpzAubz7omckX1MrFd4p81o="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 13456 )
`protect data_block
gD6l00tciPUa6pDNTk/+t0OO0nC/UTtBwLB41d4inuAUA3i/ALrNyoJVcBnAmEQW
ptbcNp5fxEUJjnOxnedyZEuEBxWRieZFQnkRdF269oO9x6CJgW/fPrRdGPKXD3DX
cOF0GOL5KtGFqfuQGGQqCwdICMZdFZisikth8EMkoRddoEpghJH0ck7wwh7xn4Ng
6hpQfcERJtnx+knoScLzogXPnUMkKK87Fi75HQjYM1RUHCUcbp1DorxgMg4svnfZ
SBVUs9JyNDZHR1iitHX2A8mtThIT3hg06dJ+ohXugfiFQgBFi75Q26VJnrpgRn66
TQrveZeD0j4DdvgUmi3eOpynS25eZEQKWHHbgTg3d/sYVgUdfceWdNzaJ+esjhwt
A1sdB8586opjIiFGY0EieC4D7MjhdPCR3E/dTf34lN3USo/pchjgpQAjBz0vNiKI
jq6nWkjHdGEvsWG4qd7S0XaJjfMwEJHD/q8+3PEY9Ll7Fz5vZy7b7vsAJ9zqNqDe
TEBu8AKmd0X9f8ooBOUpiIvb17AAphtJgOnagOIQtt2yEb8lMQiFV8vKtpc7mGL7
+oNlFXelo6wHFFennSypdV4HVBArFXgCjyjP0sfCkoKhavmW9JqY52kfPVE7ou4B
dzXxGkfuVeeSOmeYrbqS1cJIWX+xOUDNu5DNlCcCR78q3uNEp7h6dHG7Fs+PJMRh
rXPJ0yUHCcUvC3BrcN3QbEShCQ4W6A5vD5dgGgRk0FXQsPjgJA7ABRC8bnNoTmOF
L9kor3LyKD/r20c5N22bej/mdqqOsqIhUxcgJHWs+yzkcMgCrI641zu+TzNuVRe6
Vpy5A8OFDQFbwqxX3wBzFT+v9XguIFpiQhSNJUR2eliot71YIhx9d5UxOemxv2xv
RlR9d0bfdD0oxm3l1nkD6bLCv2vLB+zkXiaC95TGP704X2Nod63KR5voyQbXKDKu
MH7mQYFDiOA/Zvk3Q+TtDUoETbbTa20pkou16L9XWXmBM+lVq1WvPmoC5crnq0dd
+RoRxExBejYSkpdcD6U8UhnQq/2T82X13eXnDQ5Nm+t6QZt4ZwllpBEVBoIwpC1n
LAiiDnzG/VX4smcZFBlglr7qcyvFHM5feupBpuIzG1/nXorACxyUhxOOWXgroNiI
J+S3jz10VfYvcdFHFX64oX9n5vNwfi8Y8WKnTmtvoMKl/60FUUDpdqBhSoj5DKtI
LD0dMzTvbOrauRp+PNc47/JjGuVuDgVNu1jhIFXHXMW98EHgaYuP+YIVg8wbFFO1
G3fHyQ8sVx1Hw9momRdW30Wj319W1fiMZ0yaI/hLx3WSib9yrddAPc+y/gfYAjE3
/QNCFoc7B5Jk7gHjrZrbklDswMkSt2BUpW5wfKSI9floz2orU4vlCQB/5IXUBwPt
HZtoZZIc4fX9rVRxsntpZ/W/+hl9WWLYi+7ZNEgyOMayAUeTxkzX2dXMj3ArOKel
lChk0tPK5ntwl2DvqYIcN9sBxq/kKmPRUdBKJgQ5LwABJo2T9WfMnUiItvSCFDH6
skoMnrBXwJOEbnp9aZDkZteYt0Mhauov+CyLXEGuNQs/hFeC3jIFBuxWlxS5H+2N
nDi7c3bAZzfxIbVFhS/8bO5TxizWDywtfQhPDzgmOskn8iIb4AD1cBKv4zO1uFZD
ZvaPH6icdBxZjLWn96yzWPtApSB0vVnBysSH/iQDCogkcuu5K42CyWhcV4E9KAjr
02Ldybhe3lyq1CZOeA+SLosUCpXtHyn5dH5hodpp/PumS5saK9rmQyJMCEfaIRzP
Vi2gzSMP0jsXABKw6jI8McOG6T9o2sw7f8Sck0YGR9xaNIPQme2N8TuXdbew8kMV
W9r/+JNYot3ZgpXqwjwdXFVZK4qWZd2to8q/DXp3/2G2+kB6zzuCObaAE0MzuE2u
NRmSi5ran7Gv5ObUfj/TQWjXfmcGBnIQ/59K5TJPfAv8Mv+Lg9bThj9AccClZKAd
/i1WhiPW1YAqGOo5r2CBi+VVpsXGlf9AWMHraCMUESUcDWrQAmjQX+fAGgCLOg4t
2STlICRn1d9gZTwz9UziWm8eHfwKRFEJEDYNtFUq9RmdROdX7PUxBKMI9N7ttVTO
bflWlvSMc0l8LThTEJs2aXJjawqnxnsvU1kqr1Wt8TE4STjWM4UXmK1Gq3JCq1OT
y4hV7+aPvYN8LuTeVaw+2QR/Usjr8Nfw8mRVGuoT10Eg+Rtgl2qzQ1X/yKhOqsbR
8ihe0gX3P6edZnUU+Y8mNmJyVhalJmh001yJSEnn5Dat2+024WuKEfcfppij/nQP
lHsMjXpZ01RWPhwQqzAtcX80H9U5Zl2ORH8673xmHsxP5lCnsbhOpHJatt4H48Fc
5Gi5hCbg0wsyI4R3Yprnl5PikMttZdwBTxSCOpYO6liFO+KK4P3HsRWrDtAE46OP
UmIm4a0Cqr3lycHgIhEz1oQrG2xtbK3XQ2qH05gSy1q2yKIk+HvHNQk64V/F134B
weii61f59S+J7wK38XVQDUr+EkfYvs7YfLrrIxEjDdJTtgFy+uYUpYEdlPm9PZFl
O7oqsbLmG2gsvKzRheSpaqlpiv1p0sWoGb/088EgYLXkw/IQoeW5OpAv7mefjQ/3
CvXkGRiJXx5sCn+lEC3GCMv1IcXcO8m/Qn6ABYjZPjeSuYfPIY3frTO9t1DBO8s9
EJf/qDgB1YlkpX0x7Un6xst8uThmcdP2KNDIHmR6p/oiHyqwP6pfFPAcRW+pLhNr
nkGVv6HmXCKCH7UIuflAqTVqE2vt3robEFtMS795FasipoEh1xk0bhsp7jZPXXw2
kiY7NxrTK7682e1eW83PVNzX5njzqvKoxBb9Oty0PS2GDi0JMXxhwxRuqNC+vSZD
gia2UsDXCHdsmAwv99/8Rz/cZ6bQBpd+eBMOskQS77swvactW27fHbmqWanHQGno
TdZ6S9pOQQ/R9/44kXOILExHG4+DGfzk48CgTN6ZGQViCdH5dKMLni6XSpUtxHlo
VBVZAzgPkJ//LaJwewyZ3dDCUuiW8MuxDq8kV1W6UYdkj8jFsMNQIclj/YGHmT+R
yyNXeLLQV5D6hX63KcH3u88LRySGqPB8ePkUhRHNfqrG+A+XmmhvdA0zPnj0j8Y9
8xT/ZH5PH6TstSOvzNQifvmggMIIP3wvUMYKarZIoYQd7kOzjkWuba99neJmdqXE
H2n2Nm7l4bOhEjpY4ZzxOEvMlLGfPgDiSLznfr+DTlQqdfMg50RTrwGTdtaB+Eow
KPMNQwgmIVmavfsPdXlnK3r2laVfzDz1rnA3uAtL5Pldlmw93bpsk7qL0dpGkfhy
SwZaDvZA3KyrsT89uXoBx1oPRYQNueXRJJQpXnA8com+/odGY7wX682WOhtZXxZ7
8US3LOwmlVvblQ0i9TxlFR9nUOBMMqwln5IM6uzGZT1+GIbpkv/nhe4KpGBuBMxP
6Msdfwn61KAWQzJMCZJKcqTwwIdCiTqBWXwu1gzbMF+k3oALN5ceLvp+oPRSzij1
P+o2R32GecTOVtfWmY5sFiRjBOAmp6n2+yxHJyAjmenV2V7Tsm0EJlGPr1e3ZFsD
BRSfYSDz+G94/q7EZZsEHIvkdS5UYzaBiQPoXA32YbXs4qRdp24Bn615JhDX0zIp
VE2JnlDXoiZCBZY3Np09pfcL609+NVcMKmjXj0KnX6HIkGvocOJmsHOAJb0LUSel
r8PYC3TmRl94fAmnrNMzjz4BrQAu2DuJrgi5IZfkhuosQfSkCCac55/RoP2eI/+l
2qP/YnDQodiGLiZiJeKCb0aOJBWthQghZOoOQVgf6Iv8xOV0F9jmoPO/p5GurcRz
Asa6pPDs9Bjz8gajZIgCGalawHX/xuI19SU9kg/TPaAs3Vys6zSLSzaduKfO3FZ7
EjzK7itgE1mv53nNpxD9l+u4WyBNj745ZhUqJE+TAJNp/Vyi/m9a2Jp26DpKHdjG
nN6ey8cvy3jjsWmGO0Wemx5auqjCgKu9owOO5O3l0/ExwudZL3oWz/XWO6m8e1n5
h2qzx6lW13gtuVED6pyy9Uh2Okyr8UQ23zwiZAQ79c2JfxNN3m2znO9I0zKqnNAP
VTIzgc9ZNEXXD6FMPiPIxsM8XFHLn3U8Q307eQ1Y6PfNxqQCbEOWPNRw6ZGfvycZ
pC2v9Kkk6MEOWw+hX0Ez3jd/WKgY9kkrHtw/eevEBFh7cURFERYkTM7YSIsiJGzT
cLP38gwanRO/RJ4PNO7bUgS2k4bIFFWz2lp3yYjBVbuqYkL2SqjELuGB+/Bb2FNq
FTDTi51/FYkkJQ8Xo0JBU3wgqnPbI7GjqiXhdSN6PN4OLuJEXlmRUS8PaDSavuft
oxXuEuxXFy13MLWSK33Q+M/zgiKFoyGBU8jJzeISmR70IJML+OxzEGHvW+b/T2M6
9Z3A5gbGDGTKCWlhEJ2iPYNI5rr3cT7Yh6K75rLERYbbsIuiLensUvv3vJQXKBCB
kngpeZUKlpeHs/HAFzMxh+Zf2dy2yWgQsPKNXt7bKkfTT1Y4IyDO1XJ01QFwAQJs
9fN2+83FHlGklzGwwweQoaIyiwGJSaW3158s0DkAV8jzmekOmN/ouPio7RuOYJ8o
xv4CUSNlHp9Qcg/dHdiqimzr9FCb64n7PlGkszEZj4VCjIf8s/ulORGj0H73EgGP
aa7iazUiEdT0i4g7IAj0FB3ldgyRAQXdYLJVihLOQOEnGiB5nD0bBiis7JO4jv15
fDpen/dpyXOvi7/oiJQWgrcIKNVWx0zg74lUqit4FjPn75PXarHCsEVuO/PR6/L5
GCL/MsCeUHw3Zxb1LBiH3npEwZZn/qY6/XYM3YPCFEnqhbyGS/R0fZsM4oNmV93I
wEaN18zQM84hulkk8bywkRfpy1FRIBh+wBqDDmeyuj0bB+LnLF8u+z6vdYTdQ4Sb
oXQA3+KCVJBesUzYIKuhm94c0aYI6PAmG4kKi9y7FRO4n+esd2bzO1E3ugHbzUAX
T57pm8LAteXPljAKizeYiyScQSXU5Jah3Tu0yYJbilYjc2476uGXYCHhXG2iavlx
ItMAKgC2BE5fA7lUIkcMRKw0aKo2fYtKG+qQdEW74XnaKYoKwsLQycBs2p6kHg/y
n9OqTmyi30tdDksesuPpGlQ+0aZyBCWSNiLuMbRy02it1m94IVTR5sSODXdlz8PY
/DpCI8MRbCIeLT4yRXj1ulR/9HhIZp2NP3as6XckP2MeX2KjIcSZnIA1NAs6a3yu
DO+pfZHmSLBoRjurI+H/2UaBtapkrCxSri64ohsmL/NBFhsnlQq0Z8ZnCQ/uC/SL
y28byR+rKHRz2uMOn9d0pJG90N8fY4Lowqs4xkyEsrcDz8b+LwMzFeYEhNxBcxZu
vQne8o6Cjsrs+LUcBo3g/AFknBTAcXdfIdIEqMmFiEh6D72y2KYpFaUr8MEnhuLH
TF/UrKNkMvtpRqQc7xi9XsSeChoavP2YVM3Ik1slQosAjQGCNwtYb3hRQ15T+aeJ
AaFQkGUOAarQmgcV8TTWRDdSlgcrKL5sLSaKLOewvC65BeNiuA4/am1vd+T1XqVx
DPAwYUdVIWxi7eU4pVM1QmPtiYnQXC/Aeim+xAlyjGu3FQ79MJ8/fXMUBDfYo9Nj
iHu3eF5PGSdMEtNcu0si6kz452tOJ7cP8hAXh+IKJiLH4Pkf1v6IlmRhIdz802I9
mTO/B6RuvoFp1YBOawpHFDbpmOfgRd3LNXbZEdwagHWpHlMaLg58HVYRXzFG0FhR
jeddZbsnbwSL5m+PI+P6696SEFMXEASVr3U2CTxYsLx9Z6ilDuSNplk0ZcxqB/HL
Tcr2KZlj84HoAuvMgT9eSyUZ9u+0OlmhyPLuHczmnC+73hBelpGDYetqtga/ADU6
rkid0sgw2SniH+FYSMUEgGm/FQyZNHkMtPRVsbuEy/lN+9sv0xSfzJuHZN8EehGC
2P9Gi3hQmNhsDbZuMIpphjqaVlyZBPe5BRKH2snok9q6w9CJ47Qmi7e+wR/a/NEQ
1cCSfjItrM6dKtlnhhm+vMdGsIuq5vyOwyGa5mhMcfltzdGPHDhmxpupEfFzOuAM
HQejKOsHD0+IwdEZSFzm8BjIqyUBFVKg6Edd3NERG6E9MWmFr89LGhTdFqDTHdzz
PTRNO2BS/85AhnYWZKNg091hJj8FQijapFSPmZsbCllec9o21gdTgsZdiXI4tLQQ
SV8s2QtQvMBMu6RovGOxzYvd3/QrPyx5DyoydCEXE5z49wgOvqE4vbhaOumZ9CFC
WiDQfUajITVxIsWSEN5g1JHOta52ECGv9lq+tlU1nsKzYNuse9fODJs7PPxcDWbC
v/N6P1DB0C4EzWNEV0T93KESsIFF3vfI8rQfyy4AkX1qpg+gqfbKouI1x0Tp2j+d
80dW0hgITq2zy7hrObOHXv7TDIfP4lhd6yf8pCYGt1A3yl7UQbhf/x6TdxHNhNU3
sKvd85zfFMn58qPknnHewcXTN9nFoH/bTXWQs4uvx5cJwQZLjsCqGk+/0NNgDWyU
vqjnC25b1gWAC6hO1alUHDNGi9Cjp9hGJQsCmOasGAQDcJ9J9yrJb6xoyZu3ounu
cQG3cc3lRdbm62Q+5d8XxsMOoxW9Bdq4fHVTP6phwI0rnwsokRDa4ylcpaUXVvAz
isyr4TsA+HetUIrbaHBNqQmYDQAmzunLLAhjWAf6I4TTcC0TngFJU7Hx1z8x7xb7
DVEH+P/TD2fqBpaatnEd58P3UODIu6E/Q1MRFYy4MuttRJgjCuMZT+ulLDpfSh8x
ge2VuyhaG2eDg/Z27yZdfB490B4FaRxorGkDG9xhYL9Zns3GZdRy4Ql99oyv0u8d
HRlF1+/77NkKVhN5ye5+8iiynrIhvX6gjEQCpHEZiZ/bVEw4aS2+WIXQYSMy6fPj
F6wCHTbDOCpzNtdAsYr6+ohtJaiv/sc/JeA91I6C0j6XnsFcl1ZepUTLojOQTByQ
muWmWOCgWBtVVLfxiD8t4zidY4RnihSIoUEkkYxShZ04ng7fwELi2M/KY3B9xIbA
rruXR4D0J284kdCJGZ/WXBsgdO8OAmzfqG1jR57D7NcBa0jBppLG3bxPmuEsuifI
mmQoIPre/8txMLlAf6lathyZXqCZV3m+7G4QeVIeT6H/b8cbGBS6uO/3eCUHvsZZ
1dHvkuuVh4NC+Vc2t67d9hJlTf8utfC2gr3ORDookeuJ8A1TTtvcKUqhGWjpIfRG
P+8ZE6d03seyDVLlhInaxhBVf9mypQTWRhFrTUSG9QiNn+vwTHHOvl+o6dW4fE5W
19RL8JluVmI8wzdI4AOmXNzGoOaR/0Hdwqi5alp6OZ86FFLsBy+9LHBXH/O0rtOj
ZRtbBILIGWfKcWVWFJB6nBkJqKvsqrc4gqTelSyw2LpkOFL34gljSMy1wToRBc6m
OHu9uzBYjMJ2AFForI5R7RxusRmsFeHS+cOOlfHKT7PoR6xRP6PvJoyl9nJvmKfD
+4GaKRmQgovoazgsXsPvpJEoyXQPTOv8nNq4Sv8snPLTuJLxtpY9aQggkMJEuXnh
QvcV9pJ8O4en2X/+h1p6GTKpl2lrTEWQ4VXZdyi8hW1xoBCv1Ik5ov2PWzbdjztb
XCa4EXWbvoOUQoscBMzMW5L03QwD3Quh64WB7ee3YRfcgo0ACswYSPX/awHk5KCK
c45e0JUiG9xFliy2DJ5qW0++nBPwOlg1N44GkHajuPRvP5G87ms8g3undpd/kj8L
bWagGdi9kBhL1yV7fZtd8TExGnUA1CqQZGg89AJA3O6ZwqXEY87oPpJiXm0x96MF
Iu7GVvVoW+MaANJLAG02zQNwrAYEzm6C8RPL7sqvOUH7QgYva5m9CI7fPdN1yJmL
fHEOTqgkIPXfXRNzAUWn+dJbe8cq5Ghu7aYhDUf6HcQqj0ijU4bQxMjKSJcDaQY0
rt3MMKL+XTjvA83wS08/UJOKLkFDokG63nNiZWuRcgRPo1ddT0yC6+CWH6QqHakW
fBd2HkFpfSOU2zYXtIxStqACncnSvQllaO7h/RPPeKvo2QufKpPg8u2kClq6gF26
HxGLOJ5WoFXdY7SPPkzVpenGGMS9d68PTEdhjOQ8avmOc2ljp3KH2cTPQdeYOCIO
Lurq8uaGmDpvdkBpASADd0GAqqSPw8QemQLgmIC/4Kd8kw/JzN2J1uCTccNxKUsH
aev/UOKiMOrZj1QCdwUxVVLr2Q4FM3psLcVA2iaDNaRgmiGWirDe24/t+POCIKeI
YL0Ty5IOdhQLrEQUP7oLy5jQglbf3ML4dI6z/awYAcJoeYLZo4qfdIinnfgJpRVH
ARWuKj7YTxbBdIh4ikOisAY26311Dhsq3Sw0Ne1fgNoaEGA9wsLcIheZ8YJGOh5R
5i8eolAE72y7V4yOTPdvQ3N0iOmtgmigtNWWqU/V8ZT/IUhLeq6zVz+SiM2/FH+p
NtsOTiVv6kgbgkPrJ8Yuh5FgTNxZyv+GOHwQOejkwZsDU+pT+21/vI2FmHHWxvS/
Kpb1QqYt85BQ6+s1NpVwumwS61Bt48WpL27q0cmeC/WqsMXw+s3RRfiRGv+PUpj9
S4AQfE3dmRGJQy22DKvDumgo96mTyNJWJZU+zSXRwC7TReZFdoQnh9ohiuD7cXrS
8FAJ9Ndwv65E2ceW/rcmO6WKdQBF+QZBOUAG5Nb1mf04TBVir7DIZNZFgtevIYmc
bKaNRD+QN/0yApbVnQa80a2S1Gh89HCCiVoCh2IW94zDay2ZR6ZQ4kzgOrqd+WO2
y93ktRVfUpsgVWuoaeXPG2xE3L1wjRXr1B/nlmNMo52iUKoqtQeouTMjxPRkdyCI
8l+BsBWSeCK+LRnnxUliOljL3Y6YvZGVyTn6GQjlaATFMcg5i+kSLXPZT60iO3yo
9NETPAvCxu1PrAb6uCq89eLkHPiMKMJi3Y7qHolN97vJ2QVANTfhZUHHCiCm0H4M
KahJs1lcdMlOR9RGTXhnnXtBziUYcr/86oPHDSgxYHz/QZ6NN3kBzKHP/5gEvG3r
HDJYdUBAFqgJKuy+rm4bp/kEZZcChWFfHayZjoXYUhMXf+DIecRXxuu09t6HkpYR
6y5pk9fLV6KF121VWE4jw/W5FO/8Wv6RROGZUOqyXCEFvxPplr2hg6fmxPMCuFFf
df0/Hv3/vygYYsYjJ4lKvWmGUfcr5QMMYD5k3zKne+b17XcTfOLxXlnzPgMaQdKG
v+9HJnhr0H+wzMy+pxZfODfCRkTK3hJI3GkEM9Ov5uveWkN7MYYS2jBOXU8QEvE6
uKrjQehgKj9z1lJOztnWoQ3cBf9nJtlmBpLsoc0ZjXwWHpCb9dpVX+nKeXv4j6K8
Eepq1CSaIUNu8ofjT5Eex2ywGIIdzXZ1G4ULTXvuQ0X9pAOLFDUXEzjnE9exjRSM
Xw/G79R42FJwgwmxtx/IWTJQWoniaPaCb3Dy3hgwErsT4bZTLp4ag0FYKq4Xnk9D
IAXDGRCmr9sW9nVEH6POValhuxI1iZFxLGHVZktPmCVEPkusFrRO6V8TaLrvEkdr
gTzFSA+rbDWP7K50alD8FkEbGbW9Kqo5UiFTPkvYtS9ih6lp4Lu5EGd+ZJYGq2ED
J2zHeDj9l9gppoX4GNweTJRYa4ZzdA3ef3+xPcPStuq8w/k92+gn4YJitT+mVqJW
e9OrcS3clUmqIO/dkdywZu+TsbdUK8VJnw/RuJUdynm3w7RxRQWRq9jXOdK9slJQ
Mu9Hf56Mx7g17vi7THWYbHFgbC4F0uxlPp8JEAm2GudRIcbwgzn448M/xf9bGUnd
2oelnQe2QUBhzKd4paeDQ7UZfCrizojudHVMbMhPd1dFWMKALBAFP5kkN9zlyVDI
B9/GEFlTmNCvwcEgRF+oQOLeFXVywCw9/fpeLgkKUVmbwslAk1owTO0ZOz/xfvID
oSRu/JvUJ9vEBiQkCzPPzCuDht/tUlhMrjpiHBU01QO7B3BfyY92aVmbPLyfQhfM
iJ7wXIDe8XN9fdKPxSpOC8zvD+r8D5Xc46s+L2OOEWv7Y9XJS21qHbFaDuy4eaN/
DUWAVEtSqmeXXwnIfphA50GtYBtBuMN5V15OGRMOytXBhdNW5H1BDccLeqX1WflL
kHimMZ+8xvYh/d7kgvhq4tbeBX4gYoCj7XGMarEOz3bwNpzNnPcbbirf2i5BxG0X
OTT0l7RBjKYzewsVUBf4/UbRZWgaVAJM0QzdDYW4zNH4uPiubrbdNn+ZekZqimbd
8wpeiWZmquTKfYY1IWPI9zxYjUC/yVG6Pagx1d4wRuEVNPi7dF+TMw+rGq2XXjgH
KvjNhNpB74HsFt2VqpCoXcu5ukr40Jk7UPkf3U1X4ND70k6mX5OWep2uMvN7qj90
NCUxwMnAOnIULD+pjIw+RHhH42iZ78jYh2POOMIAzjzQOXG4QKXFMtdtgrdNVVaY
PjgcDIk+jb79ToaHKy6lW/p/auFFN5EoFrbTXzjeJwGW2XujRqhhb/YGX+8nwGzg
+mYP8/tEVPi/Xc1VfdZERIJweaThvN5bxph9Ncbw/aFPD2zFavEwdbjSxFtC9qst
tDsHCo+63d/cx0O0tdl3xk/31zxaUarZFQk+NRrjyBHaWM8ZjS0aZNKw1VgYjcYU
LUCvyxsCBhRh4Yarw88WZ/SuXe3O0y7B0M9SIrtu3XD2wDybREBrQcMW7dqP4bIb
vJSmQaxHbyVqXYMKirhLYCmvqJ7l+aRBTNev5IaUT7pwrzPA8D+19VKggELgsjUS
Xny6HG86Lx1Nviw33YxHLut6p9rA2BED+5UDTeIzBhJncpQ1ykf6Ld5e7S1/BHWf
tsq3yqVsldzLE+Rn3xGPWlzopkI2N77Xc6i7cnbCsGBwZJJTPVcwH79o+EZqac2l
yGHYOABjhApkk/VLxa07nbUy3cB/nBnSnPMTA1XhnDE9EndJFs58g2Us+82opVRI
d1ZNz5VMjQIDtR1C0eTrxVttN5WZYgRkPlrQcsiIUe5eNp5Nck7iedNk8i4zYeQl
gjnn2oxFesjsmZAmGpj18DHDivMBmmIp6pHDMIYVi1ECllKYJ8Q8l2L4kse34yzw
AYIHvJMWW4fE7FocoI//yfvVDsP20T64fbl9OLodgUvJHEaHVvoSFCeXdldXejFD
pe+cxddQX2VQzVRYBuIt8b0YBdlXhah3DP0f1g94hr+yedTPrfVnQ9NvVT/UuLak
L6UIXxayeHVGiwb+FhJIJyRoMLwEW9DNB8DE8O78noVQ7rj1m8pOKKd+D9+9Jz/E
zVehnq4XjxGBYCQFd0gBF5l5yGpTJdZ6x1k1QJBTeslbm0Hqnl3tOXmy6pdoJNGx
CAwSAS86ICbbkdh8gNsOirBG4iVQlrkPFGlY5wLVC10Cq6HeBawWRsu7rvlLNcy4
VcLdK3QBe41IEQed2dF5YLfOJHkVcyScQUeFCcKwYMyc3XwWUsil2eoCZJR7V+ER
uw+P1Q/pT4YCzA2sjMd8r8ho36Mg58JX8DEB/EOnuGedb3xsze6PZAKxbJUZwXST
JDst1foVOdMUZgGTn78f9OkGacEY4HsCTacLHf/Ymq10NayckbWMr4AsKFL1/esO
FyOZk2WAGLOEoyHueBZWLpP8VTOqA0AxhRi106P36YKmZjbP+cVphyiAuz/hMJs9
pWZ97NDcGMi+d7V/pE+vmDPHmn+crd2SGYNElu8Ee7DR8zw50EdqnAo4vO/4qX6j
oWYCPhe1P5rJ/aAuH8v5e0zIm6ndZthqHWbkAkvXSbZATzBG09IQ92zdVvNiXzEe
KZy/OnZN4G6GqApIdZtkObXK2GN0RTqsK6KIln9YIzD/hx/qTNR3clmNPlCfiiPf
GFYqT+i7yYRC1VqdTwZbrLDwlDN11jnu0/2r6Mu/pQ/ywOt5+0BDDCW+QtZ2uhqC
svUhf11FLGen3resx0nnh2mF/rxOHVMKcxPZLiMLxqRERpbVpYdMNHw/lYzhO51z
lJ2i1o210S+IkCmdvESY25XiMaYjCT0ql+9AE+C+JMcR05K8jtjTO5JoQrgLR0BZ
C/zMMccdMX4erH2tDmzPyFSMJ06xmeSSGJFRuCT+ABjEe23ltZ1+lF7BRDp+PP9y
fzMkzUpHHLpexCSm75MQ4+ZSDjaKN9be00BTFC7XB+sXOi84hey9K5RLcxnguxly
7z/MLvTQyCIKFBN/CkqvaIY3OF8TK5JxBBMWQ4mP/ldmUs2jLIoZNHTcDWnkf9gW
/eQQ2altOseE/MLqP3j87XWc8UH7yjzoVjzLkufxoWNVXuMOTHLMFiWphrfBQuR5
EHsnCmuxiL9tTFyxcRavQi8cS6c/q4JS/2xm63Lr8nP0H/zal6q3Yni1eNwVbRmr
3nvzHBNJ6vXikLDvxl/B9Bp4UY/dQ7WWtDEaUFHz7n/WuzRdPl1WAl3xFd+Z4rIx
Aki3mbq+k2i68cpJJEgNyCrxSoaqfNNmHX6lvYx90sTZU7zmeH+Icebv4MR8vl+D
GjYoCbVTdRe0pR1gU46xLr7bqbIMJd35B78AYe4dEQ1nejcfRR+siN1Lha/a6M26
AXwx4Y0xBlGuBAwhCnLD1YotJg6em9Mra5B/1XxKaTno0gy5Lp+DYRKdGPyqM7nM
NwEs/EMwF6Pzre7e4uW3hHQmp9Q/1RX0R2LPm7tvNxiiIXaffqTSyBk10Y+Xc0nF
pTD4rFBBLAIebloPU1NGrKplixtV3o5GZ5BDD1h8mmCM6DLSw5fTtQymnSbsts8e
wf/T2OBb7OZwGBcQm7azpEvhhvfsCnLJ8sB3q626SVTXh/H9BNAeAgTQZ3h5zxtg
dZugl59Q+U54cizlvvR4zv0V5FpHeTKpiHWmtn+VREqGb3b8bdYzSMInicA8naSm
uKYGwFlMsvjrjd9hNuepLW0ahIQzXkVDuWvjFzLPUiOnWFMvJSSMiPeExEro+2gk
kQA8o7GUREdvlvlNVxXAAGNZ0pmkv65TskeUGF/tAUHOqAjgMffBhJ32yu3humwX
yyMaj589k3S7VqmHls6FLnuhxxuABRJuwvq9t5LPUli4EKJ4T+JRrXdEm7qZkcZ0
bOvZW+8gRxcJY1BILqYSHi3Oy+H6ZxpHyMp/JCk/gf+bYBPlON7tGmVHXpk1tcM7
Mo04LW6VRvhidGOMzvTsBQU7uP6DQiM67nuHjPiPHBpBIuBCssT2zhiXQVVl2Y1J
KJM6fHFBEA1r6rdzwLN/zIRzY9r12LgAusSsSuxMucdYn4rbbIrTdnx7TId3kxtk
R4xG72s3dPlx3qesoZmPXP1vDsMbFehpx7qtPEFd4XESYPqFcl8+EZtomjMinUMp
5OhqLVCmRIg41Vqfm/AsRvuhEABjlbUjHBWNCtBmWanDSwf0lhnlTiahX4xSQ8f/
tp+b2uMDroVpCnUd3GU2DGSvCAREXGWjKCU8l4DhVblPmlyROrsFLCPBdk1SpmI2
jAr0ji/h8uUlPJ1PzdfQLLgkmzbLME9Ef3jf7qVycEDgLLRcq5123FqjJo6Y39za
/WSqhUo9JVexxTp7KE/uzLnfjFYc/0tTYaKFfbuchkCOew/UNNy5Ee9nMzY1mgme
fX/gPCPTDG6D5L4tC8n4RVdvw3l7SGJkc9vZF5j2X9LLVg+J3/rfYjIwzGzTOgxj
MKl8YpTgMSMZpSZhe/kZT2cBCRforG6x8MDV11Hx+NfSGCZpDnDoQZW9OdX2P+50
WG7Nz/nMK/5N7eRvcywHO0BH6kBSkGj40wqFRtIa5LFygosT/HkijUlLFy27tztj
GclIUbRkObG1fiftFTKu3aLCPnW90i2mpuiOIvP7ymKh0lCWX4Axsyyn4BVA4cA4
bQCv6UiWY6q/3nd0ZXdms4G2kraj7JwAWvnRS8uyHz0xkYFjoYsBEvqUpr8IIu+u
Zn1lXQK1hhzX0XcG2TEimCNtq287oNtyVZONDd4hPJz2tT7xXBkNiuyMuLEFCIyV
S01P8JYJ4pLfbovJLEo4n8I+0JpQZCog/9ya9cIO5zDFlyujsRk03DKQti3p302p
cx8JuZvo/38PMgl/9T0j5V7fBFrhd5aWkxVcpzLvPmge/kvfmoHG24R7sYlytZrn
spB6nHDDi5wcFycAPo0FIxr+spe8GvNsntIarP7A5GWu3NoWreffeCztlcLidcf+
Q7nP1j0DH8kqdCyj4ZbNb6ylixvjEL4osBtGZwiCMzXsqrxZW5g9/wVGa+wYMA5D
c049CYDHJuayxoWn69b79vGaLhv9cUk+c6kWzOz2utNSJUvlNmp78nh6Xf4ePHqx
J5mR+ZuUhmNcUVrPPG8t8WXVFYNprfn+taI+hwb6ma6u+ye53cmpGa0euCchF4nN
w+c3Y27v2hZCj/XoSsCk3MwmpNzlv5dOFaigbuwaGbtIHnKUOiIG9rVQoHcqWBzu
dZB9WR8RjWJqZPKosqvsC5dTkAn6kzAtbwgPuF6FExmawtzBR3tb1/hAo54SQaRi
m9C15lq52/br+vBfjUlfnfFnQwB1qgzhN77zwe/sg4SBK/qKF3GZte/AsBkwOB1h
mTCKejuhmJ919z5gomGrStEEKRnjQqgE9QM2AGn+tT5ZLpQAP45hQna2ndwvRBd+
jxAsKY3OpdyFveYrZFErjkQi2dzfHnCkorEkIaczVay0VvaweGfiWGhzEtojl45A
SYCXZ0iB5XHS364nNNi9Gr/vscQxaWUI+Qpt36Zh+Gtb8R/wHQXw+uMLgmdGdncr
itdTd8ha2p+jGexpT/iAgnMdnRQknSx7+gf9HRM70AljhL5ueekM/nh7lSoRjQTr
UCIk/NPjU32ALWGfYPCSBgXMVbcFC5wz8KyfKG0b5K+rOWfhiKYYCGyhY8ytVWoq
/t2oLXdh3Rqp8jm8Q2EwEOdYbmmrX2wjkQXltI8KxjruQ4bynBOrGjSGUyNQFek/
jL2TQzSNYpYsB8enmk02eEfiuuXcic6wzstzkUiR/NEaBcqJp5pwphO8JCePVdNM
t9xswTjEmFHywMvkHwEvEceCcneOT1fPO7PW4htoFEQ7YRX0RNx6sIOkSJG3MIWK
wMxKUkkigCRvNlMQ2GfVhXQf34n2tGkNQD4m2du9fXWFXKan4pwi9ceMZXclKcVt
BTdoCHImLbfBuvuZyJpKbtcSvZFFSJ/R3AZP8WHneMXVkoTr2UDXGd7nnhA8gR4b
/sQT9vqD+h5coaQ8nus33YofIXDFA3rHIn1W/KTc5y+FhsYXctVA1HgYU2E6pX4G
1RZtF7Msn5Ke9R+fVkQSk38/n0SI6t0Wf2qg3TbV1a7QGk2Fif19xj8wm1lAwMO/
T0NdV8bGpRNii660QiNN3vwAOJYAuB/ZwVRQbnN292FWJoZ91DLWs8hkBc81ZHos
OZt2cofuDVYveM4ivtVIrFB6zVOgVIqcd7TWrmcOASPYxbf5DK+PvGFrnIBGIdfe
oDzFGa9H1omszIzJKmQ1Lt6OB2nXrEMTq37fotfwxkk6cKCPWGfnGhFg9/t5n2Cq
7idFyOj6aBTXlzZUDSR82FVz5w1DqOPU8qFsSXCS1fml34NqhkKqF78nw4upM3ce
keL4661s9GiQ9Zvh0RpJol0RKJK7CPxnqm8ZJUzEs+euqlNQzljGZqpPb65oxyKO
mXFjKb9COyiO9M2qtvSeaRwVWMMi6j9n6VbMbU1S+p3Rry28+PwLsMEQPgU2Dx0l
mofyE2QmZA2h5nlBox926mIUV11TIWssidXaJm+EYopRjYpY/d7TnyRlv5u9jjEN
Op6xvhZzI2ELippM2eBv/+wr18bAoqhHF5mAJbTlYehkhUiFmKJnWg/2X1oPR5Qv
pgPS+gg2fTNP9y0G+dZV9zA5BWI0lAI2ZkC0CEVh2OMfVeNomoFEfPs2nz+UPpXK
PsEqOPFvPUrKx72jsVNQIUd/iYdNQYJkQ5fvQE04PGqV0qnde9GEp9UNtnTE+paJ
Ut2vrex+lgx2D3AcFG/zDSbAsxDt7THy26oNoMmNLLJDAz8Jj9+6Nx1SrqbhhIHJ
FC0ws22CZTkYF5VgRh6o1RV8twhGUF3k/iWQbwRgHF0QZlLXGHpaxbYsj1XxMyuM
TMLhjcLMpWp4V6X6674q8YcHdsPH06UmUS2xEosJonS/yevgjau+yYelDwwbDGqN
/HIcU5COwJOngd07WSG6IKU2dooJtvzjqI8h7Z7l2fhaIfE9WaVl+IE9A9aRMunA
JRXawGUqW7z+91wE5rIkepLrX4G+h6Gl6cOkyGFVCJS0hO+4CGSrV/ZOlesnE6sN
dPV4zKqc5zFiv4fC+BVZel6AtLeALSVHGCsD8s1iLXmuyQtngMpY4SQJYO3nC8EL
oBHISwJVj89kS3b6oBbu3wZgmFjRIc/C/n/jfzHYXFGzQxmn724JrD8QE7YpqqZh
Y/ae0Gq6pPlkvB/kEy2InzEgmMaDLE52n+37XazwAxmqWWsP6dgVheiI9CkR7EcW
wj2HVJEjdhlQ+PNKn4UxbZ9sZZ1o9uDo92XWZZAWUZl+WresfWfvywCtBNC6ZcwA
9+s1JH5S8Zo41/mmBlUOo3AasH6BPLCRDeNB6Zy/0zTwDkrOOCvIFC/Ttv2klpep
Mp7qsVSyp0Jy65jy3fVvgZJc/1SNUJy3RDwSJdTtPJLcpJa6fc3J7Rvi4LNoEeaN
7BHbhiYNnhjLjRGpZiluPxpcGZE/RNzKyuzairR93uQ0OqdTuvPRo/iEFZyR8HXd
j0Ys+XsR8gUSfm5HrDeqIc5ULnYWCYGi76gVcDEu0nSi/mst1BcSJO7brDoahmG+
mGDvatGbTagriVRkEuABHdrYcPc3gMnZqG2szZJoQf/m5jw0QaosyVoM5eT0XLt1
ayQ4WPMetfI83iDglSeuK0ny69ORvEGd5vo2NFqsb1VVkj8jfw8bcKCWX8PpAcuH
voepOYz29u5WIU6imFHMl5uXjrV3F2rEzt7HR58hG8aLhQzGjjXtOwW555NM7/cv
FW9AUz7ZjqV2VlVXSvwN2abY1YgJ5EmQZvsYI0gJTobX/sRF5sMNXVzJ7gGQ94et
7KuFsJD0ncpKQeG/WJWHSL2yiuWL6H4tMSUkM+MtuC2ri11F5k2y320kD/jfyQK7
LKc76/avLYb1tXJ/PTOxc+vz47Sh2j9nGQ5JrTHNs/vTL7+74Gn383CA1J3+/3Zc
Mr3+tY9DV8CjiB5U32uAqFeDxioEqGVZ1ZxZW9w7kdodhPZ+JykpEwlqoQoE0Ohm
2IsIGQCGRd5tfLgGttaxKss/dauG43efbs0Tn1NPUv7E3c76o98HEP0KVGIIYwya
JjVNrYLwGGpilgbcM9X1uJ4fgzPMzfd0zPcKaIVD09KNp5SzVLxfWyK5lQQ+Txyn
nlw1+ZOExtLq9JtPTHYUacAjuJTyCeiWmfQbzw1EQsKQ9YWEDAez5NtKX+vHXZl5
xGzC6bOsUvi7sG2pNINjfJ7CbLbB4i+9QRjrVBYSGY5CMFLadnFNT0UniNuBdUQI
6Pl4EtWzyvH21F8LSW2iixCXfYc0mbWheZuS34LpJ67joavMecsm+OsLktYY1A0R
XUjvRfChWV+P/iFDOF4egNpuGf9UxfjLQhQmsKAQecV/DzZVxPYQapRT2uImkUe1
6UVENE8573EHthmve/6wgWyRam3XAbr5fix4MVnVogHnRZGcWfRnl3QIdXIaLsaA
eV/xP58VRiIL2jysN3DLil6/76nkDu2RXqPrOb5JpZiELx05OidnGx5v2seeA/xu
PzO/lHfp6fWVg7+SO635C3BBom9mJNdk00GKjcb6ZayXY5LZ6Jxja79X8ZQBIrAv
X5qPumU7v3RSzBWOkBydwt6IAHi/RkYBcWv3l17PcTkjZJDtXkC2tixlRKF/htEw
9vvbr7HhfSipPriex6K9mJF/gQrSmiQRu9KPiLP281/Fhb9bFXJ2PDNDgT/3IlqI
yWDXBhwVTcWgxDbqbHSbNQ==
`protect end_protected