`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
ddtXksX2+yylW5zu6QL2Lhnb2d1sD00763mmSITNX595NcHTEkwn0zB1Dry37fOW
FufOhVzEJp80NC5qZ/+F0Vk7Ik02dIR0elf3clrjeJRK85K4e3Hoo4xn7YbFUIms
l/8VZSb14+JVGURjfswrIyCUotIzlzVYZ6gzoZwDXIi5gQIBf/gI+KxNXPaKV+PQ
Ufys/12rjO6aI/pPlqSm0hCvftmBcnezN2hk1UeXgOIuKZnogjOsf0iJVX2aOOWE
6pD/psybjbnsNB6kH5uFTA5frkzIzkzl5d9+YDm9OyC+k84E83I/7/j+rk4L2dah
QJOvksSIzN867/4Qt8qYTQ==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="MvBXkzurAa5VTw+1JJ70nePUfoQXBvZOku/SMmg4TwQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
oRtzZL4VJ4iwysPsC8SXYCzXS8Fw2gtZTOskLcDV+1B9Nzn1zTyNtlo6lNICRmmK
ZRVu2BmCc2G+fmzynYlNTnSa7C0Cuel6FYpxCBlOuk3OF2tzAmLAuDyOH3Z1Yjzk
a0aHuoCdIRKv7BrZCdALt03JeUmXKPdOmIlkVGFl8yw=
`protect rights_digest_method = "sha256"
`protect end_toolblock="Jn9CQpRhJt4rnzZPRk+dOpzAubz7omckX1MrFd4p81o="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 14464 )
`protect data_block
gD6l00tciPUa6pDNTk/+t0OO0nC/UTtBwLB41d4inuAUA3i/ALrNyoJVcBnAmEQW
ptbcNp5fxEUJjnOxnedyZEuEBxWRieZFQnkRdF269oNz3Q6LfFp2j0aAhShs0UUq
/5dt0MOzQA30LB02NDgeCBarVzja8H2R4g3wRYi/KR+7M39bK4nBE28nDL4aVS7N
MNoAQrqhxjXHo57vcWaZ7HKVkBjeS0Ie6kf4GW5YMw62AtI9EcritZjYYNEB7+tx
AzvNZv2eA6xskezjiIvZsfJo8f5wDkq29XQQAVQGEhwvoULY+UbnUuBmCfnjgT00
QQ4ZZj2p8Jet4hiXXT5zCuRcID7KEE/mr4T8g1OcM7ysHByH5KDgo1S+9HDLve4K
dYPnBYm+eszUxrbodQ3qZr+LlidOI6sHwKxQpmQNkBclozQSajUo26dhPZJBteYv
NQ74hjgl62/CSfEfBZ/stEm+ppwlLgOtxbrLmeXhWYkbpKMb1E9kDq3YxbwIrA7V
Uhkm+/EM14jxjG98lNCDeJxM7mqPz2+80S28aFKstAkIDQyDxM1nAl0PU6KEEUbw
G3qn4pPQjqHAddOQWdiSKzSHtjZE+yazj22LyWKStJFyuNoNlsqvIy7o730XeBXT
t9VYAfm1KIfUTgt511lgYyKY+WXsVkRana8kvmzHcWJyrH4FDltL+FZyCderenaj
3hVcTaW/4r2ctFPHlCoE8JGaZn4drYB6Poc6WRnpQUWWnQQmmeo3uVTPq5zp4rhX
6a6Ffo/dxs24260fpAOKY1HKQd4EzpyV6FD5TB/HcWDpgVv22YmqV95HaaU+6AuA
UkGW7mRmpz+XpzbnmYV0IP5X6T0M4X5Lyq2MXYQD8KgFrOQbrhoQ8ROPkotrf6DJ
7J5M6hhnAq3CMMAXz9KXBBbKYEusN4lVTBkvT9JINk9nOnQExGnV2mp7qw0cAqbq
VAgqZC534UCVTdwgyirrNJJRXXGMjkJKDAsIKWO7V+90wA2U1tu2XytkFLCmzjw7
JfWawmnAZj5JUZ1gHLgUS5iJ1ytAzIIZIBTic14tv6qmEbW1fCvYF7egCkz6OLHC
dkSFoqz1z4a4eWYJzFSt5mP2xNBzTwGussTxAj92pj6AgT9XnvIDDtGTiBuby8lH
J1Kta4vpfA4IWTki4uJdz4ILc71FuOsLlV8IEyn27PDGLbjowyGZsaC15KqUxZB7
y/jymt+zcCoLf/P8nVtHq9+gMk7fQIerAawn8Ozo3DZVXEPdXo1/IY/eV8/zSWiT
aFlXoqcfYV9bISqMYvzJtoKOiq5+M6LaXa2cx+pkby/RHv6q/RsgVCWCiz+sPWxv
0SCO8mvHcy7D0VUpWua64BA7nmrlYLqdyGWQFJo/OhJVIlsU5t0NmJLUQEoTp+LW
afQO3BYq5HaUXlQaxLGv0TDG2ur5S7FXrcY1rKtPuWz/0YKTMgLYJprZ1bn3ZZPT
ktuAFvVPqyckHkA8V+Wne5dY3qTxgBe3Fkvbh/WbpicR5u6fAbkVnNsvMtKtxikP
c+8Syd8ynIdiMJFCXU6I2SuKDPeD9owpH3/fZRBZ49/ZQ1FBQLksONug9U54fLUi
oyejBTJDc7YpAyU+CavejymfKSbYmaJTHhvuBAMT7EoTiGiKBWtqv5FOXoEv26SB
5/395VCSAc2cga9e4BC78rQO1KP9IfyI079yFHfTPszzMOM/BmOn9rOTFFigwN5d
NXW5vrSGCsCdZcLd1UqwP0PXqajD2CLtpAdHOXrrcQyrzieoErQacZHWivkom8Xt
7MVAYqgQqyQ1hPNpe+f0oe8AZ34Zu6fWiKFDnvmw39McNLOUblSNGBG/oE7LLDg5
Uxixluclo/yLeT27WgyC1Q9HKRG0LT1NJ02qA1EavTahJKrz7XOZGibrp7JNv21P
NROGS81oOz/Oe5f+9erhA2gB4FT+OKFj0l7OugTdSPAQfaTVW862DGZJtQYCN1Lm
19Po1Z/Frf2wN8G3vW5yxa8hym33f+lw3ofCj0ToTreV4GznQGIDh+etidy9lnhu
rdjEUzp0FHR7vp95Co6ti5yMZkYBD93ji10HRgSOSi4Ce20UoJ/Y4qFVoV6ZFSU7
TP666JhZYiadTtW1iZEPWpJqN/KABW1VY6/nZgyF2/bJSJGtU4Ou1juONMOVE2ZG
WhFIQCbFf6Y7kBj95ApgNMuDUOnmKEZKzgsTpXVlnM/lvSvZZvGJhOw0EkB1phVE
AUYoTSucCg6/Mmohe+KurK9pfV3x86f/wyUcyi8gop+zCVpn84SoproMTPKPCMc8
BgGh5NWdHBs+yuKx+096DR49jcEAHtZ7b5K3N38ZZ4450GrftvDisCotCTOkcvjt
VQjKNrTFJ1PYTlvO4eosje9VaILcGC6ldpisRM/fm02j/5QGyxHLv9VBDyaL27lw
vi8nu3Fcoo6e0R506HpkxERx1OM3wCQINwH97Ez68XTcS6h1lHl1Pqmt5zo5/Ny5
Ky9VB0vMSLpIA6iz8MG1Svs49rRswaqj+4K+lEpPKtY+S0WclMlS4+1Sg+b/aNIc
nsPzUeFg5U1PWFjn8+i1jUEby9wHkEHlhH0UCH6lU8g2TNqZ3Cuh/qj+WQkJ6fpr
IAXzYUStCCYvpsloODC6AYIiBphLGvYynPZdBTwNQZnOScRcL9HtXTm7a+P3eKu0
PuIkFc78t9cKqe+HiU04QBUbJudq89dHBw0Jz25odLMLMw+0mzsKGEujISA9AFWA
PM4aZ9HwxeO/6QAnyywq8LAzR0BWkj9/7ze8+Ptrm3CEM1ZV4yNVb3zydStWIo3m
hZD96TQCJE18YHdHmSwTgUG/onE63ZM84PFIoA/P63gEhfry7t55nAxjfls3nNbN
xpck1uou/SS/eOBiRUJzmIeL55JDPyDhGcYukzf/qetHFDA/mkEbpZFTCg/Zfs8w
O3jeCHVWlgzJ8C78e9dtNq2zUJISYn7iLe5Oa2zVWxjMvB0C2+IWaJx0uzuCJ1Tv
wSAZTDWSn7UZlOBtbZnKPR9BZkDoaRo76zaH8bEpeHi3utAfkdAEM8slt2t1VgSN
oixMiu8j382sBg668DTfidIQWYDsm+OY+uiT10AVrnP1/CC7gSjO+GeXAu28lW0r
RfcrC+D9gRNfi5XrMc1AiY/OwqK/lCprn+GTxYPLCTwjO7OEXlHCGhhRHn4kmFiW
hidlatuzuEL4x9eb0VaaFIBoWFCS2aVQXPYq25xL9oFTnIxFJe/ADt9OEMwiP0oc
5hi75Cfg3bf+jGtwdMEnQi2Cx3FpD5N7KWuhc8TAvTlpmQ7bIOqlt3SLNFE46Oii
NtLrlDieKG8e6I8EI9E4PnE9m9+N5FmtDpHa4to3+CvDJ2Y5iJzcCAwezP559Oh1
Wfj7zEa3k3Cebp9AWtpsgdTxJtqkW3NDCKGrhcT8BWXAo0n61XzY2xtPC3XdvZRH
kSVN1KzXCGDo3vx1Y6j0DogQyg3fMdGBI6aw4/blkHUe7OdABy6Qehw4O32ZLDJ0
xgGQdEjFLx9M2Ed0RUCxDVfhWR1MOGXTPV99/2OB2fT2Pi5q3ZVIpoJl/x/xJf9Y
HQBVNpr9l0Q4PEUC0F8oXydW+j2YZkTtsrmh9xGjZKw6YTis6RcckY741673ygvM
lIdkkp+jTm9oZGNPE2lSACWwWb52PqWV8+fDnkhSQFLq5jlBt0gT6DdIByPObLml
d3HxiywuZIGFuyqJ9r2fXg6tj8fUGYXX0b4ADWPTx9MdtGmFiBBJWO/gCgP2UXZo
IiuJu82ZIfJh1UpEadVUSmLI4iT9TA+T3CKFwLpPqPQI1jD7bHHZge86D8kmxMhw
CYDQUoK2Jre4ypFbXPF7KS0B+kexDbDBwxnxzuMh5xWsAllj74ROB2TAh6ngW2mt
w43z04HhA1dzjX9b1jY+C4UuKh9KVdCJrOU2JvdqhbHFkdKnAepNejdenvLVuf4h
jbwAPuNDg1wJbu1tS8L2CLpXOLbhSbuhQzAng5JgRoGce3Z84jBmOUjZPQcq7bZm
wWcAuJrFMROxi8jPgTsKKDOGwXn5M7wXVFhB/QY+OWKMEivzyS+2p6Gpls23+1sQ
A+VtFaDjDkISMcXJq4ijK0wEA6LJlocEjWZuksqDjjNGSz3DCzSEQAtpiQUqta4k
B+AHQn8hp0JW+UU022F1Xdy0wg9GYLSaQ2i5rB2GogMb9KqhbBJ5bCORt3jjSKPb
aIF/ybd5KAcPmAzhzKy1tB5NucI1EUKx+FNAs7k3XLOFTtJbRDfM6z0NQw2EleLB
wCDnHL3S/oIURdnLtNar6HoYM77syYUNbrqt/yRc2tSD0mtmvq6URVICCLacZi1o
y5DG2kbH9vKla6vWrgYopg8R069mfdsaE2SZQEkIxHhPO+qNMO+letv2cMpxY6EF
7xo+Tdex5IE0TDvdemWaGFvBgGTB02RzOMEFz0brRXe67TfePRbdFnD9NFhgdwat
FaAbxLj/q1nQCyvp5fMEAWVKKhlFnzspefUWc2/9UDBSU1EwfAvZbpkA8BW5wj8w
Zx7Kb1IJ5+jDF03k6NlJd6Ws8zCyVJlk3TCnvT3bA9UjOrGlx4iPWB/2dGgTxNlu
7/Jkufh/zoiINWpJwZ/LE3hCwwx03OoccjbGzpz6WUKeWWV+361PvbC5FCq3nu7L
C7H1hTe5mwIzr/Th5+WTlUdGIY1DmmChOIAsvSlGnx0tMYQzujnxYbFL7EXapat8
xkIVYWEfP+yFVQU9WvBYblKgG9PK+/yky47VjVy6b9S7CQRPTKNp62XAt/cTB7hx
CEwryRs/+ihoBY0XctJx/XW2tpw8HH1WZnAgA/RjYBICnfo8PjYWqIgKr1zzpINV
JgTjbwEOA+mWFuaosvpDem98DoxVmg22COlPktNcanRFQYQva9tq225Z+M0DuE2K
c7Y4LdJv9vELbSC0rsPp9szxNikz2+pYtDvs+GBrZ44Z1dRLpHb6NG0MnP3hQuqb
B1HrhPkFWiXZGB+pyPE3n6ALFRfxPW89wzIYaNevInDXpeey/I9TGGS6mBP4K6Dr
sTTz7DG7oWT1yN1oLbN2H6WoNGIvpFgphCosE776DoEO4VvG4RyHm1g2vd15z5jn
aNctfhvt8QmtjPO1ft+VqGjB41UOgSFk1qmyx4jHaKPb0HxDWXGwuH01gKeOOE7L
Sn0xaLF4yxz4PCIicyl43rr4BecFetwUu7BQKSvZzXBxRlZmmJBss762A4SPRrzM
rmacvH0iP4Oyts3KEOxD3CJ/FWorJmxhVb50BTj2vC8uHcQXsUXvvk3B/5IOrZGC
zGgxWpuWzVLkzkWFPLOc7uGS5PyU6SElc+bf8ASL1Y3TOK/6jFTNoU15UN4nOEiL
xPFZUqRIExMppGr2Cnw46sJhQ58U24YTMA+7dV2f3wTj/Tn0wJJx4ETPcNFAHSzc
AkiGVYMktY4wxA5oPmzjW19j4jMUOd+n3CiZP9e8dJZzP+Rovv7+n5aIdko64n6r
kCKZ7zmF310DSXaeO119Kg5m8zdU9XdPG9Mmr6FTaVLooWccSKZBsdtgODjj257R
pWy0x3Mlf/ysHCfWNT+CRj6D0/uRHviDJ4HUkgOBTKn2tg+Z9yX3bkGKon3zZz/5
35ju7qtM/A2Z/cVIbGRf/r/qglJSz/3NegTosDEUYBUWhH9IBtPu7fCDVi3JFsfY
CqeskAKMdmGBfT8kXOWVoNi9v84g55LtxL/6XY+gYi0aSYWj39ImILRAYVSfZ5QW
BB0uGVJVxYcDYW/4ZUESo6CsnmjSH5PYffaSYYHyrgtG+qiz2M/FPjH3OCgbl/qv
YlEQNSBw4UiwtABaeMRmDoaEJ/2Jo8siRiRSFUfA0ni326imlrmg2XztBIPhyvsy
FxTwgSw3USh3EOTou7XsZlONZ1IMw/Ip2Xhwjwwvk5ZCXnvMrpdDreuIj0nXDa/b
cRxgFsHSXbEtMi690UrKVO2l0H/8piwpB+nMwcMicEsqC9xB3gawBjcPwt5yrP37
NgBRQDZqJq35nQfR0K3gsbDiHJDRHtVUdBFvnPUBeGQyg7FdSybbonG8Sjs8bQdk
oGEDLUicA3mxq9cvnfph+tUU6JcPuZGnipmPcOJCVJdFhdI9nq5WgKHHN3P51QMW
Myreu1H+9uYiIVeM6RfOUrYgVJLd5G64aRkGbV+2anrWkfYWbzKLnFSCp4J0UU5P
q0+BOtxqX7GmnGxk2jA6ZQbriiEY9sIfmgsIqLVbTPERSi3pY8M1icp4Q/8jCqHE
JV3JUUkiP8qmBFwNidD5jBWWcshX95e+vQpePp41mF+LF/oKy2CXLflJGCfFT7hv
/mUvEmYi84lzl13bwTaWvjeNEYNMk2ezsXjC3bgM8vcW2pj0BTNjoiMPxAGaUf4l
MYXnJalmd8pJPxvq1hq/ZSn2mr6LnrLwFMXorbSPhPcobDeNs8u2jfJ25OhQivlZ
ZcmsFVZ4z2LGg/AhKzkiSXXDnSCJpkDdI2MyAM8AgwCSteqEiY0RwqTIR20kI1TB
iSxh3pL2uGb593chPYFtD5CTEvuGNxTDBaBYngdJQE0wRS1uFBfdUJgiGGXLY+Cr
+wcRZyC/TrdaZPtyvhYH3R69H4tJTb3mZvFZ3RvxArgR+OcLjnM/V59/V6ebNvsk
VAb9rX/ppg2ZYHqSQJbBBl3FcNISbGSF6HTOTPq3GvM3xgPF6UqG2o32o2F8sj2y
EdWOVw+G6HxE1Rcy3dUB49evZd1fqFCPiKwTNg8KWu4ELWDr1UtiRpl2ZFv5sGma
SjyXrEfhtVEcK/pD5HsbgTBCOPt1kBlTCZiAkzLSWtIB0F1DL0JT0Gvlf1ot8DX2
PGQlBpoxWngQcBnk0Bw8N0BBxycatPfgQ0KNHT74TWjft4sAkN+ZZ8c6MKhy+OQU
S8pKH801XUPkuGDRNjq752WMcwqGKjdXvBU42ixqTKBvJCFIrMUfw5d/ylOY0K96
BSvFSMgf5FY1mrKFP9nyUGYXPvqdpgn7rQkYiqLcOQ+54+tNLa4kqBkAizHNmTJo
wAMh53QBmxKi5sA8qUUBWHfpV4dAx8DSwbXyqCHofRD7i9yefyv8/cwLfXhcWxFD
ud5cNEEzhJfEFfopSbLZTGibFl1+r/AcTGlCXXmreZ40kLOFMyIrOSQV4DK8U40J
W73pK5sMLLOGx4ioz3etaqYMGXmj0jEZwyKTEfaZN32xOt4O1XdtW7eE+mydLsan
X/aorK0ix1giVHTBzzaz4dKCy7Wm8kaMwZBC6xRov+TEbkF1qWL4EHt3legQNz3R
2vaYsVM0m4qt53/GC3bHrC+V4+c49V8D2r+75hmqJ384Gnzr2kRn40dVcV4wfjoj
Yp8Fj114YmJOk6eWM5LeDjVUiTGIRdEN+fvQDRv/Fs9obiOXYQQ2vNX/SyFfZOqu
+P6UCCCvfLfvdReWxI0rXcAbvWATu4H7q7hYTIQaPUnYkJ1crboqvrzHBItHMhcg
4ZQC2PILpkAW0P8HriJVQhaXxhz1XqxZVuA+uXi8R+DeSIZei+pykPaQ7mrvw9bl
QtpMXbI498y+KfG3Z+feyx5WLRLChQmKMZ7KQWPdOaRRQpA/Kaq8OaAuVNwOW2Sd
dicTdauENmMOwVfB2V7VpfWaqxGLH3FYQq+OJGUJWGsYUmgHmpUwcsoHs4R8dNi4
SXLyZgNDWVqD31zO+kG4JPU17XTC9d1obz/9t6Kb0lOjq4v6fZf/YuFVhiItKeOU
AtkcNTI4s034Yj6FBpOsC5JkpOW4rDEpGHJ4P4trCK9M5ghZQJyT0h2ouTlqy20m
WUUGmUJDUL1hEURoApoD/TufG6SSVS68rKTskXllR7ZESLoNU6/nxkDc3zSLCcaj
unGJMIjitoJCf7gbNQKurKl4UnqKmnb83iVKEqhkRi5ExbqAxEAc4zgSvHwXAdJZ
USDZa8DZ4M9kneTEsc8xD7fAwYOMA6UTnqGg6DAZZ/a19vfTRQujao2a0LOvgTmq
08b+ewssKAhLi8CzT1ZqIUVZ34v1peIiD9DxRLGVNrrf6RpHuz5fJd2NzAiClkwb
fh/lYokQctp2nUplmyMUjEPylEJm7rV5TNy7EB3il3nTRqEiZRrYXSYTBMoN/DqT
P73lTV+j8UUy2Dng4n0N0X/Of1YfZYrPZVwTTV9/bwtwRTNgFQUfX1tH/sDygo9q
VlZBushu3SSo1ztX5g3KH2YXWsR3PJ3ApFUiwlgeq19sQi+ga/00F6+3F6T1GbNA
Vk8GTbp3SagUS6mm7XgfNx7bzs0I8GmONL9ysHw/Z7H+Hn2Z9cvJMr81dBjZznWo
835QuuIueHegHQzvmhii4pB8/U/rpveJhZXVllCeBSi3Og+kiG7ECjvzyFf8nZ5h
FDHG6Z/yoZk6M6uDPtPcBnigbDqeearxpNBt23v5aexcjMMbZDZemPgxRcOJ9bX4
SDxX9M4nEhPTupsJueKTaT/n0AKMmFyLMY/wBbBBdumBjs8zsXXlhNQ1GlWQ15as
rrDYqVsguVcVLjLB6lNf5gLRkNqxNaME5MYw7KvEJ4B/bkqb95r6Ob9UOA5OvDc2
QWggVI402I02dQWOxjjNTjZ1LRvBQo/YGVsyIxdWSJGN5x4+JB0HWrCiPYi715/3
fafc7Y1N0/4afTXovFiK561DOydTqlCTATBxYT0/+PL27SxRspuhZO4qsH61YKX3
0u7+5vyWMoscVSpzZiMw7MVTHL10aB8ifbf+ZjyiQ/IWY1z6GZz984bmJV6SAFUc
Qm4CqgPFTf4KtTkyjl0RxyWwci3jgy9tlGtl4PQDwQpLFcGw62IqjFl4Bsk1US28
7b5DNXvCqRGOitdaDtlkMrNmFcEHssXwC/jHIECNiKaDsvTJVk6rIEJPAVjXVWFX
2HUNLe3K+UpE3nxJEdlQUVmmElsKDGe72ZO8C92IOe+nbKha4LYYYwKneP7pgy3H
OS/ht0XTZUwNMobqah4Pj2mH2Lm1WMngIJ7cZGQlIi3J7iv+7LIY9EvtITb1+7IS
swVjFSk26WPrkx4xKDwAHwcl4aidPWdI9uENBnu6iRIi68DBsxdOM/TmMPO/sv4K
mP8zO9YWjglyGCIVcII8q13GzcCaSOPukUrO3X6xgA9q4VQMY1p7PdpjZnppqVX4
B3KGeQSbdp77Oji7BnrR6xMlF5dktzfaH8giuNBGq8KUOx8iL2il6nen1vg5faVP
gFPiS7DZGVrpswHOJi8bq/ZHYG17IQzrbdKXLl6Bn1qSiqc8GPGVqhkXQYgymS0/
XfLt6PrIP2LnMRN+2i/tCai5fJ13b8+seVeWQ6orW54dQhtIuD4qi04maP3rbH4H
cyvyUAAxQpZK/w/3EhfoDj03kJ66eFnkmZk91HLGJPS2comhkW3Oo2oh1ayLrMPR
KaIHy4JPqya4J7wNvqhpwsORlE7r4OnB+5RmzqZKWelSwlOLOhFl5Lh0HrcMHhag
47krtY1I1fy2s9hWA4qzalWoDGsZt5re6dSwInkIHbyXpGGLQumUvj/CrB4TSj4o
W9JMM6yCBk0yxUoeT+sRNie9nq9QXMWslsovjSsuNOuw/QgGQVO1ozN7ZypEVTqw
MNWaafhDUp1x3opG1aFCkRf3ZcGUm2CamOjSO+Z+GJOJFmXqZ3WsYbFnieEA6sFv
NpEKmtTbmlFcwUWH2DFjhiVazDbmsFCwrkq0uIUcmXdE/naqVQifrGhS1ivngms6
0Y1hY8elaNKsZZR+roYMpMchVMfJ5hcEZkA36NgpaH0V+cdWuxL0FONS7+8Kso5t
Z49BAI2uWHB+/fJE3uZPKy0H3Qp8HA0OQwN6tJyLBIcb1K9621ku+JAGLQ+b08jK
8loW9tl+hj5DdHUiOsfQxEEJimXEasEgPguOfj53ToqOO1NgwTrV/3ywlBV4EoAu
o2/yde18TEq6fc4uvl3Zp1E/R84yHLhqBANnuyWvtOKU6xIvw96sioQ8QUKmdSY9
XrTeR0csv1KA2M5/TgBhkPsYCuNfkImEqb88TNPY6bjfvR8Y+vkQsMBw3kSmZPKG
Ro5oaTG5pMENomUNKHfpcuRfMchg7Ggg8ChGVJIzBvqMRJsu+bsrLdRscYNb7qbC
olpMVWK7mjR7Ukdr99+MZb5P9aXo0juVSX53FBbKhtFDlHRLTKVI1LQkxu7LmvP3
QWTdJjnhZ/DNuYL/C3gxPPooCpBjokEifUDZa7/BKzlyKkJ/mUdpZdluQsFXJLgQ
KzAOS9b6AUHlURa306/DnMTOcLIOQwksP/ivIHf4xeQmA1RPMGlcSU3a+n+2zEBd
ZvggTmHENJZW+Sb84cVZ2hUBHcHlWQYzxUQJKfmbHA35D/IpR/9MFPNMlwmfnNsB
X8UhUMWP1OfE71ahk8537C37sWpDdtH4CEcVyxRiV2K4cwWECWc/gD4XqpSZTWFK
7KrvACIKUfgLevzjIxcRiAmXFqCrWW0J3DC5nQiXNRmGBWOdpDnscw3z1qDIFaKb
+d73WTk4ZDGy8T7xUvMwo0E7ohNeA9cVwenG3ki5+qnugsaRdoRjXB4DCilkFQwj
GcyGlOcUkbj0EkZQJdzbzjAnSGfBe7judK2H9e2az/A9VmVeFRd8R441nupjf5yT
Zq44i1KBBSlUmP/+Yw9IvB6XtIsFv3wXyO+TLEJanQMEYn7jFbZ9uqoL5lcqqa68
UvpdySVLRDHDSP++rOSnVimw3rxg1VA9OfELjcxE9m3AwuzEQp5DC1LbiBDtFHQy
khmtmLJ1FivTFE7VIcL/AtAYCIKJ6o0VDKvaqz90bVJtB7BMFUSMJtQwWaxdmZA1
TbLO0w5ojr+zW9os1AyTLHNOFXg8vrr4exsdaHMtnKZIrW0X6mS3h38zQQ+8+ON5
cI3UYDUdOPIY5eTtGpPMmRBN2IhQrODj9Y4MxzCe4/BJBp+UG3MmjGaENpxB1X4J
OIeNKYOqBGR8BizQe+JckLfMGkT8+dxJdfiQaM5+RiQhXr+o/A0mkBSgm3nBj4ig
5eIk19zr4UyH4wWPnZBoDVFme8cQnh5vnxoFfR7Kmej++MdgqhziPf5zSVIQU0NC
lD7HuUGNYN9q0A6EkybopdRtgEVqeIxxHglSiqoHJN5KdrMCPenZR8sak4wrhP4D
hnTEkfghhet74HSScgJK796GuEUEiDcGA2FrZv2T10iL5iQQVdy8I+Va8S1RULwr
5bPOI20oAhVWBp21XTnxj5l6Lqc1r/+GtqXAwgQgotLsBLt7zaO2hsdnpMdosHAC
q8/6PhYRkC9Oxt+AuAGs9/vjkH43wkb/r6e9si0fX8CFe5Qm9fhy5zDnSKXGNCBF
G4/YuV2LAmJBl89CDfzsSioCoBBFLA/5yP7zcqHDIZSJdLV1yw92RP9u+3xBFz7T
uJsd98NCcoJtDoYewEG9jvKYVM6l7tehV6ahmXlgQOQSrMqGZ7dqle/t/uuvjfmn
asGT89BQIXLdYisQ11fGxQFl/UF4FJI1PPFQ+rHiPFnNKCLtYW4o3WX3NW09H6vA
AdyrWgfWEUkeSWFjhX6QGJKew1JqP8Lu/5QoL6rZ0DMCCuBosFMh2/J/jwtAvAhr
PjMOzCXeY2rmDGzIcnSke24CYQaThf34fA008523J0ykWo3AWT5b3HdxFIJBnfVV
5gcgZR7EPI3tGS9IC0RTVU/2WGVqqs+/1RHlDLnRbRLHifJhdVjJzqDHEMhA3ixs
iLOPHUcbooDVoZZvQkJ8MCT+jJJErdNP1Y6P8b88dvmOztXoo/uFqCyLVuFKunjm
aQtVtmL4MuziyzHSqehGvJDBIe8QERUKWEslew5moyXaPC2O4H/uZjUFlLgdfyZK
GIzdnTXV/FzhLBy+ghiu6apyVWdEJFNfweO0H6vt4zkG2/lztNtyWhQpOGEBLHGY
r91wVGb/yNeOF59lMdjOVFrek/EcMEC1JNevWjcq3Sm+FZiuPdH7VaOANMqPbqSP
VKtMfIaYoqlY4X7jI8X6acsZsImSSLEwHaME3kSOWF82UDmdyYX0AXrUFjaHdONn
7jBQAALj96kaAQYE6a6UQ2LULU6oKSpcBAheYB3rPX/4ZIEjAWEm9XdpCS+H3M2x
wmfOJNeKmIsiDESRfAffDuOLRV5Z/synvT9idekKkoJWzqpruTc9hA8J2MuO6SUB
SjIY6DV/lH6rUYz/J+RwxDlZW1GXeZ4kf0zzs+JTO3iVoq2ZaGrI96GSZ767UwlB
TgMscHNwHTAulMx6AHPaaMyo7yAGMvLYTe2d5gkEWVjrqXxxmmQc3oQwS4dvfRnU
PY6FvlkhT3bAEtF18iyeci7tR7AVP1HCN609a91zCd1yilbZ/3annbT0Ep0ss32N
9g/zksLTitE3WfvIaMMdWadZHnAOoQByK6oxfkDdMoehCBWp8tuoGpq2+f7dk748
4cusAaAMdGlV8/eaMx1GGo4AmFpf4QlPtar3YvjvPTA7dCrNaAWavhM51Vh14YV/
3S2Je1Bgo+bJ+a+pToUrudq3uL5501A5PtQKR3G48mpAWMbZlKbm7yWw8SsdZpBo
us21QonmxDpcGlaTcDZdvQ5N6cgChZgbJybPfSYcbaZX8s7nNDfg+WGuK2JpG/pi
gQuf/GGpQXNI2a55ja6SVJdRdvRyVliNGvxJhwlQZjcgCtFIFJSJe+eUweb8tfv5
YR0lsFTX5C7/JJ57HtSjKkf8WSjq5MgKPRw2mCwSHQURfN0HmOB5EdChKMPY1AJw
d1R2zC9jm7Ho/dSOluFqbltxov/VF6Du+lS/BFvSM1G0lAAJokCpDeFcaWH/s2eV
h2FNpmMFmZT67cVvfRGMnK/FCl715hQm+3PZDhz+JlKsbqi3pZlUONCv03fR5/cc
FDt4Sh3XVi+LiqNl2x4/zQKM1DI7Rs9DXisX0760CC6YCOYCxWAuFQOq2ypt2B0S
C+gZEX7j52NNzkIbssKMuwtxVjgCCASCkflge1eFvIOQK71ItJFAPP/DggTU3KHh
fTdmiWaIZ6vec0GZvrrK2E8ybqQ42sSo4P323nTiucv9xvfip7s3fUkH489gCBOV
0sZ868XbAP5HIVsCDt6vxsFfIM48SYnn46Pb7aWgVl0DZJq9wmlOKxjFdSOSed1n
/StDz/TodkMmzj3ZrUdNBZidjoFZKOypxOVp67HiehBv4qr4jWRw48vZ+Ai+Ed8y
4pDSgeCsah/IWTKwCPbp340X4Sd54z2Q2KX4uQxCcE6bmYoYLIVtWQRmCrItbJ4/
F4465FANudEhebN7Rexd+gqLGy9C/FFECzTxHYKxZIkLPfKqwv+YC+yGZe7CW8kW
zzbmOsDUF8DEamJ01QtlkK1AjeiEc7Vri1fBUh1wM/579kVlJeWUzrn/YFaBiX4q
O6nf1ewkomKEiHv7VQ8PCf5mt90oJVUD2+rfEQfyXqhIm5g88oisRPgXZA5KuolO
SlYo7lnjKD7VFxLJLw4ZRWBYc27cP339nwD8UZy8URjeoWqFutLCjMqm9+sU09JU
ZsRX6SYlAFyfx4oeAg8su1EZgatA260pPMklWSuBIM4NonD2W+wsH3TRqXEYXMI2
xADuFWjj+ErKwvmqlYK9RD8QRlm+UXE+h87H15SdVDucm/cgZsJZieZ2ebe7oJpG
u0UX46OfCUbmJuTZsspV177OPt/qdSbhrN0cKlHuGqPbATVyDwT073/p1+nPSqRS
AbepSD2Dj5x78kpTu+udDaIlL3EQZ5WDWAONJcygWSuzLfIv7jlguM63AJbOIXkr
t63qrpVJj1ZBPXvM2gfxiA2fMt04A40r0XpyBPo03hWbNytxhDbJCwZR0gr6v+k8
254zmLFgG05yUOq1bZ112jF1wUCAY3ogC8XbqYRwqkWLt9X8OBdChEI4yJArz8Py
1hiei9oU4T6xZvddHUwI3dFZiXs+93/OdS9vA50xJzAxi7G5xlcrEnFIN8Q6mROR
RIoE2hiOv7oMIlkL1+BYmAElVYNOLU3vobVgig+zUbsuu2mfjhghr24wxNmKUWUJ
qrG70KHuMuR6AzEo+VnwvWHTpPryIz3H5lJGid3lL+rqHn1dqCWc+wPXd6DNoWWR
Lz4Y39Oz0x5oZxiQgg7TpSmCa3ITQm8twbx25+Ha5ge/FKEvxkqMfR3y1NLR+0QF
3amFehzED9rtuSo1DLNoE1Dxc0krD5NzCtlJR2Pj4L/VhAZgsnq6pKGOAqhttXdg
lhV3goYRUoK0Yk8rJOa+ypTVBpy38T2+mRL3KbrpV09R2qxDXV7TbNse6p8iVw8N
Hb306p4EDvmopZ6hgV5ekWJp+W5apLjFbVdmOqFrLvjxtlXSZ8qlHl0Nz1a2YYi/
L4I9+9MAhxxsjVSd/fAF5PQ72XmEPOCT3pYd2dZKQfiWfRDS/65WMEVN0xsjqXOh
ZzEfKfjo6UoqLJ2lCvgu6m/ndOvTgtSQrqAxcDI2UikX2SRaaxmw9oiAPOIDon4a
wDvnwH3Q4tYgMkxnYSYyA9i3FNz7QqM2Qn5TGuy/u9q8Q2cLESKg9XdnviKlSy7G
46JAAotMaRaGao9AtJZb5DKEldWvFWKNMqRrc529iPfpI9XsBmKQATrHkTB6ZBEu
AZoX+HZLi7QJVi2jwUdL4gMnfy3QZXxJlwOWOzb/uYZjANAnEdLE//0mIsiuEmUd
c3/hKn1oMmNIpSdSsXYTV2Wla6gcKt2xBBnRwGPxyYoEPFlZYk36lhvVEGuOmYm5
WolLdjwu2xbEFaQ/f1/PMRpmhKdnduV98KgWYDPdC1P/VOEyumVbHd9XQKhDegLc
dqccW3+HHF0xVp6DVCLG6/qtG3KH8nZz+j0T6GEaZ0L3aSjeksXFKECJEjYSzb9Q
FZIV4xcRKiAlWWV9RvrE4ltq68NorR1T7HmJeN/rjq79I76CnW0RUHcrcTzleEZz
Lc9SRm2uO4ZyeIf4KJwebmxMiUIb6BZQw5aT/Q0QRDLeAIbe+aWM3G9l3kyrsQaU
LQXzqT935OlFVl7CRipLBMmwF59vg79WJLtPynhHUpp6WO1RUj6C1fTxI0N+F7ld
JvF7Br8pRiAxBcfb1tZ7m5Y9CA9QTWlzp0Cyd81hCrk69Yrl+708Q+yFSmSUpBy7
n3TWDEgN9mGRpIJTXWwEgtwRQrq1Gia6rA29uSHcsHpjbE5H5QuvpW8IHB8xmVr1
i4f9C7rp+CypSZNXvHj0+64WZIdyJWhsTltE6Us+NqdBsPc2t5flKQJsfeC3KW1V
GhaTtEo+qsiQI9VQ/45zDZ/3X7y4ATtzAyqp176HyaijPyE1hm5phYKyCELDRjPN
ZhipW+cmO/FfQgg/GWgUHXvTOIf6kAgvqmbyIXGGKCpwIk1RnCoZTdHRSiUba9CK
Y5cVjdJRr+sp2ooXvh8PX6j/yQO0heevCMYgH/89aleCdF613DWXlfl9NnG9x7Tk
T+E1ZPzz4HmWzKGGNmZu0bBcVlQeDXvlYDBG981CFrFLeyX/MS+BRfyrwAs67odr
SavoRSdXPGFT9mPbO/mdoPOGF2rxJK0dHaD9mxE4MBtZF0fhTViNmvAeezDiy856
J1r8WOjnk0RmZM3/f9DZrtbmsW1lPbZMvXi8kp1AW5LMrsmxDFsNy2aXKCW5KXd9
1HiZxKDdTjk9xdXhRUfKx0/pd8pCxZXUw9kqvrR3ZchLZ6ox5AXMn5hOqXigMn7J
TzG2NRWvgJPhgwPWgH5mpuGIctY774HYhE+XfX4ggP8VS5DR/ak7q79+qzYG+xa6
MCZDpNb3Jx0ujymWhKOoJEYFpPZkQCEjwLk8mTRGzposLVH+kMDpNZ20wO2OVhWC
qi/LWR3jPwZS09CS8OBzMtPFGYPxtKfPwN9hTce2Q4tyEhiJR6SXFFLCuf4wi/9e
AFIy+/HGxavRvy81++GOE6VDfRDHjOMWky8VVFJoEDOTyfw6E5imeUUKzR+aVeHn
LFcF4LoDlgrRgEmlfLAx7rbk0JCfoDWhN1e+dVDUJRCXtDlEeCPdHkZdd7thrghY
cJLUqYDsLi8F8wbpeeAkHyxQmAdofDnBngYPSO92pZxeXReULXGDOmrDkir/JH3/
cuMVwQhtVn5UHyt4SQdsb2k601aO57li6Mt3ZKsaNu3Bn+WxBFFXQfRkV4djv+jU
+l2q0aNlRNULHAWnXDEmgnpB11Yv/CC7DiI29TjBW+z73HZUBxBgU0k92tHqdCmM
2n2/0CmcG7cTbFEhQDOMhai1/yRV+FP4ZFsncpyKNVIDlO0kEWmB1UiPqieqr4oP
wmlWRXz4i5kHn7qc7dooUeAc4c4xu7WGO0bqbSlr/3b0fyneSSREuGqFhO6AhRkX
6WGYGjq5tGxvAAYnznhDB5Pi/70BnDuim5PAmcdMCB5aGYJ2xtzFnfRoTuD8CNhk
TtMaKfN7c76LqmMpfmWu8l5ULcydIp6vZAgGo9jM9qxFvYc8Y/JnKgsDeywHjbNE
Tt/HxyaUZA/eAmq2K/Zh29ryn0w1wEzm3xHDmqKb67TKe7IZpKiv5KUywWojt0dU
sfW7iPqn6xL5KLzjxSxrqwABk8Vl4dWZZuPdP61PaBJoM3hjtd7A+nFsgfi45gcI
tGJWyOMTBKS7CmXEPYdF4IdtEJfWyM0vlW2EASumgGjJBR5f03YLbJTdjVPtJV44
kC+FB5c4nJN4S7NQMzB9xAE5x274YU+NG5a2M9f+6qVJuL6euFL9U7peddWRgCAv
dGhlF6/jflumKn/4mijevFtR9HtLKUsGver96M0VzsNAPX2F5Y3hbFofiR8WIMNj
Q1jRb4p6GqQ9ZDBHl2BeHv/qJwsiFvqG4+lnk+YfYN3dkeApPjSU1mZI2S/yn+5h
ISliTMoJnoAhUl2myhV9cPp8vbEl4DJHQ7mQr1hJ64ddSM+5PAEu9XQaMr/tQm7A
3v0glB4LLdruVmaUXvFD1S8x9SuW4QglBmB9i1ACuW7tL1KHV/jqQjRoyAqDN9cY
4w5bPflMNTJUzjnXChiS4y6yQn8dDc052WnxkN+kl72pTKm7RQUQ0N2FPmppkXQ+
CWpSXHMZUWpafnOHPfLOKuGYf/SfKnEccuppkh8AOEiT5k0hNusDc6TXSGWOTCJW
txW+6pZGL2Z/Bq2hxTEtXuCdN1xk8haSv8O24ZOLfe84QnUxwUbghZcKWlSry+fC
1GQF1Wn7RsZx6wNw6qgswetD1YH+iPD3PNRPn7mpJvu98VpM24WWgtm9jGwa1oK3
mtG2w9vLuC7zFaz7zEoZYHag5i/KhNq8GrmsGKxxaSDy3aBpGykdn9n7502VO36F
Rkr46chtW3lWE3rSupJ0VZb9H+5N6osQKWwE9qyEEz5aZc/+oDcrprnFtq6Iw8uA
rz7Ma4nqozeVN1DizPi4zvhWyEbOrf8+SJxuLRG8ViKjlwMAd3Kv4Ll/YaKNMXS3
pBgrBJxXK0OyqRm41wItQKwhsQHfBEyMiOxU9YDK7W1/pclbF35ZKggKK2HBJXM6
0SFDreYHQg3MPoSso4NvUbU6OOcif86Ed7X/RYPrZRPjyGWYSyELhak+QG2JyqQS
pOfXipB3TmSfojDB4opkUSr3uitUrf853b1Kyc2sHoyRBA5YOgmY5LRtmalcDncY
AywvoHxGGaR1g7qNxZwlUghX7HUn7j/ETfYe0+BkKSVGawmS+eCzQDWb+s23g1yz
Du2Uqf4D3JfXZ0tVEU3tywdG6+Z4syLPfJFxyQEggrOJqp67o7ZNqRcTZLZvwlaq
D8Eur5k90XU/XHcrNvoLr8Z09sm9D3ukh615P+ADxIqjVTMSHxTUUq4a3OZb031G
RoytxLqJa4QDFPLti607+aHdC258lFyi6oc0Gf5d0D5x1ZwBdgHQX400zWiZuL5z
q9RcNVHp1ma4ibmbzVchsZOf3dQIT6yTJV9HBZMhyd52ItA8qbp/wWRWsT2HPPkM
AIDGPQAzm8LYSYlJmnvIXVMFcTMI0RuxT8SRLL5fS5NjCoMdKi2XZkD+PS19jzJa
tXqTzweeFHRoY2HTCJJebdoi/i+UNJJOnSpAuuMBuVTlx2SqfGeRVm20XlrZgwjt
fj4T0LT8E8TxJzpRylg98/Jxkjq9WIzZQLf3kaC1hYb9K2mRPYZEyiqSoXeRAF01
NppKJZU/hZsYcNLR4TtLHdEb1yiop34dkuRVwfAs49otmSAdxQkoZzJfkp8Yvqqt
8aBqGYfiTyEmJ3jBSkQwuPfECknY0ev4hBPK0hBEHeSbQ6JhGH873zXg/4TpZiID
jtSGWio5F3YldSyt43rnVdIxiQjzGi0oBWmA4l6epfZU7JgVQFidXXRbObz4WrmC
i70oEExxc1jiNedUtI7BTkwwpaQuIsLrOexhwRTlFiwE3EEdL4EzAEKIN9hvPUcs
B/irWqEFWh/wGjZkcg6XvSDMYFvXNZ3mjpcjSOTBxzodLnLUCBz3XLRm4tA+l11k
PURcAImoJEbDJycqUGS9mqyRq4fGb7cb0wWSEobrdQBuUe9ib09j6fAOUd124+5d
9JzhQYefF5Gn946K7VPR9dnLFA3R/1XdMugnWFdK9SQCO2emYSNdWuUrd0v0wTaH
25UC0dUTyoijH/eyn30g8TmMz0YoDIV/L0hiKe1RXtj/ve+zViuMIzXTCQF4K59P
TNCXzxoPR16sHNH0G8NSYeBdRJjFU76m18JAxv7vArN9W6C0airWE7RK1HZmq0mj
WG+/b6lM4+F5dL4EivdM8cIJWqHG07su9NdabvSPEtbWs4YkwWJxgYYY41M4in4v
jyaRWeg5WmeqeIqb5DJr17YAA9CwFWXYd6FFmTs+7kUE2Y3OWyAWS7M92HOJajRR
7zZUMDMgvDM1YBALEJjBABmzCAm6JMsjeECvRIlXX4g5Pg6YlVlobOeTr4K5dNwx
CWmp2RSVI0Plrqo2U/wLsqMjU9LceDGCXLgxWepg3E4HeYuYmfqyzXFXwhCbjIgp
uBkYdqHBdNGeZmqitDNmSULfBwjXecYBurlHV2FAFnnmRTJgKIpi6B1hEHJC35R0
gAbWbxf8BHK4WegHphSHB/rtcOE7a7z1+/ipm+p+A67qOi8GvumHwBv1PAZNAnlP
lZS16/8gPN8HzQM1K3sZbTHTOQ22bFk5Y4hNCUCh0dhglCyVt9kfAwU1KbQ04grD
If5wfZ0xuyGb2R/urZWfIya7/pzlN+YBK2IavgNpRhdhRvKkR/ayfTaq6DsWWzk1
MpTUBibNoMVo4Yr/ooZ1WraQVRxeFkk73R70CqfrseTysq3c+76WBtqCBWHUi88R
UDigQJLUMH7qVos+iP9Cfw==
`protect end_protected