`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
ddtXksX2+yylW5zu6QL2Lhnb2d1sD00763mmSITNX595NcHTEkwn0zB1Dry37fOW
FufOhVzEJp80NC5qZ/+F0Vk7Ik02dIR0elf3clrjeJRK85K4e3Hoo4xn7YbFUIms
l/8VZSb14+JVGURjfswrIyCUotIzlzVYZ6gzoZwDXIi5gQIBf/gI+KxNXPaKV+PQ
Ufys/12rjO6aI/pPlqSm0hCvftmBcnezN2hk1UeXgOIuKZnogjOsf0iJVX2aOOWE
6pD/psybjbnsNB6kH5uFTA5frkzIzkzl5d9+YDm9OyC+k84E83I/7/j+rk4L2dah
QJOvksSIzN867/4Qt8qYTQ==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="MvBXkzurAa5VTw+1JJ70nePUfoQXBvZOku/SMmg4TwQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
oRtzZL4VJ4iwysPsC8SXYCzXS8Fw2gtZTOskLcDV+1B9Nzn1zTyNtlo6lNICRmmK
ZRVu2BmCc2G+fmzynYlNTnSa7C0Cuel6FYpxCBlOuk3OF2tzAmLAuDyOH3Z1Yjzk
a0aHuoCdIRKv7BrZCdALt03JeUmXKPdOmIlkVGFl8yw=
`protect rights_digest_method = "sha256"
`protect end_toolblock="Jn9CQpRhJt4rnzZPRk+dOpzAubz7omckX1MrFd4p81o="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 5952 )
`protect data_block
gD6l00tciPUa6pDNTk/+t0OO0nC/UTtBwLB41d4inuAUA3i/ALrNyoJVcBnAmEQW
ptbcNp5fxEUJjnOxnedyZEuEBxWRieZFQnkRdF269oPlU8Vx6MbEsYgPECa0rfRc
k9j3UXqARLfG9MqAOnaViSKiLGH/p7leWwU/beltWy2We6g3jYuFeiDsf/FUy96y
ZXkXjQZTlnVVho+W1MEbtiMZvnE53og73mdutuKfi5SkerbYzQA11Ilr7CBitCIx
FoxwGE0dfFeiCGSxZKcKq4PrxwCOo3hk1yljOwydMM1VeYtF6QWcZqXBhXLi+FuE
PPHprYfHO8xMFdiTnbuqgeO2HKx1lz4BT5ycg9GhGybei2gwWFJ6S0oMkMUjYTwv
Cky21jkkFvr7mP3MTmmSOV1K945SOet8hEXuVFTXOMAPqRAIZ0yTh/SAoaA+UeWf
ba3qmN42gZnqyjpiG9m2qJIZaptOZ70RBo6VhpqOFzwOvrIR2rCS27cIU1GneqmR
0Xi4wg5rb79EA398M0Nw8B7Fe8CqlqnVszysv621bq/sPtlR4ds/r3IsnJWKuUM7
V3847wP2WnRzbN8zRnvC2Dam7T4wT+uMZFGkCnIby88ZhzKQVcTjqVChHLonRcS0
qQYoMIjRN2VPq2SNjtj9wUQScTAIyIun0VOGNqjFQAsDt6IzEHM5wQ2O5ukVd/X0
Vk7W/rsT0lrhDFsNymTMVXDwtLBCp01eyCtK7mduvG2fhRvs2d4q1jc2ZIDaBdrW
YJCJR0zVUbXOdedOokYLgWmenSP8gEUOND1qX79fMUtBpKr5OoWEcCluLV9vmZ4J
cUoiScio/Z9h9FC+oV1aUQrKufAZvpPTKeJ+gbYpuykPRGOwQSNDMjRsJvxKPDoO
miYoJHntknFSnIFZDyzctWiC8rKPQR49mHZEFi/HWXcBO2IXYiidZjYSKQIoE5Aj
EqS82gMVSXDzthSEpk3yOCOlEsbGDcs4PfneMMvDmutTeZDhuPyKYzfbMe79x7JJ
jAPSGwwerPtM5RFLp78R3DYUi8CBN2p7Zk2GQI8/U9dpS4+5mocUe6Sguum5UnvV
LSZMj9rAwfhD4garFTSu/4r042i/k5SOd6yq5WDch02yThrWz6rcbSwQLFIS9I5p
6zwxirz4pBAoOwYyTNowdYUTDF+9o2DP08cYY4hP7vD5x71jY+lYkIL2/PcuRApD
V1z/eNJE/1vDXnOFjDZ9+HD8xFB2yaZ1k4eOOmMGENNtC/Ud7uwTpxDCmSRbLKZ4
OSjAxGK3WrUnUGdRuBAs2T0pg9rA0GptYmx4BOGDApAR0bSy/+NLgwiSXeYEcbxD
U9GMB8NVPDcZr7UYfYmEf7GqL5I92AATlqOrL7hBFjbjKKlIGsKlRKL/jWDdBRc2
+W4yy9rWsq0LOQhhE5fIPPuP8ZEGq9HKMtlOCazZooGkmGcujyGhGT2w7lvHuK00
7uW9X6oKmoTTdcTxLzEDCSzyJxr6aBquX2c8fT5nb9oSleyYPNdZQ9hNMPdd9oQN
KctgsRB8GAI0eeyXF7BNQhcTyggyWIRA4SjBiyXsgxdNI1h7vtdj3L/d3DXe2Pcb
A2JMLvdMccwffuQaSr868OsiS8DMMyxkvLdPrz35JYvWrmBFU+hxTcB1ugWB3Zne
m9R3LinheeSiROfjJOWH083woKaq28nK/WhjVldLBJmsNxgH5uE0L5IgauzZmRUU
1C1cywcWEtmyqxqFkfCrBgShNGCcHSkye8506cXllHQTndd+uFdlwT6ZIOxtDMci
iUfZfIxKCFGfVEp87BGk3iNSCalpICatQxXU3Np68xwi510IbBbHvqbAgEyI7Isc
KW14djhpRY8vYK2mrL+4tvIx2stBF150v15HZnrnCtAt4FR0SQq6GlYAv8ki9/SM
9IzHFO+p8Alo/HjLbOUdscekdcvUwXaWiQ1udQPAxaAD8tRa7pVKxaFgVmPh8ISE
p7TJwg3SFGxfPKtXswhfTjnQJTwKt2y8f+NS2P/aT7tevXd5rQX6kZFEqAlAhxOR
UNkXGQPhBLyNboZXCq/NkixR8Y73FMpPk+XWagFSmBEN/+D8EUYzzgPTAy0NnMs9
fVznkHx223CdC//dFLhiWl8VL7P6T4GHP4pnatNQ1ponym6IXTF92M9IciPuGKCf
iBLP0eItwaLpiVCxQIqrI3cCMW4kOLD6hSThh+o2hJNU00S4tDiJCq9It9XxPt6k
G2kktRQ7f2Mn0A+S2KxW7c0Dau3tQb3FSr6hjqz6mKDwGSbPRsi/D3X1asYwa1Bu
ZDOW6bBsDUT0OJngcSMjmoL4MJlACo/ucxyhBkQJ/5uxk3bTrvP7CN4zgfzLUdl1
euxWIqQVBHWB3/kIE6pEY3frmEC5lpnbmt/EmRdYr0SYS8MnI9bt1X7myugazS1/
+/N35Zewp8goInCg14xb6lTgv5L1l9M1C6g13rhoNd7wS40gLPlrSroSEdfxAryA
h0+Q6cjr6UfL6/NvtwvFstnaM1xYUPJoLL+NiuCVobE+vBTeJg4Fh4YBxu0ktA5R
sNfSWRsSQiQ8zUBaM5W26TbgakWoCTbNvI4vodSnuSTsgslg0n1hFliN4zNccFU8
XlxsXpNYxFo5F+fscCOd5BG5CXZIfn8Cg7gYJx3DpUGtwcD3aD5UkN5giRRTjtVJ
Rr+6LI+cZ04fvuUHCrCDgv8p7EvCwupPiuhcvGhWKuVrBK7M5xf5/SN/2n1iP6nQ
5YEl/ZmJJUVOCBg+KYWx3UakY0PbPqtdCXHGZuBpkny03X1CX4O+26ldq/HPZkp7
DDZhV0Jyay323RhXw0sn0WwR2hMjldpcnwcf+o8OBa3/Ek/F4L9SjNQaCzXBInul
Yk/ZDj9jvOIcLLFtQcDch0F/ETwkdrUgz76kp0vhy8TzjuMEyfQIv6tCE7EiUmdR
pk2ku7ttA/+O4UIhtRB7bzRXD34Mltl+EQnmTcczPiO9pYXLIPC+DGjMYvealrno
RszRjgPQomvpefur1dNUbAYXhWHyreWwipIV14Jr9TFlHJst5Y6l61mpAVTRc0UK
zT8+PRTC+W0vpjF15cJnlq/bOrkwy2rCrCjm/ZQaGu74EDpFIWfm90Q9YyxxcXTy
OrXPOR/1yJjC7gL0XAtca0Cdnt7Okn0uxiz9gZxiRuoU7NFutWvVKprwFOqy7vQa
4/FTXgAV417RAtC46gKt0OV4PUpqV1ypSp9HmJOdlOyW+ZGE2atabfWHkFdNbb/d
hA82N5yDp3CGxKdFJpD8TVd9wHTu0FUBCUkuRUKXvNVK+IfJ52wAinik+WcP0B/K
GrT41XCabvn39lDBHbaZcPNinK3N9LighHsJdt/j+tIPhUsUGd4rEbMuz/jrAFXl
FFGM1CcpDG2hwl/GYmNnXYGD55FZTC23vAcOCwepAsZhJQdmWbVnSkbyWUZcm/f3
eHOzDtGpsTOXkMUxRptRgb6LpaSKMOIemjV2Q450g0rnFWJfZVHYiL4AfbTkYzrt
4PJ3VOFp9iXdzQ2e6LTVM1LrlxtVgvdaqH4HFtIiCzqJBkMWaxtyAMObCJ4WUZI5
eFoPrrrPA+GoQpgLGwnwxZCP75iq6+I2uzKoJeSD50D2QkCW9fzHWaUHJk2GACUe
4lkQNL+docnhZ8Xi74toWtmRW+Xb6eAm2Zb50yfH47wQTlS5uzvF7l7LfH4jgPOA
W4WtddJ4+sh+hYE7ZLOeYMTEkBd1ZfavQcp85jEhs8uaJ78FfUCXcG4K4VMlOXb7
aOG5uQudVtcIDrh2CJCSg6HTg3xb1kRtyxuszXLH44998m4+5q3UxVmOKmCbc0n/
8mr40wSFNCNg/RyyKsFDn8Zpa14Lk3Zuu46AyAU5j429oyV3xqdckPTExDOBDwWN
9fBh1Rm+rFLgXcz34meEHhg0WrM5CI8B8i/UXvm9nxO36DhPvRQ4qGXxOkqcWri8
k0OhIn/j0s6BreiPX2nDA92nWI0aV0mMYyn96W+2WRgH33tamh8xfU2tKGYumikg
ljrASSjH8C/nYV7sIG5Tht2Z6BEN7qfspGUza4EhuHp3yDGRIt0eENUeLQ2+r9tE
pLxM9HiLB7P0AMRrRTHfbx7860mgNtjwwJkfXI1uMlX0HvRuJysZHI039IduJgOY
RWLnPXH/mYrri1wql2Wi1/2hZDnXUFS8TWgruzHCrw5hK6/RrSPqKXoDeuryLNaM
EtBDUlBReo3zJbMsPhxEWT24ctTJ/VW4cUv9nV5h5gbk5l/k6GNygtdgwGPysXpN
ddXF64dpp9eu4jOaQgf0hALOQ8pXFYY8oHtaD8/Os/PPrroOvkYPvP6yzAEgqlKs
5FszkC9BEymMOlE6v3rw1USmrYl9qekEJvSJWAWtkYY/5J/j1qxO97MWhHG/2nFA
M8Ype2+HnzmadKK5wtPQrYNBHIHmkKXnJJ0D6YhiRyzKSwD8pk9i8Q+Ca659NAys
8chykJGv3UjJM2VVDR+rDFynYvWGeP68uYZKw2W2blVnp7/WluZxfyJZU6w8iSqd
tx+LYaRzfUbj6JTX/ooKNrUC4kKzpBI16v83ptkeEembk7qBe1F8NgEEy8dBIFbG
jy2B46eeK4OTO3bMOdKbhEDScHefpqGBny3tnyPS51Zaw6I2q9kkm94UDeLET8LL
YZY+TmXrxAFrbV5hvaIvbd7Y+nyxTLe0o4Y0boIHGAmVaGlRLxKi/HujFqOUpyRK
aT7WOkgx3u58lI4WqiTPSghYAw989yCP0OOdRE1OooV41H4635E2oSni+Lkwxj4S
zOOO/SL6uh17UVec2Zh5nA5N0di+3o+WUFzr6ntKgNAmi4/e17Z3lYkhZd93iuw9
DTnqQoMwNlTrQ6MXYs0JDQshuMfmc2vNAVbU8eSNXAbso4w3joMM3l8q6FkVVXMX
ADpzVUhZ3Cu1Zc3cd9ZP/Or5iTSRno0YgB6PtHZL1uYgJAdte1ZPHv8j+74fLtM3
pHKGbCxtQcs/scEek5yYhFYHvj++4m9Kmh5fje+99m62shTkoR7I4mRP01udjSk7
OdNMk0HCCikXhpowROmmj7pFjdYxF43ro13wS2VVgTrEs61Ik7PmboIUmSktcJEQ
0Lw3MWjQI7w0mhPhWFtLRKUWBwxPZlTBIJjFwAG9+UMRpT05qpx86cJ+Gz+p4yrD
2n1DdFCiH79Hs1iVmImblpLNiW5o+lqFRjmO1zxudVKVEk/FUNYSDu68S84oz9Lq
cxnXBMmgmTVPRpnpRii3UWN8TN0QtlyCjMw15GoD55jTGp/6Uq3PfGaAiF2yBAza
NPoSt6svawOr4sWBV9UdtBWbo9LDYhjycishKd67rV0lD/VtEnvzqqrj0GZjBMHf
Wr0wfn6+yy/xFL8RxpjQM8XZ+JhbsSM2xsKEt9cranFdIEo307Q2/61ZhSH8Lykk
2cGLJ9mZukaTwvHIkQjQzIZfFPAEbxmzB3/i/ynRiBo7o445qyHTE4RShWmbLkqD
I4tK2GkdwhzrW4MNAY7hf8ODEGcv08JIPdFt/4vMDZfIG9eNMQJy4Ys7cjS3Ogce
YcZGS7iwwBIwtabFN7VvVxFE4IQO3/OEQW/zj1o1ZJrZ2cQRuHoSX86YICo9KsJT
4kdP/Kl49qn1DPTtrEJBj1ZoKnPSVKnlKLi618BsKE43+BN+ATeybyhN8R8gie+R
B0pRDJUPgT1QnaYeawdCJxO3tEhNFSlGVA+K/tHMrn869bvV+MEHwzpl/Pqo7EoF
zjZvXqR0t5OrOIcpjLE33oAmnB2zO21YOQbw7bjZsGWuwD/M/KNAd7gMTLmoLg4E
RLtEeJVd99pDWdh1lk4BtblvZdmYq6Msronswf+n0WJARAm6lyuvUsoLInPSHk/8
pc+YZ9zKak80lAuX4ORD3f30Ar1l3MxiFDxssYCKN+uNEp4kJFny868W/wumxfgo
3KBfkL6vtxwESmVfX/ZwLoNX/Ha9xl9yPcrpJUQSy3gDWFK16P1OEoteBNzfVpRR
PLNj70Pb4v+CjpADI/Y/aKfOHW4448XIe3sRsWYaafun8S72qTvRE8A1SOiugDee
yzVQMwmpIjhFxfX7eeOHmwDcnFvU/eiSjfn+RQ8QW+Qj+0e2yL6q73tN5sRVAMTf
RZEpjIFQILUSMZcJDYuQXT8z7NUQcD1N1aS0pHwT7blI5sVNT7umd5rrrd5M2VVd
tMHbkUU6muONA8aaHE7oypqmPINXAfUwYHI7VvLX6u1F9AZsEG4ROrWxZYiPHLqs
iKiTbzIdmxi0Y7cXYvtEE6WvQVBZ79sk+8+MXF6C/jz+8bK1UbPTLDk0BLYOc/hG
z37QswD/JBcqyalew9PXdUapT2/sl3gRe1XMpu//M5dvgGyZnoN6FBlUyUFNtdiN
Za0n3tT6cDVATv5+HBkjOlDxY0nesXn44lnaePyOztznFu8jHuKn3r/vV+6H4F38
PPassiAZrrsotpSwpMe+2GirrQsMFli4ozwGnRWZnkQn9EKJfxAZW8gGbhhyudLK
lkGTOAiSR6uWBmbTzxxmJxi9inW+fEtdpvgkzt6R/z4/uqnkaHUbw0ZDfb+rYsEV
Pr7QzeiSsFmP4zcR7NI3yhti9DY7OGb4mWMhyIodxqCm81kQBtei4un2zMGi1ZhU
K8cmb8ABrFWGVrG2O2xfb/4+IWibdSAovhhkW3twysl+sRODfeUxacgnmWdtytjQ
eDiJnhnuIB3wAwS1f5xP1Siz9DFojRVdM+YXRji7q1Sczkyd34qn1W45MrDk0j4i
026Tt08Ui31Pwm4VEEZeUzGrMZAXWxIEdWT4YLkaqktp5T8VC3i1atZ2gLwSS4Il
9bh9Izn/rIUyoGRVW4xsdBeC2uRkGDYZTPnCCcpR7eK+te8ZH0d1mFJPpOLJS5kQ
IuLWRg1awyVWmf8k1PX8alSlyAzIT+cW+K9de6p/3P1QkgLEJ3bzESlY1fNo/8oB
WoLnDGBs3bXKeTWcoIxa/1hSOY0qk6wZYk+AVLqaNznzhcPre536rnlVajCGNcMi
l89ycqUYb+UM8MQQXaMtibem4CXk0Hw6y/j1z2hrLxgb1/4n1AQgZ8KI1d3Y6tEj
8VKCfOuNqhptYNQbQ2A2Iz2YF+nv9Oy5+G+B+9SCXs63Esa+2Av/TnoQ+7qwWV0G
B0VnrvbUkIFFo2wWFg8+Jh2SH0+TGvx25MeXQI6MdYIAr5tNQpFcpw6RROXuJw88
CZU8iDbwUVNMIHPXEKjgUfjqoWk8wBlyyDmPHBrqc4xzyCxSbqDtSjhJlRUC57FO
hAZnmbYXn0acLSzRffnXhN5sAuOCxY3uhV/aLrG7lBxrewFXROQR8B5ihJfravib
ZDPX83lG3n5mhKLW3Y4HRxcguocLXrglFJHPJOr0XGN7q820W9mDnzM6+yVRm75y
Anl22Rlf9Z2PNkvanKWC7iTvJ5opnvKXNo0yhfhTqkAQ2iU+5OpG7zKYJ0Ph/bCK
+jyce1gfgYDevjsfHS1+z8BBuiohHGWvoUtaNcvsHzCF7pu8ubgp7/EKFsACq/pX
P5ZRY/iO/A46Tr793xms40eJM4As7ZiLrMad8whKT9faulx1MTEleD1hJIzChd5Z
nZlhu6n9+WC9eHTajNaTA++GCF1k5xw/HWA/newuBbjaxjuB5lm6NfsKZ6c4+4pR
EpGJphDbLBDoQnZykv6amZ1496bqDfyEHMjoomWyHDJBbDeDZtgTXXnN0qXXH6M3
A1W9ZmI3fZk21kmVKB5Ql+7B5DukKOke4PiAnCWLF8lfLNYsKCG9eoOQappzSTZ7
YAKMkMK4N59WmG2H6sBN/HDmfcAfMS3tnDtQ9weZbGQTLyUASCdh4VF1pyK+RK3C
TLk94i1IMFJIheOop+n3DyxD0Qiy8JHmFdjJQ0YP4hGdnpIUUzYoDc2Ucgubm8vg
`protect end_protected