`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
ddtXksX2+yylW5zu6QL2Lhnb2d1sD00763mmSITNX595NcHTEkwn0zB1Dry37fOW
FufOhVzEJp80NC5qZ/+F0Vk7Ik02dIR0elf3clrjeJRK85K4e3Hoo4xn7YbFUIms
l/8VZSb14+JVGURjfswrIyCUotIzlzVYZ6gzoZwDXIi5gQIBf/gI+KxNXPaKV+PQ
Ufys/12rjO6aI/pPlqSm0hCvftmBcnezN2hk1UeXgOIuKZnogjOsf0iJVX2aOOWE
6pD/psybjbnsNB6kH5uFTA5frkzIzkzl5d9+YDm9OyC+k84E83I/7/j+rk4L2dah
QJOvksSIzN867/4Qt8qYTQ==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="MvBXkzurAa5VTw+1JJ70nePUfoQXBvZOku/SMmg4TwQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
oRtzZL4VJ4iwysPsC8SXYCzXS8Fw2gtZTOskLcDV+1B9Nzn1zTyNtlo6lNICRmmK
ZRVu2BmCc2G+fmzynYlNTnSa7C0Cuel6FYpxCBlOuk3OF2tzAmLAuDyOH3Z1Yjzk
a0aHuoCdIRKv7BrZCdALt03JeUmXKPdOmIlkVGFl8yw=
`protect rights_digest_method = "sha256"
`protect end_toolblock="Jn9CQpRhJt4rnzZPRk+dOpzAubz7omckX1MrFd4p81o="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 4176 )
`protect data_block
gD6l00tciPUa6pDNTk/+t0OO0nC/UTtBwLB41d4inuAUA3i/ALrNyoJVcBnAmEQW
ptbcNp5fxEUJjnOxnedyZEuEBxWRieZFQnkRdF269oNw2hN+b+yILES7EMbvIj4+
GhyWzBVVMaoH9W043LnqL5sLPDmY7smV4Zr8zZCxw6vHeaQEX/o/7byD2BSYtaXF
qj2Grc8qrHeDO0etXl1/eqC1nQL7ubUiXqQEZo23EMpjKSGM+kojvab559Lz2uby
9G7SuMkxeGJ4F6yw5lbx/bNka2dfjRrmGXSa4gZjfxapOP9Fvps37Hmh5VLz5W/K
B7ae7n5XwNXxiL49haTExVUZ4mFPtUV6UkF4TsjORQLriLjD4TUjMwTCGWXtKUKz
+APpuoTD4w0sPzaDx3mEuDD3pxhLK5UssIUgi8LRMHH0/ylWMYX8rRNS0km8bdHJ
YLg+r4HmhUnPvXh8u2t7d6MM3dkZimnQvklfY+ieACjdQ0wbxATuHmd7wKf31ZKt
LofU5VPKaly0rEiKVpsg+ZgP6vhESn9qPMbwetH5Hlgqb0ZbV/F9+jXPgRVIcrDQ
eDL0NAYm3c/Zj4+jE0P5/Npf9UjkIPorghW/09XO/2M5zCzA3u8sHqzOp7BuWkmV
tjJlWy5PIyGo83AXb0VPRtRbwXCMACwwoZTVjxqtCoY/IPlUCsGgXhZx+xyZdy/a
38Liuny37Jqs/+9FKZf6DIC07VrBEnUaVV4BsQgvZ2vmhuTH+ZxC01vqLq8JQGyr
pu+YWQGXR0iTCfwb4pGlJm6WtC/DYKRnIyf3FHkjvkXJqZR70Or/3HcWGOwjDAn6
UQNjlzqzmiHt5JIs6izJ2m3W4b2sr+WTazRhjn8PeZhNC8vNKPqP/NwsnNSNIVeQ
dgdqBzJfc64sd8/86Wm0JnuspvQNX8lCXHO8QE6xUrAl2hgcz7G1pEjsMSsNh1wz
eBChGXVq6V3HN9/qdtdn3H7GTG7Nhg9tb7E5kgtwaKbJ8ARW7sM43zApwl1Z75CX
bXWxJI9DBcWu2FGtmetA0aw549tD2sCYCnCZ1QvL66D7+/VyObJ1Z9gYIdcd9bll
dNgRKmhmrrhqU9vCqv0hWCH891HBawf6CZL+krEzFHYagKpZbMZ9yKQAx5/G2tqA
m8me4L9zkXqxAinzg79UrJy5zAXVuvrgCI2KdmA5tZDa5u2a068ljE3HRwyYXpeZ
s3gc+K0ljru72kRyvQZCaybz5TnztjQx1gS83Tkz5FH7YNRrsj2xq8UnZY41SI/U
jH82T+FHHwwqYId2u2cmtMs4aaS0rmoSNwMEHGD1HbSVddMsfXypxS4GnXQMY1B9
2rXS2ke7v0/2aWMzdYx7bntBP3QS/SeoU0Ul6bJnjQx3ir2szQi6wpUoo2wU8440
NrLjJxndYfL9uCF1ppaO/PXUX0gO1JP4wrJHNZBOtHjffgbhYGX35ph57ACgeFk0
GNB9XkVA/ydQz1CCtWHE8Nfoa7aQRnuVMv21pl2ltYgKViISiAa4EuRLBraozsI9
tjW2/QXTXayfZWv4TbX7cslmz+S9Undp4J45uwjRgMI00Q5OGChmdMEOuOB2FpJY
gKO7164my/XgucRS83aRnXzIAzZRLcK/0Z5EbRFP76iGtOyhWRvvwiflJRf4jcvt
1QPFX3uQbVEW2mzM40HZwAHitwdkC6YqDcgh/IXoo3xnJg3oUq2M7z+h8LGKxUbS
C3z5slTQnUwE+1Ocf0kAEcUFAoeMtUYvHbc3kOhfPGSy9dYvOEwFwi3x9o1RghT2
qYURI84oUFAAzgb1wjPycAWRmd8orEY3R5AKHj9CkvjzMecms6m8pSZDgt+gmmgo
ERRqsOifpfiK+XpWT8pPW65tX8jubwZuppD0p3QQ6FQiNyn8ygtSs6j5guxKaCz2
C/BDxOnDLm8Y3YgyCPQCMnutNEQYm0Dfzq053pHvo3SlK7XtnzBfp7vVjZpE0xGj
GQy/rWM+2MTz9ejNf8BdFF3Lmx91k/LkhrsqALqykzwEukCgzyA8w7sgR9l2yzCu
H/vwTwCkRcEuji9kCOJ0TD2BRmxRtF99AFWD5gNwl1BsXxzKT3ktcGmDYQozQvzT
hNQnKJsBZD3I/uLSrK+rPM+z+DTdutlftzspTbn9FDXuRQgl5boy5kQ8jXyiq3QQ
K8Nk9n9EVnDqPIBBJQO7M41zOqlADTb0KPHRVNq2pHVlygxI0O8jjpTHhzOwAbzQ
YDUdinx3crTE9Q8sgKzWREDQtiK44bnCRmQlXMjfYtCqAUGt86o50ppLXhhZWTlg
VKAFgCuc1ntjG42qOI+tespuofeW0+ES6FKqd1OwBl20mzCAy8js/AFc8HQaLfyI
mYFjzf7Vk3q8Z41+f3lLEePzpC2Pnd3inrCLmyWwvEKLF2bE3CrFkWGYKpA4lzLI
pC1oEn+O8K/66sq1PX12SBoOaFjBjZYgqp8sQa6sRZ2pIyAOVVfv1Si8aOS0Aqwu
9grD/M/RyObperCJuPdVcQZSUZ/wZuGj+ywibT4sRzOvVpxEkQHeki3Qm3DUAWaI
NSMiyhs6Y641bmqt3XzNAd9lVi/CkUhVKokr4fPBlPovEtWj2/haNVjY6zkvKz75
XmXXD3afT41xC8nMA4lca5Zr+iE3NgK27O2umHQt2QonIDkuGj6Krklh74BuQWW/
5aR5pOOZVIB2qtDMy1Tp60JSqeSAbe61WMksvP4Az+ulKrUqHVcYmIvFVLmLFcRT
0umZOswc1Regdf4G02yBs4d3/8yza25dQVIWRYaX8qejoJx/3aAHJJWrtTebmjDD
XLpcAcH0OzcECnZA9jvED7p/pN7vxD8a7nDi06sFXIH51Cvct5ow9NOxtN/XOngZ
8DMOK3XpCU/llN0fSS2gGVUfkE/HcKXYwie1Gauh07112dozevMoDuE7eDX3eLn8
Q3rMJVTIQ8QTKsWMZrcmK3BXfWVVsWwkhi+MNEgwgsXqSwKCs9qdcwGD6DYvVER1
JE8X0nTaml/nzgKrwl/N1F3n5FQDg3LxV8hOBWzhm5/UAlmh6eH8GDsqgDcZQ6KR
QGiAf7hvr1YxSc7w5tNqj1R1lNTo5z5gum4wuJAN1mvqut02YF4YhpEuLlEAov/o
pNpQBrrZE921NNncljBUwh9jMsMf54O8cUuj3Ungnp4tPe+pX37PU6JsrI9AUIuc
qg64vf+XeywyUx2qPVjLq7JDjcM9dNLkNec18AKTgjylnuxdPhXjBX9Nc2PsaHaq
o7cHL/qI9MCyF3umf8M7fcyCu1M1UVzxMz0zB/JnKIzNfTWDbCcJtcE8qFJ0KlYV
+N/tFWgNuQ4vLHqTe+yQQXPb2Yam5U3QyG6+fZCapvuzcTm6zeDAdVtwlBb0GQCF
DO7V00BGf5JR+/xfaL9q8DXKN36oZ8C0d+ZFWwPSBqvoA+hsd8CF5rPL5Xrrh50L
z0+dqs7b3lPPca74h2oaWkwdrXqfaFuAmbPM48WA/lukQkvvJYDHieMdpiHgZJzI
IObzmcKBFmsq3KVE0m+DrP07TuTkRfShNk5G1SA0DyxaxNDnM0HriuD6k8F8O3bb
950rOlpKsoxymAkIgp5HHXHh7a5LWwf5+Tq65i1DJJE7z4gTO97t5zUY/5zyHcb6
AHj2S9a0X5lrErcluMGeTL3LvWM8/0RbF2bPI47uVkyxqIsUPHtROVvjZuVNWt7x
f2fZF5E0q7w/SYlgfRhBYU3a1XF/Ssj3uX98XmQICfyRumnquYjrP6OqeTpJMr88
PeKc0rWzlEDLGRJpqr0bxYwV+WqfkQz14dKx8OIHpet75aTetam40RFbXK1RBzk6
Fgi1CICXoZQzpeUc3r6waovlGlPAAgWvmprM6CCkx1NHNadHRZZ/YJmbVZuW/ean
vtWYRQBgFP+/88C2ozpEPI2lcNnJZkf2qh4EN15hu4ZyHjbKL+XoSnqlaj+XfjhM
5hMpUeFUDon/TPuowQ56JJHg/lHfKJMUgUVSEQaknKPw9xcpc1WGRYQa7T8phNT7
JYsLrtvvITtI6S58ThdJVDmDI6a7PoohvRofDlaFp5SRJJc5cgvvHRpJXFgiAiNX
OqRYuYQibO3nO/29FUD/VBUv/oei21XWiIysmT6ceMBAYgD/dUuO0BufEmULQ6lr
MtTK00CH/V4ERCWtRv4VNqXFhGu2YVb8Tk2rrD2qDhJDfhEklGN4wkvH3BJ3E0fS
Rfq/IIWLdHZ1b4n/5C27ik5KQiqF8V4l//Fp+kOTpK7GE7Zd8th9g4+LVkOlIy4J
6IqO+lKOwEtxtyr5CFW45MSdsTd86t6mKz/NthJe0HyNKpYzOqu1+07qFL9MWYls
aqcXXa2T11fxZ9r78SeR/xTN+2nZ5i13frJ7vZwX5NV+t9RUI7FFlKOstmJbi2iK
dNlbCUKr71KD/P1c3bmTZnRIt9eSry6BG5SPpahGVRsx7XauVBexlbstSSdahzve
uLq5zSiALVL90678+5nXfvn+hyNzfMbzGoRwTUh5xpmEQzMR9LxGV6ZWSFhXzF0L
8lYvnqQGhsan+/ez0cVbjNF4HgLyOV6cY3lHE3nsaFSS+/nw6vha20sSGhv9tzWc
u/tnhsakqpaJdXmHgDj/L+eC+igGvOrn5kx1GJaAwLpGdZLSCaqVkmAtARYdvl+t
+CUQkvnFsHmFqTE1A3naxwcEQdZdyBxkpJo1Sx1UenrjnZoIiENUoL61JE52gSIv
R5lmssjemWVB1QkeMr8pXCwMQaFNHtUAmUd7yv/GTJLJlYdkrhOrsVHz4vUEdzkH
9XIvAfU6JBqpfWDzwGiejLBIStya/iI7iBYB2IEm8R7qAlWtT8OEcexOH4QZ2g9P
vx451/hbIfyj2bLYvcMAEk4GBKj5YMqyNeqLGkm0WJdjbJ5l0vRl2Ga43n58fjRo
4b6NYcIvnssVvOFfCkunHH47Woh4jXqnv9ydx/oOumJfwhNwykrpUBiifm5/OOsN
L+H25ONexGciATKAUQ3W0w1J3X6kxxOIGRBxuswqGksARGMzMfr9qLLdZrJBOtZP
rymoDFJxkzhW0Q/6Z76qafVINUAtafh4uPDvnlLBdkBs5xzr5CYpoJVsaPQix9Ub
2nqeTeew+kdNOvoldoaVgOTX7NVcxa1xBl0dF0pYPIGA4A61le3FRxf5HCOu6HKn
KlNheE9tBlGu8ZkP5UEyIJuMIw3yDqDGs6BBihe50H8IJ1sP/uXjVZMPS4nKpGkS
m5yKqxowqo143WehlBQUUpkwe4NojkDf6Ugo/FZ/rfW0FSiFYTVJNIU1D8K2RIDe
kOEUFbl3L7bMhB94UdEVZO67COh42rNvGOsPKNpHT+p9cZTctJc5NpBwAVbO+1EW
kbSi8V9PES4QYpD7gx9LEMqaq3zSoQLTR4nj6S+HD7rxpHZoHzyYEosgr8QC9tLe
U8u4abO888LdYW8xRn7E3BCONnan1SjNKAQ+rAL2BudgbeOxvPQYo0OyptTdInNi
s4C0M2vEDz0NdrpoAHianWWv7oFFUbzI8akw8ph22LTgz4kJ/nAOrkdkFMWXHzQ2
`protect end_protected