`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
ddtXksX2+yylW5zu6QL2Lhnb2d1sD00763mmSITNX595NcHTEkwn0zB1Dry37fOW
FufOhVzEJp80NC5qZ/+F0Vk7Ik02dIR0elf3clrjeJRK85K4e3Hoo4xn7YbFUIms
l/8VZSb14+JVGURjfswrIyCUotIzlzVYZ6gzoZwDXIi5gQIBf/gI+KxNXPaKV+PQ
Ufys/12rjO6aI/pPlqSm0hCvftmBcnezN2hk1UeXgOIuKZnogjOsf0iJVX2aOOWE
6pD/psybjbnsNB6kH5uFTA5frkzIzkzl5d9+YDm9OyC+k84E83I/7/j+rk4L2dah
QJOvksSIzN867/4Qt8qYTQ==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="MvBXkzurAa5VTw+1JJ70nePUfoQXBvZOku/SMmg4TwQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
oRtzZL4VJ4iwysPsC8SXYCzXS8Fw2gtZTOskLcDV+1B9Nzn1zTyNtlo6lNICRmmK
ZRVu2BmCc2G+fmzynYlNTnSa7C0Cuel6FYpxCBlOuk3OF2tzAmLAuDyOH3Z1Yjzk
a0aHuoCdIRKv7BrZCdALt03JeUmXKPdOmIlkVGFl8yw=
`protect rights_digest_method = "sha256"
`protect end_toolblock="Jn9CQpRhJt4rnzZPRk+dOpzAubz7omckX1MrFd4p81o="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 26912 )
`protect data_block
gD6l00tciPUa6pDNTk/+t0OO0nC/UTtBwLB41d4inuAUA3i/ALrNyoJVcBnAmEQW
ptbcNp5fxEUJjnOxnedyZEuEBxWRieZFQnkRdF269oOePeGrWkWAZztkj/liP+Og
FIkt5q1amscNfMSi+pbVsK0BwYEJwbvu8eoD9H/8eqEep+jywh10Ns9Ry/Ah2Vrs
sfW7wcjSkTEdYE5/ZyGNKNFWgO51ixoV9xMFak+TDzEy9gq8k5AJIbsDwGzgwv08
l2MSEKhoZghMzqy3hlBwa9oPZHq3FbHSPyrz1CwSe2ngd/CihbJ43X3oLzNRyKPu
oP+KIeoNO9fJCOHPcVGKRv/mhQ8SjOAtrJw95tPITS9/N6Oy7wtm8Fw/ADgZpoNd
A2qP6dUzlWESqCGbjo/HpQMq3Gn+C6LroBRe9CZC3/XD3j2IA1esbrv6w2ONjaa9
mb4f/Ax0uYCwmf1WHog5n2Z3umXrdv37IHv1TMpuKwb9HxYamC2HFa1lfY85nj28
xmJdHaWA49dLIlKLRw3JF+YxjsM0UzhqDdVimA3LTDrdtvbMgfvT5M0GCR66oHGY
coOS4GN1rhHiVmvtwQzBr2iJa0hQDt6OLZ3s6Rlsn8xYZirMrseC8QsbkFhTYmF4
mwL24ynsXv4lrQGHEv4uJ8WOhaM3KfH+4chMNxZtwID7urLqzyao8PZMsCks94ek
ECUPTR/fahztXZo997m+mz10Tyf9NXAhnUOCf23uQqdGo8axzyP4k8/yOU0S0G2D
E2DonL4d7lvEngYthazuA1kfEkBgVirongVYOqp5MKObuUYeCLTsvNKh9EbkF/XJ
KqY56e913zaheH78nNFk8wbzG4qAl3urW5w1ntcEp0c0pmQ1gDnzPoiP92Q8r8Vc
Ks+EzQgc1TskFsE7ULTUmjUQIihthFtu4+wJYrQAthRF0b95rLYY+Uo6ZV+dSAh/
sb/VTaL88r4FKR+/6W1JqHKBWi8tHUnBNwkcyHPnXvvkgWwW0v8WmvRrzjLrLliD
xGpDgtL0VT3SfVUNpV+RaTlVuUf/5+i+zcSW1bUtzvchai4Fow2uHJ/WKwmRazBO
IF/315gHmgVnid0FgLG2t5H0wQVHL20Tt3dwVAIEON71tSQIq7K2I0DhEl6V0WDV
pWePyybbGJSfkITqVQJZMFgl1aFEpskdBuiRDl3ZOruK9uSlI3nL2qkXceag+dFc
rZXii0FVTDIP/YX1YDZPQ/N9tCas+vouK8fWa5KNEnxhaOh3mLmbBYu6aRVc6M5n
ZZs6/cmQfAYFpiqw9rBRcI6q+dv2VOtd/i98ixpiNienYORYOzi7TEvyJk5jSgyV
/LRkm3Zgsh77JotFKm8y2Xwf+B6R5zgfDdAfS8cHRhrZO5jdNH1MBVSJ93VnAX7L
KYaimjKW2y/w4PMl14B+5UjOIa+yVyvaCBFACPSVrayZ/cEbwRTpAVaJ7ZSJU3lJ
iBgjuDtkY92uPVTJc4C2sHr492U/B9+FbRxDVye8/QIZfOTrgi8n1xGGRUa7ajeX
eTnPB/PCpHBP33OIzszeJ06vnKEeNOVoxS0uZ2d3qWU3d9JNuq7AcPUP/GBEBlAG
iNJXJEMfSgNqD4oCv4RLNVTlu9NxLJyYYJ/Kigr9R4t+s711rR3wb63iyHFMWn/S
4X3f8C3gd3gjbkm1kLPoOt9JPdOAbpDU2pv9lshrXuLcM85swaGiRV7VY0Q6E2oO
QDhPvQHpNx0Xe8kj14LjMnRff5pObyqaOQp9ViCAUI3kp2xpEPRO93ahXo6U6D0T
/kUv07dLr9Z+0y9HzlP6mIwRJ3ND+qPussKKPVP1/Nt7P8YPOVHE7Ww+98qwTiCC
TTT7JHhxRDZyf0cl5BsARfKj458FiJWeyvP6yS8Cjg4A4r3abyF9cXMK9sjP+8L0
jgmSb4jHQLKWVtn2bFRvXwP/6YPtnpi4AIb/7KeKyKDvEULt2oAGUAf+N9ysejdR
FfhTl0IZGuUWS+US8/84OQu8zxeZx6zIX/GdMp+LHcXgf2E7wt/8AUBpoardbLe4
P4EokZAE/UZcg+DjuXnm9mTnMuUwGfDHnN9QfyBgUJAI0ADb+SAngTwDjRnnuHQp
v25FS8SZQP7SmrKLwobTyDOHubZjs40xMLndA3RuKKicxQeC+66+FohPeUIMQhnU
ME7x2qTo3qDPdElvvqa8YPJ1FenYaiQuYzMYU9smGaCKToJBgo2vJP7+m2iAPZxZ
g4yTzgFBG3x46N69WSqUN+bEwIFCokl1ezh/VMnXY4wWV0TeWDnDwH8NaITEcGCY
GPMfW9B79w8ip4IX/F3wgHguuZ80qqopqsY5fdLBflp4JJ1MoaYeiROwjq/jb+9u
67LES6Vile17oB03shuikMARBeGnzLRswnbbc//eYnOeXXjEhhiZ12oCdfn/860d
jQwEQUgx/x0xJbdUstSCK28WeVJykE25N6l6Co98hDYnS5MQ8wLW0VzFYKhfRz+2
RLymRjXOKqYYMRaldx8bxJtoEWKqwammwdwUy7DDe8k9X7MlkAt1qHOQdCG7RZGM
TQte5CKEWQRgMQS1TMgzaGufyXEIBGh6W6Pq6aqG/zAtmpnh4H6hTfiV2muxNQai
M5clfUPVZwKv/uwOKToezBy0OqWBPJSAsv5qkFlG/EPnn19Z7jlx/QUxtgZfC9jb
TROJILpNFITYqThTiqjVyXHyro7mW0ma7u5B5wnSFGFiHOeF746n/kts46wtlksR
x00Vav+tkrgrmDKheLKrcVAjVwLO9MCtrpPqT8QOkHdoOjrZ2+xSJyHn8LreOrM2
xxHagFA8Rum3M+UMTdLelZWbHsV9ibfw+i/Gv9u2iW2kzqt4G/6Ae6mMsxZnrJcX
O7/rhPgdSJk6VzytzmKJ28zJs0THZ2W5Vjb7l/8Orp/w86glraCzFRwgNQ8jH/od
GSH6okHK7KqWByc++YDoQtmkV0ED3gBtQIYN9X2pYtvtgW8rKUtQIqUkOmr5bMUf
cbRyRer0wcxCqn/8oFlDF9Ho6SgtxIi0UBToYy5e1p4VjlNj6lo7+l/bNm4yFp0v
1v04tly4YFaF0tnGiW2M1JZcnYTzsv6P7T7YXNVYw4EtSzlurHX8mO8PIM2La5rA
8LaZDf2ECpYRE+50YIVCM3y+lfk7Jo+RukfCZzHbU1JMcnxR2ZkUWAuav5/n6r3v
y9gLOVmBqCUW/aZF440dSm6XwkigY5sTWYHWtu5ELK7CjyhJQyXBkAiVVkOGq+F4
1v7yAlrq5mZhZyL49+EIMUbtcFexS3OTu1ZSzjPz8m/ykdUdix7Lu5glC6m/thW7
exiXtj07viFg/YR/yu32Gkarl0eYNTHVB64AFosEqHkp/H/l1BHqNZStPcSezU46
SXNHOLu6yHuFNIaPBrewSaqTMe93NnhE1DYPR3eWvwObnDYGCGBZoM5pXcKDMUs+
lvRDMDgFdss5ZalPNrIbUgeHSo09+4SMj/xxwD4mqKgGGIlaWztMATp5IK7v+Lmt
90EybYjvOiD+CYFXyp3PYZCF1AJQNCPGs88MvbuLNIMlI7HOOeawhhF71rY7GH4n
jyaYeP94Syy6TttXkgsVBIg8pyUjNkYpZ+efLQHPEzIQAqrJQxZCp3sBivLkbUvr
KUasc7t0Z3MILHmp6ZJfBlGmyofq37zmTc0VylmC72LAzQ5YTmZHzI7lXOGjxS9K
0ngw2i5Jj9v5KFhZF6Ds9XosB2LUNyzs9/0jSVyz1WT+h8Y54bK1mJUJMTGRKWZf
ns/28NXKHnGoHmyTRT16fdTYte4VUcnITscXVb2Id9T1Jp1lZx152otbgf5/HXfU
YfGnQcBoa0eHrXzRz7vOHPph3kmc+FYovi8Ea7T25bqBvKLgH9wGRrqgpKU3N5ob
9eP1DWbWr7wHSWD3g3ng5yVJ7XGJROHqtWeS3goYlFMr4KIF+UXFLY0J9kQk/dIZ
jPuupsq0JDM2RTuNnpT77aqYyk08hw9EEknX2u9deFK3tF6hUbn8v0UtfBHiE4dD
d+MN4GNgwDEC0Bh7wpIIQ6WmCgga/y8VIhjW/fiIlTzl3foYiKp5+/Oi4bXpAsvM
mU74UWdMgMiFAuvdVFN/IKhh9F9nlnoP9l4idhzwchi8dh1lupDg2/MragIvcVRq
0WktSBW7nF6KNQAcA/kjmapA1PQBwkLmatQyydL1jjoFygurE0TS1CSuGy/X4Gx/
RkdvHoeCqiA/oJ5tIabofDRKmO4YxWf4vWXUxhpbTkFR/aSok6ylthGlepINW4/H
NHWXjr++QmzQx9G0VdGjUDttlASIiDsLfDif0ZPsnBfUg6DlEre8e6/539xvM56e
wr/WIfAY0tWfe261aQzHfBZ74sQsbkofApeLC6jWnSzGGqw60Gn+nYuXrA1jVhVH
nY5F8APja3Rz2MuP94biHQGuaJwWgm3j+4vk24Jm+uzPJavFqf5aU6DAgeCj4kqU
+fyRUmct8ZjvRwWeT98dYUhQPK2OrZXOoTgOmOCjR/YH60oZV7PGGRE9SR1uu6A8
LWjk7yyArdZkrFUa1+THrNf56cfyYsCMvBJbpS0wI+DfuUlJq4tARRAZ+jkeWF6K
WTROBc6qXwrga7Km+baJoFjc4szpazbz8j6+ky9k5U0UrqhuAw27G+hzvKIWHQyu
s8HqTawdLLyZNQispwybFg9y81Axt8AKiQVmwtDjqcF+siprb2AWhvMrStv6WP1+
W2xwSbETnUXdR9F81HwrcViC3MGtntvutEk8seJfMQbnOBtivpbaSnwfw5LTevxW
240fcFItbvsJK77mosPa0lFZU7bEqZqEN0R7aTpjR9NMoSs/t+FXy374hYMspRRG
PIt/w2Cia4v+vzfcxsjr0p+rmcKFULFYQFVAwmBE2QmClag8OhNfHv1mVoeaYZ46
owhugo/GQ/FJBvmmx1Uf653s1cYkfr3JK5SQoMdeo7JhFdAmTwTY+4RWcrUKoBQM
ZzK1nAREt3VenPkfiv27mDm8ApKd2amR30GDDwVE7tdh+Upzfj50Fg5QNlz/lrcG
T71l7yvzvwTktTXxIu1p/3bKZ3cjGUQlP+4Wss29jnkAYunCjB16FvSEfi+0rPU4
6NCYwVh13PCcMWSooYpanG9HgqiQI/Ye5PpwL57ac9/TLWUAWT5T9iNQ1/LRNeIl
xbMl6MC1R6K1w51kYEtZVVzoFU1qRTy9Eafi5ls5nrE6N4No/mThQP6DgO96DWJi
TxPDSCNhEw3ZITfGRb2VxqxzIgjpQsJ/ekztYJyK0DD9LP2IO92dyynbEGZn7O3f
rEzpt6MGtTcyqCm1gN+PbevUJ4FaAElw0peaK8OIryLmkKYkpVNExcAb+ydaABhg
xjYONCf93iCEFDj04Y3DUbF4mYI0cXDwPdPUCqMvwkM+MwlpNPbsfxQrmO43+Ms0
4d0JxuMjUUex5FvY8bsEliKUIgtFftQJxDCHrlXTXumDOmPdif3b9Vn15AD6jfU3
YKJXDWcNzY74nll9/PVTWDeHkA4mt5Y8grO2t5wvITiUr+cfKmDeQcZulrhaBuiX
Gv+oTCVRIrPIawgfiELuZtk+NTY2KgvQZBfuNfQIdFsRd5Cgxop/eFBThnwwKvNc
GFT7fy+bHybFdAK5CmRK4gOd7NLULaOD9AaHK66fjXhBfvjK4PB8BiYwy9Fi2A/R
upvhF4QVI7vEawTd4/XRt2gAR2eLmL6BdpBSOLZnx7m02I/DTftq7w/nNUGcBoGU
BRbkGjuxZ7gvxRW5jjIYn9k4mX+pLee1sra/APQ+w+JNkEvLcggmJ0XzYX8454Fi
3uD8FwM0gJLIk3v01/IaN6PePs/R375d2XY/7K+9b2gnYLrPkkjrELGf/1gKV9rt
zDsZHW9EHc7+yeE9w4E54DuDjHemUWL2CCc0AmQdwsM4Be/Ipd7kCUgAo2PFJXUe
rtUyasjeEcsP9x1aJBfXXOGFKawTbLO0f/+C4gBZyrSdZLyvJRpl3lnOkFeL9fxT
LKixPePJ1vZwR3T9FmIFGg7Q7qB1IaYzgb96cEV4ugMvRYCc62aGLBzJy79q185a
S96dFM0lTV483i0rSLkbZlRcM2i2+rnsuNeGuzL2U1ZWOBOP/iLvpBne412oqTjX
M/IYzscFq0E/jsMs8dr9UhlCpKDuXsmbHOuiVLhFX8nAZqt/g1/Fjjuc5+97OSTf
A2RYAwbxoqijj7er+xVqX0jjmkewx5r3xhL8uCP63ZIgkNxLZD3E/lZdsXuR6qBP
jvgKwD3uC7eodr0js5feIwm+YmMLn8bcTHtsMuKCQFtezPPQwqRUDHJ4K0oZYMgM
iWpj+Ik7dFJ/IXDsK1my/XkDtylFI4qfl7Ew7ecOafikmHkilKKoPrJCgBbQ4Pco
MKc9ryNY02+cS7n0DSpvmE8GATMVNHIgFe0GSeyDnXgbwUd9EM6ZldNu2B5RzWvV
4I2oM44aeiwCDOtVAZv2m1Zres5ENPM4wz6eDFbReQWwpSyyw9AeEpPbkIsHdgrN
q+S6dM1oX1Y0gG5BL3KQ1D1C3ddqIb3aCnpy2CR92y7qsc6Qc8MwI1jCq8TA98Sx
D+G6RgNkO8PChVZs2833UNClHw9AjGLmNFvaCHG6XhbgBHpHG3pMRBT84Qpd5K5g
+gDQidyDdirtsDVMC/j++48NTwCavfAYWlwhJW65/9nWtq/tKwS5xSJv/3POnbJY
4nk+CNHZGBJ8OwuXEY1AISqCc7hWaffJttPSsxsz0wy/fH8+XMCVB/VU/zb++c6z
IbPlD2AHmU2s/9tADfU0h3NMZiCwfnKf+HC4qtaoYhIMCXPbszNWofCgsu6rL6WM
kmVyOuf3nzam8GjV3s8TUmA7zuSSUa52elEKI2jI1Hgo0f5D74YUhaNbJ0xnbcUA
R19Dv3srUpx8OHqek981pBJhJQSYWWEvIP/FkBNiHSREyLemW562PPtf31k6IYQ7
33Mafp6Wxn0RjRNE3V8ItmFJTv/qNYP2KINk9u6ZrOrTXXVwYp6bzFtOpE4geXVU
xMDKQyjGf9fg/pqWYrBTd45sft+ctz25zwCHM1LHxqWZsVDJHb9+2a+Bf/tQSPla
puh7K2jRjus8ahv8Rz3R2E6CiUeZWvhtATzfnPok/ZMoIkmhpKRIc+/NIzFISqrV
zZ5H8pmy00Pr9DDu6QVdqHaOUNiTj78AIbpkr12njAMWJ5H/3uxhhXcIA4EtCeKS
vK9+O9Wf4g9tJ/3p0Ebqn0nxXbwt/gyHYCNB2DZ2ZDj6n7sr1vDrHlFJNbsl90RM
6xi9GA9i8GnpT5+w+4Uy463UWDyviDbyJaemq6plaT4i4mOXZi3dF8MmN1tVEd6n
KLATZgcBcUu4bfcrXVSCzhKpuyjF4hMWKlLdHZ0fC9WG5bHNOULSmk/Zq0KeAd5H
IEsgjGjL3GyQZAVqDbbmb9dHFHQrhyd/QIfQkaG8EWyH25Te6f+84jrtznp1H2e1
WgYn7YmLFdXnrgs3GCDf/jEW9nHJuU5WDorrzekKfCr9eSfvlW8gboDBouLClJpW
ksAR5Pgwi7nNDO4WXT4suMk2y4OTGoGQhihIFQYd9HC7vGRx03g/gL3+w1fTDfYP
9AvJbyEfQYbeOCnLC5bARxeEiF3LHXAHll2mXf8YOPXaZUlf2U9fs/Tn9jRFSKgw
E2qNGOZzCs3h91G6WvYV3J0UAAQYoEarxYgQ332SHsntc0+qd8X4FnAp+oDmoPVn
gvsYDqpu2CPghoNpxIDA45bDFZJbVrycNMDyDqMmY6xoK84Pnf8Qc5FiYyG9cVbc
O52voJ0u9Nzcig9obIPCwNiNkWIcfumquhIAzm1G+GzP4Y/FolrjiTtD+PNydPEZ
1rr2vmJZTHCrayheW8fQGyexDCySmQ6kwwAuXZgb8Q32kgnrxWeifmyPvJRK/9iI
ngBLKz63RwoLovqSJN8QyHWjAU+vl92wC0LXC1YCUGr0qBpdTLIRmNPNNYn8VrT0
YXlc+qu+U7HLiNpozYoUZzCzWREEVCZpz68M6GBvlT9vDdBkznVDkKvPnikBXh7U
DcHT3sNPHC3D9v69MK71zdgrhLuVi43H9FsmvrWjTsm8eMZHPviwzMqPqqWBWR70
A55E9TLiZ5WHi7hZVuBZf0dyky4MCLO6JuQa1LPF+SJSmyNG7in+TpVF9fGQcMvR
OhteQv3iC3PQmjqbc895oZLwDhtlXOMHcplzxdRZUBiAyopyLC7z3cAuqMnBU3YM
jaK8Kjn9GOXTrPmvHIe1KS6MBfcSSZvUzH92bC6Kji97LP+dOoED+WbnYvXnJxbz
HbVqepAhV9amfXCQdRNegBsWCBzX0TFpryNr5VNKKKR+W3uTF4loyd8IE10DLBdm
JMh9LKN+A5hw5Xgz1/+CWxnYub+pYhjhiIwNYATeEM3reepZeNYTql3X7/NgZX8f
mQxljbDqkXJRNVSwBwcP4/HbpJdth4Ps9MuEQO+jZ/fIdWqoSakeqvJbnoG/qG9e
CNH3LaF/RAtz12YoLtf2YaTyAUQDu2Qr3Wrx4G3Xhz/mcnU1N+HVGm0h7qbvsc7O
p9LU5GSCYwBHHQJBu50GfZHLlj1W1UvPUjImknA7ucleTLgoXZBqSCg9aYLykG/h
0d7tkw3j3mTSQBHXdywiR6xqZOz7h9xVxAMiiUC3n6dfDLy39Qe49HLG42OraHbV
fBd0puiHZN/hK/381pd7zpqEiiJ/FAZuP5KY2Q7xBLe4Fqq5BVcr5UhhDTEOTGII
A+F/vjKUWcdWi7MZPdzxuNHoSLp/7bAnuxxn4PRBvinNr9wwcY8mb+/GvL68GA3m
uKNyLLlSF85OShH38UEneS2jIsJJVMc8NJmCviU9d2ZLW/ivS7osAX82gLfE9Tm1
T+cw/S+A/df2fBM0mo8d3fIVJ2h/MC3B8Yp7BsRE7PIEEIBafiDWEjmlEQkeejow
xLwtZbQIq9SKLkxf6CrI/PXnNviVNDWG3MQDv7ABkuheu2YL8g0vkn9XJ+/2ycUd
FUCTw32je3UuMrCqrugnTfszFAEooi3tx+h51oRPVg1Bq8paC71QkRpaAqg7osvt
tNsB7qfGzxSk2rtkFeht5gWkUEODjPqqBF622SJkwSPmLLYJ2+eQmBBBoixB/mrd
PKFifKMOUBBpltKURTMt5l+jziPYXwK0PmF58FsCq4Wc9gmJiQCLVaJI2ThJUieR
fryZMWQtVEIfBmNeog781ljh0XooqruaCIRbHQGlMOxS4k4FC9vW/h/3+kyh883m
7cHB4KkZXfjlabewdX8qev/LROt8XX44csQIiAtLtkHQkef80YZtGMqQh7gV9trR
W0wLRuInj+Sn4AoeS8gnMWP/DIDQp+7SYeXNZsov36lVksbimn+vofu8ajW1Z7Y1
xy5OVuZ5+UvQM6X22nb4kub/RKUEMCApfwGwPU4A4nNkwJTYonXOtZr7WYKGjaD5
bUvtp3Z1PT+vRrrR8F4kzMr1Jh2C13z11y3kOUYzGSaN1Lcqh183tu64Un9d7BpS
NoVp5u+PKpYJDadR8eQLESHtAP60icyxzxWc/5k7hWiwrO6g5ip49LSUh+nJ+HBH
Fu8u7SpIHuvGQAVWCkHeOLWkcsXFnwrxSKBUq7c5DmmzjO6LIaP6xX7PQ0y4/Sgp
kT6utSZIZTz7OUiVpBIq9Th7UloIAdW97lqDDv4VB9HnfkwwDYH/yqVNsfuLww7e
d3+HpdtAVJBWhICxpNynEslYXVgPUaL5QWEIwE0+zKVaPTTuRGeftN/od8f5Ia/J
K0wwP3EfRksO94SvDSoa8eIpZqKo8Tfxgs4pkayFwwqyNVC0p0ibalUD5s7GY2Ui
vM/awgbHqMMVmijUdYrWbjVKaEU9vJRtPC16Y/ig7uaW0MGk/qIZqnL5BlSeX9ek
6ogN4misqlmc/94+jxoroWhMhvLhciFDQ6XAqXgBqo1Wlh4W2awQYziyy8gSMqE8
XMI49Wc/6ZQ421Jhj6wtqVx9wiozth/lYWhBz3IRybkrIdl9B559SH08bEDFmmkq
TguKQRrboJs7oj/iA2p3rcgX4C4UhTBhLBITHHR2jA3Qd9VggjEcoP7cjA1Y/gzr
XTx+OIFHvqiD5kaHekR1RCPU/Wp2PgtK3lenovFiRq7shpJyT5n5rR8XyM3RSsL9
5WjPyhDnuVWqgMYEzrzUD5lzJlyVANmk7eMR/UTBbQNslYnBAgB+o0e7dlhSqoM5
XD9KX1CCpQs93B/Qvysq+idlqyYwJgCN+eKW80O0bMdD/l/Rhls8/+KCxMoniI2G
iP0C368XGEJw+wEhZOi4URTKvYmhADd1JXf7OF8ozztDgXRlGktYMDYKs3UerYdJ
uE+219LEuYx5C1aV8G3Rya6s9SMA5CvN0Mew0Aoj5XaO+chNLuz87e4I8vz2WNgl
tFLwFaPTEXpAkWsfTHwn5oY2ktD1PprkVxyZNEJzQ9HXkVwS5jlakX8eLRK5cgK5
D1LM8IHrSJJPuSUCxYDCoIahjQCQidGg9YkVHyXWrWeVMo2+JgGvPbs9f46vIZHv
KO4YE1AvkFeaFPintRXXZPzeHcnB5X59KU6lu3R0Y0fKiBiwrl+tbcyfkQxnFaHS
uSXdUAqj85nMt8gVW9Mw6CDDMbuxqt5Cx0ohWsXypfk7zYR5DcUVbJJGEav2BHcu
jAe/XnpzN0BtJgT56oR1TchJom42xdMRL24pO3ejzHdd/3UXc/cRk60DLW9IECch
JLYVcLrSXkbuLgfFlmqCwxslx5XiF5oGsp8nLagG2S8K5l3RR0FOjHBBgfWBG9hP
lMb5HpCElrpKdDhNzm4PaCQT/D+fLv8WN+nqDSwPrasKBXqIkF02nqGdWy0PQaCr
dZi+liiYWHQ8OeKXgqy0S1BTvsKX62eq6pJ/5AjTRB1MFyQGMhZPxbyJyHDGCYkq
k6+azNtiK7dfrJwEgWiAO9llskG4H4ATD2N+DAkMNEL7n7oLgxrygj1nNuikC4u0
wpfaIJihrEnRoS2c0WDK7xGmvZhHoBfsesDJD5gB79k3Y5IDi4piQI5t6qwKmYNf
ZkwwPl2g/bqEoz6NvKVbOfp0bNqNyMNwtA/ccVVnLwHen4PXaZhXfNwgkTc9DAdD
d57ibzaCfcFO8Xn0gUN9yrkZmruy0ETXpTcbgyNqjdE7jm/71OzO8i3TAoEJ6S3w
IU33TwRnw/iA0BzLkFr6qZeos//fZkDv96FW3wGvTJikG+6DLl4RTOo2e9/WDTMa
rtxT1dJ3alzKmC+CeHzjHt3Nb8wTAL42pXV0jlkwwpeKG+7ldOAVDYzwvIPeRcY+
aPkOC7fVg8Y0S/mzqX4DBEPEOKSVgNIeX1AzLu6AnMW71Dx6voWMuD3+5Flh6f+d
+crkGWz/u+k4nQc9uzqnOJa1ml0L0Y4Aqmxo2APxl/+XflEO0jV8Bmj4dRccp/3m
WD4mOwi8q9z4nfxt3RkmCoJqtiGoIUWnk5wZWWJYx7Exn5yzbexIdFJCb0nnXdu1
bQhu9LNwGy1WII8Vtkl7H6sGX9s3+HJYaaq8yi+RPXYjhMnKfLjBxYNlHT638Awx
+95qqN+VfEp9TaxNXrRDT9oR8Ef6kACTxdoFzbGqW/yWXI9dyTQMviaSuctxAd+B
JLhYzFEwiYCGnW9pFUxkEeI7T6kkpPMypE3VuG4SWqjQJ4x6v85aY+GVH6d3m85X
h+CrPA6w5SnVSRHstaYIjJHf9wi40r8DK76ItYQdVvSV+XmwLsiDi0nTiyt9AESJ
w1RwvhFYCFWzQ9Qaf1kM9oMzP8mHI1jVfw302Rzd1MePfXsSVTbymzd4jegPvWFm
Ut+LuHhQo9CnZXO5sN76sKqrJ+iD28/6LDa29kY6lDHkDNQWlf1UuhWYk0gxSxCD
WbcGwYVw0VkgDNxOPL8ZIswZM+bjXy1IHIioaOmBu7vhWJwMxYGqTXbMXp2PI+C9
psarPmIAjKy71EXHCVRfULR/3kaW6dN3zLFbmFCEu/ItwvuaF4bkS3iPYCknrxiO
ockdTWrTcmq6mYaCIhceO2wNIeNJsO6JAMqmLlqnfK6ktwDQm8U5GW3zvo3ENHt8
D3Uifmmzeo7CJ+d3g6WagxmXE50cJJqORTz1L9v2l+JPaAd/ADyCOW5KWfzOCwoi
vVcR8qUcNATmuxxhJLh1NF5qaY2xLlK6pE/wethgMyPYkTK1FNM5EaZM86D3/PnY
6e5Oy8tAxEnG8OzZP0LgLsT/tqfzbdztg0JpgJISPlCZu73hoVgEODAAP8TUvIAs
hey2Jz2CSlJMARekGXwHHDWyrUvGyEf2cFFDSs4FcM3KZV1YLLNL4V7zYubdrG5a
WzwshqAuBzYW3hXApsuWU9k6cYMYH/X4Mn+Dz+NmM8ZhVKdSIPA4Iwa+tARDtI6v
8JWV2j8446Z7i5IU7aRgzJJ/jJunH2ojkeS9p7r2gezZTJDXTnHvFjgVP5Tcjjxx
DAtssfVRFlVCAOmL17FaPTcO76g2/tBpnVFJY7cUaDehYRYQEv/3Pfe5FuMee/9/
qD6kxbdCIFfEU5FtToLHX5QR90lwBTy4mEI4Hj2qyPvvU8mmdpEaPBwGU6Y1PeOS
sAlQ+Or7/2+F1LZX/DiZg4Woylfg2+1mM5owapALo94xKEKxl2oJUTlaf0Rwih7T
Npv5SY3rnNMsR4lJb1xaofUSgiIQKjAJcm2VezaIIbtXN/6sQWuZ3yN9VrgbZjxd
it0sgi4+gzX2gzxNqAOIi/r4QpvdCvFiU7bjfKMwGXZkYsht9Etcf0+0wlAiNfA3
j3fQIHzNWKyPylOcBnPM7eDYP5eUVss6JTtghohvC6mYFwGdfgKcKxlDxXSk14ms
M5E6nBToGoIRrR96gMi7eZZIWS4QnW+bwfUv5uN3v3jdjaao31Zziw7ykAbA32tJ
vDqZUA/B+d4OOADcOwTV8+5rHS/EfM0YndPPwxP1z12Vfv77Ts4glJGSqQj24ayT
47plVBxbSd0V+mZ6K7WZJWP4W/WR5UJHU8/mwwNjxrhjsMUcYbE0ai9JrTMvZ3lY
PEQEMcPBkOhK7LUzwUiM93yMwQ+GdqC3uUpUA+rFkkMRvgFDSRQjRuKtMZsLpVgA
4GLHm0252JSgduqK/KxbNDJcVNxHJvT4z52781fM1+toqXwk1alzDcQWf8OxaOg6
DN875Eh/vVXZEmRsChkJa5SyzHxNO+I83/a00fwQveFCeY+LpqdIybGv4tW3Ic3y
88Xekw8RwH9AUvHzf3Y/QdnflkSOPCxGidZDxwa57dNz6TNh3e2+xQqZDREPt4vZ
iFXDjmKBHacBfDtxDztEqfd4RCNbNUN8TzVunKPsBP0u+iXHZHvZUYlKkP3AJQUZ
5nnH6/g+8gkEu6RUZBGs5LnQex1I3On0D2aL64zBTE5QYN9tDZXo23dgKKE/sgxK
3/a1sqYNj3JiSpY1/AIZF9tSLmUTNKOZDjnC3yXHL0Sk1rYYNVNyBKQ0BN7e3nnv
ulaZWRP8z4ruDGNzPoNkqYg/0arInbn+4VbWXDXBQvBo6jr7cWcD89f1V/i+c9pe
KsGkJjmPpKRIntXUOAvIBhQr976SAxTSY4dptE5axNRTZyMeteD+NJY8y4uDmFS2
6P/hLJU6UkJVgeCsg+p4qHvQrICt5uMiytBUNpZwy5sIUVHxSUGnTGIZyobpRnKd
wU3ivg/EpvvixVOBgZuuqWSCYxo8loMr3t5bAXzJXcZ2gacWBategeqrRVxry7FF
BBRPrc0ybegyl401KjHh8ErPjtO9o83QCWyIc1PbfAC5l0qPgru7GWA+15YeEW3E
bZHsUhW8r5CpE06y3YChKZ4B3Z0Jslryt15V3c9a15OfsO/GY53gswuvAb2wNOA6
ARV8TCmkbc9VkdhfeKVdYibNvKJzofucqkrT5O40lFKdyvSu0b+Ja1LLH5UYNAZ1
G+8JdoFSwIl6YZv5dbL5Ic4IpXZWp7g1lBrOseQVORrj1PqzOvc1KZzv8GpgwN52
umUYrqCjN/2+JTuz4Q3PkGK0YL9C0fZf4S2M05ldrv6+FICb0Hg8LmH49dxog0yV
deIHvvsIWFO2IISJrEo5GbJLZ8jWaxObKuHtZgv10ew0NVKFp6+QwJL9MhlGl+yK
0UdM5X6S8c/+3SrgJuECF5pOaG5yU5R4hTzOaZQJWkb1VV1ujSPmPq/yYdEwQNAu
gjUBzPmSgcm4QH9KoByxivaZwdLcPWQeh4XdesiLDQQyjvUS2iUi6OorKlEwxlAd
U4pkGn/NJtNFdKaBEOu/5E5Jgcv3W5+ZDI9xIB2Vh/0qUau+2n3rmJH2MwO07tCT
a3r4Toi4yuTqfzsJxh8y3ZPrzVBthJMhtidHPn+ASBT4P9O3xoIdniYipW8xSO4v
WO4RYcvf0MjcgZcAbuSJo/SWcNaxA5Usy8toBULpGP3B/DK5Ijw0Qz12oew+4Tms
VlT3GDKTN1J3CUQLlrQOFQzhKRBvMjXXVuv8ny0RLKeFpBdF+kenaD1KcvwPSpEq
qIXXwSIjpoeM7j4GkGfII7YomKRt8oyeNnj+Q2GzhTv04cXcfJaRUfvEUzeTep3c
WMiRFg9xq3mogxlmmvlWoygEXxaUoxqC+/HOdbkZYzEneZvtKdzgS0CM/syypdkI
/BLV1pjv5xDZ23Lx98DnedXoXZDgxgGjMvxs2OD6YWdUSHoPtNmjCvM3RrKBMjLe
rb3n/g8exyJRlgiLiIvzRWk9hs0AhZWYN8IjPxEYsn2N9WVcMLaNEn2Kabwq5Zc3
KOPjLROTRR/nR6V+8Vk6lZafTiqKRptVHCRVzENUSrBHNfRtBLgq9oMuAmbz0u79
UOObx4U3jtzRQmt+MHyOwUVyQlVgSiqdeQlwDNuv/fDCuOiIbBACXk1j6ex8LkzO
Z7z201w0/7NzjhAO8EKXXzfVIHgzvBH67+L1dibnSYZtpuQV9sdFIIHqeEbUsVIQ
xtcSY83IODyGfIyOKWHRHryKontxd36LYKulMp88oRzZyPIFDy/QIYaEtFc7FhKP
0FNq8KXvO7gbfxK5arTPgISfXsHhwjo7h18Q/GdXsWSuv2NM+fmQjajreuATl/6A
5mzOGCG04v70qeTfQsw77d9jAZIDzFEmRocW0V+Ri/JjpAXIPR2A0EowaN/CXyNO
HBhHZvlB4/taPz3e6QjMEa+is2gDrMlxTAgv5OD1zjapFWwcpIk0iHvOFcvt46m4
/1E0Ceqgbbi/lm7TV4KKsJ9CLKIzN7whjNZJwC3/Z2++PazcS3j3lRoelHTG7yR5
+VR7d7DnbX3UUaN+Iowdd/gSGvsACO5udRbw5LZYquOD//qtbfvvW9+WJwaAOmQa
Vih+TC17m5XFl/ZG3hUdkRKBwyF6CNqwsgeIbQ+EwY5746GgcT8lx7X4nK4MUx7A
bB+9ukohoPBgj4yEKlGZKIlrxHUYbuZ/6u35HXfrQuB9WFHaY50B7y/wBLRRt6Rz
+UTQbBPYVvMjvwXl4BxoZghRPqQEmynzF2Y+MflXfxHtmn7WoU9t7XxDXoQVruBn
ZNBAv0Rki1nwZ11xLQabR02IRsVu14nKw5RgxkG6jyDmH6IQGNnInCqAJx3NqqnW
G0Pm7C3HMScdKXBbG4JYls+fs7PPHakPrNCFvkhHjKuwFXJ6hRa0BBjM+ntU2nWe
hjuvN3eCxTi6T+cbX+bhbz61OxDMERk5ZGTjXaf/X29OdF8J0HYeT0D473SgytHb
oSSc2YyTszToVrsIGXZCf6kJeRfszIIL1b7a0F29wZSKmfNnVzITZCaxr4QVL1+e
DXnMH/dXiLninT2RrlgE+zly+/MiIdR7DfFTZRQ1rfjBc+uzTwZbyvNzc5avx00j
eItFlovNbMqbFa1gUA46YQt4QfmzngkdHJFK+eW0WvRZydGUaqMkMDqvXBWLZEbJ
KqxBjkh/mvWKPnyd2q88Ljds/KkuuI2a4/NASqNrbGCIntt8FulBprMCoKqZdaVu
kvfVEZpBu4rAqIFQaeYgWSXQLoUiovrS2Opi24/y0f6ZFomDcXYYXbppIwUkQlNr
2+OMro66hh/6Fvm9PYVlquOzjIptrMG8BTkh10FiPomXN3GCiPM4jt6zDIS/rR3o
qJ23OoEMVIjhPV07aO9CPC5/+eeICzLp+PoFffwEm3/1ip4QHOP/bedeWta32vAZ
Wsp0ttYUJv/9QuZuZwpyocI1elQIUrQjy82KzV3cX1J/TBEhaNAb5RQTD/kR9N8L
XZyuQXh7Cg+iTN4/bYscNNcX0h8Bqq49SuiRCT0shcJRbx9PQO+mQm9fMQISPmaW
pjsoE1j/3Gix8JsWby80rsPUexGFXtAka8s2vqiOE+TYB2SgxRDbwTEhljJU6Uko
pnBmcrbLCz/EeeVOy+AOMlVvw0/fVWFrLYFzyx5Z42Znu6FHtXIUAtRPsXcPq+QV
cp6pcTrULrPXGFMhnX9S25s01+QuBRDIba/vOc2ZO4OLKZsQOC41mk5agzF/3ALY
tt9TD+H56PcE+3U/Ruc+/5x0WVgJZMa2iclljgaT2AkYbLn92x9ELgJl9v+1OEba
7b5PbuyqhqxZz7eJPcUltp95XepM1r8TMS84ekZoRlSVAtbAiMQfrM/iqYDDkwbh
hg0cYe8c14DHtVKzHsaF9CelrfJOu3dkZy1ECfLPZGFwKjaU/lKek9rnUzldkP2m
RtL0w9mGlyVkyZ2Ug8T3cZ1HrrxIvT99l9sLHovXJKUxQvRisxxt4NMtJ/yOZwvC
aDLzctWpWf05aOy+CLBEsbVVaIDnjpiSMmc9KjkwjWk0iMGRS/GQDbp2JsKT18V5
/4MEGpe2vIWVM6XBBRELJhf7t3V1NyU9F7xAZ5oCIHz6vbykOoEWBKEFG6bRQSLZ
1S/PzXCjqcx5dX62t46BeeNB9G1jf6b5N0zvrTslnmAdUxUy/EVsq7MCFZMFLw+k
34dZsED0ybSNKd922a3EUrIojyJEE4fw7K6h5ieUp0CgOIgqIoz7q6PVRGkVatAy
MKTAsaNfCKdJqmK57iebJ5uDvCDqsK7ttwGNMfGtgvulB4V5NJwdoJtRizWYqaa+
8kGLOma33EwHN+1vuA4EqIpx35GuLoLkMC/wGPV91QDYIEqiHFR3XPbfRtQRJKN6
k1h1FV8q0ONLbGisQXit1bkf7SgHs6o+53oZ/zxrEr+msPBN8XJ1dqWVlUqhP9Ok
4jFajcIoYLGe7etwN7pc0Nqq9nitHUV3R6BIcfW5SsK0+RgVMuCkdq3XuNYP+bec
JP8JGDv0VDw8FqMrika1nZO3R7Qr2Jv7XEUf2Kjug6bg1SQhlyjBkuOBOjNJPi4I
95QXALReXpOo75/vTsWUEpCuEtC0lqFs59ANqVYM6Bfw75UfMiTX0F7ltkCx7hbi
9E168HZFSsjRoU8R+mpqkEwQEAcbFUTuGQSOtALFYrCaP44KvEP5jzQE3xLHRpgr
6y2IGECYJ4XEgfaWV96gDGjCKRHTWABjeliGOgCQs81so4G+El9Xyp07LDL1fi+2
EoEhB3Z2nbm8Icrx9pMwq2wd8uEH+u1NKoTHqGMg+MhcC+R+4W8o14H0cxvGGC1W
U0mVHkIO7KWIcftet2iQzfwhBtJkIF3oO3sGEihqUQBrg1ucfuXzplBz6zvaw3Vb
N1Vnyqzd5cJ3WYYEUVi0o2OSI9h2K+eSMaUt6aMovyAWha4FCAU2E99zKVsJU1se
oO3q0DYmj3q7GtUnGGm4ODMSVaFaDtvRjn+p/R+fg8mVm//hGHXwIVeEmTHyMsw2
25ommNxN8p1R/0BC7oImXvJkjAK2QqUZzf2+j5qmGAaIkEGfpKKgiUdPt+qw8Xlt
1GF/U23QcRvaJdl/IrKJSOQIfqIn8NFljbvAsRtIQjw2BstXOZhDCYmwbbT2yp68
co1AjKWJEWEnlYogVtLLfwH2Mn4Qc1DbCH0/RzaBdKhz4345kopqjq3exKabe/bH
y4CxfWuCA6mldwGJd/Iugphiq94PGLayFB+OQcpureel1aE15s+9auRVOXR4f+gS
rhmN0w7JrmwjkW+zpy2KTM6ouUKRo0OwEtxG6bFbuT5nTEuE/Ql+ek+QGlRIi9DN
6XAnpxqMRRa8DPYDAqcR5MJWws5w+A5hoQI4np8xaq3dqk/9gHt/oLGQR1boMA1L
OSaDrZW7yAKSkAK068hsNmI56aiOMvMUd3s/2qjN5zqb3ITkT/PkMuW4/0n5VfoB
NLlU3eT8Y/k3r4bQqRpbTBzrbv/ma0VUnIZwQhDpQsVS7sKfxzyMT7ciVmAoW6qd
S/g/U+TtJX37+KgsrEYnzH57rOC2MMhltu6hbEO50zaiGRBz0/BfiDYNSO3EYtJk
1WpcAYOCzl6NcLeWXDUCUSGXfzv11+UEJ5wgxaXt9xSNy2WthdD0/L+U2WqY+L1Q
0DEeVN8pKmT74pbW6S6gemMOtlRqEWjYCyNRgXMM4gf3EhuvJQFpzefrAx5pJuLt
N29DHoFq4ANQZE8ey7qYuHP3REl2OJzXw5Dng9ao53XZpMzSy9t4SjGtxqNNYeEP
YgW7+o5ka54KxxVUgWKm4wSUsRHeLMPyToHwr8ddTU59payWvnBjrJIPZ5uB3mM2
MCD6b8GnxKjqhHFPLh5kmof2GCJWikQVip9YsKL+5pMRfw4cMcHXTkdbsNZpnUss
DDxE/XKgU20GhY3qdNOfr3pHUlNy30pyduqPTc+8jxNuku5DlEyloFzHBRmErwJY
K8TVtjiof8HQByozFhPwbVplrA8QKsLIekae/eI3YqlROSjdSxAzyvks3pGD8bN2
DCPxmlzmFEKalw7kuLA6g2uwNcbqoxjgQvPB/gIVcqMG0e3gKFeVW3n+uOpHZit+
I8FcP4PvEXmIijqoYRK825OWxVQD/PYjXI/Y83m8ImEZBCftHDJ2APR0L9zzn34H
e3rhEC6zRhKhIvOGsm3GuboJq3Yqo/2HZ83ocnY1kkLtCEyIC487xMQZSzVCI7Gn
abv2GLqb0hytyqou5dZ8RfBiRIj5Y8ktrTQ1aVHXQoOeiL9/osgm/7MNLNKhzubU
9zRYwwbefJrj0rzX8pp0JZMIpzDWHdWqnx74taKxjp1zOOd77+4bzuftxr+KtAXw
pa1BZvZmsZLjHsBiqhm53uba4fXFqdgSxgscwk8pbEHL2UryTluV4Fob2bFJ/Mr1
pDB8ocn0ryi4tC12c5jFsHyK68yuFJIcgu9Ycdsl/m9nPLrDhwmRUO7yW0P0tQE1
/QCnHy5tpDkRN6S5qCZ532pqiZm7EO5FGJvJWgDEeptMeAv66MApNYMrnCAJk+X8
bDTtE37YCXHyI+nD4qYr1KirN5ib2lEFdUuMXxo74/FjBNfJhcdn+j96mksZRjCs
A45hqwliDwYH60zLE5xVwjgGab8XG1jmoEf4aS2lQYz75qM2+neqxylRliEg0U/c
fwBd6qWdCPAKOuK7KYVi7kuhbSk0aotehWCnD3+sak6EXBXosDfn+CvTFQpbtqwv
jwdNko8n2SxzEuctgJdBe1n4N6yx9jzjCq7sfz0I6MncUzr/qxDnJn8BH1YbhkrJ
THhtEQEfFZe7LcmKxUg3kJuQrVtvfuwNjW128kZl+RUApx7B3CPtsyBm62v1UM0R
V6+yrTtvT4id72FILVvn32FgSWeD1dZpkaq9Qf9d8kcoCzSb5lPMU/jz08Ud8dkO
uA46xvqky+ShRc2KcntnTykBO3Ay/LTkYfxq57vCAwybDakSi5rOKD7DGTOHSynu
g/yqvuP1p8sw+/binaH+4bPLYBpG5lT1nsNMH2FRfwOrwZnwVyZN5KhQU/DLPVan
i27BNTs9Qzu3TY8h7uRd4fLrSM7UMKydVYwHippX59xUx/l1JtLP8SfJwxim1gbm
+a/IvGiqeuhSKXYPWPRJ+d6ZTeyJmm3IQy0H1URLhp5YCPFXY1vcfhB5ujWACreo
i2gSpuBHXhHUP2lAUZi0vpkR9tCEzR74gzn+Y950OG9DdCqq5QEDbgKmY1+4WTdy
VSaTYqgmUCnl6ym3pkoEj0f4V2CZhqYraDdmDLDAeiscx1YF4GFS9bzsBZoiZ2Hx
58HKrBBVGIHcOEeDhUPeG3LViKNG6DLJ3imyXOvDiiIhx+qqs/cjRNLLYUx4m6X2
zaKZgX1SBwZB+yLJp7bGz0WM/8id1NwiqLD/9RZanRR0bJtYsOen6zyJx5oNTfUN
6/GVmEKQ+ICDW2J7En8ab5++FE/7LeCp6JPP1Q6ZzKVikuOs4YgohRXTFTxLo1j5
ifb3eGeQdNEl/2EvhWBX3i/kdp018RrZRqcO8kB3H7iO2OwPhWKV5bS1OkE83FCI
xpIJxdWUIhv3SWW7MYdTIApHuQJxh49xq8eZwaQnNp8nn2FValOMBtGIknQjy92A
mguiAIP6Z3uYjco2avkmE4mXtq9dj+hMAAjjuPel+H23wSBxk7I2uoVV9NHx8Z/H
hh3PWm0xpHa+4ITmYbI6rBECIbKbtFmWxEq4cMTSHbv4SVfulpWjyQtSdjoKMnOZ
SnWwA0lYFqvAxa623eqX7OS40LOKQcelRUOmMJPJmuRPYkHSxBTZC7NH9yaDgjP0
LcgqCpt1v0j6JLu7GhjC5Bcl0Z9TLxL1qc+/IPTO+vDKo1GaQCgtpPHyw+xRSIle
Nvr+8M/8TilfLppFytFP+SWwfXD7jmhCID40hPYCP8dGl3U88N+Bfkxg+797fQVC
YhzTqAuxU/zJTC/WFAgAsKOrrHhQqkc7J9eqZOLuzLHfISCIum9iTUBtTgzLESu3
pwpCQ9awTYv2dtHIdi1+Wt71Lyt5rOy4PgskLW1u2FlXG4EcaBCyhKBVZhlJeNEI
ZBO7ff7ZFcaKRbPQihMNbMaWY6kqqeoWZXFBo4Y53qxxnEcHC0FXLxFOz5Z+E2l0
oeTzaPjbLq5KLeyLMTAOFAu+mAFmuHuArVgYWR54MDREj7LuU2FORM8R2UOm977C
1NB9CEH3k7YXYKlfitZIIEZ7L1gzfn3ZTwEqdxczxH+cec40i4RrehTjzqE8aEmt
Es6/6MqxtzBZmAkG3TWlBQ8IeWmQOOx21HvzbBC4EOXz5nrveeOQ9m82v/Hkk9Ou
Oo4irx5qdPnWCuSEdurTSIocQMO3/hgZ9Y2qddJgolsxK9ool4ub0VmNxyx8dgTN
Qr+PZawRGMIn9zMdD6gn3QGnaZED5XYW66mLhK9WIDXXaO2e0dM1OxmK5CvQ9CYO
JPmvGfgeuYj0u6phXzPRcKvoBshEctKDvp0VT0ymjvqUu84RrSHH/D1s4QBsZaV5
uX0mkXEOHmb0P0QE3iA43yKZc8MOdqErMUm8GwwqHCjivF0dAHWt1Px+p/kdAS0e
/l1S5cduIlIE7HEDBwguCYYvGG85RGFbYP0/zFvP5q4PAhtggFiNuCnaYHhxu6Ev
EIxp6xcTnNb610Lhr4Ea/fvre00oU4Yc4r+AdSEy2VPDQaoFngyViMtuBiT+j7Q7
96KzdAPn6EPixrSXodlYEvnznEgwuUMrX4RkewEYCfWIBaI2vSoo2ol9YxHrbdGy
BCoKFyOjUV+e7j3qaudRLy02ixxZjb1WNO3iIaceFyNPovX9fSHPGvihrmWBcIO5
cRnfFnu3ryumuc6zK4Ytgk7uAqkWqsf+RDSLLe9B3usT/DyPpMqujPHN9R2+79fo
S6R4X0nD0MtSNDO9g0Gbu1p/hAPPJlRGnTY0H0vtvYi/2NBE33oTArxpfU8vurBE
BVAS1P1fjc/0gJt8CbpxkPCXxPNUYQIYq7mnrp6GB0A6gisDZFepr+m/GtCkVp10
OzMOftXpB68d7mhv4It+DSwHp9/Q9/UZeyJkPj+Z2doDMN079v394Awn1QPe0slu
fh64OzGWAx0mo2P/DSdMLysjNjld43CtvVm84gFUa63twd5Ibm94uGykPUmz1sAY
uJYmoR/L/1hPV3+yyg+YPEYcDAgi2nzlHlFetZkcHuArim2/gNsRgfLeyg4SBPjD
8yAHdAQpKZhzQVg0WQptXAkRoqEpx8843/P8PxXJdX3iw3pmsL3yMGXOfBUn9c+R
7ys5lUlhWYZZW9suv9D6NlYCN147Yf/E8omJ6EUSj/JvRWijrUN9V+CKlqy0S62H
cYKdu8fRLO6ADMLCvfygDjcv70b2OfqH3puIu7EVIDJPlUR91avbsc2cNOI6W1/w
/4Anw854wjAnqQboslH3iaNmTtrK5xrUaJWyPtIu3bDdKUWOt1Wl73H/M0/LnD+I
zJMsLdDunzvIIFGTi/w9LQ1C9Fn3CM5p2gp9PMbHd8rgM2Stttrf/b7DcsVhAsV9
HpthzTQQM2XtMxgSkSgS4GdA1BRIvYwr9NLQ8iBtOyzgEgnYJGGZsRRp4EwPmEjJ
3WvykZnTZLNt1R+TCQ5qmNKAMF6MVcMR57063ZFCyQPtRni7ovQksJdxPsbdy4H4
oDA+I5KbnVy5EbMJ0swXuQBsHg0y9fhnqgDzXr/DZsRYS2x+VIoEbwhEFslqy7dr
EiJ1D9S4Uaj0R1coGWmkzonMLmEOCBQ4I5IXSkBC8lxKAmnD5N3r6RYT7p6Q5Kvf
M20DldXZsMBvqwifSJZ0IVZiSpEqEtBRsvF89Od2f3gaotAVN5fSg5ehVMdvab4i
lK7EN5Fc7WiY1zAozGLZveCsAQMhkJx55fKGQtZGdc+DOmZ07S6W3RDQQKTfXFFJ
IvF9P0JpQDKeP2pthijCDB9BA6ACOs4mGiYjDga2PuqE+K+5dVm4JJpckEK0zT4s
PUZkZuLQcoxTARi4wP4VLKNB6XCx9pkSgURkOmrrG6EtdwKZ99w/NtnS5Ifiw2jz
bj0g0bTnvQ66X6CuezcVMObtsRe5H61HYidqzqISq6JAIIHwkwyyqVJJTjc4Y7dI
nZN75YLYGrpzQGfrciv+z/+y3S/A8re47xBaU9dWbGG9KCAeC2sr/lR8dJtz1/Fq
n9ZNIp5gNPGWxH0gG1Eyq7aYYNzaEZm4TTFChLr2UWTaRZ0NRGf0nIq92OQn8Tal
Ynkb63ThLe7Ik8KyRymLxWrzl7ji/FZUoTXZq8h9E2OEgZTNJ4GVPk+gjGpdU/Dr
w3hjGux/QJ6hQjGOtTHw5vchgWz47T+qpUANnD9zkA4tzvsG+GAu4UqEbfC8E6MA
eVNj3BkglLPvqOdeOOh7stwUpWAkXbhLEG7nCSansupguOCpBFoGCm0YGHU/oRgc
mmLM0gxMAqXg1VXHHyLiCe7yCVoY5SgFyEzC3D/MIRmSHwU2G+5xpzUaoLSxNVPT
EZzWETCRCuOtEBcr0qt14ceIuGJGsJml4uEx6XFXmcxckpbiLqak81tz6JUyx8tt
yNFtcRgi3EHO9ScNvwxZUcIN6mgfvt15X4AgZO0YpfcjJzFo8AYrwFPMlHbBb3tA
VSGr0grGrQaUwg2DbEzVhDuc4VoHacrfLzf9rPpI0gmNTm9cE8tlpYJo4u79qRKj
eVMdWf/r6dnlsMgfLvZave8nebCitx9dEB5sUdPXdTT+z1wQXXS1spqx7+WTyjrG
HA4bFg/VfNdJq7ubXSCCbiYqDZknU3pf2/seRA0jkYCsgUlLD+NhEGmJrG5uu6jM
EOEIcNxHJqGDFs48SjmB3Bu11hdQjcgrsPhwireOFo8CoqOn8Tq9KeEtrmQtgJ2Q
J0ZkLaI9BjDRf9IcM3j12x7eu5l/UPF+t6z15RP8S7ctZCkgRh2m5cGRMvSMAh1X
tIkFhL581PTnpZbVcpuUU9+MYEkw2wRDqtq9Yjw4cl5TNisbuz0qTLo5t/mpCZMD
j+orOe2rOmw2D/dIuJNUQscU18MfDZARlKSGBUOYGVC/ynzqM4tiQaukkbj/6GFm
ScaTNg7X5PR5P1/sMzTLAVPQw+OCKWya9JADpPI53eEQKJxdECjIjJHN3rzKh60O
OJw3t5Fz2TY18uKwZLDACiOwhysiuw/bpyMWMiChERLxz238xSy6Jg9VO8Cx85h7
Cs7olsgm4O9wXBxrYv8JEuI8w1MCk3ilwkB6+vqm4hQxRN6V0LahH3cdMyFiu7uZ
V13waUKAXig8a24e3W/iOMjEploI8ifQYKeR8xNHokIYEJxZTq+FY9Zialsky7lG
BNCrMSqW6kHekSAZ/ja/Y1uOlvHIf+6YONn3OmAuGV4tXOU+BAmbMsRUVOQtpCv/
sF33emS6je6zrkPzPIAalGZLwoV41Plx0uUofyudfSPIcDz20LRBmM3iT/1Wn9f1
TFjMAT3x4oInFrWsvT4JzLQParDt3ZvuJbIELMePJ4BW6JV8SDptAg+i/J7yt9of
Q9zSNGYFDLXRkoQ4k4tCq5GO6/SHVB5abNnqdqNymDrKpL7V2IAgGXJJACSpjOun
sp5VTDoxrZ92wD7E5ZoKWZOPhY46CCcc4w3kaA6ts2lejBQaf3PuUb1szGWC1xul
KB0ksOMJbsLSHcbK+aUdlZnIrAMaLrA9kd5NAbQcXw/WzMBdBBpJW0JWtgB+xft+
9utvu55iCdyA5UE1dp6L+XZSood+COIWP+xTUFLYZm2+tVwzmWRsiAVSTzWoj8N4
Q5g224c/fe61kuJyY/Ciq6boqfEFewFRRkWjn1SvTs/pG/H63DG2ITBkFLqsCpPi
uBUapM4LvZLdEcKVQc5pbbMVKFPV2haCogQyr3eOwYzPjLQWJTpqDuqG41fUEj8m
6Ggv2JQRyE/tbaEfl7EwoesNLNNR83rSQc5iFBzESRHuttXvV08iDBlZYnKxD0pg
ustBGhUcSTgGRR9RiBLDI+stWaHm4asd4i2JK8WP8SwjpbUuZjvtgePIE41YUrI7
BESt87MWBtizYJBHm/zouOypSn3I6fk1Vko3wBB6nPhE7ie+JmunQ0BA6/jNsaLb
xp0/AdKP+zw4LeHSsrpM3xZm7nVQjdyrDe1Jkpcf54c1Pmk47buMatzEwO9eAtKd
gLZrSz98dTPamuX2uMvvr5gCpxgp56qMMgtaAVwdUydiCzbraB9exOnS6Rmw3z7j
GvM7KvjRG/MNM0pZhy21yhZKdqx81jaofCjhqPgu0Azu0MKigHR4TEprFHh97djb
TrROYYeNiTunW8VSZ9ifs2a5aTVLSkKAKFKHD58LYKVXgjNLMYbNpI6/vg1Drn+C
RzHk7AqD7oCvslqdLrrPGSpFPaq2vyIEv/Rmi7sFu6MqEKi1UNTv6Mc7EUMOXczw
V6YN53zz5lMLTKPyi8FFmHNJb1QtLkuzDLEIid0cMVktr3Iugr8ez2igH1VPEoiY
M6RUd98StWReujtXgx5E7u1HHp1x+/LzhbcsGF/oYDqeehFYLACGu+tF93Z2J3g1
qRolKEXvw/RdiBIPAJfmR9DgBU2W64cREArP/hrFFsanIPMjqTM6pDGFjmLSYdRj
cD1FuijYC+K6Z/IcAgM2atB81gcU7UdwZo+ceLC5HNsdDu8MyCWzSRxDF0j3PiCz
CDGAfDNiK81mlfhH3o/UXRNaW/cLHtHt4UbnPbcGhGPMpy2O7MEZX6XoNOujBTYf
+zLA+1ZPzHnHVrvERsnQNiM7j6v5W5tFiLUmK6TPATk8C5amo9GwQQ1uYLIIstTf
PJTeGvmSDGVmVFaxjfnVnuH3S/Y5eRrWgUKFeWxvAoDMPvyYr+DXohFXNXE2qf67
aXfunEapzRXKXTlYZdg2yGTIR4bXiL8hp6ZW5RNNIx44bBWtLfUVWSFQpv5SdwhM
p4FQV5uWAWZUq6SrrwEdIbNaILFDXZ4k2DJpCiJN89jcQhT1lI3eqQveh8Yg7ZFO
GDNkO0dgn+DxY+xMk3VPI8UZ0qpJVSwy7qWtQUQT4LKDOVz0CnFXbHE5daIEQWV2
c3UzXgPFxgw0pD7W+lC3zkrY0cKUn17QK04oeccpVXvsPqQJz4hwwWiOveIfMOuR
wmUCO8TOV8U4NUXr6VbgDYUm3U/MLQdWpz/I9XYW4r15wvcQmoDCuA7NzbFbZK31
8E9EMC0BkPo2I/rw3xgdp8anx/lUK5dRvEJIV7ig12pG8o7ylRgieW/2ekzdCZVB
+wfr1JPHZRr9dadEcnqmEsKFgDS2DZf4if6mLBvIrUWnuvtLVCWth4iwVFsRaTg7
FcLsBzxaUnODeshyaxmJYRSTgIZ0a9viWqwuQd9UCjLmUpIui1t/u7XXrDk9F1tG
2UCCC1i1APasqPh06bufaf++ktPCVrHo7Wjbzq2BxNnDPqAKo86AyAvPJG7vx75y
QpJ/ncoYXHOju1k7jatPegOThiNPednl9KTjYA8WYxjnpHJlm6D+LowON7eC3KcM
BiK1+ItW/hRfAUH80SMKgbVzIpkkOOeaIhIxsLKTiwRGw0zf5ibVxZF7QNm1xPaP
oH72s+cogp8pXocqwab5tu5nXCO9AW6+4fL+7nmNtrvBsZuq83Oo4mCv915p6L9W
SOzNb72iuCyG20ekEH4kXM57d7QXoaGIppRktpX2HYaGhKdr/zgyHqgeDeZnbTA+
HihXbSjx5ZhpMo1cKFPSfrLoEKI5X4IGcMmraT5jjur4X+HlNfxKxuA3uKwNjNtg
qrWNdeETqxH0OAH0e7jmv+hByvaEPW5oqPNCo1e9U8EW9dkcttbw91HsQMIs0aUb
ZHaGzN7CaFhxas3lgdf7sTfi5SNXdcyqIEzj1rHJX0C0LRUY+DN1ky58FzrBxJoz
xm1HOPrmGTHxFVCVzaEIF9jiYQfIKUHDU/jcjCxUGOTpyVio/mTWTCG68EPlYaUJ
Xb37Crf6opRfI66zq+rg0K0YR3vxRTqCgFwXM77NGe+nv7RKOxAJ4f0Am6z7oPic
eLRsXepa2Ps2Q6SLnyiIqO32rpr9V4QFV6ZIDvgDYUh39D574ZZF1IbRp2cmvvQp
xSlCRL+dFuhRwFdBO4DorfOqtvGUPGjRM20K6L7NUy9EoAJli756YZWKWL7wL0Ru
DtK6UAMVZWyj7f/Z0a7GioobLTmsAJ246iSt/PrRFUvP+wTvfFeXUyN7BWLU7/sn
l0X0QPevSteaiyFGQ3pc22xLJ1pEeyQPVLzV3X3DPDCfW8wALnpJw3CPVUhNCCdc
1opGW7NE7eeERrgIJrZpf6yvUuqSp5b4WJoRFizmDz6HIW2mjCnyuD5Bgoyk23bH
Byvs0SEPwp+FBsfvo0f7awoAaNNGGXiS3TFQLQwQE8IwV7kl7/OBbXNNjKKz9EGa
fSqsnvNvoBKGIxdNTgDV/xRGC5B2T/syS/1cpZftKfCRmQct5r0bVOwbkj5aQqV9
KlTasss30CFxH+TakOttTBPMPlX39vA2kQyNfX5cXqHbA/E3l6RRleisU7YKHxSK
m/NDgX95fcEC6kaYZ70xxUT+HA8TBzxNgcW1iP49xxvtL2zCj8vsEeKT2dJqCwCK
MqYSjPmhxggulsW4UUw9Im0QPbgUDddIsSwv4jN+sQMPT+luFmRNQycuIqMypxHl
6WWDTUCHR4G5e4be6xDQikrgH3jN5iQMNK2PBNSdJd9h9F1iJrmXUG8+FPld2FvY
4mFnuVAetqCb/RjdbDM1XIswV11QMWFzj8dqSWPoF16RqAegOCJYmfT+9HJRuD81
UUVjHPWft6SoizcMOs8g4T+Z9D1r0ZCYWTEfnXGPVgDgMdsMYa6TAFR4qjUKRdKN
zVJMo4BIFB7X75I5zP2Da+A8wwG8O252bgeZs7SkVgnUlX/wdNUa4i26dBeQG5xj
sYNUXxK0iRxUbulGzp4esjqLKvJET9MFckbXflZp6qCgoHtT39xiojFLF5X1HfdD
Sij8AWQsMyqYPnCb2Y+Zg/WSyRlM/N8w9mJdxvCkgizBmexNWE2tYl9exRgWewji
6Hv0Youg7vU4NnV7KdRuZx4TMY7K/khEMlgP24BYkQZoiu4cuXb4oA0Wle9Uopj7
F3xE8wUWoGjB5ZE4czynqPvUv6ky6gdnxeKa9s9x/Rvgaet7+KLKzCelbcQsIYpS
gn4wGKhjimjN600y+/VIP5nPSbsY/cJE73fIDQKJcJa/PuBy48RAiNYGOuYqT2O1
TDTcFlheYRSHs3euvAtg9tltF9/dkp+ck0s6Gwxpfh7X3fnkY0LqxOoo+3fKrgUA
aWrV56hzg3Tp01lLMyhzNjVi7i4bbi7GeyYaZG5HiwpfQ7B/kxQV7wr9m3zr/8/c
3pL+Dl4nJoyKBjzJY1PWE6Y04CQQYIuD6OMQt9VLs4iH3UGTa4Le3DQKSMIJm8hU
TSZKyxMkvy30ywPX41Bl3axAwVfkCDL0z/RAxoUwUBNfCPPNnO1jJBgRrV+Nzcrj
kEwbsPDtbZ2zanhbyDWHZ6ACIpLbTYQ5TABvAnGCBQX+PCtUtBJw/hUTiAEqERGB
YkKjMmIaXMY5pCRiieyZFOEDYjamPvW0YDfCW8Cqw39N8y9yn2CUpSbxTJnztuXE
bzU376qD7xtKHSaDaiP3+UjiW9Eoq2BRT4BEeK1txXaAvLxzqWnaAumjmKL2rXu1
2GroreqLTcn+4bGX9le0cheVAdHp36cl+8OTqmV3DyHU2DxpgQ6X/MZd+O6Mrnnq
OS+B3Rj2uA0rIu+gMCAPJJTj5QgQbawuave2CBt+BqU3Y5pFDypd0Ua7cJL9/sdX
XypqR/ZCFAGyqJVp2XmasGLwNxtMgU6ZcB3SWydvshgjHsso8XKBm2iUmtPnih1A
qPkhCp84krv4Fu4T1VVw8u5NQBLnx6p5I96Tt+aKSBG4F9PKPMEKKSh74rheCJVy
fbAWpryzzLEAmbM4tPkqsB1uK5CODWLBn/U7OLUfjzGj0FhyMM8eKXqxWq9E2H+u
lBwHk52aoCKBYLac5lAH8fWRFaukD858Xh4c0CiKykVlcfs04u51+jYyCSM8p5Dy
CEeUxl7/wr1pVtUldiFm/OnMuhlUJyKUhPv/fLdBFkYieD+gH0dM/tZxKR8TsxDu
MpDlFHw7Fkx8lU9dIYi16MRaK+BeAHT0Q5erKyq/IjPtSvILhkrQ/RHazCFsYurC
EzkvdpLCiRtxoChDsa3VpkRWrVZiw8+3aRa8OOZutMFFQbGSu/PCw4BUCf5VVFux
MWRIV1/rAcSjqGieUi7hL8NwGLhnK117PLeZ4zdYRaD7S0HH8vvYK5w7ElcNwoIY
+wVvapITSB6dXVZSu+rkHm4gkJbI7qX/bY7QZkDrKAcqcOq1+BYdyovRq08N0897
hEiuZsDXx17WvU4ZmXok/jFuGqXhvovb3Lhaw/UPlxGq2+C4O86k5SPIpo6qXNwo
PBkyIarcQrDgayqD8yA3SsWdAfliPZ7Y5s3OWv8psllT5sLNNsDAZM5J3NeauSHv
JC+opk9bFOb+zHrmUYXpQVn/xGHyIBuuw6PbhdpzmQUjIiNg2xqU1DdIBoJC6gVL
rkB7yW6dcLv109tURdJD462qeuKsamaWEgsLMsYhXqeLY7hWNa8F1mrYoSiqBM68
5MSsD7FkZMbJbfdn6Ofef9Kl6LFILxhgCh7d8hBFAs71ZHgUpGPxitOtfRhYPXBi
O9Ti2exNUFBUWXn9iczdvWVXk3u5w7ZGjjsTYBtUmRZi23MygMhE4DD9ijz6xEMB
2NK/gmkbK1x7dZtUhHmCcyl0bOOCRQpsgrHp0fdrnhtWiJxBTD3L1fsll7nveEWD
WF4dX540i+mhJnhTc01Fml8KzCrQKdrF1aUMpyTzNjmu02wtuEZA4wg3ucOQdzW0
/yCR+dAiTArFr5r1YAatZiTOtn46VaRKVxJplCbD6Xe1/EmwDP27pG3iOTKKk9C1
53Hhd8SLqfV2MFB+MLuJWsn5cO+x4xVh1farBfa9AZkze+Lww6IdJjmPHHEUQW1k
KgpR36UnZKnnT1xOZciyv9970fsuzvxvcBjB8gunjSapVmnC5Zq+xnzY1meIlaVI
GqESVeW11zTGD120QLWO4kVUFzmSh/YzJAvWXvi/4Vw5yrtePFEpt2UcbQj0+tP8
YZe+wjCkgH7sa33V2iibB7LDhNIdAY3cLmWtZMxEwb8VMy0la2Xxn9USMLkmLGuI
MGL9J9bYEjfLa+w+sKDNTyQ1Igg7MtkcakTbOfKo83zBZ7j9oWnfiwRgIkUtQVZc
r4sykes8id942B+SNp9TfqniWpBwBPE75wwLIEbTZrWtssvDdxI/aeH55K8Faux5
ZseI8ukXEHd73iDS5ol+O+isn1etdvzmk7NmoHR0Xn19iEqjqe1Wjj64Nta2zZe5
C1hODsL4kFrbY5E4muOxI0lj7ZJwW+aWFo2FhC40zFnfn4nKBEoHJDPfoRM8WHqY
H87tCnrE41LIQsdO5+zYRsAa1sFa2tluEf28Dg6m7GOnRW7allDJH+5U08OrKCt1
uRKKUij0sytpnVVAB6aWMTvEuMcqgER1FZBUsFpsAS332O2QCHTTzpurBSabAalU
jC+HIq0rNBry2dL/zUJgYikjeLL+PkZAUjK5T1WuNb3S03G7KvY2RXOZgyQ1jlk+
b+LABxoSjZFKDGmwsxeNm/N+zcU20KIeCxrzi/ob8A0oO8PDZ8BRS/eoWL5JKdf3
MX7oC2qnBwvF1XzerM7Em8hgiXlxpGQWTQuoJVCMQ8mH3jLU7SPNDsU/Ri4aZrln
OU2A0aoNrDJNcmQB+CmniXQMfAira1JTvvjT7nTCdMfmbWALVQ7JzO3PaidV780N
4ZCRuL3aL/5lYxzeFRhh561CPm+clan1pkn9nGaPmi62graz+OnEoZ+WbmpdZAXC
obwEqcSrvgXRbZq7aa4tu1npJW/uPb2C64DrRjpKjqYSgYNUXhP3I0nq4GNcAOTw
aEMuxKdSXpwH0stkPDDPQfgqbB78cwwms7V4HHDaDZK9uaw7PMuP/+OMMSKqk+mg
oAOhlfO4PsBC6rupac0WTo5BoZFYklgGqABqfX9pRBh/ohwkKuXZ1bgFlBmKUwpw
uT8VS7X4XuEuD3DFMSt8wnXv89o4ZlHmQLg5mhbqyURRapL8pa0TFVjcN3RF0LXP
ZRouOFYGueokIorTWgZiqBERggGvtKaSsb1blxaB6GpAzjiVu27UxS0PTmZ0b3N6
vcRnNDqZ4pI/bq+imLr9jmRIeF3Co+agRcOlyNjO7bjOXvnfkGAit7tGGk+yBGnO
W2yCChJHuVoAtSQLkbwPHn+oFXdx+ncopJHMKAoub5D/WAAqyCeZK6kD8NuHi6W4
C+za14mMv7qKZuqv9finGLUYuoXkfsupbztnXfpiknUFP0i5v3O4OpQquEa6I1Jp
EgrEeZqHz4HODgK9kmEUceCYZnFX/iEGiaWSS4yhH0vYjrG7ragthwnrg3O9bigj
hfp/uFxA2QBfHIeiKVwnLQmEGs6YP1lCBLSnKpupVz1VrDjsGNwHk7epgkotKnkr
+M758TENkDpp3OUyvvXG5FWjL02Col9bl7MNFJZ1vyNbKk+WAGJyTQVmCuDNwula
AaLxfEN1NvZ0Nsq5Ys5TFu4SrHyBTe6bsrVf+XvPAdXzJ6De5tDPvut9Fki+xEFZ
42J4ZxrqRn7ygCawD2m9VB4Hn9fWagKJGekAEgcDTq+MLu3ivcVqTuDkZob/yz6V
wAL4VtIa/ERz3/Inp8MW+FmDEmlA5nW6d494BvP59mrg0vIoNIyLquM9Cd9AsHn3
OT7zWpmbh2DKO1CMa5wdx/OqBYvPhfS9guc+0S2EYWq7S9h5FkRKzxz1rsmvAiHB
ocJYybqa5jHNH4aC8xXPZ3lNwFq6tAbOGjiAP7HHBwhujSJZLJV2h3wvLpaGl2ui
e93DQ7JpXEIOe4pIbL9Gh361EjpQwNzu1+dMiA6AaRXlzsCtiaYuRmBNfBw+cL3i
3n0wQbuwLGwyeL37rPVkmwceGL9VYDwwz9YBDupQxQoZMfBYqEkk+lLDBTN0jF9V
8w8DXZ8rpoQ1XxC4mgyek1lZwxNVGopIoc7lCxfEzlb/u86ZYnmsks/pX9Yv2ZwM
l/dhZc2mm0K4hWanq3jY/0VM9ExXj1CrGJk+uLmeaAT4DTnK/jCvy0F1S7mvuHkt
tijxd5bnvpOUZwNsKz3VgQcICA2xkSSrbzRux4VepKnlw2XmSDXhuE7OpXL82x+1
lvujgsIqnrWBZ67TwhKsGbs0Snt2lkNXY9zILgrEyZrzpUObVoCMjyqalp986h8Y
ugaBZVXcN9fpkjVbDHWHHwk6HEW58MnQlWLt2yFte/N8XN0ERgtm6+vKV6c65xIU
t6vW8TairNZqalz5IUcOfP8RL1Vn8NZKxpvTbT79Vq4q0OjZI+nPKdZpZS9riRJ6
a0IQPzNksVbi5YEDvFmTr0tDZokADsy7RL7/nkg60+/R/ZJr1TSleAgwo5qnw5Ia
u8EvfBeWTzNUjmRhdkeCnNPOF5aTnIMyXe6hT+7l9TdKC5ghubNh9i6DY7zR/2zo
bQgofYv7d5Iu7uF+6xfljfh045yrN7EkOvJGV/4LvFrix7I//OZ88IT27Xh9IGG6
6Au7czMBjsxqh9KH9UmFtic18OI/aMg87vKMXrrKe8gGZJLLk/Z9fMDd2vGLUw+0
xqtKU9MHLiEeiYrP6SW+hjOzGhzm/xzt6H+FhImudAg71ddI5nFGymqBiNXhPxNj
S/mP/WrcUC3X61PMMHCB3gS7r7/2KHxZL1wMglYxskjU3FRogkEn/sH1GFf5ShMR
/BfItOO/SSMH+74jjDeqnT8ngVsE2vPKNM/vK1BJlZYiQV4hPWSCfLlaW8gjvYoM
73yJJygfi2E9fv2OOcuwFj9QTQjX5I2wXY6JJmBlDSO2d4EZAb9oxD6Wg8ERKjQJ
fTloBQ6s+cNekL9v0HXZmvGEs2wE7NiiO+5ZCf3P1gqe5HFhKgWH12nweMQh3I7h
FLUsL92iNWEpKu6BMVWbvajUyz3NJjtsUOaVdzkkQA8KZtvXiRC65F9AqEyF8dnG
MPxr2zSInAX9ZAYd6Zex7kN+29cuQHBmsarrxJbhDaER6hBkxS7a8gujmN4HDGGq
x9mgH2Ln2MED+Dl/CMY7anwRleA7G30Zlmy39jX45EYYwKdoV7TSajYR7h04KrhH
rICddZEmbUCiH8Owgbp3+tF4GZwotFQrezwlxlBsON+TQX1RMTQ4C0odqGQTaGBi
EldiQJuYMvN+ZFpaoh18w1XSm6cUkbgzvXTwPDFPxPgtNEAIBsehcKBLyNlOECHQ
J7lAwEiFmwB1I42jj/5LypivkJOtlnBGbVkawvKR3hoWnh4+q5RKxDeJrO3Yf3bB
1whTFGf4Q+XHI1ez9z9/bq+XIkWzLPteh8+eGLyb1BQA4im8vBrSEtHZk3mdY3T+
rxMeb5nnCmC4c+2KFwUuh7Jd1AI5gwTKId5/fw2whwdjOKr0GGJzlL4ibAd/7Z3a
HZBTY1ULGYVIg8muOSGn4P2clKuaRSquwQEANGorZEU49tkfKK2Pazoyu0yLQ5h3
NKy7WoFNAJGmfWyxoXZHUT2rxAuAhBWox4xjV99v0GQLmH0yPvi/vL2tLj80/+7m
3x8/eBQ1hgo4VrDc1ampVQfYkngcS3UtjfVD8YzmJpiLLjiLFDgSUPmZ+teApH2S
rWSafRcG0BU5CG98tWacS9qwyNi63YJxBm7MddVgGRKVrp27m06sTFdHT9A80APc
kToPV8OKYnoLKfmo9VtL9MT+cRCyr5/pJl/dpeIXEDjMsEOJbiSwrbxd9yf6jjW0
xHbqOexP53maiUp8LqePdzZp3cuuf1rHTn6+YwIZ2jbTDiVVx8X8iUpUnmUbKyoU
WEUDNu2GQWUhFJwZ525Yc/jYBl97oscK0jd95GX6lb3Mu9OBcf1Eh0iZpKR9UznQ
9Z8xwSUqUEhiyFbKBVMuG0hbIXVEkm6swZv/1hn9XDYdpWI0DM1b+y26pYJBkFle
QvtogQ17Og+UfqEwWig0Pj8aXGIexdVF6IuZ2TpN9O5Ur12mzCjLd9NULbYKqFt3
A/2MmnZKZ1mlq72XCvAPX75Ty1RIsKW4F63luT4PhRV2pGX/S1bSRy2jQ8g0Z84h
sg9o+Y/ta+zXDoTHzRUO7h+D4++O3zj23aW81D+LMy7+/cWdbNpEvOuas2zhF4R9
F4zGI0STJoGsi1yGtSPj6sciwFpyfE1l8kACtprF53/9og+Kanofhvk/VucXl6aI
YrmQT75zm8ahJWZQQQaDamcirbc4PU6UITGcPvkxGU4zXn4MhiPK5BGh1rqvzvTn
iEkO1q2pFnmEjord7lgbNyelGqNTfuckQFHJoYd/u+SYABlu48yMgTntXN0dSMJ0
iTaUfzEPbIuIsvxPazQpTwqV+LBCnl+2lTZKgQaAFWkJN9TvU/D8bKolLQXiFPjL
4sR9xexvfKx0BkpSAUA98edG8wDh5CkxfuSTlxwqJdJPMG3b6XbQhZyfKvb8GwVm
qJMOjfyuH7YczJjfG99IvI59xaM7gywptnuv7Pbp/ixEzCzya8bZdYrk3XcTNaxB
26XDPBqx9Wt7Hfeco7cNJZWV4AIqdksKAPtJ6YVF9ryj/vz0pMQJD71w8NRx/46j
Xt7Xo4Y5MVqreBxhbDrY5vyffUbAh8YNDofhNunSKdYO08q9/5AtdOftpZSjF9EE
lDV0GA34cfZxD1HWPa1ZcYWbHRZNUT8ZZyMO88L74wXf+rN0SKmi3vSDm5Mu+QqV
nFSkzjGuzD4xorUiViISdMJlD7Y8QNsJN92FovISGERqCdvCVHQ8oBWm4bGt39aI
udP9vmy/oL1lbKow3UksdYSbTFs0H0PlkEuvZ/LBNYEy8pCmEACjrkEpKFrbpZsP
1/WMC71HMMhJbKNzesTtbm6mBJJJJDBAjLACVphX94pvfaA+F2i2NwFSX9xcpQsO
UlqpnKejPniH3vZFdWcRu7wcD1kEemdto7JMNWZ9IcegCbf3y/96iUVzPejfCyUw
ObFfQLrmxXl4N5V0BCuH7jwQkqzoSMT/97/grwapnNNnVNENGuiYklr9EKjdgjh4
XITSyMp4AYZIMwfiJeXIlRg5AVE0NBFRnXGb6nOVCAM7xZFAJSL8H2llZ4fNxubo
1e1g/G/xejv4RWsY6hFEY7BnrhrMDedxuK/jK7vvTQsWIgcqmjDaWMqtn+ByPEuM
DXNRx1S/o1mXJLAZdS4qABZQZ+52NDQMK1smF/X6ZXyscWISVTt4xHJhrnGndDYU
1Pbp++SdJ0y5xPPomA/DMftiFMkLDIF+4DK5qt6NKaaD/nNfXtR+xq0zB75BoD8h
ispQntx+2YtKYukkbTcS6NcR8l/6rY3NgjD71OOIvO5FrOrp3EqieBLvZdVn6IMD
0edo8oa5gj6ddN+sVW9e6l5ZqejFvSnuU0e+ajLkOWglaP8abnRKLhMf/5Q54Yxn
xaYPrhfbwxjgiV3PzoJI2OHgO2HhNodyg9/IjoSZITNyLCJ18QO+Q686ebS6RqGE
6nA+ABdvzsqE7SuDFOhXVgNKpWGoC+sJ7ff6hTQdVvcHtgOzQZqeGvM/oahw2CHR
hDiIElBLp7Kwxqo6p4ofMA9nCaQWth1EQRBdJhIJZkSFfafDO64WoqwHsG/TgUnK
UhcH3tSHaH05cQHj5ywkv7gBpeWNSpuPt8XiI5p2gIFnydyNf0UWNdAVrnHAUnU8
YlXE+bs+8k9SDAHwX5cC9acHe2DIA6RrKpfqie2S3/ZIcBcT/WPGqCjyGKt3Ioad
bcaqgfq6p/xCgeMmkcblGUxzEztr92BEsZ45JnanXQJVBNOrCw+OsL9aqCz4Ve7i
LJc24iPGROFSpjMFDkYcaEU5YPVXolUjYHHMcFy6fTSrNFhCkD5rufGzAWj2lJEa
uN+TrBJ3uKl5L08QIZ7P2baqg7fC5/4pmHqxPgwXAbfgUbo0k1NpDCKK8Y0k90Xd
LTCLF3/CaAL85Mol9EoX/k0LigKCJyXKkBluJoZe2NQ=
`protect end_protected