`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
ddtXksX2+yylW5zu6QL2Lhnb2d1sD00763mmSITNX595NcHTEkwn0zB1Dry37fOW
FufOhVzEJp80NC5qZ/+F0Vk7Ik02dIR0elf3clrjeJRK85K4e3Hoo4xn7YbFUIms
l/8VZSb14+JVGURjfswrIyCUotIzlzVYZ6gzoZwDXIi5gQIBf/gI+KxNXPaKV+PQ
Ufys/12rjO6aI/pPlqSm0hCvftmBcnezN2hk1UeXgOIuKZnogjOsf0iJVX2aOOWE
6pD/psybjbnsNB6kH5uFTA5frkzIzkzl5d9+YDm9OyC+k84E83I/7/j+rk4L2dah
QJOvksSIzN867/4Qt8qYTQ==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="MvBXkzurAa5VTw+1JJ70nePUfoQXBvZOku/SMmg4TwQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
oRtzZL4VJ4iwysPsC8SXYCzXS8Fw2gtZTOskLcDV+1B9Nzn1zTyNtlo6lNICRmmK
ZRVu2BmCc2G+fmzynYlNTnSa7C0Cuel6FYpxCBlOuk3OF2tzAmLAuDyOH3Z1Yjzk
a0aHuoCdIRKv7BrZCdALt03JeUmXKPdOmIlkVGFl8yw=
`protect rights_digest_method = "sha256"
`protect end_toolblock="Jn9CQpRhJt4rnzZPRk+dOpzAubz7omckX1MrFd4p81o="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 14768 )
`protect data_block
gD6l00tciPUa6pDNTk/+t0OO0nC/UTtBwLB41d4inuAUA3i/ALrNyoJVcBnAmEQW
ptbcNp5fxEUJjnOxnedyZEuEBxWRieZFQnkRdF269oNsNdDovdW5ZxL9jmH30FiB
X6VGrrfRRy2Cg6joO1CXetmjFzouIWgD7FnPZ8tk6HA9IY/AtKR7xgbJN901od0g
/IjgJUH446Pv5DCR5LFaPRdAJIAbreibHkbK2O1HKWA5zd7783Wpo1fp5Ol1IsE6
NIanlBKlYkX+czlijVtI1+fZMwlbw9rV90yGl4o3mh6aTjdtfxrsS7FCs6ipPYuY
9vT1fBKPsTIn6JfrslcxE61jyPBIhILvuoIOOBZogOITMMI7sXJwBfD86/qyHzOJ
R0EatEPjOIGm5gwPaoZP+PZ2xZzXuxn8bcGlDPf9jkeLx91Lw5QZSP0fplpCjUDu
uQL2SJkMaEj/IEFu1LHxyNQB9Zg1L8J8ZSoZL7Io2980rQXrhYrl3QgSBJiGB27Y
HOBJQ56s7/Z0dsyvkxecJTR/nxOmsyx/24sbKZDJdSxVC4eNBiqzWaITjrSU8LMn
l4YoC5CR3ADMsDWuL7sGIf8aHSwI5d7wqf4wVGHGbJ+LozRCZfefLtQSuejkTtCq
7QE1R4pA4uheCSp+jMOojYsUEAzLcJNgV255XdShvyBxdEz0aCUPMpKAjA3RJV6H
awMYKZUC/DAE6nmtW1vfEBiyO2JnBqMWs2CEg5P5NeyKuBZMxVhrg6QljIhcEUjP
byUdtaHPUtB+vbtG4H+3UHa824kI2FsAofyyb/4bzdwjO3tlH1DvBO1HSPp/7oDF
vJYZF3Ai7eNB3lFESKktN9O1wF3G5XgiuqDsHfeihLXClG8VmbHK/13ADFM3Q43n
hX6aW4tphZ3EJ74Km4zDfh/uYqd1HdIMzSBNJHqfZ588Hhgw1CNkYJzIZwmFxpPJ
CxgcqgP2eswNFaNH9aF0KjR8kb9DGKvUtsJ8L69qPP+UfbIbpXqDfRSUhLUlVJal
VQt/WHkmNBqanrkYF3DMslmwiLCZc0gRgJEXEVXhYg5B705sp5swpF6SGGUXhQj7
ih6JCe0u3WC22dnzC3j+g28ohHX8eMm+Nethrz91SX/xvycuKPnaZaXoUQOdVDCf
34UpWqhanM2kpD7sHtwdHi+nLJW9Z3amciJIVrus23sMWmu1PfWSy7tGX3kwg83n
d+CZdSmyx8BJ7dON5oZiwlCch/tux9XMcE7d1E32z6hcqPBtS6Janu7qUucR01X/
7mfJ+Kyg8/3KaDPcn70C0UV4EBUBiugvgBYhTInp5osPppGR6Wl+6PmdHf6mVG+A
EVTRYPb9okpgH8NBFVoaNO60ai5atl9jy7UVpaTd37ahVrYsKgXr6JGyeLiipxA0
Id4F8qlPzlcEjKXQThcSwPiruJcbduy8M5Eq0O5rewzfBINxH50JoQ+9quBxcE6h
h9a0N5kTcEzOabep8iLxvjR/Z8JlM3VlPpWLirXyAosUpaB+36dkV1mBTSPSR0cF
eAAN88UCYqLE07oKus8v1qQCpy6/Z42bG+2qyEGEhr+1ANnChx0XssOhQpKdHqvn
um/nhXZ3yJUW5Wax0I5BSwDuwVMrlrd5Sm10g5dn47t9XkT1UMzK/KxBpQR0ENxJ
Hy/O9BWI8rlAOlilQ/yB7jEUZ2MXLFxgtduSgUUmHWaxE0FMJ28lCT2bNC1oWwah
Q/V9Nv5TJIvkNfSg7V94SDvYM88b3hzzUPIiHzYmCnztJuvCf4bt5W2kwuRCfQbR
ORz5vZaXbK/Su2u7S/tglniykJpmUgq3ZQUxaCZlI1T39Ow1GXQlA8718plrFHSQ
cMBafc7ryMP585nB0iibheM04dXSnh+Km4yn3YzRDB7A/TeQZUogxduH8Xmy77Az
cJ9ldPU+fUAaPyIXQ3jgFdVk72ET8OSDfUHkdSs4f+PfgZCG4ED5s+u48Ijw/NCN
q8OyQeNttjaivOKUvPjh3/EDT1JW+NeInpCKtck2eYn1gG/4FTiZOQe5SwRauxKf
dVMhu0z1mj14TBSC3NfqDHJDq/aJ8oQJaNRW9fq7ZwLb/yCXAAcPbi3Oy4nm6iLe
rttVtAus7flUCHFWZXGvRJ5pvd0aRuSmC7Rvd2kcq6zMKe1v9hjeJ0k0nILdLtYL
pjU4x1rUR2KOy3TVgapiK+jkfaVL1ojtKKAD9gHxQ1yQqTgm4GCrebE43TVN1pVF
XVquIRGolX0s0X7/nSQuyAPqoGnSjX/6AHU9d49xBiE2JoktqkQ9zJW0K8STwb1i
u+CJ8fh4d8ivAyJzbMfBJvLlfyeATSIthr0aWCK4Bwke6x4mZciIgiOCvehLvl3/
dT5nTpJeWhcE8pi3xgKIcIa1eT+MVKQpo2oiuJUmIzsBXo0mmxN61WR+bf0aahl9
XvWas602zS8sDP9fpYHyUYPSHSApXDnyl/Pk+9uha19vkpdW7X9l6ms5Zigs7rDB
w1j3v8kSPqa7QyY0Z2VSbyhtkrbYDHxLxw+DlAxABGiBCS/C2Y/XIOXWAwTfHvrH
vxOQ4sTlSghhvnboKF4t+HXk7Qq9JafioyqLZqW9d/R1RyUhhp+zc+V90FQTyMAg
SuIWRXxPTw1S2ZchomG4nd1Wh2Zo7t7VsKN45Uypk4E2G1ACCy6exE/QPdgB2Pl7
U4VgkT4qAVzSN+BhyAa4s/etd/zj0NllxXDc6eUwToGUy5LY327CdK66GcneZMb2
k1epEqjq4XoV0ZsNw02Rl0tT6YMpbAYEoLmXSHdYHylpP+PX/FaVW0aUriXdKMQ6
Pl5WFwD/XLUvcndLV2gYLWlzgWv751PmQSOQVfF1LWbgRCcKKhWC6x/jIbCGtSEL
bRWiVRD2zXohze2V2I+BW1MlGI0BG3fObVq2Iq0uQuX8dno36dFtzxBiZqr0ejGy
VGTzK32kcQ+jdxRvNSxUvIPrpqaN/iWnUkW0O2omjnY/VPgOcstgKiDELNmzz4y4
ZJRiDiqKaFrgOdGUrkk5xZRuNWezeJI9t5RoEZ29oDJllnlGdCq+z0ZdliuWPQnE
3ecv9vjKD9Hh1HtcgqKSsAnwAO1W/JZY/exbx3nSWLn/5rXAlg5dp4dlO6KFz+Yo
HMqGSdrT3gCAf3rzqNKRB2i5cVzcS83LdBBtGoSP28Mhb3S2xqOr95vdNJqDzwQr
hR/BDzGr2DW9dpVd+yGuAUGXqocVv3N2urg/jhRX9NJ8Z0izArDv3yFxbyMQylK2
pJ5YZ84RpFqO6KTn/O6cYHoAbaVr8mkmSYW/K1VR2djs8TBZgwPwDgmzvJS+Tjj/
ujA0IgN/psg628D0FYvdHEtVm5yjL9EoOpQo07mTByR/dMvCHaO7eIZLZWo/7Bvz
hexd3Vhoeb2yDKpQiN4Q30+gyIeDeGCZvuutonK6piH+ISAgj26PbMM4lsX+SvQz
AHWqa026ZMLSivJrlr3khcCtFXO7zRrmNj3HMutGW/II1zjVDgiXLXbM3xwDrehg
BnrTWFpsjBMEWrK9MCMfg8KhqehoClA5BIvWMj9MHPXZb/cTi/uLE9lgOZ5pedki
fSeNWwg4LqEpalztAu/K2FP7oIAEiz8uPmmx06N1CKFLt/eMB5YLSjWmyM4SsJET
3e8CwJNnXofvC311nLEFHd6fZPC318X3OT0Qn/dZrPNCv1JMKbP3goYUg9HAg+9h
z7s5OP1qF2nto8e4Q8WFlSlNopSW/hebtKUqQmcfcsNWIzL2xXrYvTDoX9m+Yghf
iX85FL96GIaToJg3GjPeML1B8Wzm2OceIdXLmFdvW44pT4rAimESHNPYpTYoCL/N
rgCLnVCLSTtWfp7ljr3qJcWy8rqUhZVPMSuaTUSl4cApvlT7ZxPhhH2ul8XKEF2T
jftJdcGIT9GIAdevZ8/NJMxmkVA++NOs2FcHHM+qrbBhtUCmahh7cS59z6wTj69p
PWwdP53Fl0anFZdGblXIykyL1Bt/AqgfrL3d/s2ICJfpd+eOm/G0WWoejh1ObJDN
k5lMPwyyU4Ohs0/cnXAP/jQE7EZJCXJKwHWL7feUFVrD/Nk8KY4eDAxHb/TtLOHB
eR330sLxstxXVUF7TPq18Qn5PwhOWXvsPtXaApub7xLcBm/F4bOWfUy3Or+j/uXY
1xhsvHj32V3j2q8pi+PUHQY5i17t1vpeCJWaNZZbTY5xK9FMJ6/+UvyD3xOb1qe4
DBkWx6pJdYxUqwHZW3c2JRtdM10vPxdusqW2meg5oVPlBPFoqW7naBV8qdLd2Fb8
LmDkMdJO+U6bmA4J52+omPp3GM0HOlZAQ6Zqfhq6ildhOXfzha5vm4oWsy+n3gLn
3itXsKEP/MO9DkY+0zwqoxWI5GLUOsJyK14JgufDDzuKybsAFFlJVfaR1XrPAGqM
JKoPH8o27y2mhD/nXnVDDxwBgu2+6jsCzIBpu4c50NAX2P0qi3pXglRMXWglRqLq
96xR9KFOv7lqFCnsIVi73D6E3fvnVDaxK7O0QyETvaV65nvtHtuVOyALbGt+WMKN
8vsbcf9ARGNr8vRMLjOywYJZnZDae0qw02bFP6m0UQFjkUdgcV+1fSs2YPsTChaR
LC4DFZWpbcLUW+qK0Z9AWXCKMJdMzC3mq38APVE5e6d1l7mVG2MAXDAvIXdJ8bWI
yjFyZh6h5qXzMlsX1FwgGV0wpo3Jv0oRM/8LCa7yjcazlDeNlD88H1Eo5wMD4zgw
aKfQMoclfLjeQznQfKjAnYnr1WsOitfRu2cwgruMw7Syeejl2miUyeLeVq2bHGBc
Tvl9/+BFbWdpQqQPb5AnBn9m/dHAVgDVuLxpPc2c5chRLfiikOmhNkvQXlwK4UBz
lHzienPW8DwE3m6LfqfUXxiOXdjEO9oFQSgNycu27YxCDQlTVT6/rBS/Y6fCGvwm
oq4EW3GWV+GERNdUI+PVZ40dvVJ8f1UiB6jWUFQHNNsJfo7SOESK99KRo+cM9NNm
D4C7mIMWeaMCpJ//I1OnuhnX4VfmPCjHvmsTrhewsMI5sRI1gfNG1Utd6LkXEHS3
iRQtOT1FE51KuBnU+1GmbAliFJDF7aY/szizX+3O19S4zpLzUMshaeZYasqbGvh2
TaPBKLeHqMjPv728gRGXxJFH8Jxy8BuJc0/QRJQSFvE89AmS9UZ9kmGZYsKteBYt
BK+xwg65aA9B4f8OpSThzcrm0ujaNEtRTd+a0wvQu9IwF53LwhB3QwyIzjIjwC7y
cmgrbRadPs+UacqCw3U59rKEeGaX7fGJOY3jtqNTgr323nhMqbbrElSn0W4jT/IL
KG6qbGOxWyeZ5jK0bHxiYVHRjlNm/neEPUQojXrYurJtJTi5bdZEaRWHsQqozBNm
DvKBK/LG7ssSU3LJaWD7mVIUE5drDtZEvBGrJ5N/KyIMAI56ciSX7ZDcoqyWBX8L
7VzFxa0neKerwk1SYqoyQFJndjUM4sUMUo5Rpi5pl2+BCSp7Wwe4TF/Lf5PlCvpP
wCsZcINGaMTWf7Nin03zy5RVAQLUKqkkUH1qByOnyTG2TrKKDETdnwH8mtcvDKLE
Qzw5h4V/BJgYaLI0md6mlmu4JZ7/TxZROhDgNGo5ei3Kmk4pTLM4H5sTeV98saxr
VL/4uT4ZI3YnfZYUZPm1/a+T0IOO7Gtcs6s4SB9lMkTZw1lQKCeRuDYpQhtPFo2j
RYuD+aWhUYC7p+4F+vCM4w1M5nNxBqVarZsCCKMC+IKTnLapDB6JKKHy90j6b6uZ
755YKqOPYUxCsRPWaN2R+73zSiDrdTZ74SEBCuoIxpaMlN3vZ9RHMyiL5/Vb65np
o4dvg2kg0wHnQaypwHdC4XyD845vMaszvLJtvAr4HvooExfVQPJEJxeaNdqYfvGJ
ai/4pUmvduLSc6WhjBcY+WBnV2RCLxiRWq6MfMzaeaCqLIJGyqV90AO1YKHHromT
49HNDeHajBTSOdTUSrTYYC0Q68cmp06YS+MULSUtOU7sWMk2chf20irTg5lg2EPC
uO4phQ7VVatBCT1E+H23w+tKtfJriidrpY9ptpvNfHG0effas6j8PlycWd4uizHc
/rv6s2vJm1ojKfMRLr0dFckD89Q1mlgIx4nrsOfd9OokrD80/PKS9jKxeO+rsYZe
paF6TZqBRNV7xtKT/VK5lw8HoO3tSZAaP50dQFTqXvh1Wl1XXl0WpicokVgbIy6K
YJc7TPPO8P71JnrPjz0Zc2hP0Gb2yzLwCBkFhnUEGZXP1Lk/4+HrkEtSG47/eXFR
HivXHoGzVny1Jv01bHEFGzoYtHm0Ey4BtwFpYR3mNDj7tqqxfpK8sgmhiIpqXoQL
xXybJtZ4z6JPQMLdBv8BRvEgafvu8hOEsbVI5TMQCZRXf9X0OacSsr6/Xnc5expg
2mYvR+ku0tZ00PKcljkxgCvhVJraeTi2+oTXjgeZk3iS3yAE6okhDGXrLlAshgMm
mcahj5iO4PG3TTsoNFXeDPIOJNXpRn3b6sJaBcoGAgrIrcAvOmGzQV4Y4v4urr2l
Or8apcq+NiCiymv+Nn5DoxaiRFC9P+huxux/7uBXghQxrf7TIo+VY2ChamRvntdg
w3fo9BeraBFdgfn2AZdTdA61EkW8ug6kxXKycCxfsqV2i/e7bdtYKmpQR6+zfO/K
5Fnn9QTHX2Fz5MPg/HNJRIrI7mE+8q2w3aTgaGUsBfsFONJoF5xr3kAvrKXs4f8J
Hl5Yliwhc8R943sNKEVxLE23Ak7foKRk8ay8ttFdXMSINUmIkVh/z796h53kEmw6
txBUpc90sieTG4JA2HaiRytsRBZuqOhWQXc/gNEdJMNTFrWO7DMFbBUCkO8h094N
4pDrX2MTgLRvvoHlSKSBsM1L5vHrWDcUaykOkRUqlzjxzdDjnrclIBSVxGhYu+Ks
+keiaXPgitNze/dklA98wc88MplD3J54nRwQnmqFmKRrG9quA8TKTtdPvmyKbmhq
s0JaXxE9FzcEI3mWNHu2/bNFa5h2dHkGm3H89qMPVXUAJlEpMVkjIsjM6aX9aH95
Fvz03mt7yEnQ/fAX2cyOtaj7KGjmC9SR/bevnGOv/6e/TaN/093Oz9fnF8Zxi/hD
bp+MctNrhi8zSGIABEyLVZU8uIFbOzSa+hMG9iZq6AkYHdl8BOEb26FBZeFsMi/1
NYzT//zVDTa+OdEDit9NXbwE4oHjZA5MeYpFRCKpX/5yKf/EKJY3beGVHr7d/Q03
9RfSpkYFoMTpNV+zyeyZGCJnlVGE9p0JDiK3m0iNUCObe3KQMHetO1Kb2vYdJm/t
9K7Y0fhbfFbsjT9dIuKl9IYSl6unNZkHv5uwjg9cC7Rha2EDeXSbWOwMP9Kc3jCu
EcXufhWc4xicdhSDQc0p1NKR9z4Tf3MChmZM9KbwmXFbpvbpRchyebH542xvSMpF
SV3A18l2/q58I+U2uSuk9JAViShh9t7NiXGDbm8WUBTqhwrMCJr6VPxPdx/mz3Jp
AfRKqBvsmXBU/iWb0JYRZxiBJLDgFBrSmBeghZqn0B2ysKCOzq1j5C31vkUlyXJ5
6dCsaQGToQ/593NLFw85b3N7M4JC7FZG+1l8xu+teyREzMJq3gzY1cScthk1XHz/
0YSTHkO1VgvnPFZ7tKNzMq5/uuIJC/1pedDdQA9F3hSMcF5jMfNs+Bb/54nJY/9d
lk3ddW26O6lgEdn0DAkkk0jWL+W07cYxIhOeZDBhl6fkF+3l9PKo3M2P0pPA9XTM
f18ILzU+roOjWfg/7tQleu+o0n/Lg7U4YpVWwnNPq/8lzbmn+lNPm3iZX6fO6axr
1u9F2okCq0oFLwgGbFzGZw7UfAnTKrrPHffZYOrl5Y8vX3xtocXbXxIG/pzvsFXP
fPogc6LfIpRscwmCYTraKWXLbSNgq793llk6JthB96BP9f/qW6fVLrRFGQbZJtAZ
Nenxo4mOtnuvJtB/ryRWT+BGBQ24IIeCPS9Hn4xqM/YfSiyEupdIPeOIOUggM/b9
KSYrGNkKyA8Nr8bER1wiFbZBnj9npRX0XUkOjJgvyWakoCz5rN5yTupKiQqeeVF+
LAR43LVphE7v1llKbWIY44Lkl1zSJwq923h46lq5si5E+JI5Y4/cGYCWt3wPLZbz
wrIKZzSmAOk3a4TW0sELZfhCxkxbxNNyumk98qxmo34fRYa+8g0lfM9A4//EQDAn
mX62C56391CiyjsJrPcmdvDEfRcj2KGDgbGZEeIwUKfpkBlnQFlx/zO8WXA4YlP9
lXag5YcnyEuE8SeEQQp0AmRWVyCCmfspYtqDpbgLDuxOonpsD6loVQk/2fn+FomS
chq1Dfe9jcklkGTG6ZVC0QCgiHrY9BFkau4lFs0SED6RcLiantFN6NoYE6yd1Joi
C3sELaS2SGwR6c1ZCArsumJLrarCRfse4pfnq4jWDFaSYZWsMxPVg90ekW6jmWxo
eavrzcp0xIs+IWAxx7kOHFm9mKu0kIYJDUQOE0142uG5qKFd0xX2Th2Brt5S/vVa
iCfy+k6bkxWhtUfsHRH7Ao9Om62n33UhO4LS7O00EIi/iPZthil2SJFlDS1VgZFx
bDM9XOq/2RTDyb1W7/alEuePHDCzLLqPflMJJUugqZ+DsFaQvqnOQ6WojDT7jmMl
7V8chjz2HLKVUv6Qja38/2xrHAqgJUOdXCBR/qqAjh70CpuTdwMnrcU2/v6vmFgl
/DWRRL/DsCfQcUfJX0oWUDTCaz531kz872f6sMHLt5NNNHi5qL2qlkcF6KCtddSy
2WVrks4157KFcUWC4DLprs92VXrbs+RIu5l3wCLG+NWlALCzdhbBO66inLlErAdx
Ne17xmGV/JBCzfK2aRNsPo2iBLO84+IzRyh7oXL8zMg2PacAM9h/7fTt+DJjVspx
2BXIEf1NoxSx9mqf+0UX7ZZ/L5O+kVz+pWZuB63dUDBGzaXXtfgolax+/6HTyMBj
4GHxKzngPXvvI5t/RTGaA8dzn5GjlDdnk4t0EejFhH31c3lkMerq+0Yn+CGKhxml
NMTQh0rj6oQTkLjjfj25pwx6uG+T8bXmQAse4FgKTI+xeW/x7Kj0rzFwxKafi4Db
zZ4IA4pxByGqmPfAX+1vYAeogs3HHohkSNA0mwu0zRy0ySw77NEoW8nJfxLjefwn
zYFPiKLYoL2kCgG+AWBRm6gA7H2BBLWxhXAi1C/AbdwZhw85DGligFDmUS7kV5WD
nNl2JkSwjuKog6CoNHuABopgTCSY6Chj5S0c2+VhUEvaT95ys2prbXDcgp5SNGDT
09QjmaRNxei5HDXVZHLiQsQpSIsob+8+nzXpkd9a9Seo4TAuQm4EhioJzeeWqJgf
DcUeiprH7kKs0uznpCTmp2QeVLHVWbiy8UQcQyq8eHtf160596pZphIwoJP839Qs
Wur+WnbduL/65So0GAked/KnU3xuZqGMUF+5dpz35RbNKTSvvJOib8GN6sb5ZkfA
GeKz1GRJBlRZP+4OFG/jnmLIbjGrQ3+y59w566OL4sbaZSa7vmEnwVtz4W4bqrMN
S7vzGiCFSdsXHWyJx98GA4Nh6sa+n8AKGSH5X5gpb0ZsbtWCCRq7bR7pN9eon6T5
+Mhwa8fqD+fExJXyi6vPtdwYUMpFyN4fQn7MvzpEm0pelctSye09HwGe8Jr3m5Qx
dl9ISDxhOuv+7BNWaji0iPhmS3v055zWH8Yue4mJScK6S+bLW0hDAKXOEAyCtN4S
67L1SmwikWzFnYPX7oZm1Hl1BrMV6j461LNuq6kTyVjv7jqQHHxCQaiyjM4UFH/e
A2/calBjhFgxszhMMusuhlaQdLvoOk2PB8oklgzlzl/s35fx3PHdaYWHzCU/GQoO
lMMnB98gLNoCuIJAQPKMU6ldbsdrHzXxt0MwR+gOSMNp/NLzz5FkxD0sCljA7O0C
7USAgKBrO2s/41PsfMA57uX+1Saop5Skb0XxReEy+3Tnh3TxX+H/57XIvLK1r72L
WYaLiYGUO+sE8mLgEbXSkDaK9FBLwWFhVxr7DGa4oFkf2aGa8vX7AvFKjaxiDvlv
rVk9IJxBG4Omqt6G51g500iobddhjiKY4a6kFVHiy/5QH2/8EaO0gavSRSsJPy0r
n/BDUUqKlsI40XDfmmhW2baa827Dvu2UxCauxFY9nvGaDu9uTkH2TcGiexsUxy9m
rTYCtVO9z2Xzr3H/SX1uN3ZjhOVlF1tDzQMdpub/mt8LDN1M0s0GwHhxzgql5OHT
dTjfSDo3AqcHAIsrYbwZZ7nvMtTopJVE++dhRaYciawlUWd0f5mzOlfCZhIiUHFI
baAWmGippREGrMK7RmLvUNySaVaWGmG6E/pjvtH6n1XipFWciVrJ2IXihwcAJhVE
sX1+C7vIPvAW5pGRtxMhl7kr6q0O9UO04nZFkpM39EObHyYD9p8H6ZmeTiKojG/y
B13lOmD2xT0XuVWpKwmsTRCeE9j4n1CSUZnBkBU4HZRRoIY2LkZIl+ngQRjje4Q+
chGFVee6JpDUbwcCFgAzBxzAfYeXB9n5jtSshNyMpMrn081XAPzBIhPANLmxgZCH
/hBotObNv9YoJpXeIwtTKrr06XzpbCTAvehZy3J2HH+BnwaFsAGMQwC/wFICJP0k
sDHoiEmwMxVJYOE71u8/CzIZPgBrdZFy+4E6v53Aw40KL+P+1ixrdEkcaMxjhxJM
REreiF/VlvPjPdcIY1x6EXmFydN9KvjMS+bRChn++owFyHpEVCA6k3MhAG25hFG+
WvhWT1XTXjVjHffIOOFG5+zyu8uBrHlPfmTW34j8j4ZoXXVngfo8W0oQ+iGrxpth
P9/nLy31tTrIcfJNIJpQGGTw3iACr+Wq/WoRbf5oITxus+K06K3m1gAZgU4bwAna
TyvEylGsd5pe3L2YebbcY8YUfDTX+lzOlveOR1nFnFNH8pgrC391FtM7LW1U18xP
12gwt7YYI0z5koMY16J+aGQF/joIi4YQszIhYKUAjNtNy04JBbk861HT6EQ7ORSf
EQoIT/zWccEcV+VelMeTlfgepNv9k1FBr7VbPL4tF4BA6a0YeVF6hYx3DsAGmccD
0HfbXZRhXKl3BmPXHc63JBQu7Fi2Cyomr4UL2uhAh8lyukKkI1svnPwuVJHV8cNw
wLSunKwBAWZxU/VAni+RhHZKFKXB/9F+jzqejT0B3k7fQDYbRLBRiCy7cxix/oSW
1cFLHxEKPXMlq/rskRCSbuWoNHCIEn/5driUHwR5TdQyNtLF88UNw1JZ9UeI0iS2
Ydz2LpjJf1UFvNwtS1E7UHlvWmOCoQGqZoe79phREMkiPntH9kuh0pYbTXcYJEbU
VQNhruDa+DmBQvP4XIwvF1eqC/YYC2UZQIfrMXS7ZCcC1glYVxltkTOYiAYaptU+
bleSr1YnpoymrzEP8f0am5AMEWXoxXIj+uHHF+bDKV5nLPbqY89cUTeKFEdFXp9S
Zo7JzGoTXD6deg7gygX4yiAfOAsC9Vb+Uvaw/UCkrhL8w9GhKl3nKErJUPJDOUzL
ifcWLQX8km1Bx0/NUSi8/xHEKjqdzXjX1fAFpfNLeRCW+CajJ5eCv4lpsQ3+W3bk
WSvpTC/Nfao3k6IOyv4dj7xB1L0PGLED61d5l9rjtn6L7CuCKRTTsfmdoVEoqX9u
r3E3JQ/gctMcFHCjjZN+07veNP7OsoQtZBBTipHCaaqB5QJ0tWTv2UBcaU3q5miT
uaDTPYj0Fwv6amczbw1dbfHuuYHspGPm3ysh99vPSOM0DaDVFO1s4w3mU5dGOwoN
VrZKo7eLFGOinspnvMgOBUB8POeHVMU/iTU38b4HGtTgZD3sOvRzMGMV5ntV3SVv
jWbglR6nBPCo3rVWOPC0X/9A7eftAIImCI994eI/FSOloRjE9uMuy/9zwfqzySFB
NOX3BB1K4blO925H6JzmdNnq29eBvGcXY+5RVX7QUTySOeDClA3tICT+lS1rxig6
FnA1BlM0Mtca6XtSdPcy8+kZAtxuMUDFDzIidIKX2DtGiKmXJ1b4tdBCvq/XPRSI
w6cS4UZfyckRkxwaHgYLyZAQEiOeuJ7vd39ZYN3fuDqbifTBW/XFpwa8Y8f+/zr1
EJ3Bx2PTHoAAqTNk4BeTBD+9Mpk7kXC4vpxkJOrA0e90SyfY66N5BO21myrN/QZP
KZfmjm3hGmANx/N9vuD7ZAkAsX9UUupI5BYN7MbHzpLEmF4dQ7EpBgtiiqMmB2RE
IWopn3L6l0Xp4BeRNBJRMXHNn6IWbr6GSmeXD23VmS4HVlOqZvRN6bEc/amO+TD2
vqcWWk7M5dPH7yvOUqDgVN74eg8cHQKGGujeiibyLJdOQ007XlaXfJ4Iu7r4ylTj
+sleQ4uG1/c6q6YO6je7tI/MB58i+0/uMZ1Br/tuqQYbZJTeg8w4P+FQ0YC3+Rr5
t0NQO6HRbUvJhKj9lZDS7rZVaip3KSBkgjcWc0/lcvdjNhcmftwOrJ/N8kc27JYi
/0ncfjUbJxrQA6qyDPHwT02sHkWiCruw/NP0IGrHH3HyBObGfjPrfUnJhRL8W7TX
lE9QLCTXhsfjkuDjkfM6tEadzTiEBU4Cq/9Zp439msk66n+kTS2yrQKMwM5UPAbj
rZyUlWYpbuUNaOzW0K0eZQFNmonCWBv5QGLya9xJKXlPeUgQ1JOAB3OdylvYYvK8
eVQBzWqYhtUx3ZLs3vat7GDWqzsZYD120qdOW/2YVF7l0Nj8V4Or0dhrvQ/bVxHv
QwiCj9Fw48AVB2aUHjtaUPogFizAXlNQLQ4GELECGt9YPIwFg3hKqmPxOp5Zu4y9
X4/qAl7X7DHdKdjQ6Fr66TQjVqv81o3vfA6fG8JR08Ep2v5ETVG1bINNljAx3yLr
GPDQfF6kU7KT4Wx/vaVjq0IRPS5P58lw0c89OWwm7ejwcrG/O+HfwyXGf4zQmX8i
5xHCwsCLw7dNdiktYP/OTHSx7GG+pSd7R2OrHcD5zpUJgmtmNMO5OJ1n4zPYd4Qv
BSpwwulNPj3AcAiJlnPlHrilYeHBsUid9MaxK0JG1cASwRK59hyynuUuNQNb71AZ
NAot08L/BP+NrxvMBikLXy3LEyY0eIx+3tqzL/C3XxeFMFiAIBNgOOG9NYqMHrQ9
J7Ia6EmQEPQNLXWmCDmRwPYekkl5yZwNVn/HFnuSbARYii6uoHkYAR84vV86jX1s
0BKDMpe2LNbRaf5Aq+OzJGYjGaB0coyyYtRz6pUFLCugnfeuRYEgQKNUJMMKQOjV
cVuBw7COL9IEvIVU+w+n7NCpKzSI/intI+r9KT3eKwFuiDmpmIXk42MKssle21yM
hDV/SLf9Rg6vcFHNyvp+65TKLWVfXTTL1BDUCj/UgD8Ib6nofZS0u5D0NJcpV1Dk
1yrVr75zIWGLZ6lh2uqvm0M7EbRQNhtkwpewIWIToE2FaJ4UOvAfrurE70b1ZXUS
/H79bnC6pO+zxJHaju4zhRaxmrnnx+1e9UQnkmC8EoArSkEhpN/AXRDRQYBQL7Fy
O8d2xFOGLZzHx+IDWwjP6DHtcjPN4/JKgp5WkiJh5uPr4Mll2G9iHE4Z6LO5bN96
GhSZ/5WGhiVhUILQFMN4B84gfdGpNu9rYHTbo5ILCE8TQylvNTYM+LjyJ9weQ2sB
BrRYgViQzvTU9cgIvN+lEO7qf/uXLn9MqBcaw/huaVYSVtWXxiHG4Nv7aicffq0h
UVoTqDbMVevCiVBi3o6FbY+Uzmj3iLd/mYs1AK9jyrdrn7ToUhr3lT+np264AmfI
NLRCjEsFOwt2iuOm/0BMA9Sr6ddpBbb82nAXykZtL28s3Nr5pzKzAKaeMOwwPesT
LLjb/tytkbDb3h6KkPTmgcIfLmre7eg/1eF5icWj6TeuCxd3G8iuAboPi/7on5Ad
YxdZFKM0e0Pjyms/uuS3WVArAAtFy3McSs7SgS+Q1XL7xuAhuGdKGgE1uWDLFE0j
WR8dS9YJgtMjR60mFTMjclGOjAX7zUthor9/mXCgKEDk4RZmyeh2qko7UnvDYvby
Ft2Q4gttLnus/aYNpElK8sgfUPwpdk18YhODulNf+RhU3ROxq2C4kwH/HkQEs86p
jxrk3I1lOZ+k1+cIpAcqGGpkPgOKn5wQYt6iueatQTOWVASTkD3pX9yoXHrO4JNa
6oYmf0S5VNHA9zjHySeDyGWb9RYPymQ8JN86Ndr9AFaq8jG3b+CLC8TAGLzFQpki
s6ivvcN/Lr32k11vKNI9vBn7aw3DgVacLHo/BLSovJGAutwyyH9Sm//tBUgygYFM
Y2WB9MymoaZWAWhDciG2lAwXkicypt7dKWjLXDook7LwS7JikobcAC3gQJD2eN2O
elVowF/yxxdDligzpV02qxl0seVedYJ8aEfb72fuRRT7b52M15dAffAwkTAAX34U
O7XUjPpOhHqVPlwE+w61u9kiO99Nts96Y0ZOkBGrB7nt7tKlIuXKzobhmCaMhzg4
2SO+6xaoO4zND552gH467uwDdrD6ennzuVVQ/Dexnu5Tt8ENG3/pEUiof2FjXl/A
UC+11USZiX+JYsuVPvWhTmPmhJSY1Q3/Jt031GB3JeK660yWQypbzjI7pCsoQ9KU
MvSsF5dwPyQyrQvMTrOarna8svVwj4aEPlfnSUEOQIoipWsCJUrU+aCG2M73m9U4
80h5X8AoPjifHXCp5Kr3s9LU2OghfgcL9NZnl+aDJHIpUJ5Zznj6HKqBC6ib+3f/
XbIDosg2q3a2GRe1f4Hzvew6VnOo0Yq6wBcRyY3f1+YRNtfEsYfg4jdSCLjOG0JH
HlNo1scpIR1uNr8LFRBN/gy/4+7LijuKgIr99Oee5uCQqUGkhA4mt06EyrGUFikp
xEYpxcmMKqQs4xR+94T/uwigi+B5HkbitQJWS61+uy8kndswl/nzJlAFJtWI6pt3
FbLha1epRqhZIJb1P7mpNkRs0l0rjJcs9GzyenevxSSjhASzattk+WwIrVyUpR8z
GQ9k9SBqEIns8nslkvSLEVmlsrvuiNug4g5P63hyQyA/73wAWIIKsqif9Yz4j/yn
5LwX1DX4fm/V7awC/SKFbW9qiWPGLsh0pdFvskQAFjXUVx5H0oPUGqX38hoPoNCe
9X2/WA5i0foc8XwpmbCXY4bCpxl40TM0nXCIbBUEw2ZjbM01T1qp+osvepmeFLgI
jgvJ4+p6hwBP+aKZ0+LxRdMjha/AJBX/qouXOosbdaW07Q2hTHyVxK55SKpELmHD
zsByL+SdaUHbbg5k4o4T80KlEkc3xA86OxA7+mFu7l0QMdAaKQqqwFJLyLd3dm1B
Bi0KAKACXv/LWt6W42ttcEaBZScRbNjL6cGwB+MVQJyIdtxeAFdLKMAtFDlMZ36S
HueJ83Ots2ZCkmB73GXcXrsJJICeh/Bi1k0t1G7J8oJTwI2vMQA//WXErKZM4B86
msc6+WD8m+w2Tk8sXInZTxPe62TKz8fFrX9pPcpo7SJvv4J/9bk5GBW3Ti/iE/F2
nPxOHEfsOluoeyHQBuM07UK9ToxertdmidQC/AoEcMzxTd36q6jO24ddVJ0W+upY
d1S8b4TkSxi7G0NvmPq1jgNX5WWETBcsMdycWMKmOIdtP97+o21nlMtm1+cpGg0G
T5vXPLZVg27+Y12+5PfvYKwqV8+SDNxw5OnQNwUP68XQSRN+U6t1puNWdpzhCL8z
YQ1zZUsgoEscBVzeeeno+K8lYmyc/eiZ97aG4atKU20bAfVEYL6ikI5JMkmLzYsP
F2oGXdxz/DE/uB7R1x/4pMAUoJkidngrk9vMq9Cg4LbVBSO9tuQ8n6KttaSUVzgX
1ELvcPdClJ+P81Rm4abJAbaMijkbmAzprRQeHsODqd/qNQV5zcWuxVbNsqAfa5eu
4fmJksbEHqhAlRP+7agdgHOuV8lXtZw6bf3c7IHQeiQXwFjIZb76MBErGViKOosj
FyLyz49KSlBPTEUSI+syAWWwomOOX8/5WgbTSFNoNwCrNJboJqpwD2ANd6KEzALH
PSWGhL3yPHzBSenMj0uPSruDammVhwwtmSZ/Iw0sBgzaiPah4GcFMZdPV2tveM5r
Q1/9x4eW78thEzDqYKX2NCewS/K4nvag7G/qyeJQuNMvzhVBC1nRRQMGXjt83z50
syNoA5Gtw4moMmmlltxIMyndf2hdlNEnAWx5uWXRYsoERKCOqaa+rC+PixqfW0Di
GW/SBiNvc3VGFPHbcbYnEVn6QeTdt+Y2LTq9VsLicqWrCsLEVyEO2EpLHDq5kyWm
jWqx55WAowwj6pbzImFt5ab//ErKg3NxzpB6Q8BqtpovDy4kJavtEJmJoXK0gUFq
BRlYZqPX7/Jw0tdZVKHTBQWJEcwkvuJq6WIa5uJQWxF1oPfKSmINJq2IYiB1F3li
I8oUp2Wn74cQQ1s9ttFNwfK/RYTSdvp4C4crT5GohRw5zruP9oBJpsBTYI9pYHrG
ESY4Hndo7IRIr61ubkApTcWdNRs1RKuL8Hbq9u7nCmmDEQyEz1riqeJQD+cqO7j2
i+M/367fv2rhnNKDFMyEQKxIW3JXEU511GtywlhunC40Bqa4kIQTvlBsDy8q0YSm
BS68zCNKwN8SHDgYVZMc2+7uOjvpODyCTts5S362k2fkRM4OsEc566LVMh6P3CjJ
KjguRWPzACsbjwtQgt2GFg9Vp4VltukRHJUPQMGzdr+gF9J/wkJ4fYE6tNkqT0N2
gGodMkrGusc6MJKbJTCVik/Rm+Yzg2DrUVERkjJSIXkK4U1y9vAWYr5nwEkzag2N
L6il61uvO/E2CkVzEl1mRwVtTxQIUlGKeTKwMP+t/n2xbmh6/GD6Jge8QEar+HAP
nXZYlCVf6qxP/PNmWxG3tMdNij1tvd5EV/DMue66Vn2jV5lhVJdn+nDNR3NBhnjp
4LIiF79//GPcv43qw+s0uU8Xs3JBJTmSardWCnDbt7jiucIoKSyOweijaNHeI/X4
46iSOAbdn9llEmduKmyTAQ8DYSBX+5BPMvgzahx9nr3xGZR8wclsLk/A0eK/yoda
ffruy+mL5IXJ9DEfgiPrBJvcaFePc62ikOGZGk8AZo6VIf72QNJkPd9OtbFyrEk1
Hk6+dU/s57dut3zUsSkh3hvo7pPlfpbwLhGQEi4fYIWrAcrKEuSiLiEbDnU11E2j
2MgOnrlMlOGgCoxxddpPGwZ4PA/91MdgBlUYEqX7AXpEhfyYrhBpLvc1Cb6Tznir
59SdagKN4LhWUZc8+X8ztHw2jgHXy0iVjRH73u2T6neeGgguR5zdohOt82xyURzu
RS/9po+WULxcJPv0LPwvWmIsy+hEHGa1ROtY7Liy1cd6BxC/LmQaPciWyjU2AwuG
0hNkBPucXW9BIfez3/t8E2DoMexWAsB9/mk0ynINNRHmtwJKp1/Pm09wFt00lsaz
zBKPygfC6Jge3OP9FTwcQAIF9NoU0q8m4gmoyetHPjYNoN5MpKSeAb3i1m0P3lhK
Z1xgjixdBMIx7MgeYcjKa9g4p3zF6o37YgTPzVe66qnlUfGmpjlnZF3KK3ZYwjoh
Ikm+IdbxUh08uXjtBgzUr7eyw82/S+gKfGX0rZ3b0S4tDoeDoJkCbXv5RhpnwASm
z+dSR9l89KOzuCM1VKS3uZI4+ZH9M9l2QBfcUDH10cCzmEvwU3d+0GTzRyseQqGw
qK7yQEdWvwNe3uMker2d52Xj2LFFvVseEwBcEGfD1IIuJ6qB8k8IW6GkRqZxt8vc
g1lEjs5Nm2kVhLOXGh0nB7TQl67bJCrhJNSo5D4UOXXHRPmg3daR1zsIsx9xDpIR
hOn2ekXt1ZOPBJ+kxazRt4hAEp2FOE7ndDyj+IokdodNZynz39jcpQ0RuYM4hGWD
/H7K11hG9yhou1+x5xfFCMD2f87nbUG2U2h8gFHkoMIqXS7778YbPp1kxYGp5ecl
7xn7TthpxGPW94QVKDG/M2jX16KrhRJAwIwBUXIcoOIPD86ued9oeWcYn2pRfGvX
0vYQ5/B2IScYELInqnLyWSMBJZg5d6Q/l7JTG1rq0a5NCCfrhFofAC1M3YxL/F6o
CZnQYEPHKBpHSmBR+eZeAJDnSi/JUBvOGMLosPcwTxZLxW88vS5a27po+117LXbB
GKsudYrOP+dd2ZcJ320ezq8nNFfGsjTMsaQiOrC7S0psepuw+cG7RWhJtLWG3Qld
BixB3v3Gte+QjotXqpmahBtpZ4V7MFGQSiowraTV305yFtv/YL5g2DoxMDDiIhtQ
s+uIt/qIKzN+bfeV8D7SPwi82W/jlcUipVZ6TeIUCePjMNsuWj0SkXzhbNuH5RoB
A6jDNXCeLjq+aINhW0DAXrTd5bUgh9RFINOMDb9Ci05PVQ/8sSHqDiXoR7Ic8Gjl
X/ys3TBc4ptiJUjLk0XmpsxLl/uIlMbIoo3Ul9LEwsCuz4TawK0TfsL36xS6dPt9
VHe6F4z2de4bJm0bCr+bg6V62sisqjYCJcNR+EVqvsuc8h4wDTsyeJjZOKBcMyT/
L6DWd1Nhl+GWLcftCjx0GW7WwSPnN/LQMphbcU8hC4s55O7//JD5VBw2Ln2aIj+h
fppPKXouCgPdGhRtTgRO1UaUh3hkfwp1RU1FoAXC05AtwXikKGAuFOehRDh9CY5N
3aFskmHcG8yAM0AkZdwXYiFEmkONhs3RF6PpYP5L/9+5wPiBSUhtWLiy12M8dP+z
mnDxpMQRo8ym0228a7uH2Cx3CwNyCvzsECmjzaJO7Dti3bOKtrDWIFK5Wel6ivEp
pkNJ5k4jmnBn7GKn81ily3sceRFsxAVIeSPA4s+DAOwgdl1hFOcnRYqn6Qcl2lq+
W0pcHBNuMxNP9Ov+vHBCymEeTYVGKbyGtwACSiQVIIXrMvksXEb64k94KN0UQxFw
A8NAsD83Zpu7Ndds2brrdZ3mngnyfVcXW0bXdzckFSsHt/ArQIx27aVd0AH1DGhv
W2Ymrjf62QwV96ypt1VrCFSeOjPQgURsYEVBIMksNx0YTLbKPjKyaa1wiPde4mV2
UxBh04l0/D5JwpPDcOYRILutuIxStTt23rqnNhVPKqdvtZ2E+AgYQEdFk3XkOb0/
OOnj4MAclapToKS5OAmEfu3DKsMhNMiyjkhaAwp9WYa64tIf4TTJB+l1MD18eix3
H+KaCbh+eyI7rF41MpupcTAYO3/rLa1wYHw61+rPQBH0qUGmZK1Yfnet0vYYYTn1
bFhUihUPsZKslyU2PzxwW3QLet7miASHWP+jc6xvOExcO+DQLelANFDODmPa5bqh
haICQeakVV0YElwh9eqfx3N2PWtYV4srjEPnA2fw8niCBaw1pT4nhoZ45TJ8wiNp
g48lGzWCTKTmiKbfA4tLbvBV+lpBBEy/VX1ShvcNoxXnqivf2oyE1HCq/FxQtaLH
u13CRP5HV+H6Wog32yDRWmbe+fz9eJ3r9pYi83kNmr9oI9nolJ1kw3k5KQ/FY+B3
+B/8msYKSL7Ph33rLG58XXiZvAfegDtu7Go+4WtV/tdclcZhfFdxQo1Ak1nqM/pP
LVZucvBJb9eI9HMp/JSyMxCSiR/TDrbLk1sH49SeIkl61RdZznQNRba5i6Ag4s9K
260L9/k5d5qm2T0bcXvnhB3yuCrTf4IFuRJvBAgU05sa1iX7fNSeYDyHu7FdCzlC
WqFkG9cECchAUpgMHz5yBpnu4/3sugSMxTjhnaW5hnI=
`protect end_protected