`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
ddtXksX2+yylW5zu6QL2Lhnb2d1sD00763mmSITNX595NcHTEkwn0zB1Dry37fOW
FufOhVzEJp80NC5qZ/+F0Vk7Ik02dIR0elf3clrjeJRK85K4e3Hoo4xn7YbFUIms
l/8VZSb14+JVGURjfswrIyCUotIzlzVYZ6gzoZwDXIi5gQIBf/gI+KxNXPaKV+PQ
Ufys/12rjO6aI/pPlqSm0hCvftmBcnezN2hk1UeXgOIuKZnogjOsf0iJVX2aOOWE
6pD/psybjbnsNB6kH5uFTA5frkzIzkzl5d9+YDm9OyC+k84E83I/7/j+rk4L2dah
QJOvksSIzN867/4Qt8qYTQ==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="MvBXkzurAa5VTw+1JJ70nePUfoQXBvZOku/SMmg4TwQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
oRtzZL4VJ4iwysPsC8SXYCzXS8Fw2gtZTOskLcDV+1B9Nzn1zTyNtlo6lNICRmmK
ZRVu2BmCc2G+fmzynYlNTnSa7C0Cuel6FYpxCBlOuk3OF2tzAmLAuDyOH3Z1Yjzk
a0aHuoCdIRKv7BrZCdALt03JeUmXKPdOmIlkVGFl8yw=
`protect rights_digest_method = "sha256"
`protect end_toolblock="Jn9CQpRhJt4rnzZPRk+dOpzAubz7omckX1MrFd4p81o="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 4720 )
`protect data_block
gD6l00tciPUa6pDNTk/+tzLxvdHE2s3DQL3/JqqujQBC/Ei+vcAB8wM3doqg5vTg
mdfn9XB1bLOis2CVSfu295W2DNwHfMSTc/8BhCDRnTlLIX0UCJs9Za0+LoM0rMrV
T7EjVWppbP+Em6PkVKCwlmIQ7JKaifJ+Y+kjw9HCGboYo5074hY+K/CBbfsBQY86
NbkSLCO87IQEY+0Q2aP6t+beUiA4f/kKWE42x3SbCSeVV8dzAeuIHiU0G/K+WH8a
Cz4nGUVD86ljdZNccxGtdfHXOc/ZK0kAM/aZi+fevNqrZGR3hd7GH/ZOor7bSkFh
JWF5XCALQAnhInED6ZZCZ0dusorMb6spYALAdHpaLl5nD79SqFJnPKlT9+CUdgME
7AsZM/JF6a3oEMSBEpdGv4Ok5+1XGC6+e1VS6L3OiEeOB4hJqI7KoJHek4OKS0DB
lo43fzmiTFvd2lOr8MPR6lEkInxg+q9oZ/lxl8YVI0UTLtSTf2xRXX4C1NLUKJEp
oTtSgCJOHFiGEfUAn3OAtTQGRMukMAvpMe2Jp0O/Wo72x31wyeopX+1JVwQUZMG/
jfjJsx+r33PS4ees4SXM5JnY4Eb7CBrGu5dGCQ3w9Jcwv1dCB2+d1x+hP7CocBxH
E8IPYu8h9FuuaZ6l+PsUQ/0+XsOlPJJrblK4YULTF8805Bg2WEAyjIbjvsLhb8oo
k9uikhLxtFlsrssqg0ChcmR05mOJzgYoYMvX2CWVIkXlhAS/YXhSpduem2+1wmaI
TWQ4/jorXst1tcd5mzwnaHxVMpGovVbvJza6RSAge1L82Lml/w36OfxGpG5VTffL
SR01c/FE4C962XEunvTon8LSeIwJKmIF7XQpNjbqfIgrnQ/gmkUZ6xiKZG9Ddb5N
EMaPWl+jctjrUd7ohDJeWvWzgIoC4LKwN+PceGsGOqzafCFkQdrnVUBOkXnaPf07
M2evmUmJ/WyZ3CG0gT6jMKDuBvygdeEiq4F1293PgsnGL0G7kGCS8hUAnRLlJdUw
SeApBFwNv4IuWymlI6UbIDOaThFpA6JyPQD0Xpy2uX82VTZNGvt/v2p7GFdXmzpw
IOvu155bQP3m8v5jbZYH3BHvsdwyjerpphnQE40399p6K+RSZHepDaFiVSidirrE
wZxBSMKEHnAGGuSua6AqXy89lYbRzZmImYNlYpN/aGBNkn/QDKGK2iIANoNj4M7v
EPWX+6c9/70HMGksiEDkKGQLDpBlfUKPRQ/dleMEFt3q20ap3V8oNXm3pUxBehVM
zc+AAj+w+nGu+voy6Aq4DVK4rUXKpg7ra97a33GN448ulEaE2OSrd0Fd409UDUOp
yNQ6MjZR01Pg89JviRPBNwANiXv6DoT3fZZZpTzex2O/7u6sK99fGM0cef6VzWUb
AQ293Q6yNq4KEU23QzcOnFBOL/cQzZQ7bkYhmbMudI8aj4ynJuDDo+1GE5xlOmd1
b0DQ2lJrOSi94aCrgK3SPyq6urtKRy7Avk2e+51ObaA4IPvhCOVSVyrbkT6w/bnR
2Sz09Tox2DTGRlT2EPWXqqBhYfErlqlrfSaSnEFUY6XirC5VRq9OqJ1sgua96ip6
rBhtWr6IBLvPh+uveYtoD22inWCmQuwh9mRYr6xvvfcWpEmBj6E8PwM+7Fb8mgGf
CUBKgFZ20aRh/WQqAONlql5vIwSB/Ms9apPUiJRu7au1eDfAR1KsyBnGL+zDQ0qb
Et5XMMu5YasccAxIY+VCKo/VN+tCrIo+o1PD+FBl9COb5Jm8RKxkPpSGOKdQkUfK
KQDEuA0fChTyXzKlRR5GQay5AJVaBArMgw/+ibgYwFjPnWd+16Ir9e6uBoxYNrHi
AmqD5YI8qbGCcvkak0MD+dbMC4pxJ7eflTNKJKciACgWJrL0dMstnAYOXuv3bOpc
hy7SH+Nf0WrZASj+YEaJxggdopeDtx7eR37TL9v+byruDb/VFexleCfias6pz+5A
I1Jar7wYOIDr/Mi2PFMCHhMBKcNAd5xQyKaG2CI+WS0oELx4y4fOXL+3tiAKObBE
nA5pvxpo55HVCoN4r13YVj9N5UmgG8nnJBs5g2pL8H4TYxPUkBU0Vdj2kbbBotEc
X6LRbVMbO3friCJ+YV6wQ+C7GWdwnQiHNufJU6MotY0X1eBO9cGr0O0h12pB6ncs
QfN21rWFu/pK7Yjb0BMDbBoefKlIMH9Pw24GvXBL76o6M9tnUCmCxhM2bI/lRvVW
2so/VlRyEMcEkw0LcOJ3tsM39kYNXxdq9sHnvq9s4I9eEq8d5XYBDws5wCxWc/J4
7udK5vAScu1hfJJ8ckse5iJ8WQ0BAi0/eXacN0mCxMIrPaFTnv5VQfj1ASNQs3jh
uBpWKGMYK1AQICamkYcvas/T1wGjQT6Onxb0GvuEf7UJ9v7OfIXy3XtiZfnf/flz
htL2XO8ShRlbCzb09Uj09LhKX84vJXF7Y33T77Al4i+ZmVHiKx663I4V/vx4SF5E
PNumIdq8Sc88H5zzidHoV/3QsEC77PprHVmttt/qdYOs1BMYrp+VlKprhAPicLqZ
IBcljjkoEAkqcimNhYzDMMWoZW/cQi7ahY2fOmETZPVVzWhjeZLqJ6QQMG3c3633
aiefG9bHm4KvAxE6mW5Itj+TALwhmLSHb9BjZwmg8k51yzHehlNEWbV9cJ7oxLr6
N5MYUs68x4W5mRIJOJr4uE9OhAUd5tCt86Rx6HsWs7t68vH7GCpNXTkNPMX1z25a
Mmnyo57v3KH/zbkkGT90UvnFt/EeTnUGSarFJtWvVH3ba3C1ahhYSj/hbIAvwHhV
5Rxl4vFxrhXtp0pgEKPR8JUKq2kegPfVfb1QyzMVKx1N93PX6+b+jI+QTRSlM8gY
T9Hb4ER9I7mlFrOqbd9yoinu+n22PFbuaG+sOkRQP7x7UleI133GbBOJ9dKE0Hlj
wkQVZB2Zj1K9P5MbwWnRjdU22qVG8dOEnjrDlkOmh4xWNkOb4lKQa/JugxcdMYh6
lj9uqArn/E1sNT9NvBj8KqfIt7ItStvnV0RoEWGTW6TU2LlTbvGHcELp/3YYmpVF
klLdxPZKgczeualZsKCeWLosFZGvDxZb1caKT0CS/qVhftYw7+6hxuWfeZw8aR0S
k2vvqPKHPaPQ5jBWWiRya15r/p6GDru4e1pQYYOkMcao1wIuInUNUuOjadvThyJE
JHKkDA2vjcxQXCmFhujzHOCe6gr8EDEEr8XCKLBXw6+3mLcaLSr2U/1Ciun+RTXv
/uKlG4vFr8z7IKx3SaiIPephTt7Uif9ys5Nrpy4BnDp0tXyex7NV/MFi0COLgTU/
99KeNUVPH6Af4zNEuNtUZeh9Kty7HEZAMinhFLH2rf4S9SNmvnH5OMPRbfGzbC4R
NoXhoGK6AVU/FKF4Hrsts7JcHwixO++GACp3u3rTsU/qaBd72e64T4mUX8J/aM6x
o/YxkE1+d1RO5Mn0DYTHDrDv39mOzHTHrObEZGxdiQEY3QHBmBke9tlzZPlGkfAj
I5ukEVbllhEy8aiK3Pi9qIHuwuX+CB7CnUs2mqKMe7zzjHc+74wY/y5gph15Kr0J
8aU8DsP+xLLobop7xgGordFBL7Fpz7xG8FV1Frkk6VrRP2+9ae0nffavvFiK0rEB
wERWz9jMAYEO8zeNGqhGbIir4zWNkbGZsM+T8FWN2wjJAluw53+7cQMpgTF2wqjo
f7nuBGQTDJoMoETqmL01WyllQ1ySRQgATaV4SBGkQ8zMbzCSfCbkmmn1H383TkwK
738KxoI7tQPitkFvuLmImgc+VrT3xBU26RRm6v3JJOjU+ZKU4CC/a90TR0uAv2Wa
g8hvU4WLu8BLFm8i/cHIuYFbvjneJEVFyy29nmyxAN50Rh7tzW+IYhQog+LbIfjp
3dg/uvU4u5bwL7NP9jj6HJsf6bNIaODX3Hk7uem3fltk6JSkhQQBqOuGVsN1DRLw
6q5d425Peg9EAubYXmRfY0/Nwa5XQRBxKiQxCbme1s5H9PDL06Ds5WvTDIS+zyqY
LvuiSo1Abwoa3bUvzbskJosTdrzHy7l3nwl5mLkQDwmWRq724BcA98nMqUQttWIO
Og6pFgA1yAiRc1VjNrWGrkeXvbllKJv0Ha9TYqX/0AvQJybNz9IHQHHN2NwPkxfO
LrwXJYRkXTOc7PU1bbbiuxC9Wdv4LcGqEMbQsjOQqaim/zyM8DwBMd1Ce2Qr0/Cp
Tx2e9FLURhaReDMJmCCJZlPYgwnSFw5OMPEHggPqXFZYTZo4sl8CylXptm+FzeK6
FpLF9qX+ztiOxgWz5tqsbnoeNfewRofUH3In3/ArI7Gh2dX9M5wUOYFDyIwQhWev
hlW1amaeknB1I7QlGJtG+HudQJNeLS39a4HLUeg3jWlMY6bCV6/E+yLyfnU3Zy7i
xUTTcpcD5vIqWzZxJfAVaB4Y27lpeqieDKnmpi5GUJFmYmb+QIkjWNha2LCQ2SNj
QVuJLDriY0wIsgxbmnDPpeP17klGQ5DnxQzpFlX1mMxt9tkAFBOlgmQMea6T/vW1
DRly8UbJ8dfPnnlYtDFnCXRo1lGId7d1mVnw2U5/WxclJ2XrlfSxBCVCuU6fTSDL
ZjN0qQACqHCO2XouMwfZ6EfrdTfxjG3hUDmjHhOQa7WpamX3e66hChWiK/oFfNxj
b082EJuBHV8Z/n/DrIJmUqotopZkW81D1SKRgnTpLIzgVTj0DchS23xAc2iunw80
MHAuO7bpu8mih/ECRXpcm2eQJaV0dwo/H004HvHfVmC02iVB+/I2RfJUH08aOP8L
BR/AlZMtHfHm3Aod3FJbFPFh5ONKnIKiigbLKzV8aqMOh2Te2gbtpi16etAGsYKZ
M7hH7Tvp/LDdgrFj7wAVYkbE8C4RUIa+7Z8+MGn5oT7XkVfTDNSa4ewoqPyS5e0J
1yBC3PsGFxvqrOLU8kNa3V5jP8DSdlhkvZYMyc8FIKWEmhVye+9M5T1gChmkotoG
cH/ApKSJyte++TiwYquN6qb9OOYrAcff7yxAXo/ttOlh5HZnfRsmj5izx1jHB3SR
9UbbLPEiNuxd9af9x8PWWhkvRQSCa+Ddw0stIY4zZ0ZaoDZZiopSzWOHgv0dUdXT
rbOz+DF1rZTOxTN2TyPeITsCPgivFi4A5YcBJFvQKARN6OSfXIDcUaEXUxskuGAu
zMpZatvLwL/Ji39U0Sa69slbkc7TWeWvbroZFT4mV4X2QUi7CHa8y1siqWTObPPj
sH/IdhhUVu4zEUTBisHWnXxuWvV8gsxceEn0dJ+tVbcs2ukjyXfB+iQdvaDIUctZ
I3VN9PZZ0NQaxQXhf3j/r6rKvEN7ryXyFEB26SEWjTmp8dfJshLYmWAkZbEHbH9i
hWkAkXXJp7tDBH/9RtwReuySz68YN/VooY+4TY3MqQaismfqM2hCzBPng4Yd5Uph
sPBHN/TCNXVfrkefSK+RrajOApyAs81rq+Z0L8CmLPLBcEXXF6CC2KZWnTAD3r+E
4WPhpCRj5IqYsmpe5WkJwtVG/QWSU14DZ/mBEXHCLu1fH5g/nKMBb6oJvgv2qqZ/
JTMB7uCXGFB5jvWGnoHT/9hsSoWiMjeuZp+3g/4dkm6ol8KAZGerpL9HOnbiDwgb
YnHjf65J5pzxLyfAXComB8QJ5j83sgKO9o/cH0npS5B9/d1y3I7lUXrsV/Zv6Kz1
HpNg7QWuArOLCvPMEgcJ2nr0CSy5ZEW9LA6Kh+gD1cks664kOOkQ1/bTu8SROwkO
GSe0qeZaXqsKHkvTAuOjh9C2G0hG1YxfjH9/WKPpr5cx4hWOEA1QaVsfFK87RSjt
yIJWsdOn1Je9AsaixwcKmt732PuqrRR23xtyVlRzVTux008Zc93wzEYGYLDuU6bm
90vkDsBvEcwCbmdHLZcM6w6nN3ngD0d5G4WuEWiaVo++MB7hbtBW1I6CeO0izLR+
6TafEODP3ienZ6Wzf2PLXU1yF7T6qUl3kx2FQPpZJBzXasuNsozPUU9EqtsNQSX9
ue1HKiD+GVFgUQSob5ZYo5PCmbQrBO+iThFXJ2lwUx1qrpAFZCaDVNIgw09KaW1d
5xuKlywcBhgwAidvnCr/yo4KT8e8m53jq2cUouK+l82HFsve0ho0GPTgLnQEAh7k
1kDsXwc5vKAvyczc+8J2pPdqKpX0s6RUQG1jR+6x31OvfE2uUJaHmqXlsxS4OCY2
d2dyCh+ldtrpLdI+H7cAeiUT1uSEVa//xFYr6/kMWcbnGg982OqtAdkx+soFb41D
Fyq1fYmWIRHJ/xxjqn3BRg==
`protect end_protected