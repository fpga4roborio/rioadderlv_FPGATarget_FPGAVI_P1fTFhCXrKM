`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
ddtXksX2+yylW5zu6QL2Lhnb2d1sD00763mmSITNX595NcHTEkwn0zB1Dry37fOW
FufOhVzEJp80NC5qZ/+F0Vk7Ik02dIR0elf3clrjeJRK85K4e3Hoo4xn7YbFUIms
l/8VZSb14+JVGURjfswrIyCUotIzlzVYZ6gzoZwDXIi5gQIBf/gI+KxNXPaKV+PQ
Ufys/12rjO6aI/pPlqSm0hCvftmBcnezN2hk1UeXgOIuKZnogjOsf0iJVX2aOOWE
6pD/psybjbnsNB6kH5uFTA5frkzIzkzl5d9+YDm9OyC+k84E83I/7/j+rk4L2dah
QJOvksSIzN867/4Qt8qYTQ==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="MvBXkzurAa5VTw+1JJ70nePUfoQXBvZOku/SMmg4TwQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
oRtzZL4VJ4iwysPsC8SXYCzXS8Fw2gtZTOskLcDV+1B9Nzn1zTyNtlo6lNICRmmK
ZRVu2BmCc2G+fmzynYlNTnSa7C0Cuel6FYpxCBlOuk3OF2tzAmLAuDyOH3Z1Yjzk
a0aHuoCdIRKv7BrZCdALt03JeUmXKPdOmIlkVGFl8yw=
`protect rights_digest_method = "sha256"
`protect end_toolblock="Jn9CQpRhJt4rnzZPRk+dOpzAubz7omckX1MrFd4p81o="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 3168 )
`protect data_block
gD6l00tciPUa6pDNTk/+t0OO0nC/UTtBwLB41d4inuAUA3i/ALrNyoJVcBnAmEQW
ptbcNp5fxEUJjnOxnedyZEuEBxWRieZFQnkRdF269oOxgolMPoci72q6u4awUYGL
n0H6orGO/jyb0Lp0PfDZlPyHYa9s+mcTeUsjYLCmlS1IeVqgkKbwPiXhRo/iWo7m
RNaj9GhLPNPWPbU4ykC9GT/XCkQ7zgUR8hOW4a+br7QF/LT+BKDAw4f1BPHHu8ko
V1+bdMedsYw3KiUH8aI17s2rUDiQnnFrxmVFhKm/AUU+e2SSoySEcmFOhMlBMTCQ
GK/sXZP5pqblIzBmA1F/z+YEoPk3E5i1LqzBOU2SrngtNIKTfdhBuSOfZicoJpJ2
d2tFuD6u/tl9xteuGnHHf/zXNeSUsBUjQpWDxvgfM2ycAuOVF56Ut8hqA8Qaf6wb
XVIwu/ncndfTHM3Ld/fGVz6qSVl/LC5hdFUCMREDcbwxYg8SpIc4HeQA4EvMPn6k
5Z9kX5LS8iz8C7bKGcapYzL9i2QPIqJO6NwPjVlwWZNsanBNue3VSR6kEVdzdzUC
lDUDJeGVOPZoxGkc2jvZbnHGnpcEF0iSxAz+n3igFtkZFb7Vldw4HcYYgjiH4KKk
UPljd3yvqrFCTVWW6w3iyNDPIEbS147v7R49W7q3mMyhARe2jU2Rug/Jn+Vh0wAq
SsVM8Fv6NAYvKy1OjeQJEGVg/GxnEfO+Rh/Q3qV1ltR921OPgs9P0zLeCnn4x8uB
cCmoJwNL2HLMDQMh1G9e/CG156BKP4k4ZWek2veKj/3qgZ0arnBaHWljaOiEl/nJ
/3eZIGBdskm9HdA4e2lomkmbPGPRQ3hSgCj4kuCLRjylqGMSSq4adM6+g9jWwVCE
m+fLxZiuK9NthREFtZKR8m4Vpe6jVFBS146aM627a1xtfyv+Ftc7z4TyLbJAaROl
eMt4IcomQpR8GfcZbgPKpSrGo4wByG3D9efC0GYrrj8MN2N3pgPNB+yeoHHt1SoT
lMsh0qbFkAc7may/qTabrrRjmDktENZLDfUWKGRtig9Ixtso1Gb4bs2PYjy/dNMW
OTLEoZcLKJYBYdueGrUHmE0uwHCGi3qDnAk8adBJPX0H4ttnXdw7vP/DNhatoqOQ
ZUlHqZWZG9CEZseC4jpufWWKAuBQTzWpPEi0QcsdVAq8Ov9Qev2ktZeHD1e9+OCF
v+VBax4CNb2xzyWTkCNIbB3hzAuY51PDGB7afMQteyDNtQPg/A9c61ZtZW77QoZs
S1OIrP6kFR7Rv35EKVbabw2kmQRydbgRQT35FtFTMoNbVm9VH40Lcm/lDYPF2BtE
v191nayyTf1p7KWjT36JaBczZlT0wLXZr/i/1Ai8IUwM1J6uC5W7DX7KkRwez/iz
Il5naYJidAbOBzSNfYuTirg2ZqtEv+cOPSoeehgqeFYPbp/1bn6N7Nzqi21UtZTQ
irX0AjTQOviJmKbt68OjIkR5qb2CbX/2/5eoVeDsgN+/OaSXq8XEsadYjLujb2dJ
xTPAwCGVP7jLt6CAIgmM2X+rjr5vg5jYPj2T/c/5WeUVnRlVjuwIFkZUGHSxRdqw
O1qHf+KBVysY7IHgroMsk4ukDCt5/EBaqCXvOshwadCqkec6/9XXMCceMAOKQ1HV
yUajl7roLkvpLB4MAbPty3s4v61cXS0alejuBRkZq/TQDAtr3DE+2hDQlODs7lJ3
jL7I36vqdG7cL6a7FgmXoO/cgCQ1Sz17wfFijKFnrPkA6Yw52DB7j91wlVHRXyod
4BlNv61MVsrlVXWxJkAy5wP8Jmrz5AlLW7X4OmXRrNdFGPn9/8ExdhfOEqZCDhA5
bqRL1mh3iIAnDhwE5TR72SL6/FUyAcfpxjUWArjkPKdxGG6PQCx13ljvlOqE8TuJ
F9Ena9Ae1I8nwNeAB7lENSuWYWlMX+y0VA6rgkV6aJ9IC/TGAFoYLnMfLOO/duCH
ziwuMAHcAV9eLMc8aGAFdIgIFqPsxy+rMK/LDwEt6FprS05Syuz/H5gkAUH0vAIZ
IWUeq4ZYcdS/B4hFzHNraP8D4mMkG7x0SNAqvRUAtxuaoPFIxijgC0r3rgWaPpXG
92gONeKJqZ1TEjJdpcim/NMIx5kr531MC6jycqSug34hdtvk680Utq0OrK1Swttc
pVQzYccsL+tkHAyH7Q9e8ebxioXSgOrCY33nCGTaD3TQll9+aRcM5ZRbRC+WZyws
KhZ+tLnaLvUIUb9PO05tEiJGtIbtVzD+qxOijOFsSlaOv6svuRIc/A80XL4LEAh5
aN11ty+BaAmkW0upfIXpQVbEdz+EEFo8LVI8bFVAYA1HA9JzBQnGPvcTT0SDKjJT
7Njl3CgUXMijpbVjsZdha/Wucz6lJSsrpm8xJ7cooxIvxzcbovjT5x0tqv4uZaTf
MyGqqF1S9epapDfI590NRgH30DPBC7S4jiaSVmqOnaDSbjIvTOnK+KNbU4THpsbI
dWPFkvxcjxIsay+FKYs3d9Dlnyb6RRZtfw/Yrofl8U2fe97dr9b/7dKHtC8HkJcH
wbPvdwOqilOOP4OpPzohMiYIm4eDE6sBcIfhjwtnxDUpfIOk9Li7sUh4Gy4p+G+e
lB/yqO3LOJNN4R1adI1B7BjDEXrrvj0Q9Cj45MvNwT7ev4kMdvpxB29nki9fjxK+
Is9CB4QqrtfhaChh6Nrnd8cyJZ82P6CGiMR+oTueND7YNQ2Cusa2qqMnfsQMbWGP
yDhNwnVnwCWaVE7ezn7Azp6Ek9VSN2EX9wjzfLc6eNMhbuVyizvbH6S9ok3Shb3y
/Ee2QdTSaetnUnxcunS4ayPs7DNjz2hlLvCV2AYIJ9XsQtQkayuUMEcZJxNVOcWD
78uZ2t6ABdWS958voypGSYKFB8ec1gxwW1yMHdLeGIJirgofRFgmqVy3NhSqZkUo
qj1iHVnHGDGcwKYDGX8XMtfo+hGTvGPGPSakiQvFJ1gZ4utjfY+A4GSyPV+0figj
qk9oR45z8x2Vh7B/7ykp2wRANepoqc8Ikxyn4fCGHDSJEANZnv2rIxabQ85Ivt53
iWuwZfUvVAw1SpHBCTcGKKPbMEo+VucKlZ8nNlJYRaN4pdCB728Bl38sVLRZJXD7
2GPbmPhIAkbkInEHIJ2gm+nXVljqgOHYJ/1osbtAhAiTpUvqGlqGRSkKY7hsu2YR
4s5bz81KQAthVbL9sn2NOOHoLVj8GrvY09tKE/oGHF4aKQrhdwbUUqkt126g5Kuw
uatweoLHK1fGad9hjb0Efzqczk8Q9OjksS2WXorpF1TK588ZHGIHmLF5951vSyna
41BzvixgMOeC4MCT8/bL0IPFdheQ3vdjrdH6Y1jUX13rAbX/dErxLXd+lpaiCvDf
REwBuwH2siMFn24wVVJkLSF1fwxoGXvukNe3bsnUiOam/KPUm5kC1LTWGbOT1VoV
ArWcIPrff82BXqOIhupXXyiCPw0cwLQVE0/HxmztrmtdiRuqkJLdqizVooii+f2E
0+R129pcbwyMGu0LNm/T/ivZ4sx8185UCbptBnUHg25wPgh8GKYeVfXsFy9FQv7q
Fc10cpY0otFAIH/9ToqTFPLBFYfDdY50tRn63w+vwPVxfzN3T++QdEMn+HouiNCg
Os9lqYvpmLDI/dBOuedoPSIw4NDSDcf0ZWlUS6p9Bk8/aXlJlNGXHGZI+APLh27y
S+gxJXJe5vRVbNO7joPrRdOQpMJe4gPIo5BKoiZUXm4kjVYBBoV9lsDa/yYd7SL3
67KqceRgdFjXiXURJy7cyFGpgji/JDxUX11hzDTUCMIVmxSAA74gV+64DWun1LLr
N84bELWmCjMsgDeJyKP8Qc3uTxPLz0vHd3uTkZBvLufiUpiuQN20Ex+/1Ify1Poi
OHTD7yTCx5OcdDOF/qaWruGn9PMr8iv4GEjncAGzxCaNYZ5OihbsJJcBGh1wPgF5
pD3OW62ORzc5sREorB/fVEyvRUmUOr6yZ0Jbf0aUxGJJu6EAmgIVtGi51oVaqKtE
ZH3hotJOCojHsHRmLT5sMi317FPymOgKz07V4Lmt1P0GJjilhZn0cwCez2UZ1KBV
j3YYds+2ygzqz7fPuMsGB10mwYC9mnsaqoPzeX2/2V/kTrzwO0lw8K7Kw5S6acPZ
aNFXyjWK/i8BPJduLGER1jxYWt2mIjWB6jmMI2tIm701n5S+6nbb6IZfmgL7VszL
`protect end_protected