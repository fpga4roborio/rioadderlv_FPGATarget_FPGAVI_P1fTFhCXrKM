`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
ddtXksX2+yylW5zu6QL2Lhnb2d1sD00763mmSITNX595NcHTEkwn0zB1Dry37fOW
FufOhVzEJp80NC5qZ/+F0Vk7Ik02dIR0elf3clrjeJRK85K4e3Hoo4xn7YbFUIms
l/8VZSb14+JVGURjfswrIyCUotIzlzVYZ6gzoZwDXIi5gQIBf/gI+KxNXPaKV+PQ
Ufys/12rjO6aI/pPlqSm0hCvftmBcnezN2hk1UeXgOIuKZnogjOsf0iJVX2aOOWE
6pD/psybjbnsNB6kH5uFTA5frkzIzkzl5d9+YDm9OyC+k84E83I/7/j+rk4L2dah
QJOvksSIzN867/4Qt8qYTQ==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="MvBXkzurAa5VTw+1JJ70nePUfoQXBvZOku/SMmg4TwQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
oRtzZL4VJ4iwysPsC8SXYCzXS8Fw2gtZTOskLcDV+1B9Nzn1zTyNtlo6lNICRmmK
ZRVu2BmCc2G+fmzynYlNTnSa7C0Cuel6FYpxCBlOuk3OF2tzAmLAuDyOH3Z1Yjzk
a0aHuoCdIRKv7BrZCdALt03JeUmXKPdOmIlkVGFl8yw=
`protect rights_digest_method = "sha256"
`protect end_toolblock="Jn9CQpRhJt4rnzZPRk+dOpzAubz7omckX1MrFd4p81o="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 17344 )
`protect data_block
gD6l00tciPUa6pDNTk/+t0OO0nC/UTtBwLB41d4inuAUA3i/ALrNyoJVcBnAmEQW
ptbcNp5fxEUJjnOxnedyZEuEBxWRieZFQnkRdF269oMl7QqQ5HVhBtoCiVOuXo7l
aV4HvC1BsicmkVrjn7GYt75+IKVzAJlbwjhoc7sYxZ+Jgy2bvfJyIKkLnrUauo9g
EI9eJQFr81grkmE+khlx8Gisdb7oEmUJEQ+TU253WBNWDv55NYKqFaU7aiL4SGdH
Pi8xDcrZWkVuF7FZXqpJ07z6JGQOuLmvVehxLrr9u7CpH3cByvXicmrAdeaA2V2k
M2qo5NGlViDcDjjily4sexJuJbtYXFrGA42cNOY6/vBdLgCk2UB8C2e2UR66CkNy
ngWFGd9C1FpY2Pe+LugiAQghIimlS6p/wRwzpuVK5eyl4b9I60hTDTHHR0gqZI8r
qDHIXX1tdCEskX3EP9vMFU9O+bRcSZiFwxsSSCwKgUa38+Bg15wfY6uKNqvx3nOG
uWwd0SznEixKOBON9ZBBledowroGsRQLFbCnrM9zrjfBrgAYk0ZKVU836HBlzJ/0
1+bKX6q2a25WjAsfnOIrDt6uobJMk1OXMD8NquGqD04gPLXRRpifdMRPVgpduUFC
PbTL8SEiHV42CLZP/qIy5eFjIxJZzXphtpiSFnZEsvV4ipZUmQJ5EeOOSchh0juB
mFfGE1/1zzxmGNVguXSuiz4zlU25cTszreze+CFiwRRCQaOTwO0nnU+0FJSrBmB9
Sw8gPfuAmF1P1aBFfDD/5/2rFCJ/+1pfKDyBOWPyYFWhukUpPz7xTSUtK9P6Mctl
VTh8rFaYaEti7/Bh6QdtKWbqkEtU/heSNP3iuDM6mkoLzdIYAv1sDcC/IY/orkyA
LTFFtzFLW5bVOiIo4T2jJ6jJapRJOMcM+f8qSS8yFScGD5jN+b5dlciJ4FzbDudE
Z8s60J3P0gOR60JYC83XXz9sLl3u4kwdX5nNBg6avYRPja3F7wybTONmBsZjBIb/
WCKiGEhecUuH4S2pgj3arHUUa9zOzWHdrzS/un9ZMkffckCJHYu1NF3+IKgR+QZT
GK7fArMJWwnj3HmcCy82/19cUGIRVMtiIxHqpPL5nqYgCO1al7WYS/Ov8ZxcwTtW
SiorH0z6jee3NvfKYHxX3CKwXTgpzzjhwvJT92ll7CSiB8F8Iw1iYp/3UTxYQMoQ
P+YB8wALleXOowENJidkNFaYXwzSu/i3ceTvhTssWAtUypj4oUSaF2WgRKyO608T
hr+2dKUgBlrh5nKJIEETbaNPxwghNGbsd4GSXiodrgSQHlSHjBvNWXXIaS7YBpNo
L+vdkQIoTPYOIVghQnI7pS7tV+3EGvEQGeqdtUM+TIXWA3D9WCw7f4b1xS6oGXIJ
P1Qaw8g2y89/wjb0pNgDBBoZ//H6XjIEcJfQXmeRXqmfkP0pUtJ0KXrWQsay6gvP
N590D7oIFAYxABYFR3NEI95hC5Lc4Q3KTKlplhVbK/pvQ+deO3V3BvqP30R+xamA
oxyx0Ub8vJWfUYWSDaRCf8V80EdsZXeWpi+6+ieIqUwG5vdTy6RAz/CZv5gU78on
StdA//8i3NSGT/LL6OTKNAidauYqYzeh4i6U4jV8KZf0hYPBlyWZjirScZhsBypv
YQQ1qXCGstkwtyFCwjxbhJExkexhK27S8FJlUCcJwM329ZWj55V2kFa6D0plvn+/
mbQ20kw4/28zY7BmOzA3hsbaq2WZZYubSZcsF0vBGI4Vo6MfwCA9U1axmQtJQu8V
X3mlqqCGeLJmMB/D0U86frBaT3D0tRzFD4d080fmG2fc2B+JJWgt83KUFzetoc4l
jENfL320YL00+dJNpmje0bkd8fJn//Jf6syVV3um5bXL2kehJbtpg5MBV+vbkphf
W+4UrQgJG+zon3gc8ytHutzExweEPIlkszOFLLT0pVlWnqMTCCcEmOhqin9wpi/O
+CmlaZPVhAxSSXWAlPAMH+TZ1wmDnN28u3HoFN2S16xE/hTq2+IwhRtlvNt1zTwJ
SQ0BGsqXWVPj2v5BImWyU5jXgxQTY/WeuUYHZJ08kvmTmHckt4wWqZsMrRNJezrL
xvA2NH2UCmzzuVxUX5YQ2IutV2k/43lisyRdcqhZpjAzBHhLgqGlndHjIyiMixYv
kIhH+f2Fmaykwy9Snu54GPYTSiknIL+Ys/IgDbfoLusP9iLK32OzErIsA+hsXGkB
Td0G0YtxHbf2X6PPFPfJP1L4+Zb2ieErLK/TNxCkwlHs2G0q9YkrNvIVu/NlBLev
t1AZFby9v2N65YQuzhbzPCSQPwYyaEybDIh12LbEmPUiQVtD36Ztjx/S5WiaXtYT
fPPWXh5rrUlrfdKSTeFGavHl1mJuoUn79NIdQA32vnCFuSjJJeXUO3YqiXv/2tCo
PqIROQeSbR5k3aEgBAYR4FHDTssgqSvMiJC1lACv3Y9sTGlbFg5iiCRkrso2e6O6
oNimMQj+MuJp4TR6Vn/fIzDRWCuyLNnkyNIDnFzYfF3Ma6RpPzvhTOgvRdEvXQ3t
HSDHCAxEvY8MgHI/Zsw2Cgp7JPsABXAcFLtOHafwm83lgiWkHyqv7HsFiktuxT67
UjN6pnq81HWS7fEh+1b+IxjafJO/u7NP0GpkwZodIm06KtFH8/pAFy5V7Fz/aVaJ
mXrzmoi00Fms3WoKo7H4RvaKGSww9NMNdDBCjg/9UTy8mWfLqXN82FLyhtheEBhb
U3REUVPzO1LRtbgO7VKVVw02DFeDjjvIZiwqTpZp/BVqh4TwQL+dwA2PEK8LoxdO
Xk9we1rXAjdvuggTdnz6rTv+MnPD/dthDRY41evhnA4S16+QI+licj9l24Fk6PC6
g3H1EKuLd9HMZIrhyx16Uv7G9pW6EzNbAYfUw5mi8mYWrqY8Gh7DsnPbfbezx7SP
xpB8MSO4feXzVi5oyO2suDe9HXmg2XaOhdu5l9V6DAl1iedb3UnmWDmrjJubZOiL
FQ9JylBbYdILLuUuchdFh9D87plDscklaClBMpvss1mJlhjf8FEraelor1xjXWQJ
VNCwVSOjATfwNBUD17WFIWu8PFYiSsJ8Wvi7fuzdfbtHkmBgbCwkDr0GBfG7iwGD
xvdWzbW7WZMnpQ5G7pUGAbDxtpHeBXywCzdC9VQVXVXLd6PV5NU2qFmrd2bErhPw
aCgN1pTLZy9jjI+PCs8Na6PH+PLq1E9r1ghVkII13/QaxXVr9CFrMIH1b6n8yU9d
jDZSc+QIT7QjGZycRRSs6ifthZW7DQn744r7PF7/RzzWoVOdzNvM/IW2rHPvzzRt
OKxtbkpY+j+emSkVlap7JIYat56eWFPk3s4CM8dhhupQ2D6jcwTeYkFEUiSO1VXS
efGSVH5QaWtQsd62b116h4je9TlVWj1zrAQWY+twIDDTBymfHBslfA6JELh8Tzn0
h6LhSLMyqELPsuy807L1bsC9EfMoFX4+Ye8QB+YYTr/w5CeHvtjHDTCKI2/ZLB+V
52HITxA/GG216oaBEY8oxgntfm87CvTbnSaIb/QebhqzUlNh/bUotbfaTaWKU9ZR
e+QPsShbCVJW8azmvafKFdE9rcyqJb6m7UKarUH02i6HH/WnxEqt0MuH69X5QRVS
Mqclil8Mpt00/YBtTbXWhw3IaEI/7qjNEyAOHBso3fT7VGO2SJ/B9wUF7aRWSrhp
hqS0vPFV405TqbMU1TG7vRLmvtzzjrP1VKspKDsQA+VZyVmkJdqj59stBSkkvEZT
wtJtxK7Cb8T2uGqWmoA9lEvvNv6f4ExNIW0ceB7fFLVBspLiAkT14WulHnpRj9qG
nIEk5V2Wj/TGtrN7GJ6T9chxAM3zZDOzlr4qdz32XaA4r+6SiUxKJyVS7GmFBRBr
WL0v6tESxHNeHRIUZjFqWW6s1LVRJA1Pfyz2Mt5c9sQ15m1RmBGyxhOUbYnXsmBJ
OWg3qa3n8NEPMWq4VKkXrRBKWFdDapUCyid4RcnPFHXe0Fbm8zS4BCa8GBDkPpar
VzSvtuH4Tijpc8C7TOlE5unT0DVRgFMLpk5BymazbDp8f9rVmPwYSTsisjaMr4oE
/RjIDMJJLC9exKXczTa/Pj2kes+1D327MwxApAOmO/JxjOnvc2wC7grZqyuKRzUK
+FHJfiyAhLBhly3XSj1cmSO7NVFj6jceGYJ4qxn1Hm6n6+5ktGn9pJU/PJbfFP7V
3NbXyOLbTZYRXN1Ma4ppJi23jcFKkI0tMZGJurfZLTP8LBjv3Hop0MRgxlJYZmaJ
Y9tCHaARrjwc/pYKwPeTnvVROSawVCC5ttM0MVzjoz+8inVQbwtjNW4mYv9pMIZ8
BAAPUyN2HOPVTMwhwxaFdyFV28wC80p0xDuyA3Bav8rkNnklIZOefBvbtqj66kn/
OiiFW0LImPTLv340wJcbcMgBAqiA3vJIRYAMc6VZIFDEBSvdprPW/pcp1v0MdX2X
W0Pbks4GwhdRpy0X8ekXGHrlefeps7iykdOPUimpsDY71Db4SlElpAzCMg/YMA2H
3XwJk6BFdR430ZPYrknyD4HDrfU6G75FH6//3s16Ok9nmBr1OR19unTKrxgtRJ/a
6xttswUWPAGnkYN0LJh8gj0AdU7FZHQTR1XLeHw7wuvph5fHMY2adTYLn7nNtGfq
8qh5MeH0gTC5kT+R41Mi9dGeBkUW2g5GHq5OSNN4nVL3wiYELr41b6rEkPawlU2E
A9lxxlY+cRbuzyM/e2XqcIduGhfrfvOiywBBn4wGDI7UW2tCmml7j61bpBX6VweL
aRDXzryCWYkCG0bCqh2dw+gSkhCobmzyOAqVWBFKC+vIV0anW9OdaEfH9UDZQ7YB
han/JD2GSKJkcJ5mB6nXv02qdirkh5j6CZXKdm8xrrFNSP/mX5MdPfyj8gtE3o9G
R1JlemGeREYXlfsnIsZcS9NRoXHBjp61KpujeSgx50lzy6DmgPAXXbI8MPpT3sIV
unz6w/EmVxPSeUWrWSDQHmxENnlpwu3TEL9a8woRDOFfUM7+93v/y4Uhc6airbym
rEvje01v4Q/gdYUIyI+FwVIrkskQ9lq1+ZXN4eVLqvDaMpU5LZ++AV4SdrVEwGTV
7jdg70RjIJUl29NDPkVqKPpa4tu8S3/zTmfxnVjDudw9dtNkQIzpgh+/vq+3p3G0
5Q2KYO39G/7AAmtj4A3Znkuitfh9TOYdYFBf55EDOQoCwYHM7EZjp9pjqN5KAYEL
fGqStUL8jszhFX88hrz869eU+Pwl+hTEgl9KFfpHQNVRKCw49lp7L8usIYbri1cK
o20QLV6hsOjnsBCoKYx+p7ETwbBl8+CHKjs+qtd/S4YVP2aPsbFWPa9AclUPaTqV
6/r86RAkW+51qkZzmJ13j4sOrkuywXQEjvkVZvwbq+dUCUZTEjCfs/smi44ao4Bc
QBtRN0XKr0iVQX8TPvK6yjMwQ/DVZOEbhsoAJUwunmqVK0macVpRE4dCKVHuYEsa
RiNg+yfwjs1YbbVCp0YgI48bmLqcntdNNnhK9ioSXClzsR4Eg2dlln0l3QVxLRnV
gjr8gimO3TEy6CybHKcij9q+CHcI5IDCdtgJnO0xBKWYKp4cb5mTgn5fJL2Q2QpK
pJW8CXfBYNDu+qghdsKg6+mcZFhBWOv9BgQJ2LJTmPYm9X8jd04ty21NWnbvuDrz
xZ9llFGFOEiF9Q5EkSbx+BMxQe9DWSKSb6UKxsICEUy9DgZAMr1ov2dAcLmktvjl
nh1HfmIPJrCjvqs7suP31kfObeg1Jx1tp/TrD4LtCT4VB5nRGEd35PiGIqsiIAtC
roqApKjKT+TZdpUisoEexzYe+nj87g4kVnOzhx4xtd5ajZE45OlaCFODPK2P+j3f
m7ifEAQVcaNaY4AZA10IyrqLr5FiXB+FF4nFpIYbW6CuLf7QVafaOzrR5VcxesR3
vadbhEAGLYsDzX0hCccVZV4BUsR6dS77GUos37nGdOse7xs8YGOHRuNgcGuw79YO
f726j7BJ/Df/b6FYBnXjd4a35LhMEqkih3r+2z3JEsMo3eYXr+nCuTjYxb85/NaI
HvziEkMmUd4duclZyXO7TUz+boZX4KLCHZ38CUxNd/y3D8qNRPhxOCBnU25B60QN
+NQaWhDQRndN2TBFL10XkB6gpf7rWPM1gRxMYDZK5MpNBKAErHyLJIOe4kG91Vi0
wO2ZN59E7NKHG/L1k1NKy1ExadyYEChNe3916Me7cR0VIuc84H9KqFcf2OST1dVu
0gDqGz/ZdXJyMka9qLqvmsjhAQ47FTNWBbZIFavV04hWF/n6XCRP/Na9gq2ti1Pr
8bL7lc4Yt6bI/42VBYqxRLa11nYB3Fbx/4httfLWbz5Ycww+oxUCz9bpAHcJAi5/
xlVgaenWb8rkowBodCGYqAkuapgZ11sL1C+Yba+NJgJv3KWgE0Dr767e8rCHR4aL
6x2CtoYRj295WAVK9uy3EQn3GrysToynwtG879/FqGKm6Gj5/ZvwDebfxG8ElAQF
1fvApWoDRer0jIT9tOzryAmsqoGLxxitVDMotwYdL4TNh0sON1W0XuLw1xJJn9Mw
nKFmcNArvuc+PdeXH3AnK6W2410X1V1Xu0kAKiPVQTtkJmcO7T2sEXqbBlMvKK2Q
p2JMpJkTvDGlL/9FWJWDGtl1AwQaqZm3OGv9eT+S5SftNd93tZjq6MW/FwrjVVL4
/rtwIsmlqQSivYcVo3xrK6UjuNiRN2Fk1mt6rs2eCtP6r92QZGg4/t5jkIulFm1i
8USLXnnbYcyDJRQo0b9X0GmaQw5uF+0HyoNRWp7J3vKiDaTz1jFMGYfljNUKg9w0
Bor2Y2AwBrc+yunNoE7/q2vXFiwpSLzzOpVEmwMUG3cPNpMGVwTf7lC179mIT1bG
tm101W61xBe5dZEbA6DPeQ8pHsgR1ucH4vRwrrSD6aMMtBiJaVxMHD/+SKudd9wu
hHQa8GdOdKWnTSN0Yc26nP5vkOovwvCkK22hmlP8rELvYw9QeHxFVpQMwz5Y0juZ
TWqmY7r2VWyCYLJ3Oyo1+refSWcUubSzq+9bjSeCfEnMO4j+BA3x9oC7md+LPvu9
aNVlImpedQOU53LVafVKp6ey60SquYj1+wvdfw6ueuxgioIQvF7kLHlRFIuBgdpv
yf0D/TKAB2uW3SB0uOB1CoLqtTc80FdQc68YH6Q1GV67bDDfJQAmHhXq0NkSekE1
SQ6S3UmTLGuQkwn3nicLlw7qAU5PWhszTaWRxDjhJV+/cFw4Y/Zg78zerDKb0jDs
qtag/HCxbGRqWgqmSS26UCbkZ4McQpxkjj3n6oOEfNePAuWG3jXvniBsVbmWBO0M
4v2xd+jhtGg51KinCYbLVPbBWMSmRIFdgDjkd9IDib1FrKuu4QaJoSQPecJRP2LT
WhyyRFGnZEl2eQ00QcS0tLVrAIgH0tdC9qnTuV6nj2S/CJsV0hMyIU65OZcY8MtI
cjd6OotVaFwUr/vAxdorWFjoZIDipf74O9Y8VEzby/3a1oCymBopLKh9oHxTGPgD
53UlcDRFePSFCi/EGGWxrzGJPqZj+WR2hIxesSZYphHfZ75J5vOXSKrUwGxPww3D
m5aDo6/HI2l1MV1xgGgyuPtYymMgWQGZG2aYH2mxuCE2x88Jb2k2sR5z8eS8Mgec
vdgi0no61RrnShlJFk1Kxb6eoSwCpR6UbMnk5SjcaDaYQssIsbUIswImW+GUqccQ
7ez+D/chymavEcQscNYCBX3EWEOtlpS4LRACR7B/G522kNOJ2JnkYYU2SHN2Zi4h
R56pD27VvaVaV7CxrI6iFp6296R0zPmsthO1UXYi8fJoxgVg5Su0RX20Lk5zvBAp
si3eZoJWlXkHPB1Hj0ArIAmt5tHsR298OCiHDMK3J5SUqz6CwXgNWDuxEiVbYmiu
4Ld/WQt1f3hLbOhtIuODiNsia4IpKgmjBJfszSvumZW1z6MkiebLvZJi52K4P2WH
gzHDFBKocRLRJkhqkpPgkvMfBRyjuXAuxPj5E51thBFC6fxgX7ZTBeKQ9taj/aGo
OLChtSdUDwOgXk31nYdlEmsj0y8ITjJObSG5GDdOmQWeyfKSsUCqyX31qhIMVMSU
wT9gyVXhkSDkZO/Qnd1dp5849KTQycIKB457Ni7N/CBgqXDpWId/6rXuwDGS2bEy
eC4huGVr8gEDQLFy4ZZ4ws41JXitujfc+7WbIJOzGrIXrMj4wf/hrSa+sUYtB25r
pcQB4R3MNvcGDZOjvwVJ/9YoZnw6Tdf9G89PFnEAGjwJCVfJe+OJi+bFJPo+WT2X
SVbit2pnC9+kixjVYIVyDIUuxVFcAtwkgnMr7OW71/z882BA7LBbZaExsFRW6NWo
MENwpcrlsKsrIYzdk0RSbdVNuHHXpW/UGKrYOvln6rl8Ywqhb+49o64CpQFwfyBg
ZL+pTlq61Ieu7/4Mjy7criy8GdZOKaNH9HZB7mJHtuMcR2fYspdWm2UyF7zcCpRG
5spZRSWzJxkagTC4ZKWDvXEX9+1z9ZOSOFYxQhVpfPvoAdcOnpyVyXYKSxECcmgd
jtKXsnN62Uyf5hW2tlRyCxzjOETuMrYFYYAfIT/IFAMC7ZX4jweyoPHTZ8xUFNS+
geNVZcbSKjijXQDkia/nlvPdbKB9yXaxDRfkW8LuY5D7V0OWYfmPESs/ViKubzBA
Hngm0zDm0V1ePriHNAFgg9MlW3rc7SRZZPu9QNTEng6K+x2bwxJXwr/1R4hQje0+
/xEzczeqiSvBOIJvymRFSGn943K8RjELxQvW7Da5DPWwaGCJzhl/eYsqYga2urel
zrURDKix7C/BJXLzHPER5C/T2+PQO6TRdYeO+Euc2uk5AD4wS2jEJQ82wuA4X283
4jjnl5OUjh4Kuaf64eP7P+iFvJRlBKL49Ul7PY2Wte6cY8y9gzN05xqihuj9EIuF
FoJd4h87YSFjC8YZ396cdR/f5uyhhcCtj1DVHn1Y/OOzaOPx0v6REEJS33NvyOBt
KBHjXpg3uws/zlNrtNMiRjgUENweW43lT2nJ+lOopJMaeZtXL9PCHS3jvX/X7/qD
EJBAOVJi4TeESHZQYytlY2jaigbt6J7GTEPfOm69HgCDM4qnLDC9AMmtD+7KdDr0
yc+8XyaEpeFBtS8N3o8Ugv8sFuvyfXuXOs7fZJE3rpdWFXzCFy7LNv3HYq5U/+jd
09dqe4EMNC2xFmNf8l99jtjl7VXMFcdbO/d0lb9TKHfGjn3xOBcdj3hM/Wo9kSzn
x0+dJq4zIKlChb92j+nI5hYfP0bxpcs7inFkU0HSB9cmMsMD+KYDLXI/NkcfQmql
5nUIpX05BCfwKOTywVYq4Cq+GeR+EPUl5cKS41WCh5Y+RY2gm80O5riqRD3CqHd0
XsaJxffU1XdaH2LLH1OADt/IR1Ss+WsBJRe4FB21q2qMhR4MuI+fkUYfFtnjk8OC
AsPO/hIH6NkSP0g/zBDRHgn/GfG5sNarzTsm49uS8Fikr5OSI60yAg9AF9Wd9DGD
DpZUMoX5+CTGeXkx+fX0WjkbkElA4P8vp4HUgjOezEMp9wjtb2YndX+umUArF9PJ
6cXmufC1zC0IGdu72YSYkG4w9Rl0dWd1QhOzmkXnkYN4WOGdGT2YAj5ISYHxo1Lu
NUi8bDhYkDTpQmp2FYWeZWWMQYtjBFVElpRW2OdW5vBWqdB/LJVX5ZeDW7y249eT
IhNr9n39Hqe9igrz+1EuQDIPW8803EXjg/OH0Cf3W1g1fWkpmYqHzhxXcO+vE7xS
oYjlTP01cyfk/E49ho3yzmUFYWf8oyF6u/4vF16AyGSuKS2zg/oaf0GR7/Qx4n8q
z7P2nlQCZfX6aRZifWKauFchOVVTE9GpQTCzijcMPyNRFifURPT2DOjBHWgNaozz
l7JtMOau42a7TOlVwLd7wDWA7mQ7zdkWavJtXulXabtjhmq3QqesRRP5xR2tgKQr
BGfWJU8s9kjvRf18rzdFGUUwnVOsKqrgxTaIabRJAYglVNuUIGRC4lkSO+tmzViD
pKDtDs+JL/a/OtrlrYqg0Uq2Ku0Mmnu5lhW8sItb8VIBj8EmG+XhsTzjw39my3s1
cMdhpN0zZITyczTgPRfW2UHZMt+F3DfvUC0Jzq8gtThU1iqoNVceTBtjUualr0Gx
qVcFaViXUoCHMOoAnCgV2zMjm6ZIfHHJtKwzNYJ9Hx2Avv/mUis/LMaEv+YOEc8B
FFPGbdDh+IubA4N+/ixXyRMQVp7u2C8jlx9gtggjst9i+XGCVTwOCrg+n/y9ejAT
37xmPsDnXsIjSrUS+JLkmDIVvIUpCYRN4M9yNAtlhkBfcjShWC5WO28ghphpEUgQ
sSXND8x4XVMzZ7iO7M1e+IV+Vydhjnah75PK99Ph2RL1bA1on3HLtmiozKj15+XU
N08nE/r8Ip4D0/LHVJndhojml3aW5i9Y5yOPQk9RgjEwz6lZLEJUMHkRNtTrc0ZR
TdSe+og3YbXP4qf+q1iR5zksO6F2NfJqTjho7UGWJrNwVXvDo4Wb3coDfleughOA
rNNCxVY5g0kL7hUMNlK9MyWltEiTwjOOLJ6AonzCAlq/LOd7voyknKhcVndYdAPS
zeMBAJg9vUdK6NwMlxJ0ilNzSMKuWzCrLm432TTga3wDtEXb3Fx0mJAIOu/81Yxk
cTKR0c2WYpk1hD+g3vGd/w/P7Jm1FglP6TQUZ3aP9Ui9HHgcNcimmtBpNWrAEW9u
i/ick+PPKW6JLczlgfoMnaGDRcLf/1GtpHP3Ac6x1k99LXWRo/Xkcijzwknn/RoB
qxGF5+0QRo/IQzLO6G/qIa93iKgaI9c5Ognj/7OCrqCBtx1Ws7sRXdbblYJ7MiLB
74yI/kUtopT3tc7JDMyqWw8KZ172zVaI12uyAL1+TwPv2b84myHIO2eF3Mr5BxVX
KNmGQ5weZigYsl/jPUshYpBlH4kX01+58mc0TDqZMM9dj6PEUet4PTrH7nOak8Ca
zfha6iX/BhRMSWDev3cKCdZmnEzpYS9i3hcUcym9RSPwyXFFaKeP0Du+T0jr49BU
PGqKNKlAnWwMXvWpWAPU2Ed8jEVkJ4DWoaDxadW2UXDyYo0zDJrhFqBfoRHbQDQA
UiUAv8A6j+AkDVPm8mPmc72NgPi82SU8+VQPNOMwB07Nqlj96cDAOJD5v7Dn6y59
W5+UGXkpvPy6C4V9uwIaVWpnGblGdSnitTM/47JKtp2BHXHv3hIE+2BJjt0kjq11
2j+P7AT6C71xFCKN7P/s2P3hPwTGKPhJytjpxPh9XXa7GFNWhlzvL/L6Hgy0wkGM
rGrIAuJSkT+2szlR8Hr5oITriPycIoyM2M1FbmfXu5XKoTP8XAu4azC1DuJ48hKL
xca/vuA1b/m1x0Thu80P0lUqEJtQzZ985SSNpRbKO5aMghgLPVqIHEKkhPapNuy6
crYkcRnY97yTcBBeHNvP/70lnOTmAANZ51nZK2SMG1g9H/Jo4/Bg+kAyosrZTMdY
Yp2bIJH/OzSyebF9PaMME/GN+aB6M6jKb3Dv70g2V2JrEow4qdFnq/6PeeBZ0ukz
mUc2WOCqM1SP5w+hfzWxqgThuBVTtKZQSFeVOUSdKQs7XA4yLpvv2awy/tu/X4NN
vdB9clF3iukk4uGRN8wVHLTG8dghNxGcx7qpBPRl6sa6vUm//RQqk3NcISHVQ1Nd
0A9q1vM4XvFMS9qW6YxyhrUt+J/bLG9Wkh6HUc5dcGcm9NAbVyMoLoDjl36yp/55
QWe/cglNYzpVFlQUqY//WGxqDBQXtbGN9Fqdzz0SKApM2CLohldxYKLxJWRhpnnz
KXYBfY4IavqyuGBgrdFziJEiwnpy0UIetpNzN0K9VgmCspI4xFCwajWkYAb3nq7A
3cHMAqy+psNiIExNGg/7kqOayafotfrFmzg7DOkQ6vAU/rpnSHKZ+yJqDwBkXZ9Z
k+vaEkN567MKUjOKRp3Ij15w5OVx2Km28NY6ikJk0G4raNTTrqb5gLq0C1lu5XCA
Pj05VT6oM2CyRPpfd3dhlbiWppJPDsNg6MSqC82t0Bcg6q0tWlV4DyTjQen/w1YH
+dJnQkgVp4c6EF4kOdXVhF9vd0tynIZh1th6xS5FnVg3bSyMzsVg6rU0mS8CVNnS
4IuKSZ0/Zy5qSPBgwsKr52E4Uoc/2xYxWugEgdnMJuXzrMPhsGdJy72i4uRqcHTD
LpkDVuDeGQakC+7u2Cda6JWXxK951bpOrP1ub/SXkRujm95KI/6dTJEi+U70TWkc
qARkKf88HKR7m93Uq3qDN8f8WzOYLxcK7/nq89WOvy85TK/SC9daew1SZ5bKwy1m
M7eNoBsJfuS2FQLKjbYkxqBXbMEMJ0d12uC8dDAmsZNcZ6QXYiKwj7pBvSWWxy2I
kTGHCiOegnBJj/chdLc3Bj6/u55GfAXLRBld5/fRr2bzO24/he2LEhF21kRlyjDV
N2IN0SRoMakBSV4YDYgTOdDAcwNR/i3i2ZL1D5NOMloHNDJzvEWhb2GDUDKPinYk
yL+lIb25wa/GX2tg2xztIEieQscsef86uZIcDGohLAk67qpJDw0lg70pEANuQQEs
AjDHXztQk8wxbenmekvUvDsCncfeoeUxcB+AcUDgAHmAaZk1eRZ/laf+cm/9ccaS
WjljsFUor5dupfiL2QGP2D5eEBh9dSpu3p7AXfqiYjtd1a+jOHLePjL5LM8W7Bw1
3Hq8Lwr/Z52IkXzm5XN9JjHITO8RwVisBrhWoXFw9MiK/hh2c7gaCy9EvhXV1/7N
7vl59nrxLF5NkufJ7cSq31XjSUfewdZ3/iJi8U1BH1hD2VhYQgJaCwEU85uGZEoW
kjRXHj/DJrMd/CUOhYyCwvTPVwW6CuhRIjeVlqRe1bIGqD8YK3hncKAIKEWyNeR9
rLLR+L/jgvT5q+hjckVDDHhJdi4ik6ORbfDhtsQKpxcWKt9CVyk5t9vNNxsYhVnX
RWO8P5BUJUQPDdzc7tzW50JCV1RcsWCH5TZjiogJzDYWkBwCmgyuKU0LRPQ8r2As
gYh7ZpAVeraOjFPOOeiClbh2DKBnGoB4d6VKR6+055J09YBMc1O7nU52kB+XF10d
YGqglXLwXn1hPQrb+emfAGkXGbMjTyo2BhIysIwG5GDM1mMdlInsGjZAFV9pfRsP
vV+C+0XAX67jcacedqaKimO1QiARXGDGDIT2oGmVj9T0w5ALS5j8/o5K4RF0NiHa
xo7xE8ltvI4l1tcgNk7jx4fz532rPoKM4ZWEZHZE+MidqrCVXqTZvuLJjBD/aYzl
D4qnwhD79Aei853s884MKlM1xX0401FqBsKw3eNYWdR9c+/wNdjn3gXcl7kcXmGG
neUPItqIBlY1oU274//euJiLD5/v5PoAEqdv9MpKz5rqfH4jWvJzLL+0J5H6Tdab
qSyBtl8lTEmRsFklMoV3guazY2uvxtYCu/UOBQBYLr1y4u3vzHQXc/jeMoHJgnwL
bwly9tp4yIv47K9QTWK6hNlNvCsGEEx+8wPBh++SqyiFVv22IX8tLJWKfXwiOeqB
aetAipwez+KSBEf6C/nd2cPzaRhrxF17ZtSrSMDnqYzdkiwoyUqlYZLMZIhEdAeS
JtEqLLbH0la1guGcJcgYsOP++PFFGOb4Wo8oCJnBa38TAVLqwl943zgfwX/9pZ7E
LxCyXWh1srEAj0jap6zbMTJCkTchiNfUS3PnQKHefa4mCs8bdYiyD8zfLy49DG3h
yt5GPi6pOB5V2zyDxe5BjTfG7HhikVXQObjrYndInuLw9dfiOa5rf06Cqclx5d8y
bLl+vivKmykF4E/7qcRvJLDHjteydn9/dMBsnzXJEun1KbMfig+DtAsUuFtsrHhj
6RhamXoBstnWU1FfGLnTVP5bSSz7Aw0Saq4YD3y6eZRmcZAQuuQVOfcPjH0hFRxt
JfcjibYSy3M/ZTAjNVe8WFZt+ydloIL3Q8oCpzxtzrPhYZySJefsVelB0RU5Ahce
9HcG7LlPzVCX5sLHchctqmQSH+9MOCgBSMSKDgzY3oZ9yBYk4czQDfrJiUmEaJk9
HmutPYpct0caa4/kZE0/elpvcEd+irCN8egmX5VYlqpHY9mDpGDy/2vNT+oxMZgd
o1tWroHeUQkYeM0TMbaAkF1IVN1UBzaZg7G1wWZvFp+oIifXmQU2uYqaFXle4I3i
JtVdiHnFMb4ylP/KGOU0syym7e1QhKYHjCpNxmnYwQf9JV+siHo9SW/bF7CHYCXr
R0h0C/GEJ0VAkIrjsTwCyz0tfSYoDeHF8/7iHLB3Et/nF/UWyEkh1q5Z/I5ujKcv
eCepXCCp6soeCBTY6ia+zgBTEjMm9d1B41tfmaPe/Una32Np2JmRIz1lkhdnMDML
grV7W1kfUmxZgO+Xu1Na48GcOIS5b43VxTzao4pfuS6zK/7ZDROqzCmtVS0m8J93
GBVt5rw2VubT/Rp81s9HE/3MdV3u12BP0ImTl8i85VSmzT9urZD5p/QGYb2JK4Gg
3cpN8Nx4qPewfbPUrElhU68D5jv08zU5mTU9G2uzNt8n8Hp2Z9l7Ck7vNMFKvxuS
iXpceOtFKU9s2+09Z+7drwBvQUP+DDGyawmBvjOfY9gnO8tAXdQle3cqJBvLjNn1
MFF3zG9GHoO437WL3yFs2bmkF7k8F43z4GgjJUD7qwqBy+pCJoA/KC1hoOC28Dnp
KUKMf/7lHj5ViRrHQhuuUwmmLdFI8hnqNpuG35VF4dKgC/NqAInf+46dDtTogx3F
Cm7PQA1ilTQ6q35aG0imJz6yQHT3VqUkmuPMWRlnNCYhHQfBQ5ct92W7NXHorcAR
Ubr4mnBMsLueOW0vGf76AkrzlaVeKeyWbiDhXR1EopIhb3pSqwvPg/IEqcFJlBXF
W5WZuM2Pyu5ejfbNGW9IMDoMVfevv4CXTV9OpMDw1Jg773CW7Shja1TwJ5cTDYix
A8m/8o7ZM4Y+ezl422SiyCQvbyr5SEK6sAd2V39Zi3J23CdFPYBtzet88TJfPOeN
i5PWYDQR5RwCtW80a2Iqim2ZTvpDF02HdsARCghVdxcnLsBT5kpiKJ8pDtJ3EDj8
cRRAl4n/L5OkxDHtTsCM5xz4wpMTFmTczz5v4PMoAhPlYzVQK5DhaRVI2xuvaxb5
m48Dn1GHcp7asNEPE/xhv03IsbAUL288rP8zBpqJ8x7ZdH5MNXH67gqx2Hvb9OXm
1muQDBnFPVFXDLfe3C2rhU2zc59RhkQxl7CVqYeWUpHn5NXruiC2s4Y7Ng/YtwP2
7fBdAMOykjJU/RLBqW5OA5rMh7d/Fh5ulynIrzvYZYlcszrstn32MyJARPNW68wl
8/kPBNnNptsuEDBsagjAzMvFqXX//1sdSqf2anbmA+WRqOoUzf9/E9yNM0PTEwfN
cxQEzWWmGAzN54TBbN/5qCZ5UjylI87xl69s4KyYo+IZaEDOpMdcM9F276NRzxAb
GVAKnpkb84gDHRKZ33Wrt7Sqp0tOvYBDA54tlLY82SM3k6dyGStRU+TJghpHiCvb
oY0ypDjIky3UntcwlVHgEwWRpGpG0Pdd/ulsFNlW+yfeG64J5naDxsd/ukznkuKW
DnQdvM8M+zez7qOvoAuuYER5SUbzpNlmjE7wgPRgZnaYPHDfVPzECje8Z0RcMZMy
VZNaM88lpVBrw8w6pU7Cqm7ratZvbawPhPzj1/whIEESrq5fmgZF+dNGs4YuGFJP
kIQjKR706R6tteoXhpNfflfe0DAGmApsnpO0FgGgKlO2l2bsPdlnz4mhudibNFYI
NAuKkWASR+XIKSiJLBqL4DC0jvHCDFoVNKw6Y1ePLKi8nUxrGnXvYuLdBAFDStMK
8J7lgV8M0pGr8Wq9rI+o2F95XSKRneQLPS8rbFdgi+T9DiMTREbOovWTTVVAwL56
Nz00MJWGFgq2SOtXpzVhIi2SNj0RKw+kc7NxMcgxWZvOn2gK3ZpmTxLlf1noK1xL
9txQTfu2jV3vgWaom28oGdhOH32S2RGRS66xcVlWmFQ3LHamrjJprqWGSFND8fui
uCMMW84GoEMW3Em4FITkh5G6QC2bPzjP/8Tldjj35bU6/pDS9hc6c52MSpXq+KXh
UZHQ8ll1nfQjhpYpRfPrZVNXCwrRkCy7ylBGRdWV63HDjEfoGH2jX4zz21eq1WQt
NfrytTrTVj4yOaZqmcT2V+tijJVRpmfrf7d88oz08brUyE6MG7Xyt3t4E9u/Is73
82qeUnUGp4+KWHWsD+R5q/srIIv7rs5U4IhKQx2HXd5kyi1Hw8O7MnI2ZVk700Kc
wmJ48ctb1i224l2purOYvXmzTPYGxPQeALSphdzxefMyw/GUNVNVdLzJwlD8Kq8t
ek6fKDMcYyu6GtvmXIcdTBxhGcccZDXHqpGOiDOphjOoL2ukCO55OtIiLOgVP6I6
nzvKu9n91N3nxggso6tP+vsLxnTew2sJXCKngIrYcqglSwFtuVYohX0lo6P73/9B
YOTFZTiz0zU0+cr/akQakQKvothg/rrWzBzBCDj1zf5wFpX6MvKdAEKrXwSz0Syo
UlLEYfrZer0uAhxpf7SnqJL6Uyf6qJwi2phSg90swOmz4XbgYpBZC5iZicuTlZQI
9Oo57fB5jMlrQvL0LRnxOYGv35uPNmWdjjNFn4XUjlAyWKA/Wh+umV4icemacsUm
NUTPpLRtncqxJ9LL6i4WzMtguIRXmk0kvinYHXTryItUKMzAtXZi1lum0PGjtX8R
E1jMaueawGooG5RIAmzR52FgN/Rc3xyyBAOyPMuP9+ahMblM3WWnP1yiCiiGcxN7
UTB6cLE0IbljRlXyp9UGxVG2ZhWhS4j3o57R2fsg0vrIY5VooxGsqSLDG9hwwpe2
gTeyiExFdKmFiujMrsTH1CVQeN6BBymXL4VfrSjQayQJBqSOVJNyII0fzq2xNl79
rSyQQGNGKzf9vXI1xxRMWmIwB+EOjzi8TNlSW77zcbOe0J3+kxzAuz0iagn4FPGK
NTh+4Z6ZEIG1WcNljLHHdj3Rc5RC8rLqyjITHHFswYr0++baWAu7+Igjk9wnVevt
/vj3Qec9OSJhLhDUfVn0pjC5igUJhz+35Ziuk9teAX8JUGwUg/tWspjmlfxHe1Th
UrpOsGox8y1BJrV1wQuzWB5u5CpUIeyRp1Kegktn43bWEgzaWUW77p7AEzLAP1Ak
yUfitml5GDpAdV7oqKgDnTwtCtJFnp0bFItNAEBm9hibDxDyzKCamQDbT9Y1zvcF
HIrUJTB33VygZQqvKIDVuZqcGXGFUTX3fMjUwtS4MJjoSCrv0uAbGOoQ9ZMkBZ06
i7itKAHoeQ1bi54JlccFQ1mRXk6lKg9GLyQKhrolGCuOvXklkFykEAO1JNF/KDcE
BZlLeQTQ+uXpIBh60zZjEczVM7bhfGxjrRIY96/t1v7mMGLmeuBY7yVlPHPBgJHH
qPSB8NAfJttFKyNPEWiR202MBWbwoga7PsUxLY9Zaha8riOwIkQaZM3V2rrXW71D
57XGKqQk2MBNxw4j1hnNEHjzRobEsKnoox/VPWu2l89U1Sg7E70s81qFyLr9MOX3
KPmCNxwYjbjeH+u7X/9ASs6q+CEJpHb8dJhHvkeU9v6QoQSPo+DIC5h79ZNQ1Fbr
Asjl51ffJbSQqq01fyE7+A15lb0kM0LVbTHaw0WPlFsh0v8kBmoKGBtBy8yqCDXc
tduY+kgn6fgZVI0iM4hLXjwYbV/9ktxpoWCaGgqZP6JrW/GmXiJxuTRSZdzfH6b3
ptk6oapw1k2CrF7mE5EAmXtuGIB4C1jPCS4oapW/V2YZvB/JcvJURwbvFVUYQlwL
+FI/nI5yTth3FLQQRRWpMpIsQRa8yUX2Jgb7GaAFCiuy8yUT0Rdgxvjzse6pp2w2
ctXoanWsIbsA7IBkbBp69L+NPATP9rzcUWemxYXj+L9J9ACXVVAeFEd5XLuHymy9
YBSiv2Fu6syZIKk1zC+VUKeXOqyykxzUKQIR79m1r5Vmlo/Ii5Ili+95xzu/YOqe
QeFWnm8Br8AJIzJixd9Ttgwh9ZDOEsm8j+gM+X/vcv7k159aSmpotLk1uK4KTQwp
LdmweBqa+JPiSiLhogApnak463bDDZVLK8boL9Cc0dN6Qn7c279koo2V8CTrLfkD
8bSPPZVQanujBPY5+xTFraTrX9ewNN4Gcj2v0mm9PwXs1XEMdWTlbkLf9xgKZ9bO
R3M0OAmbxH+zzCW4+B5J6zK8iYkQgYje0mocV2an+SurebKp9CO/hToH6QEGHSTR
0FEXLtJTS8gmQDqO6JNADMnyK6wCAmPuXVrjIVEom0c6MxZyJ26CBkHGyPj3/ppT
5/B7PGysQV9Ljn0jR3JPmPmfjhdhpiIVL3DsWSNsG6dbbPhsX1gNkmNkhe8mmufJ
Bi9JxEa7L9AyTyCgw+iS5JJanEs6kUrF0ufFCChoEn/VYLw4ottq7IgmIX7ojx/v
KmnXI6hX93D+OQ6i0GHOQlvAr55a71P2UofthfB9c4v+QiKgI3OwG9KFWxHvIBfY
hpwwX921GEXAv75U4t3gruyvPhRTAw+PbiKVvYIwL49QutuZbtNp7V4hTDNhi67B
YKfa3kO8kSTAWhMrsiDhLyZQ5ldN1gdeBSweeO9DZzhAfgToS0bvFCukqN3wXfWD
jKkmsjUlKS274FVNriM3fGcGIEU7mMF1aARp2cKgytJagaqyJdRzfuMavB24Eoe1
A5OnbJ/dc+/8Ey11FYLABEmecpiTxfR3FZHlA8bnwQp+8fIxCz+2kHO1VKUF0XiD
tOT+9Ssg7VHsj32fzdNlYpuCbwnrBQ8fZUrtY8lLdo82UGLyt+TR3XJ8Dj5Hgqw/
/u0p8vox+NUo2Ap4Ch5ACeTEqCxTwtsrjaAeWXU2ZWCik12QQjYfm7oSR7NPCWGf
Yme3kByyQ+4eDra6gr57MTjz4LG9+dM8ilHeJg7atxiCmWihefqK/zy8NpWmRiiY
R4OykyEm88FJN6+J1ih6wGsddKu2ZAilW0SykcLhRP5JYRqvbFXj9FnYvW6+/m6D
480sdTDOF6CbSDkqzGBQMlwFrzvZFUHq70ijab04wWK/0nLwlBqb9G2nO9AhBMQN
MTrvCFXhlChC9A0VKKmgdvUELWXkkqRo7PR/vtmJ6G9FCXo0OGvu0zbJN7gtA2Ru
69xySlpq2hIqbbGkxAIDp89446SRxW6YRPynjEvqrN4jozH4pbXkbCuXbKMwq+Go
Czo02L1K941RVwEsQuis6h5FFazkkN6KA8dXa37DlnwhXLSf4xvyDHJSXzwUcLpZ
cjJvAHeDXYieacw942d3aECZkrKUKhkN/+LT21oNcRbTKgybxpKvlo4f3eQHikoi
3e5sjv4HxHU4SEicM1blOT4IoNKhCcNnmhKh0co4NaY3eeJLLLlPJAtSKFOwQbI7
ILkJhm6NX6nL3N8+0xYJl9fWth8N2XrpOmMTAm1X3hjJAZ+IgOT+FuBhj8xuON0G
vZk4oWPjEkVjOGjLwU+anYIt2nZOb74so8j+757Bk8C+BQBZYdGupXEhVqmdTjvn
dg+ENN7eB+2z/WzzVMSMwnHIvtZ/8n6HOTmLTizLExBVJJPE8LIGMLfSlxm5WoPF
nZIt/zSIpE+Ohg8FJGvzxHcAsmudCvH5Me4hFJ7Lr9Mop5amh4zK5/hx6HHr7YSV
EmIiJYRDKT1kZ7VqCuLU7ba8zzU/QARA+X+FxvuywqUFayOJ/D0yF6XX4UC9/fet
gOxY3htFmlE/3IKyo12FdlKcacEdqBk53/1YferCwegwQNb/ZENSp/AoPS2OC/8Z
K2r37/s55HlC+s1tcADFC3A59+fiirBTMYCe4EyOVyO0/afedWGEXZ5f2P06pdbN
bvz+qW2RoqzPJPOgA/fNP9QaskTto8ggqKhkWH/mmL58PtVQvJE7ih670pX9hLP6
il5wV9FPpRuF9c3Cawpa7ufGeY73CBY8V+oTjYwWt20lBzPbRm5I1l0BYb4hHhw0
AYTsPdyRqnvR625jOeT8vjnzQ0vDw+T2FwXu7eOga1wrrTXVe3/itHtlhXSDyQ9J
Q1Wue6F6yj71yX8CeqOjneG1YnDL141k/gnZ6IIO9Y/l4mlx3fuJc+uo62nh2bZ7
q/IBOJpbARpOOfcLcEm82PDcQ+UtfDL90b80nqib6uMpBlJXuwu83DDCLVm22bMA
lan0Y8mNhpAJ3v78MgjhrK3NOuS8xmBDayJPx01wzL+zAqC3wMgKJMZfZqc0Plcm
HAjGpxLkBPGupUfyaMZNlBM7djGJI2dVJt5fYx5a8XynL1JmxOwn/B9q/O/Sdd4O
iPkto6/4hy4w+W6Cxc8Ute8RxLhBiAgEU0oTOE+LNYJPmiqUHeTwm5XG4fKxQYFs
eUFtHJQtyQegba4P07qeK6hGFTZ/XPUppToqvXfvdjE32rEVzsOhk1SbK0RAgSei
XqToDRaK7wmPnG1Or1JHtp9iGw13nqQ8pt3zdEBk3W8+s35Ep+bm3qbeWAVao43O
cNlBK8kec1621D/ii+NfAr3bh7lIUnBXEQNgpmr/bYQJ16xv8jfdIDLpKXfyucEw
2Hk8DcaoNig/aKwIt9OO0Og40gjPMsCc/jTJhWV/N6OB+6NGd5veASYcBJk4domg
lssE547WB48xa61ju7TCL8iTnK9egoHzVEONGTPwgZWPJBLv0xGPQYKDAA9J3+kS
DYWEmdo1nB2Sd/9Uou0zhigddpwuP5NLlfAa/qm5XOB3QJYhpgVQ8/YiHd/M4O8b
26taScajuKk0u80KiLYM1KhJWHnpeaxAZU63fNNvYMNrRZqPxZFS8k7TGWyN3x0J
IR0xCdmavVcR1y3Rz8WUIZaqi9+yknNpdisj8H52AqhEyarjTi2rLou3hae/YG2i
aXfzUMMnMkIUfAo5ChDDBYTN3Nf3OuxpS66SEPQedLC2P0efdmxQHMHqdUp/akwB
kWD/FMHuqTPcdGUENJzgsf8WHUe+8D00jj48+pALj/OGuu9swRDL0cUsyDSJtuNG
gEfR1MjwMEKEN0aBUviylMM66/MacpPba3aBYBb2jlDQC4G/g0/zCE653UHh0Aek
3VjjP1rEvfnssOcQROYWcWac3EHT5rbF/JrHyU40C7kJ1zwUeON7NkcfIHn1t5pj
Ufo10abt1lONVnoWRX8ySgGKPTmKn6z8sOtiMoZ812Uk1nBiB98JUxHEHQki7APX
ZaTEKsrMHYTNHi7mPDsJAOOiQgYH530RpymtLKPsIFwKuK1LLXGEhUVQfW0dFOCP
+enAgaGVSvb4QZreRCla443Faj094F434J8LfQr9BbU+Q/x6Mi1yiPV0uO37Elyj
a2HF4sLtJBghlVe1U80CDRz2dFotB3CbSVwZuV6o5R/HiCs6UQayTlQC5eMt8ZA9
ZC1pqsn70vL664XWb6ihia9sLTaezXrmgarVSAAnMQ/WK5IENxkkadqYiB/sHVOm
g0iBdePBakkanKnB3V6Y78kv9a3E4GMimMfRNbliR7LaqdstsbculcIBCduLKMK5
Aq6Knqf7UurgbXZJEg0Ll9ttFLrVOtP6SQHJ5Tfl+XnoiB5KNtn9d6EkcTq9TVRJ
vH7qXaMI6nHuJUadshpMl2lFnjPNqC8m5CPEqZEfU5BliRZKcbR/DrtpvyOUhtDD
EQp8sZSiodSWfrcrWiT1CVj4APPmqJuoBHseAS6ePVf9qRXF5lrQHOUDauTR4wSU
dPrFpIfbdxRqR0+zkaR4rLnoHEGm4iBG2oD0FHg82qM7JUNZShJXhV0DZAsWLJqN
u4xSB1uacm51bAlE3MjMK2LrvTO9ilbmz+ZLjWkcpolXAkGNbXAc0TdKYhcyf9ZK
RJ3ZQqndOgNZXz5yZAys7OcQQLnKbqZBxC3gZMcnqXHUuGIyljnKYFO+yiBCaiL3
gieWiYTxyRdI7xy7nOo3dwgqbgbrTD1FYOaGKdaM20EjbYcDD4whBEIS0dqBKozm
AGD/dFYW93mR9PpLfuJZhjcnaDynhBw60PtKvy7CGZFkzKwcSOuGNR2d/AW1QdHe
+zCJIRDMhSLyfy0CCaEDbxko7ACZm5bzzHGiTwohWLXvlWJte95CPfdqIE8LgCaL
KreOvB9l1QBxQHK2R0X129qOjSeDIEMndd9syFyVq+XiWfwUote4f6P214OF6HXz
DahnBvsIMj8uPt5dI8Lp5D9FggQLrKIxbH2DDcuvcY8LyIfKdw/pQMF9PucywHUW
I7+MHUS7IeHsfsYD4MiUH6audw5PnPhaNqs0p9mhgpiniaXl15Rr+NSOnV4P6lFp
DwCBiMmRbl8FhUp9/46Luqc4ycOTLx9f5Te+tSgZkEaKigYN/u/R1iHicuMJEE/l
gB4o2iAZvJmvzZiy1D2As5A4XRgvqASPrmxYc6AReWWrZQoweQrCPH1N7rm0xDG0
RdSpPmbNhODB1y7HICM93cFcz8HCzYFo2VZtMD8/KiAIJprL6hmRXQe7g3CkA8rH
r8YQ1VjvxFg5AUgY6Cp630UPr2s7yjscYk+kogYrnULjItFrG1tRUHInEb8YdYSI
YU83ig8zGMzHSD7UILj7i+GCWHOYvsVQ+AoddV4PoZn/i0+rxOjnrBRD+lcYvmFT
nxCQ15+R84/cTBQgiGKLvsulgoG+lMo7tw1gW46/6tozh/H5DAdLEPUb5EFC6Na+
F32SPx708YPYNgC2QzHqeladNeOip3E60zInLP1qRLguaQCAW79rHhSA+SFsnQOl
NEpdhBx9LjahiNCbKT5laZ1xpG094KCP9+0+5RcL0e8rTgCrVzwyx5gH+Mt8q+Zl
HXHju3cL+rYm30ykHwHfxNwRXxUD46u7amS4PqXGMRVO26fVKrGLmMcrtJkcOUU5
v7TaNFeddiUgWO6BxZggYM3pbTphoLBoreVIjOIi8oyJgAFLBAxuSLbUPTOhMo2E
hUXh+TSwLwK9fkM9JT67q5GWL8+nkzgu/fTKMyhcOymLC1ATAAzS1cyiyMwTvmqu
z3AMqptln5WWd862oWyodyLvtzJttSg6QlRy52wfcL5CJMPLY4idGjXTvtQxBW+9
Tr6PFjmm49HJ4bKuai/x0A==
`protect end_protected