`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
ddtXksX2+yylW5zu6QL2Lhnb2d1sD00763mmSITNX595NcHTEkwn0zB1Dry37fOW
FufOhVzEJp80NC5qZ/+F0Vk7Ik02dIR0elf3clrjeJRK85K4e3Hoo4xn7YbFUIms
l/8VZSb14+JVGURjfswrIyCUotIzlzVYZ6gzoZwDXIi5gQIBf/gI+KxNXPaKV+PQ
Ufys/12rjO6aI/pPlqSm0hCvftmBcnezN2hk1UeXgOIuKZnogjOsf0iJVX2aOOWE
6pD/psybjbnsNB6kH5uFTA5frkzIzkzl5d9+YDm9OyC+k84E83I/7/j+rk4L2dah
QJOvksSIzN867/4Qt8qYTQ==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="MvBXkzurAa5VTw+1JJ70nePUfoQXBvZOku/SMmg4TwQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
oRtzZL4VJ4iwysPsC8SXYCzXS8Fw2gtZTOskLcDV+1B9Nzn1zTyNtlo6lNICRmmK
ZRVu2BmCc2G+fmzynYlNTnSa7C0Cuel6FYpxCBlOuk3OF2tzAmLAuDyOH3Z1Yjzk
a0aHuoCdIRKv7BrZCdALt03JeUmXKPdOmIlkVGFl8yw=
`protect rights_digest_method = "sha256"
`protect end_toolblock="Jn9CQpRhJt4rnzZPRk+dOpzAubz7omckX1MrFd4p81o="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 42256 )
`protect data_block
gD6l00tciPUa6pDNTk/+t1gcgy1iCdpjTkA/bOvU9JA+cpFEv5u/7dp25hHk7lLT
6tYtR8HgwcLXTcx68BnPlzdPHkVIv0lwXo6yhFVkYlDWBcqD9ubowgKij0UjlXmV
p4anbpVt/gKvAYRDYe8Q5F2CQ8AIsxOuOcJ2vhCPchS4QF3n7+oG0MKU5ZyzxTu6
aCowB/Nv3ElMtK6/mGqO8EQJj3PCmuuRWutr1V2k8cH1xnGKf7FNGiWD6T/AuCt/
NnAo3LIedcG5XeluF3IQBnijBmfxAoeO5Ua5rXwQW5Gf/KSv1ecHGdg2QDfPvx8D
Wjm97QSsjbht6y6gC5qT43Yzo6YPHOpwanPS2sQDEgsQ/X5WDDuDikGGBb/urlTJ
fU6oZx3wPyqwAiObXmxcVXflmhqCYo5Xy1/Rnns2WvQjgDqSjKcEF6ACNQ1Iz0gV
meBMxRdzNBUfFkaEAlMwfFSSjFREbOWa8Dz50j+PqYZhvdVFpeTr6mMHBFg/iOiu
LWth78ca18BtiP1RccCvZ7YPQWfN/2Sq3fAfXQGASBJpp7ZXwQ/sFGnlDaXApY56
stGMRCMXCfgneVTIiUREujIwwO6uxV4S0mXO6VF8478deJXyKYpxL0OJ3qxwtnQ5
uAG/k9cnoqygZt5TTaBfd0LgFEqSpO0dXlVL+fBjoMxpy+a7UNQigPUwZOUX6sFx
WuHu9paCUuD/qOuqpQtjbWeZR03bfhh8JV00nMPymAKsbUE+ZFiX4O7GeImt+tNi
4/vRgedl7RZ/HULqxnOCzAh/vAlwi6xyfAUm26QJ4TuqmDJmxFi7kEghsrBIb4MA
YahcFY/tTw8CtsP6ad87OZ1X9ekrIS/brEZtduNHjhFNCIGLVdqLZcocFzt1sqZ5
m6h7u/cePnu19I4ALUHGoouo3JImqEX1nbPkFvw/SWDh2FcxX9x5o4BwaGpclMSP
TFcfqDUcHACZxCzQAo3YDFrsyWM5plJ2R3SexRcAWOIHwZHgEiLwOLkygSuBzlwH
5NkParbCfuJV3AcyHHGakjQKNOJt3g6rzggSzENC9ekXp1hz/1cSxH9Ao9t1DUEF
VBV7RO/FGJiRs+HgFU70bajIriUhcHsoaBA3gRqISAnFwF9m217tGOi5vd0pJoKj
cja2pc/37ZxNpxFaIfqPksIR5q+oIYzYFrYtxqdLFVJrYZxfNguHpkPR0BzTWXGi
zl0wClfY1dx3zW1dCgvmACT+qRywRDgN19aPhDFG/1WwTR988R9pTtUi4nBIEQ5o
kjf+mCT5VMciE7FaYT6IbcDqf4OuRngi56n0qNUF4Y6BkNykPF8kGLkhaqFhfZUL
C90ahUmd/0pyN3iPn3VFPck2mvOoqHVFQNLow8WZ8fIjI0OAVbptGRtpu6JmA1o6
c/5/71juW4qFrmhL34yJy8cXS7sm4TDWftZc9ykduFhBgdBfo53V+XiJZJnCL6cj
sc8T3I/oTk6bVzE58HRJ4lHBhkwB0n63aS4FnoDeit2N9cZ6T/WYK7dcKQ9sPXJa
PyTiptSwnU9BsjAxU65dVEnY/Yu5wI+AO1CKtseuVWZIk5JigUbn9YxsQ8Ifeh8u
VViwnxEiJmhLX2vi20QgtjpXu7BjZn6amfysjL7fENQCbPLWrIPutN+pGcXqEhjd
v+MYBD4xdl6yyWlQNlaDSre1GtU1qrOizBbyuavDhixIHRw2I4OHBDQiCjj7412/
jUx0Cs7GeemkAZdqzkX6NW28nX8iPmtfs+2132SoAa2EFlNm131i2FJjKPOyf2jl
3gain7GEXm8BEGNykfAtjuIzDGZz29scz8DzMg3pWcTkKgADHrqhzmt7/oNKfV8s
49O22BK1F4FHHLll/AnGPxRBEEDAub7110UFNyZVoKDuMwqbL769ubpa7H+run8m
+4OsNkCPq92cYkjEZIGxX0NE0VDKOOX7Bi+9iLycxmh/3rlW/2QpA8wXSsNS0yht
UPMntyzWUUbc9CxN5pc6rdBbRsAVES5Za+rxqEaUJijsLjLadAWj4hwSa6zENI47
mgOVBjUyQ1e8+1fhaTZMST3fJtn4MhICX0pkPA70CpIIBCIH043eqlyK00dygOh3
EyH+H5ybO0RDI+mN2i4JfCIq3OGNiwC1CH6wLivP3pU7Zf29IU0ZHp+iEKgF3/O+
C1UXOnLXxWOUE5CGdavbSl7yomJhFDRMIlUcS5Je05HyvWnfJKubHerRtcFY2j/6
+Qh69iGPydVcT13WI5jCRlV+yPrjY1iDiWEbafbRonglpM0PEgOLUPsxvHfeMjXs
IwSaMDXflFSX3VzrtL6m0m7YQx0ykuhpPXySsToq0UT5FYZ7gfE9ldYl1qEChfhz
r2wzU5HpNrB83MpkfvzSm6b7tgZ/fHhZFFCcgNmJ0mHn/7z1bhXoacTLRrs2Umlr
KA64G6yDLIdEkKXo6I5xxJEa4/El2ZH2vtwXRivRqMgyD2QHN564u4UV/Ye6SJBG
gJuEmWdnFqCGVGYrcE5YKMEdBDtRmPPVQURThPfyR3brXPIKSmLtoGSjttMrKDpi
QDxvMHa2dFdoOFsk+jDOgRIgQppw7awcDu9osc6lz5eK5b1AY5kAs6Zzn5Br0nHc
1uC4RQbq5ujhC1Z9SuUcrUYUb9WfiHBE++Xkx5rtP/jHEsq0//9RZwpODIrRqbV3
/UosQcnuClDlT9P3bw/RhByys89+AoYYTbpYxdGcie2y4wHIiG85qnzEY5SaK3To
ebJbsncyGn1ZJWVgMIDTD794r8TMhVxWc0GcmZCfN6ZX4P4aW6l7MvNJo52Cymsk
eXaBmg13ybRfcQVAxLIgyFGjKFbFTIl+eLU/uL6wkNeVPBt5H0LFYnfhzcID9WQF
vY9/ALkIvKqqfRwQo0GnwoU2LcVRyAgTtn8jXn+qlkF+//oV6iZDkZo1UsMiweLO
yL9VCGmHYS5D76+S5tkaD0LCXSdsXqK0xvokp4EshXzyAXFIEcrL2xWMl/Aeomlc
uFym2aBydaS4WNuhyheA6pyN/nSBRN5DRSyPcgoCGS8Yk+DqjBk/pGPDSkZfnBU7
tAde04HqtxjE62UMNQtwLm0zUgTQa64286s98nK6a567jILwowJPxZhdVNAjgGQC
/8dLZ5FV0Nq7mbNHCNfu9DMG6MOgvsu4BrepdgN6+COUoTmaiORfRzVHQ76hmtwZ
u1FV+idR9qZOPnMPkR1n5jli4jIFQUyFSNLFp3cxgcdn749oaS4CKETO/odV2PV9
3p5FWyw9YWA0uwyUx7wk49R6MJbyWSbBdYeWvWGPV3W9sngrhNyi5/weT0veB6YB
PVuBs2TnmG1t4fLxvIgnmOjxIM0HUA0VbeJXkbWZuvOyvrAhjCRdp6NZCdFcLf3t
JcV3YSmoHZ9bdZaBBRshgkT+qWG2V0VH15EVUUVQos011YecR+p/vxl++l/F/7Mq
8U4qYCv76AC6enLlvFowDIF/dEl75Ej/HVxCyOy4sBIibH4ltlwumnrd9TB8yihX
sQRJDinjEUt94bXvrNa+8HIC1rosH9ecD6iyx0E/n2j3CLMKVOI+AZG5YHqbnhVv
sDqtoAxhKO8OaZlQTpHLS1VDFrYo8XE6MPEutAIAxNoCkCLj5VTHRUZnwzmTQidL
I6IrEyjA1uPXg6NggYZy7NERU+gkJm4bpryqgOX6T4P9mm9n/zAlRr59k500CX9F
SVBRaJymTu3jYMYNBa5I3tvzbn7So6Fj+RBU8V7dYRd2/uglBMksvLoNnPPq7rAi
g8wFiGCrZsg63Z9SjjdA+FdpS1ZrhjNQHbnUfV5lzIcPzCMxSegnM7RHRZxiacxF
1V5a+ys97WWado97tXXLj6iNxqgBMFP3H8z5wMnR8xuPZxW4lUv/lShCgb7DqB13
Q1mVIfhW9wIstFl9F8PL8tqtLCXPNN9HALXdA0B6Y78khx1BC3YlbIEKs0bMVL49
I/UecZoTbdnhAtxkd67hZ3DoMM//Hm4yzbOWXqYQk+NnF4WI1UsTqvIFIW7o4o4Q
8fcyuLbR+OyusgQm6RfIE6j31XIlwyD3bnzZJV4ZVjm290Q+RZim0Wtecxl2CWQ9
ms9JPK17e88mbNGvGOPJ5Dpq9pDBp/jBTsxEK0lNqYSK+UZheAsBZmnBKHpBtz7A
RWrZPYQj6QPSZpBQz6XpQXblNfeJWkpQ4vZ93v4k6rSS4aNRct2HoW4JzTSRby9e
/wuFlmddI1xELVOP+Se57VdltRKX4a/bBBzA5SpeXRoe4scSH6i98vq9m8pK6mVb
CeUN2AsSrXy0yYpAaie07zNisgZVgLNn5glu3lOY3jMt7BDXZ4HM+lPp1BwaD5mV
5087k8RIR4wr0A1w6NlABP6Bb88mdght8ByJvsbGDzBe0b46uj0bV4DIQNKDR4ET
voePaoIADGt/QzSev8KC4/qw0xX0eWMy3JFwMRYiZTN1FYchzAiuuSeYtk8+HE/H
IrgFVCrNuUpl28l77/9C+moaJXcebt96kxyHspWoDGXuUSCr+faPvFVeI0iO02Ip
jmYpHH4pTPO9BwJJg8lTli2riDhbsAAUfl5+mRyUDLCV08B92R7wTmhII7iE0KKP
FTRWs0zZI22QfRNww9/ZE9+Un6JTip5qXxrJg6P+KIDGJ9g53utesqhJgkELA+ES
rNHx1m8eptAdkYWC+4VF4/QFmtxI9ohrx7nfj9LSSpsBFdBwjeuvJjYXf3P7F1iH
Gevopv6YEk8P/b7b69MNS+DGSyhGLE/97KK6vOOVqM4P8ng3zWCKTuL0qVU1BzUg
c6hOSUGhVldIFi6lBTgSiX6Ac9EAQCPv0IUio8i1hxPH8ABHj4KRsEDI58b6uuxE
NYO/fWc7kpvLd45OVr3fpe+zkQ+Qnntt4CyWjTTCLH4WzvH8SwtA2sYhYfx5LTJZ
ErIg4srD8dqKdT+WP19yLZSdciv8HXO3JMBA+0BZeU26NeYyhJqTrLFvyPm75XNB
ZOqMKhSBxW5m59UxnBH+qSrjOL4g0jdAuE/ZmNXGGTeCN8NZaCT0+a2P9ZquFKZY
qxENBFX2p15xE3ecDYHPnruLj8XUKdWVWZvE6A7P6IRG8rtunTvilCgyvAwrhxBs
Q+8ekC5mYNM6pHGvfw8BzhJNrTMP1SAZw/JQeE5iQNSSeGzUQfvTJ82XxucIDAFz
ZraXfzagHz4+P1l8JSu0FBiQV1fKx2bz+j7TbxULSAZoubt2NKqiq1ZKjE6mQpTT
70piyo8//vACYw9jk2DkQYRhJcMqjTlhLeAW9PaFYxAn20aWPEM7/4nXsrws/UbG
D6zZhIUXIwLx03xuU3fpa1eQB8aldywHFoo5Nt3e/KR/aEIZ3rqYXc0h/U3gXT+u
Ybv43iF+3yZF9wIXBQmx7RtJHfsCCYiP5/owIha7DgT2tmmmkaAZhkQwy4pNvJ0Y
bEWdLT1fx0LaLm9a7rqskQOUSGffz32Q/W84uxS8b+cPhTnlsSDUqP3UCuOV6/V+
hXzhlMVNxLcrhgtnsaRfYM5OEjpjKO8evGZW2Zt+zFub4GbzbUMHyonHr+YkWRFv
Mv84LLwdO15O3Gq6ZL0KSauzoain524RjawOzrhRIaKvBFrNGEWTAoyr6D4rMnjw
ymelDEuSOI4XOKZ0pQhrZXRCqexRm3duGHTa3SitHRIDg6lCgVm/Gef8QehMHTK9
TgAF1kBVOqCJ9RmmvI+SynoVhwEWcY1sKArtDWRxqu9USmZyWWx5u14XY69k6sRD
3FhNlORef4Vl8gM28GB1p6S4fRpc420sk3tPvb/saYat9jakGjTM+3/NwnMwKuaH
qT9TK2Mauq6BBzY08IZwYdUNuoP/W2FSAqPQlP/5Ju5Lv/rqSKdzM36UVjMlSFRS
2ZOIpfDcw73ih+51Axun/buOY+7w22gQxhcJ3CE73vkFWx1kiQ1ts3iB7WNpnHgR
K0gFj6IVqwz+ox6xxqdha4ad9sWHj0eXj995XuXsvcVMRwy3KODYM1TuDjGAgOO8
oMCVWY6pOICM8gp/NoMhXlrdShfoKASeDDWc7yvecRNcWChAm0V5PScXv9TziC4n
Vq0QIV/SkyNhGRiSPH82bGnTD1mf8n+6Jr2Hf3G+OvK9MfVBb5qAEQdcpIbfQn+I
jxDHSxv7oyw13+cFjr/9ZEP4MEIb+I7NLjpwzeveUiMzAlxhBB0cUbPIRzwdvpCP
OAnINcT54vV1oDExQfq93E6Qw4K2smTYc5KObHYn2X9idfSG/tdJiK2fCJN/6TAT
P0B/RyEQpvoC1RqD5A6TF/DdslEVWSBxOBKP+2W26M90ACTPByArlrvW+9i6t7to
nFFI4213RLtvMZ88fyiDYH/GAmLQB5OS+PRhDnd+6FMmo2aEYSl951FrTPPTq2w9
i9hamzR1WR8XK4/hWJINcfkFBBiXiph2maXpN7LKqY55uGft+Yy7cgkxIKHvHufn
dbRz6DfslLVCd3FTv3dyc7q90NOKmLSzKLuZs82btPPiyIIJl9AYeEHxOuMu6Cin
m/B/DF0ctbDwkYqftkdga6dw2LUJTXN+5U/FSrotY1ml0y2n/nIbIuR4VRFykVDh
XCUY/h98vgAYKxFnjrmzhY1n9gqy121Q35VMGUrN0FPpGLOhjONBJEnxJ2XpY/Ui
eOjExXMu+SP9MplBg7G6n1ebDzM6WuGDLjzEU/sK2pDMfg3TEwFpfWSVEnE1yGpi
Z2LKxdOt8KQzZGLj8lBTKm7WZbeOd9HH9PIf1X8x0AyC0cali7O8vLKLSCEV9t+L
3QIWrLszZPXBgzxHFAAQr1kj2mB5poqhewZ0zfWM7J0VB5V+nKZIvRKbiTmSyB57
iL8o67dQ8KgjmxTZPoVcz0Gsl/eCKNub0J1KpAQllssBfp5+SEy9fdJ/6hqMCm5d
5STcJHQurmaBE7Nc859L83E+yGRk4cSUSAtuC1pK8aOXAlPE27/mSA5FD1ZOmose
zreg4HSt4b+4UP2Fx8YdsMaz/cwYk7pUv+STTuJDY7lm9opLZP8t5EPVMYhrBUQO
YZ0D0g7yx5jQrDUQBD3/MrDJeGTtXc04cNX6wiM+jVSiKR1mdnman9NekmZ3arM6
CR+0q6+0lJ/mk7PUUVXygCLE7zt1M9/kCHJ2SNs3LsBFIhXeYeUnDwrUqdGx0Dkj
PcizGN6OBkpeEeAwH/2T37OVlvOP/2bGMVHjXdJyCg8f8PBPsTq7IL/UjIxDiXHU
aMxc5pqC8LtRnBdXT0K5DqmDR9+F+oQ9ryXNK5dDzoLg+uIF5K4i8T3v3wXHo1n9
gvDFYwVjwTsgWYGuUXaOCGZRh0V6Q5OpLXJYhJsrbzmmijaNC4yJXngaDzNPLd4M
sSgZRc5MsdMA16ikm7OhIaRQJ4n6fpMAOqD6RXqGjEUMQ+W138w4HNrkEIAkX4mC
Tvs0Dr07JIurpie2rzbsjyU7TzG5cypebSHwitCrlo0qNSd/jZE5F21Msb0SORFN
cYy955T6w78/+pF9ghoG7u/10DncSddpOS5vSS6OdPfYv7+tX9VGaTHH16uagilD
zHXED2kMJ9sur8mG67WLlIIYfwyvh9vDQnWbQXyO5g6h0MfP1meOFnvJZDaeExMf
c6KRp+t5+A5fAHt2XdTaqi2hZ+/Q0Dig2yfHagT3kN76G0YzICMZ2bKSlyp4RQI4
vOHN8MGlddmS3ZETGV4TXtI+FursRx/RrABA4sfCvZLrrLl52NwcRxCHg0MRwocw
Afmvt2aj3C3G7DZLr06hEhnCTXg/vmzkOHDDUl36QTX12uvejN4+QEye/qelPCG9
6NbNwOPIaamtDdpIyeg+Wigf2fov0ig4fmIMb1TSIlRJn1SueGxhp0yQ2HA4FNIe
f4SPEDn+CKah1lbdspfmz2wb8UNkjAiQJ4EcQUMHdX8XUfZQ9ejRKaAFjjWe0HPi
PPPCNM0/swbtg8BQUiyqWmO/j/N6aUHrSsc9pcRf7TH7mPqI/lFjFaEQ7LVjRZ9c
y0xQTw2uuybPS/awH9ILhAKvosa5Dun5Dr8Il30MFecZH5G8vP7WsNhWOLMZe3p7
NRIRVh1jDlwXk10VI5opQoDY0i2clP7p2ckaVeSlFVTTzIadFtsQqbBsaQ8NZYI6
oy7Tu4xa/7V5nfl+QMZxGef8/OXlBc/mDnqTDlvCKx6jarJGSCi7PDHKhJI5GN+X
tZcoZ80NY6j0KCd5CBrrPLoThDBgANo/UWuptTyZiECz40i+1nRGyH9vHxo1jd7d
e+XTAxp9tjYFgFBqKC1TwOVMrsNhoPHhKXzoMKFMC4e/aWCU/zd7Nyi2HkSdpp9o
p50QGuNIOEwd3Xr5X3Yr+skIUgYqhwW1HN/lf8CHR+llIPSttwX/un+Z2LpBw51B
hs5WRLBwAo32PlKRzDXEw8fmI/NHqzV0j4pTPsQdNKr7VS39NFc8PlHCAlgbIZz/
kFIPFqQtCu6fhv4WUjWr9q5dmwbOE1ndogYAOFRxF945ZEc/l7JIzK41fBOfM+ya
GlvbjG40666JdxNY991uA44GxZ77nNukLXifTRjow7J/4qHwjmgp65f8zWK3kvz9
qsSHk8WpJ67FNJka4AyT+X/u0vFPQLnuOgtr6XMAlabQDwr2yHfKy02TI1COY+KX
+ZvQJKdVrC3A+TZad05HmgEDZ/4WhJJjWht2JyP++Difp4/FDCl+PMt03ekUkfLU
Soat9ss8l1VdYRTbq2ShIY0IMX3ggr27IMRK+oYISYrLKnfKn/yH0dcTHsXn2RY/
qXPKe1ARHavm9kmoFoIFp6uz9HUp9MFI3WkHmwCZyHBCQdqucEPVM4bAcZh/qnSN
r6iedfMPuVETKRRtwjHDdpyyIWl9bWXICP/vkllEvA1siUXBQ6/lorW5RIjpvP2h
8vJwtkYsch2nLOUiRdV/zcfYL+YRe1vSmktZy2IMA4lkjTmMy0m9l4K1jyL/FiyI
tp1p813+q06CoC58B9K9AxSH/rebP4G8krUGdW2XedjL6GOvJ9s9oJtDoQHvDUn9
zCO++bR9x1BxFUiCbBcMUN7xrcogAvl5SKr+xKbs6SLxya0WjlAKoeF7bEPprG+b
ME9beSmZLABpzUubLNGv2PZa4X4K5Oosnikgu1TczMVovVzJR7fljidDZLph+J8J
Euy0kX8vQUOh8cjRxKUT3zjMASHsKBKM/xvck+UWMOpwSc0qVMqArs8l5+LmDKXb
NqJp52V2j7USudPv5DQ2XpolbbQ6IDqq0l6J0+Ve5amBLWrwl80EeKheXSItP0Bh
wAGDWldlOGK0ZN1Wa/5a787i10DX9DZq4czqH7+2Qk9lN3uc/fmLfHmWcB0LFI/a
Ropls2OhOL4SfWIUe5XGlGHiQn/bATcClXOdqPrkUCBrmXwfbZ+C+nZWiljiJR0K
1TQ5+2m/BE6OmTEtf/BH2/zRbCYFH43W2SbvOr2i7aG+S6V09CB/7q0o12bzk9tQ
RN9o10NTJYQjKUIAb+7/fFyZtp804Xhu64FEBdVk3jOJbolGGkgrzrPcSs8/urWa
e8S+amOmLqQuAPu74Ra5dpsRVSQIJEPR5jjJIir2Tie/Yri+14cC+edVAjIhrTp5
m/fq222Ooqlsnc2byWFkxU2b4l/kda5Oq1gZcu//3d/jAJK9pL0PzS94e++CF3W3
k3HFG0GizBsrg6vyFoepujENnO4eNABQOnBwOjWPnEBN6jQDGvDs04R43fz2QiMc
SVBBl67hk/IZ1Cuz6ovd7o/BY2EvKjUHG/mMoi3O9bewT3i36wT7yLVA/s6WRcT8
lH45YBk4CmduWNtLA3Lr29QJ5V0Y5k6pZDYxdGW9D6f+BlPXBbMnAGiaEqij3KKg
PMDCMDMCDlMmL4j0pJE0/eopWGN29cGTE096KDTq3ANdUYaLcUSqwJ8Uya0Hi2Gr
ZA/x3YorthR11hmkgLLZs632kdwChi+JHufbwmDHvEAh3OcsIQ2CsBN6Hkp7tQ0p
Da51aPbiRQdvfvgZLO1VGRp+gg5BXO079XaOPKMFpJERpvlzaB6AYRYQ5n3BfsI4
6tKO5Smr3pYGBSWtZKeHWojU5C2jmfOWqetZbF9KcGzIGMcwr7Yq3/LWDrEGcfma
0uldEX+m/pCNqsVA+6FJt1jGfGXvpnVCT60Y5Cz/Epi4kz6SDR8oYsEe/rwVkXrz
mRtngXBcQyc9XZnMpW3wVgqCAJ6MxgxRcWSs3MnRSfm4lYL6HhAm8q3yysHxHQEM
EWXS2QSInGs0fNLvL4JyckqG6bKIsKqlJ6e2wkJ1dxQmmVmime+2e49H6f0e2ri5
F9IpdDxbPK+JkMeca9FWoctIt2SHzyfUq3fmzB8XUiER+mhs8o1DSvgSbYJXV0Cs
bS8+vxN2fMwDNCbmFe2xbqVFIuXk7EnBWfk6QRGFqTddg2JoozqXYr9lqw9FIdDx
4l9t0kdmALl+QRbEHb6fO1MVmhjVCIPf/vDWlayzzjCOQW5NqUMrrFAP2wCwXZld
qcVJ3xBe5dTnV27vx9PQSoU9IkQLpE6SPnsMxGCGKolPTQnceNT9N4WHgKoaph5y
l3szqDBXdOL4vz6wRs1PN7mRbRYURu+vl+gZ3mIc/u4r+fF6OlCAv5pKrUifnQOY
mhjAvmq5umLLy9N5yvMrI0OZVgiG+pXwUMjTbLCX8NbtEQOGtuyjE++5MNyFgf2x
AcSKyn67ZRalmJ08M64yJQGzRvAxELGdyW5rGpUfmuRMrYcmzLbLtXh5bts//2o/
ogYVRwERT71Oe6XrEp9C1n90Y02tGL5/mxC1u1h+04aMgactLLE64mQc6cn9ck0l
siWRIe0RSst8F6OxBPELb7LbD/JZXs64mGFt6KbFX+f1vVatRbTB99eGJgleH/gd
GlW8zYHxIRtiWiZTr7O58dvWbprQHuE9uBgMkZDafqt+k/cFeV9H1NPqPI+ivbyU
wiwaWEGuYlDBAtpxr49bNv8mKIF0OpIb6rbPI/1ywPpy/xJ7BQprr+1+6btZ07oh
gZKBNQFkVRMzyK92XYPLyUhfcn5EU30n3CYxuxGnZ0Hd8Yvuni1plrqq748eimu5
N1dbKxZk1ddZMhnhUuHz+yvmTG6cENF62IX3ieEMOX/OQ1Yflt2iGR4Nt94+uU2S
L3QX6BYrFrfTw2lJUP0CCu5s6NXnlUMl52nj9l3F/jyfUtcWUz0H5UBLjZTitaRJ
1A1ODUk0CpU49ohbtuTRGWkrD5x1/sOjnDmTiJ3kgl2fGvzwygkd7ahdJBjvxt3k
Nh14ophuyADCKx5R4NIIErtX/zkeZ9HP5wJlRPgyEguEVlD33mjjZ/Xe3I7ZTFbs
Y9N0rGxGBZTZ2PDkiwosvG40SqYuFrqPj6lrK9/uiIh5D3I2+E4juWkzjGkZvtio
Zj1pw3RBLQhzTW3/wF7mhJgudV6poCYg/Ni0PHIdt9QLf3KHMemwMBdvFRia/Wwk
5UhbFd9fMwUMQYzZ6YyUXHMJFkwrHOM1ehzf/rQC1q4iNuuUKJUbFkZ9bh8Hn0Ge
OoHfs4bZNxZklnzW04mpBEh/8IDonQTdAzHTTB9g+V9a2aPO0PYkEO+rSTGfMY3l
dBGjKNHvNh51T7g3TXtuc0WSfYYdLN7K7t7Nt+7qJ/EZcXZjMhBX4dWJqQWffu//
rEb/c3d7Q/zU288yjxXG/3NjEJxyPmzYQMD3kNdN1QnMK+RXDHTSVmqNL5EEtUSw
aR0z+HmXYl6+ItHfGqBA1C5mGpRo9NUBEewm7B3M3hDA3DOEAMErKxvSQ3D0axjy
VuOVJytC+smxZ5YoWGHdXMFPBsqlpzPeEFC6Pa3DpX6SXC5vXl3UGDC/Ptge391z
b0XsDoKYBdm0B7BMPRwUOVSte/LBx8Kbk8kGF6vlledgqlUg9OxOXooQrNTMYZUT
E498YNPZdeAmFBUpEq155gEbeEnHhd1oXigE7kvkHw8wgyVcTo5EJ0miOH6KqMKD
bRMSKmCPVbyoJTyR6NbagHu3Lz3ATvoSEBXNwkOQLeF0tm4PpQuCGY84F7IlgcCb
oFcmZpw+NpYEwNhdWy+Jy28kFxs9cXJHoikzGXjRpFx/GjHcEVn25nvAD4JQtCr4
mH9Mjm9FOtE9spNuiN8OIFO7IexXHfKMRp7vWTeemNf5BSirS7YGkGjLwiytM49n
vxzLnam3QsshBSUDtXRP/bXveuELdfaavWbmp53VPb/U6WwTty9S9B43W3x8SnAY
qgZBfSoh94ykoaTjFxGsnOBbq4sZP5uiRjEZPwWCoWbdrXAagjASuk97U4otKf46
M4mZFMR0U97d2FKDqonG7wYtNwrRpLzpMrS0EecVc5SPOsmgeEJCItXk2uIIVVxM
qT2Bm5YLIykDBJ7nHFjQa4ck0P21AS+/Pyv/YiI2WpJJrGW36aCFLl9FlTtJLj1w
g580iubqHn/BhYxwbRGJaBqWlxDm0fmbZRcy1FAKYNOC+I3zFhION3IFp3Vt/eO5
ylrqwi2JAV2Y2KH6aEuWyP4uUGvInUtm3SlujfUCZtlOPp/S0fYEfe6ZGRBtvMAo
ut73S17GwDS0UyZPSR3ZcIXApxs5jzLAIgjX7HdE9ApdbTVIjB5ID13j039QA41j
7/Gfn12ZJzMU1mPQPscL/6IGa9/bbH/V5ch8HW5Kn5WU/9kfDqqbk9uPKOVVboNB
Ms7C7/f8r64j5vS6mZox7/8TRVjCZ+SIEiJzf5+zLNjjJaJA2YoCUaiXSwe7f9i5
VW1eyYWWNKqUMJ71LR6LUo17WKBWGkhdLumIIpIrJKuEzLTBgPODePdshbxjdejI
jwut10inFTpymYCxBmzaWws+jC8HRbjY0P/i5/apKvHkPz88j2fYxyinaBM5XLHO
dxTVx1i9M0NNrI0CFAuOVOkuqrVCQLhf0M2cccb0Q/b9n8oBO//v+AXHwECJXtS5
Np5QUA0STdUy4WHvyNVQJofQZ2I7BxFvS6bChrg/EHzO7pCdAkW5s3NVkHYy/1EU
I37C+q2pCUXU9NejmbIgXr6Hs6zjVVibPGxrRvKFKYZthhB8KbRgYOVbO+0iQax4
XFvKX1sAkWzgnKerhphjZAUUDhINcTTh94zvNcjod6xu901aC3fPCWJEDNvf+hJY
PxiV+4/8GrQ4rgGTeSgswU1zw+dK5RHapp9Fy+3XR9fLp5CZ1ahizHMcYmJ96EKA
wq2/ZGUPW+IxEWF0kOsq629Znk3Aty3IC1lzRHIoVDtTVg98bcid1EvICbPb+aC2
dKGDdUd2X0gTpdp9KT/tAgigzWS3ssMgsQDF+foUBJtaQqZpA/FWkSiiOe68XFtO
Oq/rV+vt0Y+zwD3Jm56dFj+hh84QfwSuBNTRzdkOzyHy2gQHtHOZ6Oo5w8BVnkJR
tYPiEVyY0M7zc8l/OtTWaHo66g77wRYkkGIKYSfEbrxW7m2P5Vs+eAqOy9Kmri8x
/hCV84rFH3H5gdKlbyNr/z6BWQkOlBYghAXuNeqcGsiaA0Edruhw2s7s2XxmfkTN
VpXFuvzdZdo1uE+MIsyXlEBekWDofHXEMJcEUQfmFV3oOuuYg8KgAVNsGyUiSV2D
zn7WsPEW+ppt9BFz3uj8Pi8qMkrTNIyakP0nt4bdk3ck7V1hfzi4hVo1DUcKrs2k
1gDnd/USNI3hjglZQ3B8kFHRiW2zrOAQZwR/1kxcrTuLtbT3AczGnybePqy4OXQL
WoKMXqk+dXIVQO4d9dRx9eSTNesDA3PO/5CyKTDv5fRgmFmbzO31PIjOWHnhdjjM
gri00YRfAKHbwfIuasKWkw6zkKWCvCjzjtaRHKMWQ5g+WsTwqLfH2cgLYOoQyVlA
tSrcYIbqCFCFqONGN3lx6H+F7JjInVpLI4o9lC0+yRVVZVSEKFPStRDPtVZD20kn
SM7qARj5xlCaX7jKrxSbLcASZJjpqabrvcLkRMZ2V11wSkj9Y/gPT1rtVIkaBSgR
nSFNgpIFyHBIcr/TT0fP2Oi6yYHtyK+h8g2xZYG/TFNGfQFJpTWuYivJm3Z/PnN7
rODSQECChquSa4U0xWmGaDqlGgmvn4lQmBvSY3KW4XjLlOYIAh8j01yaji7cUU2u
yTYYRxumCU2UzoWmIDGjomKtq59Rpwd+h1At/+62G0xmfmEPMfD7Bbu/QIY6WGZ+
s+rduE1hn5JtNLxpOl9/ndu+K80SoU1506/QZX9dTSLncE2nvrO3+h4KLlX1Us7B
I1nMk1W+6e1ipvGLRC4sYOcfaFvaldex+8PRbiGrBONwmFiSOiAX4qoaEF3N5sDS
Cgf2mSeZ2jb2uQWrxra6HsUNiqvb4ezf2fog6x2fEcz7azzQ2zcIqoFKoDc8CCNb
RvIgtAexw3lsMUQHEQVVIme7YvMgJmT4JMLdjR+DuNeGud7pzvHhMNWjdcy4VYzt
g3jl94DwpfCcgILti3xdWrsm6mbPtk9dSyokCPy3zbBWeYBehryHiL8sr+w6Wsi9
R/4w7WU5iudcJYTj+ioHfNHpne5IBnobtbpdm+AdHRw/kIJmB7la8Z90HemYOu9E
YhE9PsMOFxgYmJThGCvNBdzRn4Qf3cQBhDieQXktBO/tAv/c7zHM3ONSC3/5ODrI
nt6TJhNNzzn5Q7uO3EfGEJOXiFUmlB2BfLeN4/nAHh5Ey1HsquiGhvKuCa+taXuF
qmP57TJ6t8yJ91RCGcoE9nuRw8iWktor9KScW8dmgMm4oL2lk0Rzohujq3cG/9QQ
w0wskA7Cw89Gqx0rvt6TuvNQmQHe1mCb+FeQFl1YuqHLqHu4QY5wJPUg7Y2vFarz
TrL+VOsEe6V7gtJYKLRy/ou2cUN0T2I5fkjZFpC1wCeI7MUneSYNdeqNqL+gz31i
wFULN0LJmt7BADf1WB33GMmyKqyqz0NpJyHj8z1SC4C5QdgIssWc1jl0SUWuLUZ6
nLhwu3fRqvga2/Qc2z2qZa80f7kOvY+zdW6MI4gyPICl6Worx8otvlVPf0urzHuH
IKH57cYasIlMhdzBjLoTHj1+WnbftsOx9NTcFX5bsVyuLZG/xu6IkMy37i4aqNCr
1XL22GY5kiUtjs5Zyz18T5V9qBeZTQWtBZP5JNtcyg7ImZgIxXOS6NOFHY6n1fPC
64gnFgm9flmyQDSURSYncLCHNQakUP63DMyZ62/a6PHCiSb2TuSNoZ3FGT8+wH47
LlqkQudgULZ4hY0n1VJ44uSCoMOTJWUSncw8Um3NzhoV6Ccb9+3SVpBbAG2u+yYr
F9W2c/MKw7eClwkkHLsPzyu9Jxc9jDUjrccb1TQR4i8865sWsjdBM5/uFaHYa8Dp
vYgG0M/458h5XAZ4CjA1MPLN2ZK+IL0Mpbf2+hN2SJNKrVIWBM1zMcFhIOAkUbK+
uoJKJ6Pkwt9aXNJRQLHzmmHi0QFtrI806B6sNTqofdzJsJjlbdvB2d2bW7L6qZz5
LVRWAWkGVBqNz1oZxY/LUo8zrgys6GAu/7QdEOmyf6MG4wFgTSrWJBzmt4HqT08Y
KyukxekaeOSrHrtRDv+J1DE/plLZ2CrU/0jFim09Wi2K3gocVxPeatYEzdAKz9oj
tFL5R/4fy8kNjbpED8nBS11pjNkLsBilZIXziV5o7/tisP6aiNRaQi2IV0v2eB8i
0qrHA7nmiWpIYBJmes4q02JaSUJwV0KvWfcT6hq9MuOIBLVZR8FWEVEsC1YkaEef
0drB/HJb7nPLwWP1iRPYNWQ/taVfcAkF2SC+5zNP2knosoJU6gMJq07Ig+ICIBN1
Nu0JbHT+fFWckpLNdRmrNWZWytgp1/XGwq4fCD1KHYWo9fso+q9Jt3Pl9b/tYot7
RxTgIHMml/2A6UbHPXDvfd1b52IfdCzU9O2rZCm6JauXQeahhekdGSt9Ny86XqZH
53RwRY+76EB6skIv+ZTgvF1zTK8cDjIKxfbcUJ7lHm/k7+0dAwvrIcdjBllMC7JA
SBogIPGeYAV7qEDMENQIWMiflqapIcJ9kcdGG660yAxhj7pGSp1e8TrHGU2UmQhw
vY1eRBgyZbMcvwWnVfzZqXOFC+8CCd0OFzJzP50AshluMzV5R2pZ2O7w30VmzD7z
xfqqQKX7knpp7LXMm7uKCyEkUEfPSoUEt1NjHe29JpwNjNlbyKWisi7PS1i7vbQ2
H84saxDG3nkkOXWDCiodSlnHZxV39guGMojEZHLP4QJevWwqNRbywIK+SxkyZ9GE
PszmFIzuTmPxjyrPH4qLwBI+oOykHwA1D4HFqoR2EG6gyjrfY2kSKazz/vn4oZtI
qDaQ6N3t+O4+bQ/3BghcQYprcuK0/Lpsw55dcoNXDQKU97r1RO8zWC8bN8vPsMB0
PIhBWn7XOSfcBYaHsk3jSBY3Gew4jXpfz/gZRopTeF8/MbKbHWWi41Wr9T8OzNQn
66EZLV7tSSFr+ljrD+OBwSNHLMJuwpkVSCM3rPfS0oJd9rL1w583DYNmdTCU12bE
tBrrqSKDPSofPvzJ4R3IRR95V98Sjcdm24uFQhIPHmiNl2gQPSCN+plPUh1ra5z7
DePBOc3sRIKefns2y9rUYcHRDSXK5pN5LrZXakXc5LgA///xV674LaTl8ev3sX+2
M/ELk/UAwpydH4wsXqELIPc+Iclc1/FZA7TC4SXDFvLUBkOQNICHbIe9/eDoZ8gP
ABJIN4s0vSIUeP5QMMpAopTCy+llSq8QjBTHw5bnwL39/ddlvstv7EznDlob18UB
iF4IGeAhB2T89+HOSlaWoXccGo/+TCa7w3DqNJYZ1pFT1QmCWZ78UbLYX5fapd7n
nQiKXRC56PA1IiqaOusFRz+3YgBMPKTS3kAcvF5zNXhORJUQfZ2FeHJXBzbrhn9E
K3GIoqDztn2ZldgKJJ6YUxKedcUGGjE/NJbAMKSrze8a7QiO1/WILzvL+cEtLueG
pyqdb/nHmKe9tJUPDOmjanb1ydnA9Aqnrct7CxHTjfJ2CgJCzxguvJttGlmCVQeq
ngU6CQTG9ISObWcTzSuFUQdxa/98/QG8EkgBtqXxdtp1sw/3LhvvVS3PT7zcN277
tw97bJVt9tkfAZxA8SiHPffHr/OvfWbQ3Cmh8iKD040+JHOUh4xPwmtJXvOgqZYE
icAmBC7uHUEGiYVyMMMNtPsBNrBUMTbYeIKCIUdYwMfcT+/SlOxF3fsqams+3ABd
5M2WAVnuzneDOcoc6anH2g4+L5PAe5UD2oYJlUjJx9ZMM8yuEnpFJnSqSgqdiGi+
HJ2gVbsI619lEJ8cdAatYp/NsBTU/KlFC2uYYIFKXMF6boj1ZumrygbPcZfFix2e
wTFQdRVR+RAadB1goQncer31VVZmZgpngLYwNNfihOKkog/gh9nCLzWSk5ht/W0P
DamPQ2F9jCdL2F4tA0ZMk0wUwLMpl7QlXbTmamd466bSsR960oP436Tk/d95N6q7
BWpL7umAnUxrlfcAHF3T1C6CdpJVL0iHEVTqrJo17/kPuXYzUwUuRUEEmzkpn3WN
MMSOFFh/pZCw62sDcgNyomw2y0yDrMD3AGwVagkXnhCj8mMIDnsK25QWaAh7zuW6
cfBVOKAwjWk+GZp1g8vwlCDH6y4aAQvTxBywSdOtk8U7foIIX5b8Kwbt0Q5UwKxO
9CuWeYimr2yjrqWbsLw98GyBEJPLr/jChTdoRKLXcLx/UBimdPpkmGtxPP7c8qsQ
BZalOVngo+K+Pt+HXEr5QWAEkgFUDlDs7wgdNTMfOL/JlBWRpVN4D13kvh/+Kknk
yFbJhUUUlXBFViXF0nDndgEEvWPzIhg/fWewTdYvOx2rHoX1yYp+t7+67V4um4Gc
7zo81tl3zLqtP+/FCZfKOnd+3uIWPX4tr4nAWCRyCwRzZp0PChYfxV+dc9VdU9ig
KiLapZlfOBTcbCw5C0t2gxM3IY+2xH1l6l2Ye49v71poNfaAZe2c66vie6khR3LM
EDqD6qZAq2dfdbE9NoE7op+of53dkNQ3+2jAihlIsqnhJbKSKP8LcPaA4TF6Mdik
phwgi/c3/rRuzavCUOCkC2NA42nQqUwLuN2oHfXeRiM11hSVcVIV+DyrRruH7dMO
vmJxeuzKo8slEB5iP4tdaCqC5UfbzEIYOIVvOGzbWiM301ID5TiQ7HgxoErm3KBP
CC7cf1MefDxeZE4e2p/7xUC9jJagz4vhp9dDAYkhW7wfjAS40Hye8SH9ZgHf6bei
hmn20LN6umBtImMyxekqnnKG73qzhq8MUuy3gmn+dk5yPJqhCnOKv1GNsVVjUjSb
totUewwsm/iIu/wGhDYuQgQr35DlRGwZp89dfj2CPgniZRc39qAEFG3mLTy8MYJr
qx7exK0U9cCH+bXDtRGzjT1nNSSsUZCK29QufAwLyTF9lOIywYSmCZiKAcRXXbMr
7TEHOXjKoNb0bv5qpll09Dzw8KrbnRZPHkKpWaivhJ+nDT3cWIz6AeTHyg/ngJP1
FTpU6rc1MPg0FQZt1pMB+Gb/RzjZQkCYyVWMhTpWDGym+5y9I13GnXHtowRuI+0V
Tw7/h5UFt4Csjka4ofnNsZIHVgukxtUqmKxUbfzwvulZFPDW18TnEdB44upB46qB
fAOBLul+ceN7yt61HhEPaKmepCQBeUekuHIok27y6wAn/1nLWJAh7npfjvhSWlfE
ESgRmm08RDu/pfU5fKGLvZzbEe/Gzxx27KYoCBgmjjMtoT+qMdXgbSjKPuckBc8H
f4+eRqQcOcZ6GPGopNZab2hmPxNzIqApPRygqx0g7OD4b1CtyxMgsU3mcUv/03x7
FhmrdJNClbQMJt5a5VSDAsisMj6zrlfYMo/wWdi4D65INrOTvhqu3YuV1VFdgWdJ
3a4f8j8Un0LLiZWSUrehW9i2bVdb9vhIJtfR0LWr5hQAtGSaAlUmsptPVaZ5Z38T
PcTH1UGuADPyPVp400Dyp1yh6afWJXxq05llOEXTLUMbPDplL1WJfOlcWumPvgz5
jx3QTa1kqf5Ui5kykcG0yCO21O1iuOPdlpCww7zMn6B7ppJfXbEY3MczZOFotlAi
M2q3+EpWML6J3nsMmOtGkRR8oQARw2ORidgiCObrHGnx9bxbd/RwqI3eyCcr/ht/
+lXWrpf8xbsO/QOj0o1PnKw4/Ga2NWIJfVol+zeHSRDE8A/zrO38+J9gNoktgs+c
9dBV3gASbmwZ4JGMS8uLt+KzjFEiC76W40TUJRXjTkdyafnncmZRIWOr1HKljxpZ
WQoRn9GEfWor+wxcrv1ICX6KQMdO2+xiV/QhJNVmcpe9tcSZGsUvnxwJOluZ/i0e
D7UjmOTTp/W0LwGMVrAAwQVsH8euWmmpMpO1x4NTyUyIHe0SduYTuh61tLuqTlvm
ejy8G2C8XKScV3jFWPUGmUQjbwKy7C70yBBbgN1SSTg+gs9oJbtK8R4QSsEKRAuw
RiqAA8KtkNaeu2sb0JyMom4pxGQh16e4kzWDNxwpq0g/M8D1DRF6lgK3ws25LYkt
b+KW9Du++CF0Fn/BMxqZZwOa6nwnVcqKWZW9sWrc1UM+q1IDyS0eraBtydIDlaTx
j0valNSpyWCQ7AyDWmGI8GlJyMUUgMREgX/gewmHNJhoflByLZfJrMjOB12QM8vD
savhSvMKkxXsh1J16i5l5ijH3c7z+dKBcPG4FlhQnC6meBLwoY8457kDnkxrsqeA
oXPCZ5bTucZgeazNKzEHphKuGBJqU+wf4piB6Bo/jMWxooumdMswFsRBrpBKmn84
v8wAfrMuakGTrOX352ucX370nwtRYUDKKQM/L6M/xQl4JGP5tOKZkMFRRoArVpXB
iITcGhnUUNRswE8FxkA3m/NvFP1jviJvF8wjl8UXN1VAHhETBi07h41/ybGj5Qz1
y71pXahJCzoAHpvVIKXPW1W083okYby50CrqSYFVb0sPmJ9hA9CJWd0J0C8hqd1z
HZegMH61wbn0+lj1S1Dt5MSRfsNEdoHs3eM5v9n7K9FIBx1BPZqpK4QZna4OM6SS
9uzcxUfNkH5Wm4ReMpLqMc+8Ae5PyRFxOdjFMnPQhOcmEkWyAyWYMVjERmH7E+cW
+brdzFOvCPopZi1PLifJJgrfg7E5KMzcm8Vjd5EjJZCt4p7Hn46XhAM3O6JcW5BF
fABm5kaOH5gIX3Q6XBpTBYs0UfAiCN60Cn7eK9BM3yQQqPjdHZcSl6/QogULoi6e
jF4EqWFVV9Xt9dXzNU38De22TgXQHbSvFD1uOdux1W7kVKbPimGxsNauphlbuAMj
oBVdFYZ9ywZ7YGDq8xsdrWrQWaFKJ3eysHtu+Kq13bsQASsk11T7pqIKU+m2ZzLJ
v8DH3HPD1N3bE71DtOv4rlw9xdbwm/vIX31+fHAm7p9xQlAAhM8xhBPZHG7oyn+H
u5lm1ggM2doo3uSYSbiWsuEwmGeHRVyz7txRn3Z0iGUON/eoSZSAqWIOOziGFF8V
UC53XS0nsIUQU+5hhTYPtUO7p6MtaTaXVT1ICYdIClaMzlnsStFNSwcPdciKZoX4
eHj78nfu4FMowx4nMXf+5tf9SVxmUQuXqoHmOvOhXdSVqWWDcCP9cAl7rRuyXBJC
mlQHeAbWGJS+pdiEhrkzIPrbKNqH9527RyjhNjpflqnY6gZ8ZfG/G4YzyDoznhRT
5jrKdMAJeICDacL/fTZD69b05Utvq+pPsxM/uKWJqjTK1rMz/FB/0V7Okzlgw1To
xXypobbzXdhzTVmGNtMG9XOJCGGJAHY7pTVdrMa9NUlJO/qG/XWBOBg1/jK9Pvch
7NukKVJNTR3W+e8pL7z8hr58D6oUpblVcA3yCpHuyvfwQ1BtqpZ4hqHqd1+aFoh8
rNEjYiUA1/7x9XR1Zr8zHnMQD7RJT7zccP6X0hACOl89ouKpccMEwBgUR6wfDHRN
1WdB96KeJRvnltgEhNnElmhkvdE59cWvZRgOfUCA4YNYoxhOFN+7B2cC5x7qefIv
vyz00gB4Xq6HjyFaisL3lCV4aaVCEYjcc4TKAZNvrswg73nVnCNI6HoGUg1WKGf/
XJr9ezS5C8m5A9FbZB8r361lOL76FhhiJnOW/p7HhGlhVWFOsoRrKz3w0E+4yWJb
TXHUAdVjDyT+spki1qIpe0P/5NKcfjn/ehTxLbWQef7ZjuE6jV9dClLbwCKybHvR
4HxwuIxavpCcGQq+IBkTk2eO7bezh34ITcPurUuYHpevXumsJIikjaCqUcdo1Qv4
9GJFLeQJggRco+g2bW5S7J4/IYPvuIAi47T4dJBKNuZguwDCkN0XlvC7uJc/lAet
5qNHnb7ykcd7fYUgJ30BxY+B5ox+IC8N9Ld5rsjTTHcBJQxzeEXzcGiB/5RR2OaH
0mvQbYoriVVia7chwjSVctf0kcsaMlqQt+/28JNKDLRxn/7doYI/XSp6RQzw3Tvg
LsggDUXzPTbPA/8WZw+42ahoRi1uYv4FE0MYWXSlZZPILcQUguPAgXRjJkVyEzcE
z9ugfd43khsqMdgpWUiDx8CLfCnxmTyNeF76xiyxJgUyn4Sybz56ODwwWjGUgsBa
h95z/ZrwdZK0C4mnfHVSxLUYyUCf3HH7z9/XDhewx6IB5SzbCvUaCUahB7Sen2Jm
8abDgavB8ryjODTpPpAOn9oNzSBNi29mTkvBlHCUJZ4IOscsvjYfVlxYSFLKTBpW
vWHFSkDqLvXjUDs7dLkCKzYNGUY/FhZbCnYK27kkSDikaep9gJ+OG9YSTe7mSJTc
DYj5NCwe29orSVEgw+NQ1OGkZJYGjH7OTeXwTfAnCX8BWbkbYK2Gi3ZyidBTpjBO
EXR4iX3kAAilGIz0AZo1aBip2oXhCtdBOrkrwuC/GmuDaslDRbM+JultJBfy0J/I
X9ncWwK/e8oNUw0prJODoDaD2zGvHV9VALZC1DKsyJ+F/k/qa2e+nB1QspuFKXSh
mq7j3IvkNDaoHujaPE1brWtvFganPeVMIF8HIYJMhl2LC9vjCTBgUU00G/7mbpAR
tZPWWQXYMK1Y27o6d0rsIE5icthGTLCK6rMs/kLgcsveR139RkyNJq3hIKXFSzR5
lmcx+kQ2wEiagwgFkhQGhY82857Xgowz1lWa/+m/3OY7ZsEinTB20BJg8S2yfjuO
z6gs/JSG4q5zn6sztn9AybsSLXsBKG8mhFDJ1hr6nLm8bKrj1HJvBKnBGpn4K3xh
EJrOX6en2oLijiiNrA+zARA/4DkSBwpKmIW2/R9PlkzR5Riuz2J8iE8ftnRiPnSg
96RFLJe66FQHs9+/cHf83EHmBOrcL9t7nj2fj956YrDX7M4goejefFoQAkcPMNM5
9K9EubCGQKVWulzPa7Xz5EbAmLv+bNc/KIos05nCU0ktdrqj01EreT1P/ScjLDIg
CPkAAkSrnXi3nr8bnUeokUs+O+mOFVyOKMa+TdSMkw01JdtTDxpQLF6BEgZeZxeU
nZf6h2S4UPxIXkVnomKq6VIQ1KwnTJ1943EwhtlYmM+amL+mpuWtpxfwiFLO7041
yFUWVqh4vW9b6ZKenAo7/XcpmCWo1k4ecbr/vbe9z4WrOJLaJhwVqg9q0qNLU3lL
JU2gleRNQc6LaCzWBmftolEEkaEhL+Cu3kdit1babRQwfRtpWZ1iZILBXtIVKFEh
GKlOLHGjnLawN0qzz6/58hMyHnp59fe5yNVB4fonA9ojR07kyQ86hCR5EtI00jwO
DpQE0sz42rjBc5rTTRR1LahvatxbQlla6tgdrnVwz5CsSWuAav2YVm98wWkhleL1
4XZcXZ5R7K3L3D9pAeXMQ5LSjDdTcBgHrVqk6i1wKrrZZthI7wP3bNaBRS/H1wfM
S3SKygbsNoPvCbd0wA5fkLccBsd89FQ5X/wD8MV105Im2YULJY10bdfk0xr5X+C+
V9NDPzxouY7kJLv4uRk5h2QtqlDAdK4jeopWcQYcS8FXqIzUddZKnU/tpJ9z+jte
S78zfiy63zVe4PGUT1Yc6BO81G28znCRAqx7ELFXZkvIVCva64yw1lPmwiZ/ndjx
wZEtxCLn9VMWporJWm/bMlQLDTtHKP2R9EIrb4RoGqZhm2PatqDYVyZPVKnKxNqD
NKkW6QH708DS7rfdN+YRNYwuGLql3oZgoDsr2BN9jdQPpMSAwbyfbPTIDLWEQu+9
yxCJut7YsaubnnNiTIOeELmqQVLYzJOILEJyYrLPIABnArrULNxgjIkgTBo6Suq1
skwYoG+vGXLrc021asaUZfSc+MnXEaufu5qswS54Z/lKR3DXmrTLpHpeaykhiEiJ
zimKl4KsMQSM6IcQcF329XsihKGidCq0G/FPCfxYnrtoCNZqc0t6qUvNH31jXYaR
IWmg2xyucDojmhSP5BXwjNIvani4BPJuLBjJAXgLeZxV/lEnB2u0ZLKFO3OxWcWf
oxQFTUscMm7NK7/vCa/+d0jaNJh7inswjUXkPtmL9asumpMrOt6EmGmLvG2Hjz9t
1Ow9Uox3+3U/ExaM8te7HFVumG1cAyxcRznnF5/mrQPQC48My9655nKC/dQY596K
jSs5pMFJNvcifVa+6nek6Xp4zq3/WsfDqhuDOQL0IeiafJx6mI0CX2GwkwvKi6at
gWtOnXU4AK2njAqgdh5fKufumPy/uBnv8GqFP/ppKHuYfY1prD0hYt8fcibKTySd
GjrrzGvnF7E02Ryka+5GycFSGwcKlI0dve84G7uNj+zTaF9DLLEQQR8kbWpEaENn
9dOcEchJ0P3yQxRfnndgVXNxl5Ekhgr5ZYNmv7Z82bUBK/PDFQBUo0JA/BWM7xom
zUNmAGl1phtLZwANhMwb9xTNueP4WxjAGYs90uBS+Ol7IUiNKwPeT+EDRwZ2cjzu
PD1u3cf8iaMwqCFcb5cvBRUZZbODarBj13Hbwze30Mq7zCiWWOMrwQz1GEgUnsd/
oR0sgc/hAUF1DvwHSjopV9eNqwenJopFOyV/2yDgEr4EEd1bMN0w4T7YWKUfgId0
G68mLdCJpbIjFTi8LDpMNr5yHijFZUEirV28AleJmpOaNVc7SAaLe+I/4PXdM+J+
vTfi/mjVDra7cx3FYVNVmJnPLWNW2FPNHjmlBVBTnO6J5dCgclnbFS5DV2AL9QNW
R4SJt9MgS1PJyzlk7Z8p4FGLuUr8pPyLeipC66K5XHeDiSv5BwrqVNT2s5LCmZVY
TvazfuMvW0sNOdKKMFaN/IVSObhTJ+PES9she2JbyFyqbbOzSxiTEbEnc8BTbTcV
4mEvZGNKtzu47tv7VZxJiTbYbz4IfjkwlSFbUGLsJBAraW8iNLtfSsp60SuTkhUD
Sy9eNr1nB3YuwvFDfVxyxv6Rb2dl2K6J2/4LBJE0ioRMjM6A4IFkdxgUeaLSfxcR
sT7HEXTPWiWB8l22RVIFk+6o597K5z8SdjK/zCYc0i9lGMMYlLN/tqackD4IlKbW
Lku5WPb9+wTex+AwUMKbDJ0+ohoilloVJpltNrsSp/guyEe+cieUw9nr9Z9FFd8T
fEfMkj/f8yaWenFVZ7/R32RjsE174VAle+SGY84NJ9mKjg3oO/OQXOxaFdJ7p5wI
yfLc/SWyvHfPGBjmF9dG75yN0cXxHJLM7g8rBqndnh25DWXWnWUeEqvatERtflHw
v7qRYEXf9apByfyVVT2GJXkJoclg1h1kqGwu98fb5KN4q6HIFp9RM/8fnfTMPH4y
frgkTDjKqUxrkf4E/e11lUAj7F787wNFRJx7DwfZbjTaeZunM6FUe3BbzUEXYAiV
2LZthHKC2Hp/leGilSUT/MLn9PtkJXd9DgWIp4B8RjkdTrgNDOa8jb2JqXBPohYO
xqpYO5dmCd0Fk+8GFRtVg3OVKapduTgc/DNMUQT5Emvt2paztz7rCl5gaaTH7GKv
uj2YH9q5PQrOUEh5GjgQX4QUzL27Rx9FUhI51jLeqWPWqG1LCE2SH+ZfMHMq3tY7
0/4Ve0IJMo0h3V+jiO+CeUbVoiZJU2aKZZbyCzrz5kyA7f6xjJzFYsNCyUK48w8X
AlpZz3OhzzCR6JNbiKwnJ5uEJTwN3mPrOSWijdgqJKmKXOj5LirK1xzFogadcO3+
sC2dUI9aPAf8saGvVoQEI1DVTlQDThhl4syrCeZ7Ihd0olrx8MXoMeauVSvzCtA2
Ac9UhabbFWqgP1O0AOWM8GplbfEEdskYmAxe8oB4YELB6uPF+eEX9dkNj0yk3svF
keoCEcfx5KghUYOwJEqnLgg5PBcBMhD4hkrmpnB4sETwIq5ssZae1hTnG6A176H8
NXI+/jHg8aWbS6qfN/fGRhj+iKJRkwe4O8UVJSvuWk8/AHUB6AoX8Vu5vAJR6G8X
iKRkXlVTvXXx14msyRwPLyyGMw03ho1nU+R+4FNiDmG/OW83BdYGgJa6VefzlALs
KXZx1QlbkUbmzpUsaVTsPbyhqse4u1PARcWVClA2DSkefU70P4ZHgkaCvpfeJNw8
ek70PAX+S9w7TEksDmJW3Ci1xd9Szomfii7G/gLBvrurjs3PiIVE5EAynJyTo/sR
0gSJPfUUjGwwp+QsJVpnaSIDaEvg5qvyrB/xs48caPUzKdyUaNEjyqyQF6H3EU1S
iSSaVCv13GerGPD2wWgv02CeFVLMVbggVqudtgxOlpGJAHOdfhi/DIDEUQLa0H60
ghvCSgZ3xMTrxVmDlq2ZPgJ4dyGZJZ1B/zpVs3hTQvLxhYUl70ZlGwYvalRhetx/
DND2KBuY60fRF94CaIMld4/afdl71oQcpjr0onddBAFzlDJ2nxQ6SdCf5cF58sJQ
c7zu/G9OW9Z6mjsxl0cROXUxcVANVvFFVT9B7jOFXlqBhGuMaxTmEMg8OyyNlA8H
fz8VrjhMDbQqLvtUllBOOxWcnxPGL9ZILtr+ZNHEI1MicyOXoATV9SFJebUvTltp
5l6EVRHSzGme1Nvn7m+srVxBZnK5luEJJ8VUBkp2UJfjurWF9xCJBI3didWSFMh3
9llRif2Z/BAN+3VWDbybsdbNjEuGkxskjvmI4QLWtqVS38fgR84JRuhTZf4eBT7+
p0AVLNBzEYLrbWKfQkbY4i4WwroFPGRG7NIOPn2bzVpgPWfNxtRk2kItJ7Xb2zcs
tpZHc5easq1fb8UD73qCICG52xrpw+1NfeU4tYaSLZ0Mt/PCgEFhkAfm2X606sGn
pa0O3T/863lAMIi/zCHm9nLC2NUO/5jEsWeQj3HAHFoYF3RL/kx8pRh8oGRQoPJD
X8O6hKHffW6RNE/z3gzQ6XS3Uc4ETu0A0/Y9Iv2/ORTFF6ubTU8ztOLf97LVhB8i
og/5alRQcFux1d8722ovBDaf3+WwV28uZfw1Gz6e1zltXpLzDsOSPgq5tHm3bgvX
H2LCw3FUgYMiZnoCCE/HLI5pzGa4ZKHi2VIsrOqS8Jg6kESs0oD7wUe3upUe+nK7
N0Hjurlw1snyq3/ahAR1bqDUnMAEKP5mZ35fkvpr0SuygOJ2dDJVZNxN+oBBdlGt
wkQDpsJW4bC/M8q/ntU+Ar5jOPLfm4pOptUxA95GMBox9qhesDxnRhYAfCp6LaW7
zHyyoSHVnIvyz/YwlE4d+E3zJFxcxYn5HDsktaeGWzJhSK+skYENjD95wo5R7XWd
Wh0ctJ3f4UpG4bEkcXsrzSqUfjwimMvVNn/hoV+RFQTVxnnY6aiLDvH4vJgdb7b2
FnC1mVxWI+m5Hocel+Pfe6oKT7IMk443djrlDfq2IYIiN5MMIjet0TYjq6xF/fTe
hsHs92TR/A48C3F8j9QyFCpIeLid3JasrOZLiXU7lj6KvVrPOwt5vqb0u+98Fe55
rgjknductyLHI2L8VFKuFv+VvzxEZ39LzDPrlBqJe3QGMSauXsC1INHv5pHAMKGH
NAkTb85K3W/ms5Ql78b96MRqvbjsDhwfzwvaklHHft7AriyLX0bpo5rCJLVRppZ9
AUrhpL4FP1+zSoAAYrGD8N9IQzD55MZOGG5UMxIWcLuePISPoKRjHRucw7O/rUbz
mLHdyXFuLyzFXURvHocTiH70KT+zaHAiUFXHfZNoClAMox8+KucLxd7C5ldn8ws6
1tMRM6BYC3kgUzOgNq9m48Jp6NdOUqh9gMoPxPBCCR+KtpeqzYC8bdv0i/Jszyp3
tgb4snGNCmtqo18z2nmo+3vQGfANx9jU7Sb1qrJ3n1optKxWPKtktHO3K08Ucnkp
3bAajWJqZB6Io31LAqltIP4fBQ5khd/3XdPUteqFqfo6OJt+wR9D2JQ98wMtxkpJ
68yrebFt/SapAfp5AHg82lVpOhzlrjGJBCDwJsCfvp1v4jUGmin/ROkjM9bzYT/v
vQoLvdUjG5EUB0r9Tlk7KonWE+zfKfMRCPQe3fAEnrHLIJOpCtbMhGnF/bakOrSg
iutbDfX64bU/dzjCpFkR31wVg/j7h77lN7sQg1mEoeEi1+IfktbJKF06adtsPHs9
GTDazu5PtwUnfmyjR84U9zYyoib8sMpyOZurF0BsOszd0Q0pZzOF4ZwumyDC/ZGI
1xpF7TSgUx00fef9D5VojfJ3EKSlb/2QLsMntsr7adXqk5ZZFgfm8oHl7cqK4Egw
zP5idz8tr5fPDAf3Ez2/vTk+7fv52bO715gVs1wQg7tN0K4gMpXb2r4uQ11i0YjM
FwDBgZf2DjEJXy/eC5j0ylQjIZeZSG+q8UPddA1lgqMu2plenaD0X6kUmOTS2Wpl
YMaCJWUEuBK7EoZTJdQI1h2NUSqPqgoSeADtVn54bN5CqAgDc0I+6ZiRRr1NPWnd
rgQu//dsOBMZQK7/yJeMPI9SHGDFdtDNjXGWpXKKJHP6018oxpEcJzWeycBZgdIj
KnuxDF1728fnOKcPFupyn6Ftzxq/3UuKYJK4U2/yEK2uVWO0NRQEACZJIW+3gw7p
dsetQs+c26pcpqSYLuZow7SJ6fvxtnIeGDuC01KB7bc0yfgCKxWfm+qwWhljg8Ot
pKMBPH6eXQquUWDJeo0pfQHvfmuUzG6N0x+8PA7pPRCylg1iJYvRGSvYouiOZvMu
wr2BwjC+jV9Jc4n/FN1ZIShRtUGDlMoafpQMSHzQy1rpK6Oy1vqsasra2Y40rgLh
G0iIigQRHCxNnTO1Djjq8YT9WbR1vjBdvaDxd/1xxOqONm1WRJXx5uFCsjFtvq/m
MTN+Qs5VFr24u17FRBA41x93ewMvaSepqDozJNBKwm1twXeNalpiAB8GaGgOm888
pw978ZtAfob7TIS7Am37/J1dHIQ1LN7vYBN7wKk4TiX2TtD93Nxa4Q2roDSmclzZ
Hy6SOPSFax/eqYqxwmy3lVxunrIQO426brrKXZcf2rbHbIFzojpEAqvGOGFkLS/m
zNsm7vHzOVc8VfeVZBiVxkf8nAnzZldOF/JSLfrQzXxQ/JF46mCBPCm3CqnXtMe0
HOMH7efR6e5Ak2LEL7fQlSrBRAQsc0bmGHmxHOFCLvW4uYB0L3u9pWiDN1xa8Pvj
r0twhgUBH8SG/zjVVMepaHlUpJrOeanN2f/37AM+SOVdM6XZ7hY8+EjwJkHq0ogW
BlOWns+cNJ+IyFl00YKIXLKJaz42zNnmiAgZPr3YN2Eq3WFavu/+fVAwVpZO44rV
+xlKxNDvnZOQcPaUC5hsh6EiE6x1DPyJYELjvlpk9ulEUy2SLWhrsxPC4aGjC0ms
Xhscw5CEeRTWnrK/MOb+GkWmVRuF4a50BpS/qG3S34VsaabA8WE3g+61slskz4NT
DzllJg8VdMXT+/N+F2Rw2VodtzmcLsI7snK9ws9DWAEppR+rrndpGixJvvv9Otwv
xeGg4eBfFPak4BFU00aOpD3PneUsYH7nw+W46Ayktnx5sSjSSpoCu8sO7NnKvZT3
to14ilVDHkyi6lvEbLpJ+Gtt11e1QGImScuk7DuoJ0Oc7/gOqGAoGaanPkjaXE/G
FBxAjevTg+PXPIH3F3u6cw19Ph0sna0jOBOJ8Tjp6wI9KvHZfl/TQ281uXSDKPYe
mddFIav4RKcClWk2y2idH3Q3OkcvQAJ3uJdHgzZfSpJvjtePr+F2Loss8T68y99I
5MiJIHz2ROcDMZRc119q15Hgkf5P5HHbw8wcEiBjk3QOZPB1nu1ukf5Vky5I80lW
slEHK8pt96497IigLGWtC9g6E725BdxO4OqmnHIvmRFs6AbhNDUNH6LIOyfBCHlq
tAK+z9GT3DNvH6I9r/cftM3Y3M3+93dgxTMwvr4Ejwfnd0pfSnbuQaX2afnqV2yr
wRevlQcn4YP6aCde4v9zd61f5AAfGz9xTFF3FZXJ+f/n4DLfHWAIPnRKQJ9K40QV
V/ZxZZ/T3DdGWXjgGYhNfamqzxfncPMVealdIp516KS8eJsdepFwxarlfSppysWh
NqxIP7S4/+Oj9m8a9yC5BhnLvqze3KrF5Sgg0Xs3NMCua0qEfb1DNlHWEeGU4uwp
vH0WAiUlwGtku+Q2CpChcwQ6kHTRXvuovRfqMnuq7N6eBT0SuDwDwsvaXD/uA7Hh
RtwORFKDChQ4696K6JMUGIdyar6NhkmZ5hZPONsvlrETKO/XZfOPqIG6pT8bEpH1
39yym0LzG4G5dKWRa6/VTodxd7rHf4XIeWCV24RbLfzja45y4FlOd9yTRsnJWphk
FW+2Ac1q7V43LHA4Cxe45y22Om/vxywPDlznJt3r9z/kk4NZ3nuVyiO2FfpiUqyd
C3YzR9dI4L2pK1AJsLmxMoSfPBlVEsTPJsdYNdI8bEEZJxBp0amYeJGpVI86LKA8
O2nxU9YBQtbOHnK6Y6QTJA3TLySxAHqnxPtvs7LGgAZI+7xA6JwTEucFgMzBaNXi
5YbsXv+LtTFjIOCTkPJJCkYtnAqrnZ3mNY+godAkPdt4pHLgRb6arfFoGZlfX9j3
9nGREcJQoI1w3vzkkk3jBR7+3OC62LiWNLPQGHWpTrI+zGoZYCibO1yFXYVTJ474
749rr8lERH84OOdM+xbmV+wU+jehpJDxOvNMcPV76bYHRgUIr9uDfTcQyFKM+H7M
L4Slnut8LZ7jyOnSCFUmWeDPslq1BjZiuZ418bSvVGF1XB2e+x7rLh2qnAJ4AmyK
Sgo4+WQ5mbQbOrtUE10MG38WS/ttsoq4pGrPbtss7MTmj2QV/aCR0eBQAYQ21ER6
L3e93gixY454SpJ6qfGmYHfLlyDWQZKsNE238dFEdKnke80cG5T4Qq0TzRY4QY15
1RKCOtHoNlHpJEFdWVE3NTdDPlP5hb1JWzZNtXWU4eiR9mC/1B4H2k0oTT6c0jWc
NxwYxQDpGz8ejdjiy1kvv9KKcV7Ht5Z2gLF2jzzEaUUnWdy3OH+M8hxARgIIqJwR
dNcC7vFUIET2d+qBUZTGGcqdiEtI8fWkoRLVy927QHd2GkDboAREzzZ3nh/WZQqp
3QD8WOSy0dT225CJ9nl5AV1v9A+8mz7EJ28e9CZUN9rz92jb3t3bnO9AdicsJkP8
MYp5m180B+4krsbRA6DGCVaQk2qz+JPsbojjl7T1n+oEX6DmdPMPce/sEh9DT3fT
cSQkytv29gbFwZFd7c98g3vQajQ8PaRFkpU73BWP+Dj/+xr9IT5knhpHu1tdp8h2
bS82ZC0AGaQ6T0vNu2UdxFLrxH7crWD0g3nWJBtpFFcyUqfwZ4wOXern+Cf3KNF1
HBxCnTmMm9SHT5t7pMgp9QgQMZiAiEC5FDhBKTw3Lz5H3eLgdMu7y9I6kZ1Hxb60
5HPXZd22I0vPx+VoGZycbkj2bR8FLu349JzQP2rrUTkPLfNYsDLHdVS8jYOw6qDD
MUV0BH8PSj/uYXHBKGSWh6mjVowrBvnJhSVk0MvDcTfWHCWHL2JZvv10mbSzOJB9
PwHoT/3UEEaEep/gej87g1CEeQneXU7FhveBfR3BMq/WCpBj+TZtJrvn69nNxiPa
OTByfsqA2bjyQiSBkztqaGXuUdFTWjXeeuipDaS2MRhHsGZHrw8jWvSU9YcW17lZ
Q2HvajP39VuEgU0HCAh17ckoUzWjRC4lGIwdhO9UBTCixv/osrYrMPwknlj1p/Sy
YyFrM3VXQwFttiRIUalbjc5AV3VAu9R1PBBa2le8S12nKKYIYZYKy4xQjsLYDC89
vVs6CocUIX/FhxyFNT9dJ3dnRvxiZ7Iel/70uAHwD+uzP1aWSNjMvApE0XI3y3ET
Ad3gZbWNju5lnIieXQzJd5jpcbnsZsdKcx6HN+ZavAaHMkDkKHpErZiUFO5kN4DI
AMWfUbPt0m39tagXEJwwfTEhvq0HZJG4+nq3XJyb5LgUE+Asrjlbxx3RYN5jnffi
VQoJQvwxx1mvWsNLNY4xaRIFXH1lg0k4uFuxetZQkY7GZIztExORZcVm2emE1Hh5
iVW/i80NI1Y9FfJ7cD0kit6n/376/oiwFksuMXWHEX3DrLR0T0h4ww9BFXGVXR/L
9Jt8lAAo94yH5BEk5m7yc1pVQoYdpqmdMb19N9KkThSHp5ekARGQquQJ4iz3QRaM
7oeyFuTH1jKmXyUTQUeJEZ0siaiUszLqRpYPjg7R5tgrvWiqyx6T81NkvjUSy4yV
3dUl1B//tn498N3G4STI8vb8AI/onY4+STAMdlWFFAumzm75jGFbR5Cu2qVLq6D1
04VL5vvnA69qpRRI1WH/7fAWvTuc/xpnf4UNjOWiW04u2PNKrJg5OYujTc+50Drx
zLMxMSk6wVOl1TLG3GN3xD0xCYeLvgNz1vrPSkMC0kmAxAE+Yv6MlE5fnWf8npCl
kXww40sIevc3pScOFxcGOxRQ5OttzxJeZDymASspy4r+ZeWDR/hQ/t90N7r6C9S7
wpC25Y5K6RlbeJTixGXdGT7igjMiHae2TkHMc5/Bgg40/J4J3h4oG7dhAYm4KBWV
uiP/xTA6HLcKWaJa0dSD7+VwA/f6BP5HdbyU2+d5b+N0frU7uO8WqQU2C4174vOs
ebtQ/kJMGz68lKhOdCVXLitRkjoO5mFqxZHbCOAdlSrXc5mLQmf7glLdr0uGeE93
oJxm5ZHqFkf/bqfoJZ9R1SFvWV2T1qMP6uYNV+n96HsJpOQ0Xl2BR+CR/+Pork4d
ZJzxBUUaApLSDa4LuOXmNmX9J6l+CCX+ngMzd+N301rvKAATL7kSuk8FHcLzk2BW
7Mruc9UNvNJ2l/7o84dFtaFikDCcvGRhoHZKINIUWTC1H2Q8uqBuCkl/mLKh95Qg
oN20xJd1THTAOHzkFJ1VuNrMzL4nPM5yqiHhSMIjFTOP5b3pjqUQqY4qou1bD24Y
aOZPh9KyCTb9XGnkcFNwa4h1ZPy37PgJ0mdOEpg1HUnRBGsBE+b+96aNYtabj7nD
iEUrn1REzwnm5uUhsC1nSW6Lw4hmc3Pu0iQLPjD2/DgSxJWtIb9TyJI60Ynpg5VR
QiAtaMfLcTlNAoKBPofFAIOeTEU1EBgCywjn1YgkHu1mPMAkCtSGXluRokBbdl/K
aXZo0AqzCStBvstijh321Ppc3iZJatio/a7Xtvu8I1bfSDOO8EIErYKrtnHaIL4R
8H9n2tLMVuAHurWkhBbIfVPgTV5wTWhAZHze9qesEWeKCOFHVJlOXFjguNUdIhUA
eu7O34Qy6EyjzmpU2SQMXDnZA0sXZsZaQZBWGNMILClgC5Yf7aJ8u/zPnUIEffpc
apqSyynmGA3hA/DuteNM+7Ui9q7flHpBD+BbEmRs2wNVTscMmlzeJoMVBONxWQGI
6AdFJNKnN90ynory766fS68smBDAzD3Y5T4HC5IvyI/VlCVHlhnyUsNuRuLHx40S
kXKFVh0e3LetLiPhXhwkf6eeTgvh9BM959ravFqPjxIR+unGt6Gg0GUXH3yq72oQ
h3HNuO6OtCwljRp9j0lURiB++N73UWnXwT5f8ztvJAnJ4jVeR27mgrx1AEkL4MbV
A6zpgBfo8Jc02KqPeKTq6p+ouaugec8Bm1Tk3LNJcdXm5/4Aw7d+t4ieDrKC+pbb
h1RnFLCZ/g8eGall665AULrwsFYpkZ0YStvzxwiDw18hStUO1jIhuW2P0+YbpCl4
tfe7Uwz+QSCYIZCq9Ow07bH2hZ6npOFGThcGk86lnF6VOSGazNjdbh+0wMJunW41
T9NU3Or8Tc3VHgnHpNegQRHChPFl+EBIJdjkidbYAE0vQmIypZtC5+AQpdAfP64Z
txg0tgTfX4veAfcsgwGSNLFRoNsPGHR8Y4ychTL2W3yva9G2mA+lfwVBn/9aScvg
1SKBAFAoAqM9RouUkp3miVxHYnzeJTBG/TdauZXuYu1o5evvw9UCXPuHcntnB2E0
CAbTkQtAtBs3TIZEhUGr6ZUMgcCSa4ccIfxCx3Dbb4su/+xfRkwsaRvw1Lq6/km4
tmUxSASP42nBB4PqtzSbJF+ysgUx0ko4b2yduvA3AvoE8KJ+DHOj998NiqomD8tU
mQEFrcogEDCmflELirA3Kfwg6U5Q0LkieRmpeujNjkxR3I8nf/5SfAQFfUU4tWaK
gokhaoy87niqSo55jj7/SD4aP5d42tbxZsRPaGyrTtaBnedgZ9Nysvi+oWpjQoxW
awB+gQgBJCDlpe4IOYEyBtKcGUNn+jbXbvz+AZPc1hoTgvinnUIRnZ9E58CJBGTQ
pyoL17qqI1etdJN77HBnT2eoEQurLT7AEQqGLgf0dLkRPhIintY/CuPCkaOMEr2e
71djyIMKreR9IPnnTC7m1baZVU1pBegi1ffybIMTll5ZiUEzuovPsiTUtHA3wOgc
deL1pjD0xKeulMF08M2CXUCQZs2Ob5lJnaLZX2t0ec+PDdA6Wof8skNLqSolz0f4
v6FrJfbZrIyshGlhn5Jei4cXWbuRUztDvuc4JbowhWZ6qkKU/rGWQ4qypmfTAcTV
SM3uNxCvp4KD2PdMfiCbo5wn4i2/Hqk2VB/aJxISUiF8k0cx2qV8IFUX2IjoySdR
S+B0lYSDUtkggVyZQZ03GON1VsEiG7lG7scZt6/6G54RPEU0J3kuO3KF3OPjy6oS
NdphsL4kxMQ8W3sG4y0ul8JEghJiBqKc3ZpfO8U6VVxw4WVIY/P+l4IvOvFNVqGA
XJ/2gZIDRe33jOKx2XLrgaTG3Bfew6fcndP2QJh7RaTj6HAGrZ9g8yLsCi6/u90B
hN0DEK0MYABe3qnHyKpsiuD+vzGijdW4ykTZpeERPUUNiJQtB7E4LUHL6YLUNRsW
4MHGWUKRZ+KLnHRepHEPdkGdWfIx1ZtoRZza9pZeRXmuGPuBa3VKn0k9NyujkoXh
dP+EpUBUEolM3taPU0VMGEiahxJ8ReSD3onbi+4eVzY957PoZUy3Kj18+hJBiYQt
kjzwgcykuuXpPyZ6m4yFH06I2iLIHSs3fD4OpWtahdn8eTpBGTZTt7Z/eygpgBbe
6msVO5WuVKin+BOQcJ2qnl/P5XxI04Oo+A2YN4fenjwURaLojpgMMSoqtPKN6KyJ
9A7BjCZganjL2WHJQ+XrSD/zcwG0HwXIrOtkYys+c1o1tVkizECU1DsffNot4qrP
mDc6+DXXu5WGz49U1VhsI/hvsuHX04zx0c80u2kXSj4GufGBeVcMp9pxXQ1z+F7K
j5mgdrjoxRWTLiC/8o8to6levI8lfItJMappP3rGrYtNg5/blysHDt5S8c2unBaV
kDryVuMcwus8kG0a/blp3r7enUAhnmbr6azXmsE8d1RbR0QA9NAXGaNCj/JnEZdW
3Q6MUNxiu5e4QsC8o5unL+gbh3Lst4xRYNa0C6Z1PBDNNwTaVqHlKSV+2V+mtlPi
PAHx2DYpUBYXKL4sqbv/2hrjpYTNdl7RlnkpUUz/pYJV6Y6ao8yQFOTjc3FPiyYj
EL3fhKipbBnfNiogaMDK0usrlWzO8NObSBv7ZOk8pG6szu9RaNVSJSr+juM+EFZ7
PoOZpb/gZZH/YKHGZJ2RYCz55/ssNfveXBNGlztXks1Of8lphEm6q6igyim6Kdl+
bBNrmEBOJlcwJRV4aF8mwRQgHWZpLeYEBfyJLh2DxGhCePhKnjkere7PutekpOyn
uEBflwaUDl89noN15yiilxcjScDEorJ1eoPrBRCezneBz4OtOcmZ+pqHHTdiFIFR
AgLHMEP3fuNxqeOxJjtuooi3nZG9s1nRwK9D8La7QV2nZoVlgKWUxnShYwMV18c3
uF6PRcXYrPzphvC/Bm6elO/1pk400Ykv/9V3vaw942AkaCurAN6N44jv3eGe3xAO
eSxKEDFCr9vCx6CTO+N6DIc9JOEZFsLy5VYjciNGTFNvYY+Kr0RzW0Q77Gd1Ufhw
h5DUSZjvC8Wcva+aFr6LFlxA87DWeGo6jMf00Wy2yOCBTPDjzaHKECG3ZyTl43BQ
Rfypl7r+tjMcgu5PudMHzWntxRmFqyWOT/YOHbQIUpdyNHocBUIi6r7je6/g9Ftj
x6HMbZshaPbe0ymAh0nwtpB9YkR72ZG6WVT+cWSA90At5yLKRkFK5CNTi4Mn7qCy
Y9ETym6G8bOLLWr4IIQICP8q1iRjVS5Xc2kEPD7eskUEkt6frgUQVrrnSTsEt2CI
fz7pLVESTUtcWl87KdeK/nIS1TrmD26mqZS3R+6859Ta/yTaKABrQ16OXOKuLQWR
0L5YPbeLkP8+JGhnpspF/X4zJwRjCIOh0L8QKDobwhtIPpoJwsuEQ/6W7HqsCTko
vFIhrHwgGBDazfBLUbQgxJNE6dafr+ej1sIBWmg322mUNbHEYFGBse9rKGjRQbZV
DbZDRt3snRJhhegIoNWuKwl/lsJM3frDXlCzBIApadjWOladqqzSd5CMg0+9x0b4
7DTpe4oNxDen2KgAxxo51VEYSMyvdxaDY8vDkGBWwENQDKhpAoJvYCkRfIjpDygb
8lh/dy/aShcKnFka1X810TblWB38xOQr858MIyXfoKaSyYqlH3XisA43jzdDCplX
ELCTv/TbcmuvzADY9PzNT8kBGuqnXNaP+0q0tt9sizGBfczQwtCWKZBR+KlL/x/l
AqTieJzAe1nO//nbZoeTeSO6YszblENv0TD9jIco40wjFn1+LlKvTYyu/0LgUErr
W4ngT+fzhLmMZ2Gm9rJ40btokLm+0RWB9xtsLhLHBhZTkoX8H2heBk0L+qoSTTuD
XPD3CyImVSPIrQ9xjuEuZNwHb8YT3I6/dsIoEP3Aj6BLGAjCNshZvq2GVBDXv9Ma
bUJOoyI4dOIUgSXFnSVNmxyTSFG/32uxz6YoEWQrRbY1opaggdKLKBvLVUEz2mor
HEbYxmWqitgLUdhO9Haep3NO3AMAP2NL2IkXltjgoYfJZ6Msgf229Lrxnwz49VKb
nS1Xoi2jrLeMDihuQKRtYXPprw4/kxrv/wb/1+TTpcGkDLWk70N5d2O+VCLhbX/Y
4rFmR6X9M1La1JhUo/bqbBXOgAteqfFPI//PvJj+iHOEw8ui0IRD5hSsKVmXYTze
phnNwbx2HZhQcmGhw9NoP61SPypmvEjCN+KQ9ZtrX1EYL09G9Jvrlr1sTV2ElJee
sRqw5sYuy99uOgMB75VjKbNSer40jRHLDRl2/WwRfiSX9QjHtyQX5T0r2PgSLCG7
ZtNEP8M3HEDrbeZb23sojBusL7GuPg79CYnOZuTFU1GSERrYgFdw45LpOvBIlCPr
HBhmYU3X9a0qOaB4LZd1kpTj95pr2Ssf2FfbABSPu3timOwnOF7q+QJtmJL6jtKf
pjAe6N4Xa8ZXl2ESzQ3wYbe88koY6uQC0DKdtwdnMcNNkdJQwmWe4WhXiSsgWjGm
nkullB1qXxCw1HiIiJXxQBxyhNjcq2I9BIN9q6ILhHaSbwwXi39H0ZpYrg58Ez3q
ZZssB9RSSrkFZUBE3umRWR+59ytTiiD969RE3zg3Li+LJEgV3e9Zxr+yRHHVjyNq
Hl8OH3Q/sKjbd1y7rOzMlLaxP+bIQWz1YXsSlRFP6Kj1+Od7qWQCt/2UPqmURsKZ
Mdt0uNYhgs8bZpS8+fIZh9SyYMOKcm6R99nkHgbAB8n3ku1IXy+sEyRQKOiVc0QP
5O8ktqFNx0EdUOb7PsmxBC9nqxxkjMBKwvaW8s+6pNw/aNL4AjDlORNrcoa2R1mS
lP9xEs+nFC/blU5plMYwjQOiMebmh+5fDkb/9CCqq75AMZHw2j325dh4XHL4hE5r
vGv53OMqrk/eu7Raa1EaeAhUSaLVuW5JI8OX20+thSQ01DVgpgBb3LXr4i6vwVzg
5xtGZ4yiXMSAlV1spxeg7fp3uinx80MaepGjvsXkLPzVigzL78sRyZ7vXnX+mDVJ
OcPGNQ8+0Ez9ly7l51wvUBjax9b/knptESb2uqv+ex5TyS/lARu4dnb+OJGg7UpJ
X5TRxhaZoPkxpq70t4s34LmfRBDjflVx2abB5HkiU3qtUk8HwFX7Jk6+WDNNFO4e
tXTFXxoYO662vhMFcSHfmnUmJ45gbOiNjzhfWpJJ1YJZc48qgXGTo4JCfE3NbL6t
Hn1UqiOb8llBF38FERZj54/KTgeS/fZxdDIteQOTWTleQVTVCT48iuFTExkI68jF
Syfx/64NrxFEEN+liBBnnGr11IQA2SFBV2VZjZ/AFY+cPkoy45fOKxwrbZf3pES9
c7yC0MSVZsOqL043L1YK5OotLpRfYULd7epFQyGuJjjPPdCwejsAy1oE/8Jk6l+E
HzqRutsuiJdTOwdMtJ16bJuL8E31pvgAkRO+iROa/vfDiZhfMMrsOOaxwgA5ibCO
Eir+4jvgIq+y4JDQEIPI052RbnwMvf5p+TICnNeayll68gZJvbL4DPLhfEpSiBOE
TQFyRYaeq+SiefoTXvlIVS2Tecynf7YI03xfXayF+2v7sWuoy/7WtB4mPf7GsOF+
tqFEMYGFlp39UhGWCtnocXhrJ35ECCBBOAMYjTXGyilBPTTxSq1E2/2bJ69LgE1p
2RjNSU0uo3naSLfKIdZoFgkhozwZ4LKv6bm7Obpq4Gk6huS8X5tt86cVETbTOaS0
b5ERaw8Q3WI+U4KoVAFQeZvj18jE02LocY5vYKtKLfzndT0OlafvBQMLdKXxBTjY
so22jnQBmHDcJ7NEXqj/gmU2GJNz+jerBSJHFSEjSMFl4AUwtukCEsPLtcmPyiW7
+pUk+e2X6AeE7tQRshVCofcI+BovhBW7WmF46e240a2MdD8FfJBwasCTzUDByq27
zf3PxZ92w+W1We520M7iBHpdBfufqtig9EPgoh3oIQgTc2zL0wqd3SpmKbQmVULr
jhHXhl73i6f+k9zLg2xTkLqskhiLPOeysdTHVFd+Rtwz2WOZYuXJcfWJLSQvZ9fM
YTFE3xXUyH5QTIKBmXJEjLCKpkBZxo2xECTaiyzXFbOs0gHyXy7iJbaYc3Moi55W
z5+KxJp5biqJdPf1rLWTkuiU7SmyduULHLLW1I6UffbTecp6vfgJaWUFSFAQSG9Z
IraIZGM8Fpg1bwGDQ64m71nhvcSAqKcarn00FLQvCBDx63FKkz5BgFwB6QXN+TDv
VhtrF8SJo99VaTKQHb1rxJVb26itfwuqHA9vxX6FIfrQIwv8A1pxofoQcobaPXXP
Uj3qDVE6faeAbMvmmIqEJMIzxy/F14s+6is+L0SSSBPuOATX5PNEZzN4B9M2u3NK
qbBmDEYcsm24AywOBamXJGvu3OmMzfOIUxcsVQlIi412imO/FQUd4BmCn4u6HYae
ZbiElltlr4JEdVv1/B65Ub326XA6b8x/FXHxNRIsVsCR5lRCkOK/DXXciuD4BuJ0
W3UDHUYzeEVqd6t5MY8OlAeXDFGoVSOu14mxDBoD+3xJ7TcynAVfGPmwh+JYiABS
yig6gVnhvz8FuVKECBYv0ITa3ZlWF8J9Tau/ksxGn+yZqbwSstbd76phPSet15Se
Ec/9ph/tRqmRn7gPdPmptGPW2CZ6K/ePYehxe58bZP4e0jcKnRR5VBCOXKakshgp
kV/znxXXoukNK3N2KPiTFzZNA3IGU7o9qTV4ZQEMNjrErpFHiAjVUa/8DbOrnbpe
7C51gT4ICzx7q2XfDpp/qGlcau8enwgOaPh4MfegbRVA0wtLtcv637+6Cq7Cy1XR
QSepOAvpt4y0ogf5dCPgUyAQd6jmTPZgJblKdVCYvcJ629i+FdEG68sRFz1hswWg
qvVTV8RC39MFmjFDKEFUCbjxcqQhYP4d/8t2bG1wQdhciFC42pAL+DF6l82B6vfO
p4DaTqaeE0bfrpH0BhLPq2YdIl5eZ0BFtxVAukP0NpYmyau2Z2w6cIC0CLBcT2h6
vhTcFzt5vA75B/EYW7li5uR7i/oOUdo/078EUxitDeE/Z2btTLmns+pEpMckJOD/
hFLR+MtlFzVHbG9iKq+03mrK/J4NZ1JmyYAOw5l2OR2yrkfSHa0DzkDvTcWJWJOZ
39kLnpCckjQyOa6HGtNoi7fta2l0TaaqYYKw8jYlF+fDErwJxLfo8pFG7u1f9Ey2
G6W0yEt0PiDTs4bZnUj/UJvdpC3+KBDMdAhNDhXOb4nSYdu5ouyuhXsEinvO2v+7
I40xgHSuOOMk3ISEpW+hGI6XDsCTkRnYNR0s/i/PeHm65tcUkBfcaCX6qmtZsyl4
iQClFu9Yxeyg5gD0MhLAVRiB277MU2L7jQMM7KUuSRXayPaByb8O/BYwY0HpZrno
6y+zECDHYMmzNBoGGROkFoUEW9T7qtPCzgQZ0aTEZeGMjfb6G2tHLL0WJo3Bx7qP
eDFNrU+n52py9qkjVeWXYnDP8DgnECqVWOkh0WqfrBNvJceOtZYVMRf17zGrNxwR
E8UjwOPnHjBeBwWfogwm6zmSUz4vkb56VjNZ6Zu5qgBwyuOeEAdKCS1Es0xxCGSG
NQTwOGl1qrWE8csTeOpUwSElHstSZdkZPNVVeIWs/jBw5ZnmzNVtO3Y+Cg6Tmp1v
BtG8tFI75Jx/yLv6YpNeyiqC7BAeM48wW230WqNapjsJJDdPnWsaCB3clpI5VbtK
xU+BOR9ijUkJo/vI9HkXE31VIddLeLoWKyb3nfpSYwTk2YJZStK3xud2tkJ4Hr5N
WWzKbpjvYbWkFoXWfO0vsm8lnSMHMZ2eFmmIXwbiQps6HKGZIAeHOr7wSwTLYrdD
O8/ZQmWQCCaJTDiIT86yQgaBIYI5CGH2wfMWmLH0CWPt4aD8BNw2kC4kvA7cVazt
iBVtZeBMcecFU5ITndCtgEVwykw84EElpJ06Sh9GxlUNJqpUwI/KLJfUWTaT6H6j
3lS8FDgogOIftBpzfGl2tCNIu3+wt7grMIdVLogi1Lm8zfqOuv+7tqSgr7D6qNI8
lPP5icBOx6ZiNV5jpsIasmsgXmuLlnXAJQnPowrsc+6J+/hlbDhp06B9SdCEEsOa
ZNmYA8lyEioyZMsNZdNTsjc1jfkGPloiMdMPWnQyulXpVbx6ZFHrDk9Wx0ToYU3C
Zx7u91FzqWTdz5ToPOXeGY0gfbi45xr4J/8WYOsw9b8RoG6VWj4Pr7qpgAq/zPuA
o+0a1o4OWatXRZbAKJzwJid1Bjd80MO6q+4aViaKSSRN44ZB1SJVHcIJUZhjdw0L
vsku4wNTzNG2XkFoVddrR5H7ZiANfaK0QSVEV60+dxOHhb/wvrCyENwH+e1HnymL
AKyNUeymJWAZkQ+f0KeMXAKWaxJC7xjJKlS2ZDDYf4eOrmsywPYN6SH/+XjyJRUa
b0h9cysUD6Qptbzg1rRnfNI1uZ8uZFhQzMPTSyZMksewnoswU+TxzPdvZbMjTFmc
4NeRsdc2fDk7bDVosJcpYYYiaWpjSsSFE6PmjUPCrGQ8WGXUlHIfPZz/y8Ymf87r
BGhR8wk653EUQk9GFOJi4OBM9+UP7UbvQ53788mrmCAMZzvxd1WU+2Je4lIbkUqj
yKJ7zfIVUVPTVa6IvXmfkumxwp5pzDFxcWzYhOD3op4Y7+52vUodbZcvS44x2DRu
tXcLdJWVK0bYHivvpeJd/vq9K+ubML/cFEEXRyTMtvUs4uIojW9rb9Ehcj8iOvLm
sWta94HEo601/EwdBJgWC85MQqpx+enE/P89aeJyuKEYf4hKuEq5Brzjvn5AiNhE
cfK880DufuWU9VdkfigHNU0zrpYYpn7jDdFPyC5pCzjhgj/q+sq63MbjAXnwHOgm
Qilz3t6RjWYWJjnAXrctu+xPVi/b5XyQo1pg+AvOfef7631OXYGnyO6YIYhhZ5/2
rWo2eQQAQ2XeXtiNeivvvKi9NdDFgucf9al7lW4sQq+YWhRtpdkrTMrM7tIgC2Fz
FrvcZRl0nuPkK2eNSU3UmmyhR9/TYyWCNQRwDvIpjFllQxC6Ro6CNTxJMjuqorj2
rIhafDCX5ItcOaLqr9LLyee4O/PBSr0LbXYJiCc0Scaya8SozizfNrVs9Z1ZUJoV
duaomYFrb4mKQped3h3rTcHLMOoOHyg6Lpu8pP/kbLnHJu7GZ79RRiQsTwcv2gps
2NgCHHfqZNFnKRgqE36R4ml7yUjcDwkaAONEauXol8Ci5sVOiM7eXAQNmGpZKEiW
qzv4QDSHeBqt3WxfpbfOAqM2MdZqHU++Na21pRDGlQuaAzVBBNvazpo8+obB7/rC
OLw5fXhAfz0jsHWe3ICyJk9YDkJ59Qy9HXUSpUL+B6EPuB9qTuqd3uWW9dGiiKIX
bG0fn/Ke/YbV3t3T3B9mN0b32c2fKWSsoINTP+X8j7j/3VvrJAaUmAB6gvWpaPzH
GZH2Mu64xa+eZydM3vZZBS4zMvS9Jp0HqR/v75LGRYmZyhWVY8GvZebiQJ1+nF00
k4KmZStMDVnXUGgwVjdidIT3gJ3npkXae3X3lpm4wSMvcePmUGJlwKbvacZn/Haw
hsc9oHEF95YzLg2IekO13qLJwrSH+ADyTVwAFQ/mA7Y52b2nCadhm+U6fGmqXB9i
vFobXt8Zjd1GInOFh87trCJLHkzOVBhke4cYEcaSqo43yXiS9sO7eCZPNCge/b8R
bhv6zqeM2F+vMguxy2ZYqD8X2m0UnLqEAw2VCUUJxm/gPsEeK6cd8WFd0szKAEbd
k3EH5IzeN/rcAYGy3yOTHOqSpalfQMIELEuyUqHdly8619+TDOSA66zGhVszlVTt
iRxiM3onFjTmb9OtgMqqD4uTf8qNb5T/SNdLYROfa8PAajq3MLQE6/Kuw7lTuGzj
2YzI6TZrtRpUZ/5pofs1L0FKqDY10wnIdsJYXLH7SnZad7bYgBMgOZqeiqX5luh4
8Gr5sBWxOe/LGwgLkcEfwcRCZGlndQcnt5cNHbaxopC88uKuseGRLN+/eUXKSBKP
TR3czsTefI8di630eVLMgLhqxQ0UpbnOCHW+MOb55RWdwUM6n4HtMFHnLRRgxBCm
7JVdAQ5qpRalbAc0+ueqa+W1W4oRlIzHskonqgBAt1bXaEQ/WKO8WuPVnoLg4MLW
Me/8BsUcIeOV00iLox9GWaDHH2wOPHBxlT+r2o4bZrTNb3TWvVuiIBTpwxSasn5Q
bUzm7dXHhL5SDFMA775bE2F7/EmXb5ZuD8xNYwpco7ZnlEfMmQLUonzx0c7+rD3u
XcpEiLpp2WK8xa3Mj9PmaGj5sT9GgVXgdEOwWWq0iqLX3Lr5iWsM8siBSTpmxLSD
8t8aAuKnLubPgMWDCQOc8lD3FpKhWEYn+Bs9vbrwOkY4XjLWiktJ4FitI/cCljWL
rTNET7etvCPhE4Ok7id4WQZhDSy6t9ErHhv+7rK89KN1nSYlCFrMdPq9BtTDqG3f
8p7puuHWOCsuI8LzKGWcxUlhU0mtounLR9cn2JK0fL8vruFu3+gO0+RosgeG1jqy
5v7gIZ3N8gjrezcLPfky72xZ6325IfnRSBM49JOsgHGjjNG751VltQTgwdMyNCK1
mBpMMNSlof0Oft9tf/fEW7IUehpfdLB8qfNmkd7p2Ds94+/OuY3tWe3gBYDc6OnU
gMp4eANL2ceksQVWwqiVEbKRF77nMEkMdqMmKSbv1edKrdT6IZWrDLQPQngC80y+
peGif168hrsSBRSaAOSobStPQg7J886q8qijHvSsSUElh7nQ4Lx8/cGWuPdA5DOi
JP3KXdwSPAbhOBrUWXBUmTSR1RhFC0Igy0Mgj6VnRU/rIeUCc4qvTJfgsGLEt5N/
9TbckmjZu7QpjDEQrtRyaH1sXH5KcJHDoV2MKINUHs741cmMXLAJDTlXAktwSzib
L0b78kTI8Z+b9+/aaqsniLCrEEwVj0Vhv3PY8K3d3ECNekgq/xmL8n9B37sKKG/z
1WId20GGDcf8jxRKlGZMzLD/I8Pe6gJArhnuYLTovdgfgnes9f/egMB4BbeCCk2e
pDOAcNrEPZPoaRdMClVAwHILvDRKP/j0m1u7+sl+/kutoc6uVfEvaOES1HBS7JOH
sp0nI+DIMRf3XhHUQYXDzNoO5ABB8F9HXa0TlPMy37tKgzYdAI6B1KJxGFjAvOCG
pYiIQYECCIsG2kk5n5zCvNUwHlFbIk9zmDvGTKqwTTo24BLzpsAc5LPLDkOIU1X+
8wIIV0k11HEtlApIO/lXJo7VQmNm9Zxj3vjhLNvjDQE4j8ru/HW8et+2z7QWZd4U
5AfGIua3SRFBU+4cfECDUPXOPivBKt8Z2MeDuZx7qcju8atbZaodKjGkyRrHdCAO
04P5Ualar7rzeQej6eK+MLJlji065AvqN+X8vBxp/QM7utBBWJ58iAikTnKkL5OP
DyB8hRbNHSUDhzMXcXnbfS6z6Nx4Su1yzL5/gLB+dkggO0dBbRw3VZZcMl6TgkqR
IZn61bu3LZOearhAT88WxGERcXgrwasloGS4uAnv6NqL+yNwonz4T+Er0ZUQk9IC
8MOCyYcJQ/0Z1WexV4qXjMR3t8hW5a7ffQ+vol7HKELRnY9AndqNldncbasJ86nQ
2ku30gGwhIZ/rY2U4FaiqH6v2M6+6ZwTpnuX+tObhifxnMz/0/2PGCh1dWay3xmP
tDFLqpXFRkVz64uEKmkqdCdeGmZK6Tuyu1Z4UIXFdAW0SDfcAESTG0Hw/QNBhbTz
7lEBxn5G5vDA1VbfNeP6O/2f1af006uMqvwA5w3VAg1k9ecSgyopa9Ewh+TJFEoB
DQt8K0zgg5J11rCh56SbH1j56+uHSFlGhh/7/WAJFG15VkgaElli6RoX4n+YxdST
X04GyOYOYU39SyEebYwDydy7SSxYM472JrjL444Yy7RfH3cxPXSz65RuXdwf8Pac
Aclx7zKZZ/PCNbtpfg8/Lko5cWUF5mDpVBKmTigHgv9bze8ci7AcBimIc0KdlGTF
fMOMllxBWBqJZuI5ZhyLk6aTDDqmrzb2kpleA007Yia36cPrU4AM1ql0vczlA3jw
QC/byLlVMeP9utrFUh3TNfw12bZvLpa4BR1KsJOb29zWfhPtics4DR7QT/s/pgZD
2t/QQGC60KfUjVRx0CLsTfKJw5G7EKO1ZnTcIg8tOqP/0ITgKvPgyR7lmF42cuSp
h5CyNz6BgPDa5NfGTFXWY9So/eT/zgVUGwFuy9XWPK4n85HXGirRFSBPY4TH+4mp
cX06x1daf1h3/yJH9635/qZqVgQcG76fg1RTxdnw2dDsZz5uzEjNFwMaGFH8xp6n
mTmXS3PW9vNols+n/8r3SNzQw01ce5TEbJZ2oMXxjFfU8mY/k7y1Zq0FBbfxs+He
Kg8TKhQfkcinP2u6zHUO0RahYq3cS7hCFPjVyQidwjwbvDD75uFoIhuzz/b5fdrL
rdjCBh5CfF1oeKCND65ZIiMcVN0SXtW04ympDDhdlqIZkl48M7Nwf8TjO+PAhpsf
xbjz0YCO49QJ2xAjn8AhlWsRmBeRqBSXl672Hf6oO3HeNWJi0IPURxTm3YYpwo3j
Dz+tFsElC2O0HbN5oEY2DyC8uheGbR1NYcBkHdJIvjhn7TgOMDdzoj9WxKFr2qlz
4fcFQr5iev+UDMSz+qRhuann3lND1YVnsevR8kqlg4SvY/kJ18Ylcx0QeAVYALGw
THEPbk1AguDMVRTXDC0xaWtUxXhY3DEBrYoYco3Donj5fHoHlRp93ybhNLXcs/2/
Mtndjz7fqJWW3U+zaxdKk1NO9y9hA09TPCefEeWh2tzf+K4gKm3N14EF2MSf09Gt
r3DX8Vyht4bLRjacyCEU3itojystZwPh6pFwl3woIYuWaqlbebgzPBwpAg1vpt3R
5k+7AgxUZqMCXuWtPImg9vm9gB5zaok/047ZRTBV/Q6fQJQqH84QL6api78eJ+CZ
wIcw6iXGZrIS2V7HNuoaQ82YxkdBrqJKcKV4KHNYFo9iGp0wdoijmIW6YUw+29Q/
zO7UUZCKQv+tOUoT6vxk1mGt/F7WVawfb7aGoTYJSGsbLf6RQEW9ZZs+GWgIBTQT
SN39Ci+wRvkycOb406tiAEIscZqmGbDr9zRy3SAZ/Ozy2Q1CJva/2IBUPoFU6gqf
rBPjYLYmHL/38/ZafSUDrcDAHnGpiYGfwDRfNabBtTqNXRob6IdD85RL1MZLrBQG
cGnygundkRx2lIHWKAXj8Kl7pwu7j6VG6vr+DAfz/qHUTLtjdzLzuWfrB6+viYr5
WJCGMADXFc2vuwx+y9K6NOkjaZ80Us/ZITRo3djhrmrGe61MAhk4eDMi4JaIBoDM
iLKlVDz+K5nh680esk8UnMLdBxrdsOeuMTzYMt6HR4EPteji84OtWpg4+xsPzzap
+kCCGnrda6F86RmUlSufrd8VzskM6hw6Oj9GvCma+3EvLwv59WGSjMsLM8yEFZH+
167L7jswuSkpnPapbq6jB6d4tWoYc9GgwiEJXsFR9tI56Vbl2l/kV7DpwdCKFC76
7RH1Y8OjXrB/CysZBj4bmE+kOSGJ3HcMwica1s92XxMZiwqkFJzpoUYoN5uJPN3T
VOY4/18TDauPhHWbDfGwim+tETZ6msodUd/S06Mznw++ehgg0Y1w/wwkPk10i9A2
rOoAWYTPw+V+yOdXBfBhDf78hjW6hJ0zioRXR68rqvKhSOxjv1izlolYk4WHYiP5
N58Ua9rY3faBjYlGbGHuIHvhKDtyBSqfwxJAEw+8C8wSNmO2JAdF4pXxELio9s5R
F3VECxhewj8sI6EmCp7/84UUzS5VdzcPp+FFYeVU+5Zg4x6Yk9VXujqzz4H2KVqJ
HcvoJURJylohi/nC07+arqTqgnUP3A6bd6kS/R1mBCiWmOlfF7zfITuleeEfH4BT
5MhxK/cZhE5m7R6PbE6hGrKkWuX55KL2krJzqqBoOhNmSoVSY/fIXbl/ocfECXs/
dgQjjqEl9KXRu4GSelsFBYz4O0HAh0VRGKTgsmWwuNdknUaHfDhcjR9qcvXYgChy
jxX++wlktQrh5bDg2aWcv/ho2LxO9mGH2FwbKJhU5sruSdue0BpJ/9j7ivVza1Ty
v809nQEJO6nM8TEXmoM3bX0q9efp8IIo5dKKri9Rgye3wj1aZudHMewvCr5JMTut
A9uoKTJYdb/LAqLC/lYMK4J9cK+i4nts5nUBbExxkfbCWPKbTz1w+pYrzdjC2xpt
S1+3e40l7iIjbYAJBulUa+bXsKuUC9svDyRDxGWhlZ8Kx/uxY3byWc2BghbsUPgz
eIJnFeL6jmnVwACzgBwYiF/F3jMQcM53cvTXHHx+Ix94RCqjQmK7Sle3jV/Y4lSI
cGjwnb1YhAWp707mfyhzpsKLfaMUM7MjuyVcqLF+agNslrDl9ICvssyNXvRwDWaT
SzRXeu7Yb1l0VmrUOrSpPkeKi95wEVTUp7A9Gmi6UevvwoGMFbqa1Yjb2yK1Zftu
0GynDDZ88bu9vFq1EbcAiY0uaJsJVXTuPI3pIPH8koHm6nrqcf2MNo4f49OjuXv3
1P9OeNGK4R0EJiKyN5eZxj1SQIrseiG7ZozxvzGPNrLmNIkZBQxyAVunsW+vB3Mq
7z00zVsmwgU3cgrFtcAeGDUo2xKNn8McueyY32Vt7AAvk81t2lXjaMAaF/yg9O+A
6v256OkE31mW7SqU9UgHiWbDbWwim1zege9JRhwLn2YFJNmou4wp1acw67AF7/jd
9IqgvR6m39cLx2+PicZOCRgCqOsaIhktJtOInyZ2yxJuVL/zdXwAz0Nt3LPpee4i
WxLPRglJrJWFprIzxLohLT75+x+DEW2LB2rw5ToPT8Q1bKFATR2RPTXSRU4Jzh4R
32GHdSAX3/b5JjbL+uUDb9q1D+etS0uub9pHeTwReVsB0WjBneGJ+SuDTGDIzckJ
IGRSvwYGxKxXeA1O+iNqnH9JfCS2GqWiedc2ki2mYqyORwGdyRKQX0pvHUeU81cM
ai0ymQqjGNreSptS+vSood5X0W3bkTzfE4OhsF6aXdwDWKg91Iwd1iGVViH3m42D
U6yPNMSOkLQZGt+jRgCtSDPabPnwnGC9+inyIrEoEKojUWVwVeonsOdUjdso2iok
xIuxLg80OkgirbAakXpEmhVhodv1F8Hj0X/8vSKZyzw7/AgAdbfhJqqeu9XegdDD
Drg91M6cXvQSacdqf0JJTtERYRzmUBVwjU0FdOJs1pggfdH69rX32Ruhl5Wh097B
ncGMAC3qHVdxswaefLEDUmSv1wCibXd1EtQ4bKvVFzQOIUYhy47DBVwn56cVBK36
Yw4rZxPrQSQT6w0hA4wUG1djsh7mHqQdAO+x++Nw8IFn+ircwdpj3rkmgr0fThGU
WEGd4mAU3UempZ+XqgqTbd4W8CT6qzvbKkpndTaahymVm008l+8d7G4vzaZXDYYW
j4W3XFTsvFEfVdbPVNVaTBAJmaPH6rAok5ZAIJMNCksNlC0Ap6bl+kO0G+bc2pgf
ivsMIxUILVjSmqssDQcJ26NkDPkWNtq9NE1jjPX0thq+Boc7rDzhgEXqXmL0xeza
o79b+/MBOaswBDLTzD2FDdCt4lTlZYL0iEOCrt4kSJj/SNtZiPouwH4euM/AJYmA
ahfXktuh6EW3a9mm3F1QhEYz6H1JOP7RgH+p6W0crY0k4w4sn0O66zkHgFKyieUU
MifJuPFhBKSPzsaeP1tM1a+rbK4i6OX4V+HXqDwaxQTjXNW1TYfCZpjZnjbSrgG0
hmEMJyvelb9rriNw4I//JQUQkAYEIdeY3a3XzUdCFgLTvhTapf3dYVC327vg02eS
C5T1gmsf6IOUAcX+t+b0ANhcigRjdnQ/MNUeO6bM657OgXylE4FJe8H5q1BYCCDT
h/QV4H7+uGLaGCMEVcCoVWzfI7t76R2UHLECQykEgZ9MdKptHZadQdOodvofg3H6
2jUyo6QaDhIixT1tY+LmylJwu1pPdZAzLSZ1kYcYbC4S2E0QlfuNKaNZWUlDVHeJ
Xdq44FJ/Pa5JDyuHsC2JP8L7sNHnnPQjOwhREPxn5WcJqM/EFXKPsybowGCnhoKv
ADXP9IbEz/zC/dV44FRFN3Q5PAb8SYj5F5hGPNKdrjDtXJ1pn6nHupYOti713dJ3
x/dVOAQO4koPw7gIdsP3XR7BDnWJqXuDO1dAw5QoxeErNtvVuxB6BkLSpZ/XRPOQ
BfBc+A7HzU9JUOcrEVdpAfDZUB6pACxxXisfGxPBbwficDd6whfHzpH/TPmiE8sW
ZVfwYujlF/G/0iWWZ9zPvwxYkLdU0Igok6eyRfURQpjL/bisnkZMlKrp0TMx5/YG
g/2Gv8Rlt9bWGiWddUBArV+3xZtMtmWdDCPGIYFFL2XPrze7tB4aczbw6Q0k4Aok
z5hc+nsN7NibqmaQEwuuisBKT8Mv907zIvFDmQxGjDA4j3dK43IGJ2tCq3/R2OWI
WhxwJsmjI2VvIJ/ieTT1mC5yRV0fWyQUx+tv7mMyMbz4xetl2PjAZ21jnQGkNzVC
3cOWeBMWXQ22JXokYNIwU+ctu3khK3JuwjDuHn6WQRz3WxGVVCsGOdD37O4vEbyR
k/uummmOTidOMjX7e8TwLDxNYRwYUDBMCHf9YFP2J3qBJYjEjIldzH0mXr0N2Tuf
eps6Us06+o6GnSsUchNxJvRXnyVk0ok9Dig72rQp+1bWk23KW4fQQotUMxtzXI9w
wWm3rI3pUkqnG3J9eK1jbjHFjBpHHIyYfElqP/uDAxEFDR7uwwnVOxdT8A1hA6xH
lhvr5ZjcFWJcILqlrn0v7lSFnELglX1Yr8YiN15UbviU15RVWGXkCM3SSy/IwPkn
soGLzGDy7X6vCWIU4roqX+JswTC4CDpjgLIFNabSq5vdBfuFlXsmaYpcvM8zxuVV
T/uUIIjTgi6uUHnWkkDaJx26wnPJNOxD6D4ZE6OnqHOBkhdHjwHLVU1H6EMxiRfJ
bgA6u2GcDz72mpZCrRBWPh3uLCc+vEuqj0LKMUWCYqNe+zi12WaEwcEzfIK1fYbQ
MRYaxJbOrtftpT4eR+f8dNC5jNUXCA+o39dQXB9bYlPRUkCvingtFZFOQylP7HJZ
NMkwCTJGdRQ5SUjqGf96E1wwl9GSM1aNVH1U2mkxUWI6hjzK5QNWZ4q/3byu+wtS
zPH66gL3yPk4z8v1tujgrnKaptfoZnSUTqGevTNX58CbiadQCSEsLAJ400CEQnFx
u54ohk3BVu55P/PnCWkAD34qkQlTctN84FCjb65QblSCI5PRYXsg9mOlriOAQRV0
LXOx+1Te3BiNS73PHcKVXUE+rJtfWzhyPDydgDi7D/F7YgY9kNZvjfSvz8F0NYZS
X798Gk8zEFLaD7/S4ydvT7E48ivoP00mUtpv20DDgmt+I8u5B9Wfe4s+AU9n+xKf
IUuPpJ4PeOsvPlupC2ezIO+RbuOOOloXC6LmUprVIoYjBff2vkZ25/b/7qBwFNzD
veO+yEy93L8nxVlt/NRutYDpW5x/iecPNnntSAU1//jvRDHRERGRITQWYFX7vU2q
6Ja9P35bVhn9ATStRegYjj19oU66lkYYpDaVocMoeyvEqlQ5wYncKIxlc9OvoJHW
v8oN7CWyQUfnxoMbqpfkU1rr/yEGVEbipSHhT2F6DmGr235gxgt8sYTulgS02fc0
70UJLA2a0HUHY9nOmRCwAY1Ite5rBWSIBRfI076cqbHLuYXNqnuKgp12DZcl95pg
5BTOi4FzBVCltWjoev+fBWG06n7uP7xLf0b3UW4BzDeCqVxeLMP/VKELwlnlUsgi
9iIfkwFo+OWlFOPmzIzbHqbqgDg7tijWvL43YNiUqTcDBLDesXrK4yCwcj6PCv2S
reKKx89TjSu8fK2XLBmgoYpmosy8BzO4JqempwRpdizWBrgzioxJGZ2luACJj4oE
IPCLE1197G3/5vmsVrAoLhPyzvyWgEKRMD9xxdJSAo8GIrAYdilHLOqi1g3/iBh9
ABCqM8R4ykzoMQSAax9P8JK6d9XGdCYhw71FnIOeDyDIwVxAMBl05s5yGFj7akYU
G7il6LS2/64XIit+oOuuN+tatd3BTtxSrpRZPD+TvDJaJwvfe9+7ncrBDPEp/4Eo
JNCzBKE2LkF0RWGKFlQtguE6DZ/bzTkgZ/rrXzDRmI3pNSyrUfh0B0wc4yaV3V0C
0TAyXLNZxLljjg6dgJgUcmODYUHr6P+Dl+oB5rMoDorskYb2p/tmSM/phsiPUIKy
O47iX4Ho1TAtiVxnpb5l93XJoOS7U8rQHZME/gaGn67CngjjbZzBXD2Vk8WtHGVl
67QE1K27oiCsUTnygEuJiSKuTBNLsSk/aq7M7E7u5RtcD1TmxKM6pano5tQKSXUu
AJEy5llf88uKOxfDqPVMn0Au9plF55JM1LXCb5dxt+79Oxbwa+W8t3RYuH6JeNXD
bVV+E+lZeIlkW2Ey7uMZUj+FTggSkftMAquwPP9d5MUMyzf80Cv6U25CI/VrXRVW
CpGnSlnALRluZfXVavKsq1R25UBR48zz9VUgm7dqQqvjD8LG7keFvI4/d7wtk0F4
q2A6w+pKPkD9yH842oTBX8zysVBMs4NnnSa3vza700mIuvWvlTF9SmUEs3uVEfr+
89n3POnCWibjvRXtY3Ww50Gn1KW1B4SeTyBWWFBB8A7sOI1XLQU9j5iz0ER53+g8
LzhFGyFOJsn9iXjezloMjYdxnOGDFbOrFUaqghLGZKWzAdSfWlBV9PtG9Fwcvf40
pvESs74iMiGcFsolzNy9VJw2C8yxfL+YK4wKRXn+nu/WzUMHQAxvklCBk2PQZqd2
Hq99ULCNjhUQr9g4QdqApP5VPhPeoATdN52AExgC6M9PsVuVmp/Kk7ltamWd9RkG
ZG1wr9gGQbfvQmKYmrP5T3BMhQ79TG8mQ4ZLG2KOEXCk8HPHBkB+UiG1CPp6LnSc
Wn821XsMN0mrXM95OelomHI4u75iOAIGRsNvpLH7HoH0OjVyiEX33n8HgDpE4Hxt
WMOoulMPZ+GVzcKoRBQ0/+m+WnshI9Bc8Vf8nxzmGCGNKBbjZTOYP317Zyl2eIlD
7QgsbC10IxT72e8R2wfFHnVL/u00qzZ5d/MEmPCbSTAv8/HpLb54Qr/vD5p/9aDP
QG5sQj2X/4czDCmPKhfZFqJNl5NL2X3RqUy1rz5TM2wJr20BUE0QJC2vwMc0mwo4
TV8H4C1LwB5JsverhK4OjBxtBi0XZhHCG09M3ayHLaf3MemqmGE6hUwjL8im/gtl
9BbEBnuTeo8TZwlKe1L3m1S10PA7O/HBT/RnURWpX4Rf6Y35BcmA8L4wj6v+hCSF
bkKJPoNPs8ceEzPgrrSYxxw23OEFViCAQm1SPUFWFLFKFAc5sCE8sqI0KPstACwH
SP5HVs6+SzFr72jYtVP5HgBI6ZlEwExaEvRb1r6XNkDkhG7nxlzRcy1wbJpeK6dX
C6JVfH574lYoPvrKm7eJStNRv2zMsuhGQozahA5N/ABDiaUp4ayWFJmw1x7vq5hM
2QAN3Xz1enUtDyQSPAZxDN849FJgDtJXfZzLOyORLPn1iUA5kbPE1uNNZdc4zP2K
1IflnmSCLqY8bMIVvLZBl/OUzhvOMRWB4Fs+pXl99qeWk1oUoUcZyanjHfP/6C+B
MZGfk4ryI2lz4eB3OTbdbZ0zrJnQy443MuYohdv9fWXiTa3NWzsmzmeCzY5B4YwX
f5htCzd9OMiJ2uS4/Xy+TCCPaaInN4l6rYGuGROgWbsp9Q9Fx8t9WeGZTCC+OvYN
MXXiavU0btJeZXTby6aPkddJcQr74raXqre0hLsuirhMgYwVe5Cpb0/5JoSVLU0Z
j+BkP3k/U71u8phwcWhu9UigPqKE82Ce7qqyTU7w90KNn0Qyxc48FUZ+IgN2yHq4
Wlk3rCVo9bi7vnb+ZZWWNRIlZP/A+FCbbguErzZ2q8gcWLMv4RHJzUVGV2doiAlH
SIKogQ8m4T0MIsA2aaBzJn0JUDNG+3mXDqIYMSz4ksq8L/OaPiyDDDAoUWSKF6Al
LXaXHFFJ2rq/Rlf++HBVJ6/vkEDdSxP/1WPwExiAx4POnT2tPa5R3ac+l6LK56Yu
uZO/nfCvpr86F+sGjJsABR04CQISWjxdI0B9aAmXO57DPVDig4pDUSsmkCifsR8H
mVM1K2ZfzFzKzyToFIw1khlymozTszA0lMaG8d3GQineEUtBA6vwe9oQzxTLBC9y
WplZJg5Q88b5MlSVbd50QM3twFYG3HY3/KC5Hd2U43NW03GMPtFpI4vclwPsfDW9
rujQdYUlwmQy9S8XZrwJQ34hgOXgBsPZ9+et0UXfms25RStDuTRm+ci7QPm7QuHc
eQMYp3UxJOmTVL2zlez/yRE8eXESKjh432e/mAWK1wl+VGTwM9DFCj98h2zRUd2p
2MLUtvuOSxT20CjWqBSx5XVOyyBdbstB/xeq/nwX/yal/Y2uftHsmIZ3iPopE8DV
56hIFruFlHSrndVQtWxoD/wZlkkQpTaTThK2/9mxo4L5KWnQXXuCfB6P8PtFkPFP
S/vUxKE2AIFHVdIx8pFl2xWkZ4GInSrbrooWbmd9CsNvUlEgRpOvCHA/CQFF4DES
VMqKUzV90pTifHKRw62ngdG+SBZoPfVVCnkM770Omo/ng5s6BRiBHamm4GEhIJSr
ZRnuGkxDgiY33V8OPqOAO0k5VDdNdSdOYudjLFmlwKxrTWi1Xhe9RR2I6PCpYnFp
IW3WVOmKsXO78iH4+BN1lpl89uI2l7FM90joJvypdU0GL5hmQV1U3x+QHAKBrreb
EDI0/IxOpaQD1XY5SgKaCbMNuLaUngyM4qsnQj/u+AgIiDohnPL4SY17wuyXBS3w
OED0vjRhdpPEAbCvLYNeybPKVay5lO3Hfd43FswVJtcpO5Iw+X7fDxQDGF8lj4yc
Wej3DCFtsc617lgE7nkl17bC+IrmRum3A6wGPJgKX3eXcLEHndIkafdk0fBB7rO+
yYQJnWrQsU6XpMwbIrtRciWRqiaOKtqNQbB1H+0iQ0ALhLWEeniHFkpHLNhIDhsk
bEy/e3BFmYZMBTsVFkdFWNLTlVnWQ5jaFCk5NnewqnN/vSHwBmqaypJRhNR/0224
QuZCP0w81UE0Jl7K8MUMoIqO+ShIuyYTARq5DWQtmh2U7MTs/KE0x+hqcsDC5cs2
ztcglhk+JCAMYPcL6KjmgBSNHZMQGklvtC67nrMSQbSNTCab+j9QO9tr1QFRf1xj
EDooShxlISTs8cVhdj+7HWGl38KWS3vERcsKkTi9ECz2WOi2w7zHhAc9y23yQmyQ
n6xeUlDw0t/rjdBJAw65DZoyNI3sppf1tyuW8IM099YmQO4ZPAN/X9ycBD3cPjs8
QBjET6A5d1AQNmPdvXo3hQzskKGE3TEiDY27v7uSYaU0HElZ/+xMtTB+6kpPbsgZ
zLQ3jFouf8fTpPqLN0bTRwQdNh2qsvJo2L/VWO02k50ve4L9ddqwQm2HJQBKkLne
kSOYfmkUGLD/8eL/8QRuJAG/8sv1WS90bep9+cyfUe3U+iYRYvUEqzWRpAEzwITE
2Bjo8+qAuJd8W/vDYjpR+xDpp1PaSuWKJta1me44x/MFoyeZC4AxwW5Pl+MaB8lc
CNCJJO1wb/oTClSdMZuJJLwFM6KrKqJC5wIPz1eNKaHN/GhKkzElQfPCsMkXzrS3
wcKhtFAQRpl7+kXVL4AIVvOWZIpMDR9Yp6khYz9zbYvEkY7GZaJfKFlsf0kLAour
1MWtpy1VCucOlCWANHB3kw420AewiouI4xUJQGFEwuwOR6swQCsh9r7AI9y/KQ7e
yXcKgLaF7XGaz5aMohyZ2liwpSXu6mwCce4hzzUex1yU9UW6PLC79quop1QsPa3w
wWO4pMzOTBDJzpHVBVZ2c5M4hN/WZAeYBA0pa5gG0NuNfXbNp8vlPhtEUBRlmefX
wALhZOx6LgrpRoGoxXO6i8wlC/Wio0bdT8PUFWcoJ8Rfh1AQJE7GBFlIHeAHdrrg
+FFM/MsaI3lqNuXP2kfMONfAUVpNTjD1F5dAlkB5rrY3BLZuBjWawE7PW7JFG2Ia
JWphUImVxEAZFl6vSA7fPnvj5rcmq/eREQZlxTR9Doacx5p0dCFInk9xjuaerHYG
yzuAw7lYQBrthQtG22QIe9rSYHZdqrzeyUWelAbfbKUjMDOOugUgI/1JWpFVQsQi
9zjyJnCblmVVlYKeU5uYnB33cEEqmqGfBRxKLa4Dgx+1v0nSNpwTWlI0hXTEmKDm
9HKjFGfr8/qg6C9kepkW/54zptKXByUhVRTb3H5QVIz77+As0Ak81sxhuEISRU70
gCsfk03px5K0SB0Rqiv9BLLcKtBapmXit9QCfN9U8hekMsN+HtPu34XHFm8ySkNk
3xaFn/JoewpYbaulvP2OdoL+UapIYN2NU7qdYSgQ+Pc2f6v9E/Fh+X7Aktot2MZ1
SD1VXnSjYaOSRJgRzP4lJ6ypEYU8oQQCKFnxw2wWcEMZMiCL/cbFHAWe0VBmoCUo
hB/k9w3ffCrRWAfTkmHIYMj9NYo+OwyaQDZl+zI6CuDdHGa9Xo7B5zXHN9Io3CVC
4Oj83QgACmDIqvtX8LrfguuvbbpLmzDP7tvJO/yMZKMX9BpLYtgYPRiLU9UYV6wn
QqDls8gmtw3sqdbkZenV4oQynxqXNJpwlgglMqk0/9sz7/yrMxKLfS28I7qvNC7S
1waIc6FAS9MfCabGkuTJYoUbKdjsNe040QmvwHXmrlQeRm2mw/7Fv2vU4/NVIhJK
HDkBDsCWSW1XGwUlwizQiPuROKpcXhZz9d7iGUjOgBlhlVTVt1vu8Di/lz0YiW3u
yn/zWKzMbj5vYB92WyV5PdomBtm+5YxYC7lVH2wC2ox6cWTl8pNPDf+Zi/G7qvxE
HkpABxXp3bJwhyjKEe4MI/h7S+7ZKrTTURqYFXnAMRlSWGA8PuzAQZByFEiraBBb
LfmIZIL/85kE4Bhk/aaJHL1iqtPklbwgx0RBsMy9sdTGqlaXq6/oExAxknlwrWS+
7lZ6cdAX22lF0vowjm5KZfnuFTgeXC2LouNQdabKOHyfvfrXvc6wBM3K49sPOYFh
z8QjjoAR4FVAvF612L5BSWmE7qh1vI/98MrFurp9DIFPQevKcdl55puglSA2F4pe
TZwFGVhNz4gWOPsmSEhYGg/b+kCNwV7IfBd4l95bBQu9tPW6eV0acUMaKDq0hWKV
nrHAW6H6MRa+wRb4T/+INiwuyxeW3F0SuJRlnMyow3yDNJcAzZG61CLtmo55XqHW
1/d5PL6779xhhnhc7Gl5D/YbPs9FtHwgpG2t4kaGHEpFitSaNj2MZy62MTWYwcLS
iPdQmEzzZLme2YQ3t6r74Mip/wdMtvEnXZ03Zn54tLtQPvocIBw2No3ySIP56+zo
KOAWy0UyYmZbNCm7iHPhSHvAhWBY1e3GvEqjk1JmMLuWGrpGo0II3pKfx5apSg11
X3Mmy2OHIXQYf6AjWmbQDmRLbf6WVhmXulV71m2iTmH/rHlXN5IsnBdKHWig4ynv
CgwovnhGATFtrvEl589iDhuM53UXcql50F9kbCQV0qmqw5/g2+eWcpC+PyAlEJoM
AV3kamJLDNx42biNQ6pQsLtr+ArAI1Tk7DCE0LqkorkCWlh7glYfWqhLSpPLa2ah
1gY5ZMJPeOesPBbwKJ69t6sOILGvVcjlBNsMm5yUo6Wq+Lbr8LX0M/0CKDaSqOo+
+jMFCDLusVFPX6bRWT8L64Yl45K7xZV4BETuImlsRbeHO/kbE5FSGKYsBieTnweF
+HRCNM1eNoctXVF9ZteUzQTSiF2UzopjQ/p9X31evSBZm66SrdlrZMsJJrQwHP7u
S2NwAUo+RqNau18FVoC/wT0NRwc8sPKVP8dTvQsQxoo3+GkD6LONImzrjw/EhGdX
R3OkxcflkodAAlSokcT/PMutUEFHC5/0YKW4bZMeNZCC5NWXlTeZN4vLH4CVb9fD
71606ieR5o/XMeMFGOkNp6x4r+pUIfu67f1rKf8GE69oKZZ913Q7MHwV6gIyQpDp
YIZ4V2dsY6Zehn0imL6dmqwofdSqOiQgiW5evUSxQ/cnC4KH5YJY3a0Ka6fpKMm7
c2E9ICHgXDPzcCyTpBY6mA==
`protect end_protected