`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
ddtXksX2+yylW5zu6QL2Lhnb2d1sD00763mmSITNX595NcHTEkwn0zB1Dry37fOW
FufOhVzEJp80NC5qZ/+F0Vk7Ik02dIR0elf3clrjeJRK85K4e3Hoo4xn7YbFUIms
l/8VZSb14+JVGURjfswrIyCUotIzlzVYZ6gzoZwDXIi5gQIBf/gI+KxNXPaKV+PQ
Ufys/12rjO6aI/pPlqSm0hCvftmBcnezN2hk1UeXgOIuKZnogjOsf0iJVX2aOOWE
6pD/psybjbnsNB6kH5uFTA5frkzIzkzl5d9+YDm9OyC+k84E83I/7/j+rk4L2dah
QJOvksSIzN867/4Qt8qYTQ==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="MvBXkzurAa5VTw+1JJ70nePUfoQXBvZOku/SMmg4TwQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
oRtzZL4VJ4iwysPsC8SXYCzXS8Fw2gtZTOskLcDV+1B9Nzn1zTyNtlo6lNICRmmK
ZRVu2BmCc2G+fmzynYlNTnSa7C0Cuel6FYpxCBlOuk3OF2tzAmLAuDyOH3Z1Yjzk
a0aHuoCdIRKv7BrZCdALt03JeUmXKPdOmIlkVGFl8yw=
`protect rights_digest_method = "sha256"
`protect end_toolblock="Jn9CQpRhJt4rnzZPRk+dOpzAubz7omckX1MrFd4p81o="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 16512 )
`protect data_block
gD6l00tciPUa6pDNTk/+tzLxvdHE2s3DQL3/JqqujQBC/Ei+vcAB8wM3doqg5vTg
mdfn9XB1bLOis2CVSfu295W2DNwHfMSTc/8BhCDRnTlLIX0UCJs9Za0+LoM0rMrV
T7EjVWppbP+Em6PkVKCwlmIQ7JKaifJ+Y+kjw9HCGboYo5074hY+K/CBbfsBQY86
DFekqOo2vgag6ud273wY66ssqLFwaYFDrN1DYzXTvlHUl6V1yVrebVvLEzfSesBc
A2eY5KhQ3LFYcANjSTM8SXhbzfJyWNK1c2QPfMcFv/aVcAQNVOIczIdr5nnwWfH1
LIAr4wvOgfqu/yovbfb6cptPKW7ekx5FYMApNsn7kAfZVPAgcwBt3qWy4MJr/Swd
qeiuJ1dVoMgkpt7Y8Fbds2jr+uPrnlXZDixmtg6iOFzz7gGN2HXlPRHWvJipDqn0
xR4pLHNr4MlojGSctuR1F+37VTUyuIQM23EXqz/86dSh51ePBpQCcJfKNQk23V7P
4Jgbqu6jJb6tK0FHySXKHwe7KYspLXeuX7tk0mWLQH46OqXmLsPe5BaTw7viCMmG
zL7flXALmxGbegjPGEp203hOgKPxQ/+9iONtfCzOrBnQNdleosBGhG5+BCub+cik
3AJYrk+3PK1oFY+t+yqdjKMuWXai0aDHHP9Z+evhh8Y/oOqYriYszElb+eTB7k6N
K6fMExRFUz3/xZzuqbxbS8BkvNY6lNtLiSgV3RfNbeKEd7HkL/39xuW11pz/8cMZ
96L/lodFR3QyRzS0BZ4Uu25+C8klnq9IAvfot1lTu290T0ciRM6CIhal9fkTVxRU
O0HZL1cQsvKy/e5jorMkXM9i0bAin9yuMew71KEKSx5ACz2EQtVREoVQ6qQ+wF9z
AtDinMSWp2sYnIM2JUrIGxE75XamlpxNNJ3t2K7bUQ4qbN2OMr+8GBmd7ipIuG6s
sDARsAonpNi/mNSb8nJaCwyN5zEdCVbqwnyiL2PwAU8wyW4S1KD4cIqYS6um0hHK
9V4X2ptM/XsfG3qiPXlxCKcvptd2IUt5K5Gkza6MRdLUn5mYj0gvdRiVBPmQdnAW
DvplMggBi54EN8CKhCVSRkvSJxVO25zkgoiR9D+l5lZ4hJ3bHb9kAN8OxhS483UO
QXTCmQqD/evlv8VbXE51kF5euxf7MacLbIWHMrc18LsrRk+nFdMiaEtyEBwgZ0dp
NhWi0gM21FYlrJ5tnpshPNBc/EbTCH+DsYoeGAHDSlV3Q/GC+a7K6d2p+8843yoo
GX2uKWSXlQS23fRxi41ft4vF+XRBO1hS/tT6a6RxOX29k4CgKAnT8KiePsmLz4r+
kVwm+bJvfbek3L0xu/9QnRsLnhal9Gi1nsUYIgBoDnx3kCPgqu6GvEDnjkxOWYHy
PQT2EOO78STzcc53A8ulFnrlLGbQAc6VyxNQeVTJLxPIlmiV9hQ+qWUz7HntwIV4
7nCoAEXodUQeVO7+WiUYpqRnD2CghgE94kfbPtY3qC3Bi9lhjpjDVk/wyGLB3NdK
mxx7lez9EUgdYTpuBHAYfbzuha3whx7Wh6kOkWMLeNBprj8C672lC1XSosPcfL8Y
EGIcwn8sKX86tJnAsE02mOjSjvUmp1ADbwY7jvjMwHGdNqB02LcAAKRX9e7Duu7z
LpOEBA+MUlxMgFwpsn3DnHDxkC0qRWt0qvp646LnJw6eIHhW9mLECtunafvoJsaT
CpIF4yn8TQudnf7Z3ZYQYMXpDEMriHV6JZTl8IkeVsxjawfiGuwslYFwjFU2nGFL
psSKGbGs3hFrQoOJsHUr60B4qQx4uZ43JxNaMaSrTgEDIXdsek8aQpIs+VZPkjt5
njqEN/eh126DyWrxii17Z4pkcx2PdKPx+J0k8lBRgsdUcSw820RFVi46vgCgT1qH
Ww3kKIJtOmurklXidzoL6+Ed5pbp2w59hbcov+dqgqLJdKYgnVOPXDmuLexOXGGm
NliFqpegmLnpJGt321vaNdB+hKluEuVJ/NnnXq2YwWnZvA7oDHcvklSQtSh2Mmw8
86Lij3Rx6seCLfqK4wpR1q1LrZqURZ2jsDoM12Mt8Mq3Wcf9kXgNA4tV5yhFtcI1
a9UoHnXs+msDE0r5gD+WPhuYTde1GfdNAV60YvjbmvgfVP2QZs3yr5ZxDvKpMGoE
FOTHRlbiBPecvSQvzB1aIAFRrumipUdslLPhkWGgKCTiOm3kXmlwDKwml5aiF2Ff
dLH6045k0vrBrc2gWhasQSywJPnk1AcHt+KtDrfVslZK0zoGouRzyd1kK1PjjMM+
0TLLFFxSl4qWLIvFEq1R51ntoQaGqEutTyeCZUTPYqJpLO+3ieysZywEAae+PlDD
YuWBfSdBBDo/sIBvD5qKfR6v2nShC/FKNjU9T2XvrJZgMwN0ak+9wHDyejXDowgO
rodfGsVXIr0cl9Pct6i41K77lt9mmGlzJG+NMSvaQ4ki/tdiWOeFeQmcOwxzxPlf
4pBNE5iNXLedIjZwE0+KVCpo/7U1CvSmAGkJlEXc4KCMV4lGEG0aiDAvQkZeKCoY
CFWraNtuOVI1tRWAj48M9CK6UphjEG5EKV4M2erKL4/GzgVqKDL2osvVpX27sjQf
0BUw9ACIo+MAmCJSQO1lMSULdPmBvBZD4hBrE2IGiF0VgMleRCtJlISS7LxGrVdQ
rdAiDUqd+ZT8cQw3JI/ZsVsy00k0JeLig3b9Tof2OC5WViByQjWUfZD0Yq8HXziv
jFABCOL68R6S1AUIu1OiNBbVLno9EeMNlVx69GrpwNLEzqwbqouH7jCF7o8rA5D3
gPdL8Fiqf/NQXTAebLGB1jcoP+U1KhjBt3B7wFLg1nYlMNXpeIIujjrMiWJVyF67
C2lljWsWbDn73QsmX6krELEi9U7onEL6JpervdsluwdQ6IWXmn2lVPuKPt7W8Tsx
A0zKq5Cnd+9c/XRs3Wli5DR5srohuv/7XHGf5C3e4Xm34JKaAWQS4knKxouFt/Uv
+JucCnGCC2pYWE+uIR7dOX9bPVRxR8/M4Gkxa6nQms1NQhNpuhDtvUkJk1yKzyX7
oXVifUig45ZfIuj0IIRB0W7yIQerx6Gvs5ZVzlVBY6AJZ03Dz7iacThFx+csFV04
3N28iELrA2xkpFDMRMSQ57hmIjoyuKTIjQQfhfGuaMq+4nQZSC93AaeK2gktgPJF
WLoR1aXm3HvnePVxf1ei/0r8H87X/HlLlGK5TB4q/Au8khMNhL4QF0/Ym0zJaxmH
4o9r6iZJArvkovNN5s3tUz9k9rhmaRhindCYiFQf1V7zwiPbYXOshdD+aX4Zj15c
AaKioMIf2akylgByZshpIz/+breqUQGELAhtqNDfSpYSxUBTfDUanIIis3mSb2vn
nFPg5whVmr1/W7a2Tuh0nOMtnxPDxsRpptfe7nKvaEy1ozdJtHSPMgeBQXfEyMGk
f8U7piun4UEwbp+2DYPXBaJ3PoSRU7zE/ywk2f/51dOfSR3rwG2qF2iYmHp8oAkM
lt0/vJnkwDq31dWwjptl6cs1P3524YthkZ1gC68HdnfCzwuz7GqpfOdBQVd957qf
B337QcZZA+OGYsazdT3kIHQ+sCkIwW4rM/QqHYSwrQ5OXsHT0Mzs1Lp0ATo/oNhO
b3M7LbfLGKK//GkkaQDrcrbTlb/at+D21WVzP4k05f+vnTXbD92KXfQkUXLtLVKM
F/lu1NcvwLh/vDHHJph/Gv8NBekbdxOWlK7Jmi3jZoAQITrfW6WHViRVZ0/mq0Co
PUEBRV72HWS+SWCvUjdD/Q+LWtryOmMfm/iTzYlvy2Me7OYrL5T6BXd8nGMXo421
Sq1nFHvMlG8kU3yz2oO0d2O4xcmgsjlndNI+tvPqXLXvl4XcTWQUP7f5xNOqfnJA
KnRIwdkBwRSnc5iMCHa9D0lNA2Ri13k57bf6NsM4aTbhDvYAFLHvwPBV2da6NqF/
7iicxpN2smZei+zm9rVw3c/6SOkn854VcxFYW+/WsxYLoWYrZqqaeHamApbdKDPT
aBDHT8D8FaP21k5PiENuaUSVZewT7RJzzZJwQ6TzhoFwjcY7Hz9jZXDPkGBOhD7q
pZnT0j4IfarZfRtw2aBlOe1mnRfAhrKtWvdXxHLOEuRSynZk3ei2nsb4GgnU4tCd
EXCaH/Y0vuEfTRh2H5le02Kfojk6KndJsORftEJOgNTP87MdV6LKpiqJnkFRkkmS
awxC8tjNveCCzZIx+jLbTryCjL4A6iLKZo1yFUXIYnq/gYpMuPXtUigzAcptifAT
0qAPuAJ+OIexzji1tktYDJlbanL0xrArGVmItOeG/N8bfRzaZvUwKBi0aDt6neln
INk8WbbL4+rQixczrW/L835R7NHRVTm0dfLT3tkeZD+vk+qylADZ5KWU4zy559Xd
hhREr24rY1pzyPZ/A45PbnuqzkWlj9fwrOE+SLVdOvPt/nuN0EEgee4Uo/2O6LhD
fWmI3uptSEmbfDTmwM2QiZluXyhCDfEpxbfI228A9J+qhtXx72SDlhZXiDFUU1xN
vfxfEl3lLYqe+O9mhEGEtCMxJDS6xKjUYKSjK4E9oYmWhr8NGke6BoB1MldIRKCR
Sa+A1I6TrM2iZvsKNBj3uNlDkpTVIhMvQY5dZ6QCPQ6FJIwA344v0HGjShuIIiyv
l2p7h4CGPHJ0KGSHryIrqaIhrdnrK69LeryiZha5yC2/cO65kYUYMJCbF4DKAB+X
LDdp3GlRPxU/C0LytwpWmHHxVWp2rolA4nYG8UUVcX4G9mJjrE6ez1Ix48G27sGv
YBE7ONb5/LUZnrPD4xJKn0Is2vPadBtCOEPJoxopY7POy7w6N6uRUMxdHkwo0jLh
Ae6f/uyUOlWK6mXNDawkxWWbtbDwimoYL/rO8lDHSx1/lbRGxYvNjF1MxldQCFtg
lvEc90NVhWJyy2+M9vaM+YEAPdUFM+5PyABCI58hKfRWNa0tgCZmvxcdZZShQAmm
4C56IDDRDvbncx9xn7LSc3oDUU10ia51DmSsJY+5u0jfR0+rUeYxCp/iGaIGuZrM
YmTQdx6Ffne0MRtcSo1smd5WmMkXhP3Si8VGhyCslkv7xyDqYuL8cEjyitXUbpKe
h+Q6N/1psqr6+ckS663/dtfZGIXbWQLaMWdC1Cgz+eV11sXCBuHpFbIxsvLVhRVQ
sOuMd2W0fpkAc3A4XhyICZ/+kFJLHu1gWtCXoUsuxr57wE8dMbdKZQ11s1o7N6zS
MRdPame8Rp/Uh9yq0EZkoO1fJNqFMG8H+I489VLRKDuSgrYKxCZynYBOLJm1Uu5t
Q/B3GWaytH40hMwIL721ABiJvmKocIcSDTM3BTnRw9P9DSqoHlM0fbLFcU5taWxm
5Qkrbk14w2jaI8u3gPu1amTC6mUK+xnmskGkizZRLRrGroZfhn4j+ODkoD98Gn5j
YPhG4Y+/y/pxvHcmAs0q2/gyee+9r49GSvbt7R74KegMQsUM4DXjAmPgD550J5Ra
vySWr4M5PUqR27YHk8Sb0vclQkwmE8+OHhPkRLBdjZ9aL2OYKVDRZmE2Dt3bhmt6
bzMvowlmsOOe+Nd+/5qrST1BJkry2IjFhBNG0lQj0D+5hnqb6laDxFZ+1H8oOLZR
5E30dNWjzFB+ZYbf1aSoNqWjpP+feWh/sCeojquxHf4SJWMiS2N1bFDTwu5Yvb+3
q0AJHpK5kpaFQ12S3bCsrNijoUat16km+1BA+n/0KjBsjenYG6tnwrEx2TY4YgmS
P0o5cvwEkKqgRxe302tBB6ysWlL2pJxJXf8wALLbktC6FWa3homyPiTgv04rK3Ev
4VkpnYUkgRpZplNItaTNZjZV3zp/C4pVbDt7FseZMO9E5pE6MIS5CHhxwaQFoVQz
+Jd5yS3Nx5uBJPQFO1M4A6EYAiwpG5ocjomQRRILlPpV0K/44r64OMUhi675XrvA
9eLKTpUaykfqCDnFGKi67KTtweLmJbWXKuIMvRGlIRaT6B4k36zxIdSkLZ0NfvwB
Om1jw9vjKHaLAuSh3pdmPC9MXw/TmdghjLQE+X4sh7FicowuAxW27hS6KcW7l17z
w501gTteYOE+juceXga3gdVOct2Xc8VT8g6g1qFi37KM7UtEoQ4zye+R+xTWBk6i
7Y3Vlqhpf74XCrvzHKyYowoboReic2vaURvnboiIHfHcfOP81tBU5ng7LdJOQ2Na
0r4jHTktdEVMzUvSWNGqRNPdUfo0s3jnppTm95euu9Y38+C+FofHg+OJcYOhnxcb
DpGdQIMoKBkaME8QksCM5WeNOnsWat1dyNzHFyEs+NGtT+f4vpTsH9nTP8uVi/MF
sbbRXkcVfkaGrhiv3+B5jqscYMSGoRjYG/jQzfS6K/euMopoZpERohIBCDEaLKmf
2D4jA4NbwfD5wkzuAN4IJFIEveoLAHNuWBRkv1cxr0BfvET6YAM0WB4JMSq0pwek
aRQu7CCxn5e3U2FLcGrJdgk+suH7RB9JGk0fjLYjjXaLq0uDifdsdjDMwEzKVTgc
azWkXXM0a3feiBDtow7rFQoK6exXZurGIEvIqIiw7ffT8y2bA9+fjhYJa3kjDFdd
6rD0G3y9F7Yog3jL/6CdljjUQTLoxyFc/lVqKtaB3er9fJlJ1DRTvoERYv18uYzX
oLRgMVU3n+//0eKZp+pJmIWC0iHLH96WRjbL+7iIc7XUV7hAwT5zeXk3QUkquKsp
BZTEm21SZ/yJqS+fXnUzXr8jRxYSk0MCQzjUlYdmS36c3UVAImhO7cwScE0DQGm1
E+qU1OyGQ01ar2Oai+RB6EDUKGknxfscmRBzoliVCNj08ebi1yLCX2G8G2Ez6Dsi
1SGoSvKZGBmnmVSXhYxxWbcMjs+y4FgNa+LeH+X0Fsp0Mwa8ITR/qYw3x0mwMrJj
MMAF08VVSjIiedI3odjyc7vQNGXHoZFVVpf6gyog6fOuXcVG3YxKlmnJ12taamCm
7wPFcQHfQunHSuomBGJSEN5XUYa8+Vp+ydMhymAI6cF/XMA+qqWKYF/5hO5v2cQO
qm9sg7W1Sap7vyMuU582YGlINQxzA1OQf6RSf/SoZ628gviRHckFtf+hfCyZHukG
9nuCxV33rC/0Z+zXif0TUWMG2MXsrrlgKeMTnNWbW+xjcToG2nuqhC+m3eQaX5cv
LDhM/bmOLyWSPrVr0MVOlyc7VRloM3GbpBkMBiovCHrHo6RdYMIpoAXktQOnITYV
tEC2/OwSIvrColUR0zjGODM29VVskv9KkEeRczS99uYJyJWNqY+RMy9c8sKpAwC3
Kr29niNJllAw9sK5hYMO7L7XZcIdAY4YA+woenmgTn3qQMcq2fUsSvGn1UpkSuhi
rvVBphnl5CDP26kk/j79pPLTwmx1DNXqCSldP92ZM1vkSv03W6Gdz5n7i/TFiCH8
X4cAVMr9wW+RJolraCyozKSXU/vPfjgFt9r1GmkZh2wcPeTy817AJUfYhQt16Gb9
/nwOKHCNMCHk/UsW8zOeHnBFdXCr89R1yDhqIbmcXV2gIr0+1G0HRMEZUnmrXTA2
hkWcN/uh7uwq/3oOCPax7Za4hmHJM5mL+YuwVQsRF313GFJ5lvQpJOjjQx2Pj8Lr
2LytQ+Dp2EIexWIu1Ysg9Ui4KTlgS3IYBzUBlOIZe1QSLbaAA8JER1CQuEk4MN9x
87EmOlgpvEhBwVgJsVpvR5wngOIUYh4kf0xjlzGc64crqJOn2hiLmBSwl+okiUy1
YAqdACbxhDqMo2CqIb4phvRKMgSt71AyCF25fFRMILvieiR/A68r76Ukb1wE7p6/
52lMeJbiNuwaP6t51EscOoHt/A2x+mPmOzQx12Pz4iphnnOBv9g+ijKsCh2hra8d
WDn93B0Rjf/EGpy3kt8/q84pe+eW/gRY8S5NKNtn2/OZCU/R863Gb1rtXPs7UkyG
7s5Lb4ATkfejSbCaJOAWqf+L5fkfqEKLNxEo1KkWv5S9WFrty/uivzTHh2mErK9L
nxj0Bj1wZXvNB2WlO212sTvQ+M7UhmlHiW9i5S9pZCWhZlRPWCjpyxSa1AtvBiVM
1BlB1tEZy6wk+BUfCD4QBXeACcz4UpIZ3gEgMe7wbfVaieFjwL00vkJP5l0mh2Om
HReFwlTSzd/wBMREymxrgckkxb+GTDZj66C14xlxXxEzs2l5Otc9l5b7H7arZcBS
YAoaVkOfa2meqvnh1mm5TOpIKtHIT0C5cXg0fHr3U2ltdcKQhBHbdHIENrEpbF9D
dlpJFLQqagw9RWNwh34h6PJDSrfOYpoV2wCi3gIAeOgeqgfbdeCuL4Sbo6Pk+nSe
44ptmQlO78lIBDLtqQKxO5yNwzUFZJLtxB9zpa0pFnUb+d0mglw06b7ZWkEYhcRS
xDuAQHKEi1aEXXa/XyWUT8FwVAH8Amj3EA4kCWxp//24rOJC1DKCGEjsqPGmgvB3
lMReAN/Qk5A1okv1cXi9i9kr5x+oM4kRgc/QWY50uQVJtlPo3Mzy+5j1045ovqSB
dWUuBh9d0ku58s3oeZ5SmsXOWJcZdviVx1Yw+f385SupIAq5y96WoC7JkAxszF+G
KOLOwz+y4wu0tfkDt2tAUL18S88lR4+XvWD4SXKfgjaEN6jhWqa9nC305nt/tqYg
taT1fF4EVmB8AWwfoLefTxhQ85yWuLTEJKHew50ChvOVkamMc/dxHGLvfnbaGo8j
GbEbIcIuwxznwwoZqIXbjkcljvFRGF4VoYGI1T+wEnf7vVCF0KBAa1TC3h8+pV4k
xvMZHIysHvvX/pMGHl11nbg8YlRUAv25lz/eFviJWQCn7aM0XDHwlqiM0crkDjO9
wSOsjYWvkA9AkTo1QoBKg+KW8N7v/Deh34hLQ4dlXs3oP7AboKdtmOWOEDZ8eZtX
btqAhdKILvix6KjU9QhGe52LBY2B+nyMaVLYi4lZr/7W5iEX33iwg/A+nKmO9cFx
na9n1CcW80AGqExpx9BUIjQUxl5NMbyQ7TelURcjzk51MWTb5/HC86eWo4gm+eAi
sgvIuqMumBoR8mBK98xziEH1N/5f0zr8awiRtKDzc4eATL36/GadiOWQYrV8N6M4
XljAAOKJiyOD5mUVbzNKm1SWcQfZcDxlyEmbHFjyjlADVE/+DaFuL7CS1GAnOplR
5Hiov8v6SucUddE3dZOVgaQ1V8P29K+hn3pk796PpMDe9WLFouXu5oT45PTPp+im
+LBY5s9vzE5DD77453qz+KTfrw+kmB2qRzadlidMi/R0Qcm2jMVurCSg8hTemJqJ
oxGHo2Z4vX98b7wjgMrkCWKlCRUNNOLw++EzYXUPOeMtVSiYO4cCVjDGLP3Hu5a6
IFD4NSr4+C7B3SXGlAnC4hCx9L3+RUMzU86/7dQ5FszNB61y9f+1HQGiKSvsTest
cmIM/FQ6crFJcipYbEh4Ha6HQNDfwdD2ggfETXgXDQ6qNfRgbp/AOfu0/CJRJS+C
IdyPLbJbmTnXXkMDQzj37ctc1WPdzKKegLKQhJtLp232TTEvdWQoMCEmgkOHRs0R
32hL+gdye0WB2ZA9z9EDaYw0xd4lABHpGPK5GkUMBs1VaNMxPz3ZVBl2yWU70vPu
/3C5ItytKg3NhMOwcAqJaqOReqJFJ9PqlqYD7sgYFm3SIw0eZNUeBvasiu5WsLNC
1RWPhAc0l31jmW3tC2nvyieYqX+jI4RQezx+7GuCPGRFR+NF4ZiDiL7++7XQUr0Q
B5iSgchw16q22YIYtXPlAtw8oEO3GhzRjmxkALLzcm6Nql2TrQu+Y8NQ/m1mtsPX
7qSFGmSR8eTQJzlGos+he3mqrhYxKoNzQeQgFAdIkLwSHqcQBCeERr5/WgNa/5ZI
elMpTvPyF//tTDQqOayonn/R31zZ0Ap4CIqY2COu6SHIs3sIS1avOiq8QJo8+rJi
1keMZZNO+PZDLjwkiXTYvgr+PFyYf1R79DjPS19LSY0hV77p1GODHGtp9smE9IUq
hOZXceilrrFdTZKGrf1LowYVpRMwdkafG5zj2i9YA2QvXapu5ZLBRgKB4vYl9/q7
uSEWdXUBI16Tgkkg5OrU2VYDTKFxFw94JjA7zWCLl3tMpVJNFPnfUiQkXDBpXczK
Z69ACk6hK1OmgmKdrTDTUzdKhrrvbgJpBkVMBApjeHQcF8aKoXq3/HUWSjVTJkLx
ZpNJs8kOjxfF/Wdx4iXRyo585vjqmnMemlscWOREp5isF7UzIiGbHCxxeZB/unOB
FgfD3SFoxbWEhRNpj8epHapU6ZSkaJz2lucDftNqH8Bv/a1rw7EN3VTBAbHR9k7W
7pmtmHqE3HkUQY1x0kdXBOp8k+ywJ9uyyRKi42RHR7jDCwHRsa3OLuXjlNjvJTx1
OJ8b8nl2H85gQtrvqGNb62q1aH6OpnqGk3hXpuZ67Zcoyg8AEWu6xRFuBy7bSoR7
z2SP/AqwI1Ggoadat6x70m5TxtbjvWINP7xodZDR7xiOwYylP140X+Wf+o+4pAWV
sE50R/QtBRRYjRDFB1cgVFwi2USzD6DW8IaHGFUFVsELounpjbwAPtL19FhWnmwn
n+2bPeRhW/1BphkxFL4WK/ZYB0uLdxWxlZ5YRx7O1xTtdbU6F0JuRnXGn77Saloy
86O8b1zUVpYOVISDm5AOJ3f1uqecMERtvbS9831ISJKbaQ0QZK+ycgY0+RKJbX7p
wlVozR59L2UfocHVCSlelw1YWO8t4GJ/cRGyv0MAmkkBn7IUROWaaGoNdzxIU2Me
QoW4kP54ScAgqTlUshQ7VbUZ3X/9ZFy+fUfe3KA7PnhBbr8KqtI/UCXGUa6mVR8j
exrEaB7IUjik1vFllyLUTD/3sgnauTji4CbWX6ohVEr9IQ5lLAaY+rfaV56Ha4D+
xEKJoPVpZftJoeowVY1Gsg/H8ikqwsReTzWskJtgYEqwlozrJ8qLHZoyE3tFHYwh
yei2WpC5fbelzhq7sVDKyKM3ddrgc0KH2XjpgLgZ/GWZzl2hj+j6SqXZ3R7wR2lT
28zZ8MEDQb5NlcLIoauFMzbTrYDrnqc059/9urbWkg6XLLlWHBeVaNqeEyDCOzSR
yxeq6proEL+RWj72J7CRKxi/L7UVPfJ7wAOB0RgWEH3r1K9W1qtqTtrL+K62E7dW
agqLoiINZ4SV/L0iHr+k841l2E7snyB2n2+3ptfaKDQcpcCar4ze0eFn2sR4r3vG
X6khflraGlvl35dyDZoeHisAdG/KD9qNehl2uoAAqfzhAjsff4dapxCzq8ZVP9rZ
WhU+NaBQBo6akF6Qg8FwO/3dJLIeBeuMQusGyUDu7eazRNa82B1bolsfd/x4ybcE
0KOW2KLKbBOePpoF0G+6AIFO4cxPPj24Pto1EZK1tiRRNaqhw5Y5M/L5zUsdCusR
bAijlYsXD0leR4jkdkNkovy1ThuXl8IY6Zcy8GcV+36T2dwu/YXz0ad/tG2qy7Sa
Mfh/KjBIrKLVPuDFfIO7IbilB330UXzXYaUHQXNkVV/B8KdTd+AdYtDup9u7U0K4
u7wpLx+xVVYv5pkaG7K52ktRlLHWsSQF6m0fEpjw2tmZN9c13LHkIQVcTDSsoJ4k
ffDeYtWEfKM96qN0WL0Aq4qMSVx04hafpzV9eeHTLOQYIdxAJUj259jdmtHgFB3y
+ZZL7m2A2W+FTlG+I5rN3+7Ie9GzwOXvop/rKSwyMeTJ3AK7xE2pU87Orfgshy21
XH1QVFU9I3neNYITfvWUQwPzoQxuMMchXVfojlqzHO/ENAxe+PLfqDb6hfFi7RIP
VzCoVlTJHVLJluIWJ9LvjysQoYciSef5lSJ2N55wDqNEkeZhvb1OsIKh4J7FdWCh
nKqn1x1cvtEp5P22qRcRROIq37VtFduWp1aXOVPYvBxMWM0YNRKxIOCPwh1D99Il
2S8YTwF+/pzL49Hu7abZ6pbbyxE8FToxLY5+ECJTjd+O4uZAMbeswp/imWAqk8dx
NBpnIPILveDYT7GXhEg1pB29CVRHY/crsUZ6tJLpDWzQvVqa4kIrwMwdMD57WvMA
bvif8iKPbfdtb8OHG4GqugI2bo7hkQX9KhrtP2ZT4wRYF2nNmAsnUOQuyryoQfqx
uw/PyRP39IFiibCVExD3BQRAw1TZiJYT9lRBrHNv3ySn8/S88rZuJXnC7/2p9MRn
jLJVJddJAOrKb3Lh2dIxyRt2Hn56aS3LtXYyYdmFKvXl8UH8X3lzoULM2YjYkuoQ
3Bz8ufSfaF6KKQwfu0GMiM4VYcxNXS6rxLPQNruiddQGUoMbZkxmE6o/U2wHwNlj
nNDM+RHpa34ek+9UwEdy2/8ETBtByWKn/kRa1uP/Ae335IqDozyI7MYj9TAR2GrC
on9HAcFyG/Wvy34ijMg7eEhFb3583bejb4WP9Wm/yc6KXjjMRM0i99xdUQ3N2+Eu
0/RTbcAjc5ZezP1kpkv/6WOLjrmxjLy/ktb0/voOorSywBd7WF1JuKZ6GlCu38M7
tivmK9ruDv/vsuJm3+9oy8nX9LQMa7sBZk2jrOlKIX9h7q02ir6RCNFbM4x9ZZsr
3vcQqhHVP2IfuGHxBtxf2RyhIuc2fnsYc/REBiHHFj6yFWTRgRGp08aQbsGK5Psz
2QBuIwKJk7ek37icj9oLUbAh+soZHhtpBEowf7LBAOBpymnhml8zuguMhIQPRyM/
6r48PH+YgFf/Doq5fCV3xvwUNoTMHwBLlyzwTUOra9Jg+tU20Qjcecxe2kivGATb
JRnie1uJh7CABKvzoapF6PVuDAXkVjL6Q+DaW94vkIIJJqjvCfWdz/8jYi8FjZGG
oGnLENad00A4u59TRuUZxE+sIh9ltj5fV5cQ4XoEM73GlFUwhCLllTJoHe0BtlN1
oYkgzMhXxLp+B4EbgBN+iN1NPTBlSAdgI3h9y+OsihnfTOWVikdhAdFdT25n4m8+
f+gU1j+t1gWzBzEy+D2QXf2di0HM+6yWnJRyTFa2N7gTZMQzFmIDu47t+RTyjAgz
EiegOLkKPtnhjligw5/OtzV62l+u1LQ6c/T2jZVp2DMTt1XxZOj4/SOLrWXkpdNa
PcL5IBpQs1Sob+f20y6nHgW9ZPZ3+ZdBgkEowM5UzuXqD6SSmSYQh2s6qa674/ai
8/8XLZ6n1bXeSgk402VdTYnzOO6QBirk+MypcS4wOfPcF8HLok+yBKigQioQGt3q
mv2fr1pxougITa99yv9Eze/VOQ1zTrNecF8kXKoh5F/r5VFB+H7QuIULXHsLi2Pt
Sly5CR86TormWh2L9ubvgILppgL5w6rmdofS154E0WrTZ0rN5wBd76bSMYXYffrA
dolLbFEnHQwoK9H+j0Q7VAZ+Y2JN1BQHQQ0Cvvc+zsQ+ycVg/07aGwLUc874hV08
mQWA5mv6Hx3EPUXZwP3P9tqt8wNtAW9j4IfJy0bOObS/SsFiVpNtEEJX1xWbAn40
EHKytAv4gwdU4TBiV1nwWc/ynL0YziAIs/tX/+8TqZSJH/79oe8gsaXzqF31ugTk
70tHpYm5Jk/mDHMIygjLNY+5hPzFUJRNkROn/0xGfJUzBmnZXbS6JgE4OGO5pPGP
K42pK4DG0JYzq8yi+OggkwSQJP42+XwiRiBzvGoQNFdjPq4JbKTgwqRTdm13BVsH
NsODbEN6NBCJaUO1bziersOlJ4Y1ycfKo08vHGU26R2bNIgxvWESU/c7ZI7zhHvW
kqtqj1kNF9WqCYSsfpqEkYX3XCwO+Lpgg1e+OVYbHJSx8Ej0zKRRHvMN9OzhK8Yc
PoB9JvApEsFDPpFQsveV7WZO/n+5B3TiDmaUjpvHju1S05A+D2jVfumZed6S8AdF
sfSDtl/9DaIUYcD9JvwvzY09843aQ0l8QV4aEFCMPXlelEdWu1CSX9DHzxq6fqen
TdIfiESigVs1qX1znRwK2xaFYoBBGhtfoP7MzCnIjj2BJFxPkVkK8SNRlyoTRDUm
zG5xxaiSMWoyihxtknlhQusYGjSBvXYBYowbIYU3A8bykhsOKul3MoC3zpfiIljn
sFCPL+ljHj/XkhMRvkFA+UFTls2Br7IfWoJeU3C22X0dGhO26PF9c/8gp6alwIC+
gCW6LCIutUEvuy3y5yJuMydwCyDrGE5KkhTxN187/YYvo19FqWXrh7ft49QEqYtc
TAzlJ3USZx/HR2Arzjm9/SXEE4wSdaIzk2z4DmRyDLHo/+cQRLxu+ekbRUHeI0W6
Q8sCAPUH4ZXk3bPFoOwhj+e2fX+Yj+m5D2q8O+HtnJIZ98yyZ284J4WdEBpAAYjz
064y3AZL1Ocd4CkBg/D+R+KZ/LHvsLAW2BGd1rttUfbglEeZYRzV1L0orMO/F3rm
DPvU2St1EoVNPZB2e1J+U11bd18plinRx7/4K6FGDKFL0oXhc8TezwaQuphfHX/m
AgISBAPM6oygpPl3WRK4c7xBH7y0jOstXYcERv2gm2DVD71x9Aijp2SgFR/bmkQ/
UVWFFNf1wI0P2okSkYS0HCNZub7WCNEc7nvS+MiYmV6p+CUMwfZePjjbMMVv2s6a
eiHW22EkzOCL8mW0BwX6+U+aCtWR3H4moGupDVc6VRnxfABvxeXHqQuFyi85lE2F
2BDgyMyhzdKl6raUBNVfLGfuYM44zn9g52woiC+b+VAkqjxedRwyHHmWxmj+ZWOz
hAEWZPLJWvQQ7vSGPQfJmLGXAm0dpI3YOBw1dYj24l8uiU8Bxr7i677dR1pDobqk
WHRTpFVMdhM3clB8ObIuVr4b+0RxL1XsRUWnw1Zy5PNZfq7+GtdjSiEvh3S662ib
2mP+OHqKUsEXn6EAPKTSlVo6cuK/M70bGU07She8hTvukesfNE9S78FGePrfV796
eOvBOIhk9OGPFrG/kiUrUt6HjsxHAQEYSrunGvB39gzpejuxvamXrLTDgieZ3azX
0ePkkIXOrPA2YcaqMYZs2By8W8IrRI/Crn2PUJ03IX6fy1Gi2tyaGaMPNuUW4Vbq
Xev9J07P5NRo0+ZjADRZQoISlvxdvPFS1SenjDDORp5+v06InAicfY/CEcHK2JJt
61LlJBOw2ZWwsmb83K+doKZ6akHIkjtDV/Eh91XoItuWHApxklrmb6X6Q8fKGS9q
XTIVNKGA/TOErSRU5h7plnKX4wa0qmAZWYHlCd42a55A2HoVpLWf21zaIKSN3sM1
t8KPyI86DFyVr5TFKGT685qwQfKYxF5jkEf21ut5aikbk9J5QWOEmyKU/Qjy883M
PO5eQHgbGmk+JLLd2mh5eP3g6TubN6LGqsSmx4o7wxOOu05tCYhQyWazSeWQKbh3
KNj3AOC2fZ2WFpd8F8ddbg7yujHD6Dk+hfaSJeSfKgnHuojw6zClwQlwjHmUc/B6
xwPe+fm8SOJ7gmozsVIjTYqb3vqcO7SD9pjV6li0jQLaghFDZvh/dj4IBZd48boT
7kSypHEwsvwnAwvX33v2O4oH/ADsGTsGcycDufMDUjg3PCEzKvNfVJ4rK8jL39YF
23coOnsd+KMzizVtNhfRQ5dr2sRWqEN8XjuzJRVSxGkMLJ2JFPAO3QlP1sSV/JVV
XvbGl5jDVlMOfzYOJiX5Wvg6v/Q+f0EghedjexpLVSzXRvGwgbyB1hvqgrFVB5p3
xoaarCkwP0F6zxKMPXU9hfflGOMGPaFwJm8EcNe8TN21buwdL2kl7EPtCVqJOc5X
PP4a3t09vFlV1H2GDFwTQJ5pMnAVE1tFpiORDUSPBhC94NtbCHI1FxIJoC3Gcd5E
Ye3JyS9EnwMDC6LpCi/wNabEcK33Qcs2b7iRGFq8xKLdCTdTIDxduZAoEC6KpOPm
xtddbFZmP8PtQ5QbQjNaPhdc/TkkoObzbdrfXI/UpmJA3EtSeZWCGs1yKKOHj6H0
/DUtEh3D7mYQCX5mKybm0XRRUzbNVi1ext99y41MFWj6H5OIsph3paDlxQ7h16fm
udLIr5qR4WNEq+ugsuSpJDVjmRieuhIWnTsxtWOCorZKnffjhvlCbrnj3DAgbZdO
hdKbRdyby/WMLsfB6kRyxCGPvqLmWSM+vkZ/FaXuHiXg2ThuroEHzK96kD3lUgc3
AAC8dm8R9wkntWDnx6Pm8QoQEPmZPWzWO6sZtycMSuXRVSyTpBEOeU4WDiM/vG0s
uesBChQY1kRD3i29lY2Lgx1UBEHAwW4VxwK92nvL+cz3WRF4EnBMCzoKKrhOJIbY
zUyrWbmZJjS/SwBJu2P2+gBrY7DkERxKMWsDvbC26s3kSYII47dDS1B6aQQ0frct
yUMgVF3SAKPbDPXBkccc0gSPYstM3YyybdB5u6YC63hAhon+bX1S5Z7dZyLIn94x
WdvX3HOFjQ0zV2BVUbGnooCD2FEuhKgBaeyG6EG5yD2kf25k0SazWleUx/PF/Q/c
hfwWJTVAYKIcXXRAMLmZ3ZvqhwLRAlYNSvUn65XEfCjh1T0aB7yOBtvmUUcyqH5i
6NrpjWHNE0b79ZVzf+wsJi59oKS4O3WZtG/PPy7r7JdTUWkrjXmh9PZlKYVgMjiI
9jXEJoAMdSwdMjFLlgmkGkdPHzAXu1/DkE+MNFHqag+izt8OWp20UrFLQemGnCCn
s7KULZU9XHB6V4WiUC7aZyj1tPY7cd9tXar/2iJduqdfiRVFeY0dmW1p9LP3vd/z
8H1LZo4P6Paf/JFFRKbQAqGWvhqxbzkxhIdYjcnZggaaNXBgqRFbBPn6RKWEBIJw
DNLHc5ww+eMiqGFYvBbMBizDxAfPQnJiX8uukTmm79qHOhXQrzqGAJ6DUL8rTtnv
vPAVPyZmVCazFD9j08dxDfgWI279Jw5rjNtqHxj2FXaqAW0DckEODT6QBTS++vzk
vhYtxDaeMb6BuSk+0qxyVDU72aBtPHKaDoxOp1yZnOEczJWOEFmG4VV3x9BOiSHF
lzW0vElop+kkY3SMIlTyjrwKDVdpXbSuvwnF2KHy2DO8g2SbYk3HgXlaGaH91aqG
jmRMD7459tBaQ+oZ1dOzJvgHwM/spDvLLUlBEiysUaS7Jb13IIk8jFEfU7CcBj2Z
/JIUnlXDNzUBgebBtEUssNh7vknALqYhmAxmFWj4lGjpVY4w4+Qrv99E2KXb2vuH
T2E6afd1YfKOT5so8pVBlvlMX4Wj4dYCBEPAiij3G54a3xjHVkfyk2f2eV19vMU4
SNLyBYALQRqq9aXQ/0o2rn1cqNuEmgfsd4+TlnxbygUcoAShMq0gIiVaDPD3mU2o
9+RnbFvpVLMoCByX1g5uXGu/QlkjIKWTahS3J8dcmXpd7Xi8o+7da3DitCbiIDBS
18rYGn5Z2p2kzH0gh0DstRLo0WXCDTp83IQO4TUt7C0UJcCMj+aPOEy2Eav/gG0r
JF9RTRtzXRIOpNxSoAYO74zPbVGQz/Gx+z33TmNmqTw80TuUH96M79Ahg2FSkM+2
OBiwz/MqEzqNHMQYsmhJHVh6MiYzx86gR5IQRh+EgB83yxPsr71RDKYAXiJK0dCw
+O7jloPUSUQSokO9eeSfoDJMPpeShQpt2IiWKyB59cqVoFiXddgtC4ZPF9sq8yzy
dab9E1RT4JUw406wt48sIpRuxRTAgOAJJ8MqRmJOxNjo/CuIyLAN4rIP8KX4pm/B
8Ovo22SWbHauGDeSBf+5dJtFCQ2024ZKjnffl+nSQrk5B6CmQvrF8itYPOmVd9+u
PXEX+3xrwF9jDppsC6/cKa/V9/YFVcKGMN1SK1iAJJZF6/DZNckJoftgcZvZJtds
izFs3LaHliJCoLrDXrJZ8TZnIHFK8a0T8nzTwt82TkYuzOD88WcqHt9rOuSsf6Lk
r/5qve3q8nRvWF4VM0LB3hOvYGtf61v+FCTzh8PuGR97j7pDWXJTOqLX8MG/ERml
yAWgj0CQeMQPvIPZ3qbbCBPHMHKmHVizBmrBrAXQVYTDUBTjAyAKOC5qbKE1Dade
70HwElU6LNlyhHZ4Jhu1pJ1LMN+PwJcjplV8DZpQXqlGZmF2JN1NnHXR2prAD391
ndR1YPShudtO80p0vD7/rnFoXYT0wACqhjIUo4xG/7ufDgBSubtiTiZ1dI4uGhbz
Svi6XnxJ3RVRT+uHigotXH22SYK51TD4S7BTOCeaZ7r+O7Fbr0izPKFVDS8raYP7
IF6vdpJKZsQguPxlDvwk9XClhyv2vRu8IgEDnDdpxt+Q6H7q7KA98JZKkFz1iydg
M6iseV0cKU3Ctwcm/uwm6bBzm6k1Tvx4J23UYwmIfSbZi8u5ub5tv4jSWdOCJhIc
WTfzfVxLg3CP0rfDUwIqHLqFJwTnmGKFbmCg+Sp90qsdgu0jYi8Suy74ZYYayRie
KXrZFio//iFou7fPzErHIP0MdxE0fc5bqBe2q1AqO3wr36KRLgUOeGR+WJ/07Sin
d0oTjmrNM4cC0pUQykw9yj9i11AeNyWaPdc33iC+AHMK1xvd5MbfM1cecSO6scUp
GPM/y5exqJqAWftTA1rWxUe03J2UDLd1ciTjYXL7+ElunqNUaZhYVsEJlhUXYMzy
I0AjM+iV0rnMPAKRC/BhjOoUrftZb+TualSn8CXZXVjYxBtagvkcFELJYqjXUaXX
sQxdW0asq990iHAUNQWVx2fK80ChJL4HYE6+ePLx2uba7WV/E1zw9gSAyUyLF2+I
cxa9DRP+Aa8ga+IREIzQTSr8lP8q/yYku2HuRdXMCCj+xlJEAXa3ZQblVZgPAwnv
HYhNw8nlbDTmiuflwYAxyX68i+wyCUEaa6l9R0Vk4Sqx9ANHe/WWJLi4Tue+Y66U
rER7J10ZylGbAdSxvMVDwExui0fjOlJFONcB4etmrx44gvW7LCoL6uhNnPk77W3C
LmiYWfcYIYKKT0m89r1e43riXXywqeXwJHMmup7OfBS0QyjYxv7gS7m0i1DemnK4
9V8SbEhQurgBfpeaHV4fxdKWv2a7aMVrI+8MuQi1iOXWV0kzhdUopjYITVFsWwJO
LFNY9scrLUbekoFWzCdyw9fZHL5BO4ef8018ArrV+9EBFPNy9bUCj/SyHKjfpG5p
wNsv/23L/uWIptQLpLTF11uqgBBZNR3kxYbdxiZGXem0Rh42Z3vFmYRpdf2qR+rR
yLpXEBlLeSXEluBk8dAv25/HpsOeV40a7sMIoZ0kei1aKeHW+0bMIzci3KS9g+74
8LQ6ftUHsJFI9SCpEA9gjNUovTKGIIRu7NCcx6J4DapaBJtScsgHV1Sh+8rvcpsO
NMJpQjWviTK/z9sczm/aIYm7rs1hTo6IDzURaJDKMS/yU/FBj3Dhy9L+6x6n3Ugr
T0WdqweeGe92FHi7Ylm2dKK8lPdN04YDwOgSCgiAoo0EsOGqAPFCfGCSUP5C6UXf
BXLm13eUb86SI++juYSsTCXwIeohEDzaFL2GrfNobjwhMQ6Lz6p18A8is0sF+DG9
YAU2le7nwGDpLKC25uyzVYTAZMgCHwoDMzBhYXGBRaPvWr4SRsAHuSlONDMoOBMk
O98CFLMo9x6JaGhM2cU4zLZXFffl6K4yyonhIKAQb/J8wIGzI4X/j/CgMfrYJGBR
X7wxjyXdax7jM6WuJqB853JPevPcPPkcfuymdeLgASlNRbV9hDyg699KgMbOsY0z
NxdZgwsQ883qGNjJIBdOEo5ta3VZEdjT9THduPLtRfgitPUFD9ag3P0+A89HrIMQ
aJOFls/oLZJUPKioeWQAPnPOT+/wGm61dE2YiQrtwD9wYqI+6EfCIj5x0dFr3PWM
+KsSeNoHcg3E4lOcXMF/gQEQnqCsrrU2UUDCJ9/9NYIeJ3m4kfDYEQvA4EAz9qaV
Q0Ug3IOUUVn2moYAuMN0JyeEIklW/mVnbLEylDgPMryIzTMR53AGLfd0dZnUOQyM
EGr3EgQgscB8cuIhrN/HWffxTNr1c6mZQu9NPtR8aZ+dik+thiWRps08HUDGjbi/
Im9hcbTgBRin9yrxTtV3ZZoF2l1vB3SqpqvJbaYgGZa4KwCTunslUENtUxkLz1Nf
KVBxY6FhtY3k5jSxb/Y6zAHH0TqYis1ihimhGsKrTmXNgC08G9hnKZ0D0nDrRTXF
X63VsczrSl5t1wf9Mwv/MP0VgBHRWd1lPnTjrsA7H58MleZDoDrLAUKNX1hhokVV
5ZURX0a+tZAYGS1Yp6zh3LjgCK/2wG4OVtj2AMtB+1bpj+m0TMKdtxkhTWxHGu9h
DhfSs3P7U1JBifu2ngO0zb2TbWIwGDmmtNDUKBQXA6MfVQ/r1lpSyGW65O0cIrt9
u7Rfjp6+wf1LYgZpCMuDr2q4HMOqieY5XOa3ioEZyf4njd7NVN4J6xEZAVHl6T63
JCs1q8InR3b5Bs95aROjNwlg84FoKjkAlb8DEpwafNggCySzfLNQ0gqNTbYq7pJG
W8qgTId0sKUwrMrrW7n/SCHv6FqQTlsRFrq/LahXLxQ2Ba3Yl4Wgn9fD7Bi6oAam
aZGjL6M1OsqePL+DyVWKJsT/6HIsEX+OvsmCgIGFTVNAOt4zrcegrZg1CmWISbTY
R0/Z/3OTLDPKWFvOxGdt+Ri6JhFVaSxDnbGRnG304szG3LCZtOEkAZNsMAt36Bor
EJhGM+K5FS0Uawhc0kf7TFZ41/f+ySLUJ3QvUBFRsnCx3HMxlIpmjgnyf06jG3fx
iK1gck/6A8aCLWoVTugweQykVs1yFoTKLcROhP454DlWTWc4BVSdeRIuVsojGrXg
qULeVR5hCiHdnM1gIdrljoAjlEHLfg2aaPTFP5rpa3j0PSU7LmWhBELww9WAs0Rc
Zx9rF2TH/ZAztOuaY/Tk1SLpOD+JRGdfaQ04BBAnHL3CWgAvhLiDSRla1E6IorM+
rdDYvElqnXaamt4TJKcmm/N0K/AwFCYpQEe5tph5cQy8lshVBxPkmQX3R9n9gIv/
pBN7K0saPaUJc577SsoSCWkS/CbYl7/1yoMhP0IuhbNtxMihTkrQbkWRwtfRBV3L
AeF5NJvz+o6hscjRcqn8TfnKJNiu9lnO+AAJ5D/eoldLmv6NKaB7zG1tpbmL4XL1
bIoxCxNo9mu5YIo8OFgS3bmztmgksv/2aUdCOyzjG9t3vY68tNTH7UAgsAcmSCew
JP5zuOed5qlLyq6gXxz/d1JpWNofvZ4FSc5oeLFnEM2NjSQcJCnktxtb6b/eupBc
YKwtgivXvlv2aD1rGIAV7kLUYt9/X9IBTFZoYPzvnXWKRGpM7MVUme/zZbD7XibA
lcmaxBMlbaCXQjbII75rIx3Diey6sJpGFKLrMwNBXUa8yYMpe50jZv3mFWzYEMOP
9iVbzCtxAFhkFqTbFnECrQCoUVVX+4IbDwdjVKHTCt8gpd257zgVKrw/zvuo9egp
xSCCtdmcBSCx30RZKkZWWaD6y0DGjt/KJUGoZj9z3GexDdLcqzPl+zOOpsrxDi1Z
ak+7MgKttmLa9yzSkH3A0KBRKqZ5asNG1vvcpavyMGyKw5XoJ45PEzsPlD7OlLyx
eQ7vqt8nd3RP5cWg/DDNh811R5WTBV5Y+JFM2FML1GpKk03I537Uw/izzzByIvkz
WvGmO/KdV3ZyMpaIg/+KTmT4WeaOGw7e9iUPhr7BK5OdkA1xB9Ntp/mIeR7guIID
cr1gztEj2Bpy8pF5XboPb+dEMOCqfmEYnfuGH4qUrpWn6JGhgx+Ptd3OfC5EWpQw
n7f3xADpJXXFPfR9F2pFyBn3QooS40EUkTWnHCPca9XVuQPdVBZr1VrIvr8uJTD/
wlgvRxXZwr5JmaYwP5aVQKRdU3qtTxhjEphZQ99Bjy6vr1Xk387wsQ6ZVU947879
jj54PXgj0ZCEvbIosrO5aGVQ945HwrEoJrygcHcOjWl5e96rKu7jRH06E+HP1yw4
rWqmBNWWgvGxeWnWcrcgxo5pB+7eFdlWvDaAI/9BEXUac4VnsPyFlCH4j3KToCh9
dRqZtoEaDcy8ICa5NkFljU6AoFoK6kw7sDG4nP/Yi8d448lBcKGqOl47wxe8JH8V
wYcDDKF5GXC3YihgHUzNW5sh9j/7iJAGFsnMsiVl+qwpSaK1gHc/QKcY7KzbG9lx
`protect end_protected