`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
ddtXksX2+yylW5zu6QL2Lhnb2d1sD00763mmSITNX595NcHTEkwn0zB1Dry37fOW
FufOhVzEJp80NC5qZ/+F0Vk7Ik02dIR0elf3clrjeJRK85K4e3Hoo4xn7YbFUIms
l/8VZSb14+JVGURjfswrIyCUotIzlzVYZ6gzoZwDXIi5gQIBf/gI+KxNXPaKV+PQ
Ufys/12rjO6aI/pPlqSm0hCvftmBcnezN2hk1UeXgOIuKZnogjOsf0iJVX2aOOWE
6pD/psybjbnsNB6kH5uFTA5frkzIzkzl5d9+YDm9OyC+k84E83I/7/j+rk4L2dah
QJOvksSIzN867/4Qt8qYTQ==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="MvBXkzurAa5VTw+1JJ70nePUfoQXBvZOku/SMmg4TwQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
oRtzZL4VJ4iwysPsC8SXYCzXS8Fw2gtZTOskLcDV+1B9Nzn1zTyNtlo6lNICRmmK
ZRVu2BmCc2G+fmzynYlNTnSa7C0Cuel6FYpxCBlOuk3OF2tzAmLAuDyOH3Z1Yjzk
a0aHuoCdIRKv7BrZCdALt03JeUmXKPdOmIlkVGFl8yw=
`protect rights_digest_method = "sha256"
`protect end_toolblock="Jn9CQpRhJt4rnzZPRk+dOpzAubz7omckX1MrFd4p81o="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 22480 )
`protect data_block
gD6l00tciPUa6pDNTk/+t0OO0nC/UTtBwLB41d4inuAUA3i/ALrNyoJVcBnAmEQW
ptbcNp5fxEUJjnOxnedyZEuEBxWRieZFQnkRdF269oN/2w+CRwzqFLNdFc9MQHi+
3ZxPofDDcpDU/lmxR6DMJFFWCNue7nu7iTDTHjZ598ZOVjAhBhSRS8EFstJppcaC
q+k5+9LHfCm8AJUwc6iASH4OBJzlQN00Bszpxz3t4nD2jxz5H5gcDlL58LFB9hxv
Z2jdaC/iXuPUar43xq+eH+POAPRHzT5sCiZyNuARzq7NpvxkRWJRQziTPdISfKO/
ZYysNMyc5OUQ8uCeejS12R1HtMu85eWFcCS5Gg0rox44DTzRyJ3WEi9TP0KyWjrU
buB03Y+q8j1JuV+1vxafmpBtxwPitE51D9D1RR7c4PiCYwL9glZ1j/PcQ5sst+yM
Y6mF/4j2dAr879O9pWpcXrAX+JxtWY27W+skqowDMUvW86ClCTromELBHixu72Jj
pG6E0UVCK26Wmofxl2g1rRYIh7r/rK3HvbhKvYpqXeHFd4VUig+ZzEfYpChjG9sG
Zh/GYOhxC+xln3+mEY0NSHV+4bd1hKb8dYHDVNdH/CP0vfdkXWr/fuxpO4CG2osp
kIKIYnjkmOmH2aEWd8KgR+9c+aJ/8TFYHgeB/QT1oSIe7Tv+STEuEshTpZXyUnF0
LyU0fdW8DlKOQw9AT/hINdIbw7OT92TMEkEsJWQ6tGsp1Q9t772pvrhHb0m/KSjq
yIDoAN54qtmILkovhKKYAjm0NO/yx8H3t+nRT0IQU0ntQgTuEA8cDApxBkAD+ICH
vlL1zJH6RBFGjO2XTRJeLJs/mXGLxVEwv+Wg1lFXSDrxgNv6Xg1ffPt2dN32mBbf
EukHDs16Q89G68cHQWlGCWl5DjUpUChdWTfmhTjgA7yn65wWqPfUNIueQpZ30xsY
auQZy06ekJ1DFTW77wMj749Yuxz9ak62GGSuEfRu3AN7ys3yk6fnFsZwN5fjp5Yn
ww27vVCy8F6LRMH1U4KeLSIwh56s7wT/eWI7D3O3Yyl4cUxgAuyi/8bgHJ+ZmCmC
A/YQpqLShYry8qml2BJVGEo+OXWECIUFIIglCK0Q9ThDZtPIC4pbXPiXYzrbHMRf
nh+cCw9BoG3pL6EM5JqMdmLfmi+oODljf5/fkr5H3e1nfyddee7ISsF4gFDH+qYR
wU2Aae3S/7h/UVBqw03bsHayp2h0zOICQpTEp3p4Qxv8BnSk9942CfadwnbqAPES
5Gg4oug9Yl/CEAoo+AtzsD9fFtI+WmCirDmRsYf4KJOatT/bF6iI+n+qK2/anSkb
fY6DRycfPmprWJYxPoXENWA74EOfh/OZ5n+lOEpCVpYnYHMdhReHWeWt6Ryyz57l
B1I5z9NWyIH8ilg2nF5ebBgUZYpSCeTp7f3oT31Xc3ET9dF2Re2s77zTyk/0v1X2
XsHolFaUdVpJVnDJZZ4VDp+vCC7e5xu2zRSI6Fsd/jYEMiszRTARG+nyRIVG8xMF
iLbbjYOOChp/bb3KqhSao6HtrmAEwM8nwbRcFgSv9rBUZ6WuTJt4PLMNi/ey89oS
qQPbe0GNhUoBVZhu6do/ZgQkvQ9/c0aJdlJrBEkehwXWWFuSFtoA/QUH8V74cVBO
7w16KNDm6jtA4FCwijF3XFunzd4Si3Qs0P+vy7yaLdORj363jF0oSfosG/NuR/so
UhlbZr2FQ5VeT3Nt4CO85kKAF5IutiLzuYzSO6y3xeg7vZ1qgkUArs6GSZRRsr3h
EyQOAuLCknrJP2ETp1Go+iCuj1mJFqjsugot6DVVlsUHabTUVOcWs0eHNgsxVwDN
p6FrD/3OEE4TqSgH22XS3W9u33EOelN4WFvEWs8Yzuz4wd1lbNUqT5PPpB2T4f50
4MAQfCABZJFj+tVQzyb/N3egy9DoOIFzoFCyFdJb+uIUOb77nrK+A730pAqIvgT7
bJz0Yko5/HfuJZWHxdIFN/mb3iGEDcWIfrTvobUmyGRBwrI5eDZFjTxny8ECF/Jx
8HNK+v9W7R8jR9Mm9vbLe3ngLH2T4KEfZXBJI8jinnkLwBzH4/AjQLOSw8rG+/1w
RCB3s30L/u32GVfWv2q5EXrYAoxKuzfopIPFK+qiCJad4+IG9C9aDyvNsw+pKSOe
TUi+T1L7pI66wDve8bNhuq9gWXzu38+xUzVGnTzxIgM/43nLDcfO/lsKSKych0V/
SX+URoaIw0YPVqkqzVIktOgSSAhj/gl5Wh9sIpax4stC4vbSsE4yZRcMtXEeyXPu
ES6A7meIsILkJVs8bauiBaamNZRJMTv+AmH7qhiuAnlnKHjdSpDu0iDmoHMOk55p
h6tMochA8GJqkVUjfGpAOgeruf8oOKnkDBTF5rX1agZWQ8QHnKcVsHtlnhBC4TND
IKi+FW6ot2/tSUM7Mp8ZrV9G783gUbtP1XEMFDiUXiz2yYzsYR9dF3r10n1Oxgdo
TkMeSVxPzV1p6uB4ceLg8dIPdLP2HdHBx3OIsC3zws9pAsfeF/UzK8NmR1JIPPoH
vzvRKuesT0xkARcMUBhCb+K2tVLrEPQAcphnMTAPdDZmc1eNJKEgUuYN3cepKoSA
jETOalfnwX7TURSQn65vq3BE2L5ilafe1/n3QEJM7GzJt3tuCbCSv2CaMGSqhTVA
S3r/JM48BpqTJXAmHk2WxT2sJ2yvKcRni4J34xhW2DumzKi3ONO1+JPUxf+adWwa
aAwqNRuQaJEiTTQRgx1xM1Z+t0KjNEKnMkhYUTq4+vkFv06HIYr8jxVfNcCiOpQr
YUM2ogfz5vmleudkPLHx6/SqhaJfXJp/fnSJsRvVBUE1cvF84lCsWSqXBbSfr3Nq
og/MJ4sK3fThj7hkdd8guhGRR6tKL97OQKPkNCZGcrAemr9B3dinmexrNW+7JT+r
fEX2RRp1iFxbmUBMc15BVlMHtHwYC4xKThYSglZ0BewAl0L+P26ZgbfwhiEdDqpQ
ZrzCND4yc0SdwN+FK1ncd1gYLg80tjQ33XZ+rVbxZIN1LubZxaPn1n53B44WAZB7
ZGXxTmYZmThrCkvFuLK+sems994EEj4T1PUfGeDDbtHLRGc/a+UkEytZY1F+WRcJ
uCmpa2VP8JIRmIzZZFUmrVhTPcHUJmrGWQH5RdCuzgG2jif9rmUZbzO2M8cDL8e3
7iZnd1YlxcmwEKAWHBO0JxicGLIiBvdF49NaYj2v4PL5FLXGTIuyqoWSE+F2wsja
OWjBxC9jqotiidXWXthIEITNDETPVWluB2BhVdRJRpAhtnzfjK/dlyRlzRGdjf4B
I65NZNmzryxOzMU9DJ3fNjHOLu4vqATDKcoO1BGvxiE9A3Edpii1YfOugtNG/7X9
qGOGN9W8CYYlvCpL+zoMU29n9HPuTnmFOpJW3H6KaoZCmeK1llG5NGBCb+OaiIBg
UZZ4UJT2hsYr39ytdullHXn7OFQxMzRE8KNenmy+/sI5vt74796JwKMXxSvGU2Pw
LOejolsgouc/LcxVZV2VSQYbMIYOPzIQDUMol21ii2lYbeEv0ApFyIUSsTsNN7CZ
X3o1xt6DaE1sHE+qKMxvFUHe+ZhxrXyj6+EJvhP9KGO+TKQO222oPtghw+uq1JiD
LSMxFX2mW0RgUaoEu5QDPNRmy8mmoKniWC9fh/yfXaH3f1IjAuSi+GFFLPP5kZVp
o0E2EQ0QQii58fLDUI2Kn1welMcspJQODx6JsRM5uBtLOFeTg+eIoydPq7UsOW1R
Mkd4lbZaA2i0f5roEBjzb7dZDGr/tIO1fC/6xkyccm9nUyjz/+bAnKRCKtNBkztX
EywTNkC4DnFJDlLuTNDfwjbMEHhtPH54Fa5qpfN/ELlwAEQf4OOUD1r0srldEFXe
3KTDKbqDCZ+r3JbXBxtokjQ8gn7LcvC8uZlvuLuW/dbOdSfxNgEyeEehIjkGh07v
+XrojuE6r90D8h4LuWKXW3XHGW7XdZ0zF9SMLVqBS0mkdLQxEvLUlX78e6fRewaO
hNZNuK2H/8kk+kpl5xOLMs9KQ9ANW8TjKZJw9mXYyisfvRKanRXk176QLS8xNqJ/
rdKu4cXU1wk0p6SiV6HrOLdTG8z951FMiWDxjHS8svzjkrlSdIix/yszZUa6BB9t
72QeA3ZvZvYkkSF6SJuHMRuznERCmYJvnjtQzcpqYpJuadpQXDeoq3jU9N1YMJbE
sKxZsff/YS+qdPVBOEeHUeZF7UscpeBZ4lp0WKMQSU6A6bsH5qbPAoEgLfw2WAt0
i218p3uTv7hMxaQO38lnt9Qeh3u8sJu8C1A2rxd3IVHn59v8pMHVRA1f9lwTVgKz
wtrv2I8Fawg8SrBXfGbJal9CYRSy/A5Q7vJrWS5jGMnwBYiN54VsDW1asCBaZW0b
k3XDneJ/m524AB5Hw5yk/Ffk9kxdk2YH1pzxjcYH49AWmgGxc6KdIUhQEnuRhxT3
NkMP7J9HjECn06IUSEudwUtVTJOUeG9BYABc6Ac5+3j6mzx9ORwpfsVXfZpJMmSu
1/abBIfPJpusMj+qUS7iUDgdLRD+a+YDmYB1I4T8CD9z7p8H34/FyA4k2ZVP9s/g
QbO/Di8xAt3RRxpu3Ro76qwLkZb3jbCn9g7X7pIyXlz+fgldJcjgl0B22gCiKVjv
r++16pFbycVv60EAE/IIMt3ydWAnIDd/x972eY/XBXutuJyJDtjXkqjTU5oL8I9D
Z0sbF69+C9fSuROotkQ10q00QIIgTfuEznfzT3DD5s2l4ZyG6hUO+3RScO0zwukE
E3n8xnoqnVBhPmKac51z9pEhzsYsrbPKADbGHBExcNew5UI21z84brM/gGC4NNs9
5ZGXVo9Fkbw4CVZl6un12o+e2fYoLcNI4x5noEJuZJ7nSKhoVHl94sY8zzwwG77K
Tg4NOHXdtW4Xun1YtL/Qkiv3BHYd0Xu7SixoJSx20oW9Y2nw5EAhq8Nqfsp312YW
bR/2Do+tpgo9wUVQVeoBdY/MnYwkcUTgUOh/bVdK5jPyNj1aQI2+j/xs20tGd8zF
4/DuHrMI5zc4dIdcvIA8W4BbJDhVPDEu7Di3s1POlYjkhFukkg3fXG/vHV3j5rMy
t+1N4bh0YhgzPXWXGNisnjRM0bEP5ZS+1Tsu4+VKTdcjhnJ6VJxOTElhl6jO5+Es
HR5TjNRGg5KQaHEg4BMGnFBBDps00WAydZSGsbYYTWq/9c1nuwwn8EvdADKBx7EV
rGe66INqEVlYjG1gRdmY0SfDtJJ4sLLWmETPg7W9dHh5QwtiQEAefNf7uMTMLxRJ
D1pSBysnU6xxkaMwP2O85fA6H9TIGcvrX+yQcqzHknuJGVzaWX83Ob8d8J8gzsBl
Mnvp35ItKUBbVqR/YKaHWd0O6EraECgvMiYtopRlWEfUeYUeuSnlJwUqep2Y6k6x
EOrwrcxRTlvb6+Hcvl1i1zHxujzWkt2SuQuJG5ym7oR361z3hlIbCVofvq8lt/t4
57r7nSeomO/KjfWSAcX16Btal+izL/vXc2k/kGKyruU8qlnfe3acyRb9Pg0P1+xK
xzKSrFgQDEWkMUnKkFIZ7DGXkHy6p9nxCbvmktrwMoy4FoXbnNoJMWZqHVdcNC8o
ul2bx8brCJwhYeGyHeHY5HlEUdx1fu679WhxjtdMSeECql8NhU4kRfLAF/9JtMaq
N+fM5YgawX4X8U86eJx/hfLNr275eCh+ZgtyrTEXfzCsbiMobwD+0nwRrRwtOB+2
3Jao6c1V5ydgUSw+EOiXRicknSmI4KLS6BrNVeR0Z1ZbHllLQRYxR6gr5VH2rs4f
FQCc6R076jo+15knTR3YvU2J0BZu/27gUAbXDovRn9+YeaG1v21pTIaPEKusdqlb
6FpJM+ntjH2Xu3rAzmQ71Sy71HCEWqfoYgTZNokAVFtPjASme+xEpPiw1yq/gCOK
C3IfRvoQXjyx8iQLIETuauyi2LULIm40cvwvSMGudQ71U8Xxc591lxX4Mwuv9fRs
6WZPY+Xg+Lemw0M1aEuAMeaz3bzTz/adQDAn10/p1N+ZjAO11J0ofFQtt3J56eQL
n4nb4nr8mfD0AgApU+5N2RyhjzzzBI4wIq/bJABnLjx8K9l+6XFRCL+NgUrpLkKC
gDzq2m0LOKPASOGtyCY4avEQOXziAjZ8o9seMXkVk07I/R5vhdD7eGt09shjmpea
tSJFHAjz+DcyOE25rz4+S9bhIm+G5jrBE0Hizg+G3zP3dP6plDrWF0exFjThBdzz
666NZ1eb3zrBbveE7Xs2foY8CmwOQmKTFzo37mpKKCJBqXYVhMXbgnJqex8cuDeG
2T7mJo6pVAChqzUXS+8UBZjMxRuSEgZ8pFCnxXD7m9jjjOWNgneCYOdXxvZjtSW9
mIo1C6r8VYRmh7i1y3N/OWS2m45YaIAVMgWJK5zMJb4w8QxlUEj0EdKt7ubD6j1l
2gwoj01SuNADd+81swkhb8FhxOKZUWJY31Fy150fnMjYzrMnYhKZv8sgTCwugP8e
iTfoys2GwttDIbV7mjfkyl8o9ckA5tidu6ncu5rwBtZGt1Wvq6F4InLOvKCl7Doa
l75FKbPfNgBfuuqsPlilPt9YGoMTtnSxju1BI/MdSi28NlDHvQljfxKeGeqFFw7B
jSwlOOYWVLk+8fRPFOTLj6w68ZMnxTEqMsBdZUhyB3DkazScruvBDnbLGhTa+69I
xcCweZ1QlRau3UcvrFktHD5ebn0iMDs2S16Ve2tL65PW4Jw1lh5RsbyRcwHVCr+J
1p9BgGi9b51c6xF9QXd36t5KokwFbFgTyUbADXDpNzXuN11D6wO0A1ciQmnUcKCb
8i7AWLbJngT2ZN5W4Cc3L8GFhAOTXdjStIoWqIE+nQUNkuA49H4rpvd3VUjPIMK4
M1uiiVHXiZT/EtIEGZZCnxnqBp7JfehvjfdyV4LWuATHRTH+edGSNFZdruyQLqOI
Noo9wBd32dIx/iY4teiNwR8irBeXbquZmqqyxWwIDtGSwlv2EXGtbo/5imMSglOD
2gN3GyhnxZP0H99K0ZF5uyHh/C6CrrCIy3SwKnabZLMHsyPaeDx/AETQDQbDSU5S
Z5jxJuDXjcRmBQL2IXxyvToBzHEuKnTZIF74L1IdVxcpa7Ujey8s95JogcGQWyUY
+WcbQKRGCVzyptBlisaNhmH0+EbxLDqxF89b6xw2inzPpXdzmqPAkmMb41T9SGkT
etdmvCk722e78VNVMBO7g86f4gCs2ZCS94khFjULSjd0AEe5T+zd8bBELXfsQN9h
0RUWX4llKK/aKwc/9wROjlliHr/xW3AKTYaU4RssQPB2mI0u0FY1MKStwYpyJ18L
GijZNODVYCV3rh65pLwVjJS5KSUI4lAZRSP+K/DUT8Phw/16UmjFqxIiVPZkHF5a
SWa+iaTeIrFBcMeiaQWt91WnBi2fh4MA2QHAkgT3CcJ+v/7HPYk1xgo26xhpvxOM
Ix+81UqkAAgo/e/aaIUX1E/lqP4Dqz3QUPkFn6rXQZmEpJ6KDVdvjzMfbzoAt/D0
SXJfa2KuOJBouSMWoBcMgns1/yZaWRKGlPHiJ7a+Y69jkxR1c2wen7EstsUBcvMD
W48KHId1zMkCgnL2QfPtPcq3xfe47npTqjMtg8s0VFYT7SswQSZUikvW+cLEBDSs
izKJ7xqxjCEsN4CJWLIvGRjazqNQsF2RXl9C+kmy5XqbR4h4w9/8PIEuwyi/jw9t
ISbkmKV41GKGM6BBBp0Zq1c1JL/nfakzrCOjG0OExZnSqlfy2VCaon1Ky0f8Ccm+
20SNmU5N/0NBrn/rYLF4AQu8ejUdCm48VNMQAUujNDSvh4nWVQW7GF30Qpy/+4rV
aaht8lLhNiF1ZQ9ye1U9VXv7EcXusjr/j9HQPpHmQcv1+gBCntUngDeCsOtnajXP
p6EPU4F+RhhR/GgAQkB1F6xyImx7oWyXVtQHXa0Er0nkXK8luUTB/XgpgQYRxewp
ay5DNCMHkPLtDgZsOhPS2mCHsDqCV7TE6fN5SWh/DdHBt9M33gpvdSUoFe53uHs4
rUpWq0aIRGUj6f+5kIdFF+f9Y8COHJF8iwGZFsB0mMG/wRg+mZHLX4JDuPrkdQQE
Qe2adjjjDtV8++FrFcCrWEpyzv/ZHxtz9mbXP20kMH2c/X3f0n0Lf0bMXt7oR8SD
uio/GF4UJiMMzCOAVAL7eDEYKqu/0iCqAvUhA83FvyQaswxPqrix/GoL4UCRweIs
pepl3Sd04OgcpB0XkCvV0a7df4IfpB0pom7ZRgFbBtGnxLBtVc4MU4cAnqVrOYrR
UqKVYSh5geHN+KgBSYN4BxeD/ZA4CHSd9zkaXXC2WBQHdQgluJQ1RB73jbWVSg0B
k2Q8WNmTuOS7Ji5yHrV0QJTjpHQNBWV0Ioc7kjTtZT2KaQcRHveQQi3dthsct5Ve
PHkNUm2XDmn+0Pg0jI91cwJ4bKwqARPk0AgBe4CoupEdhu6EuFVC5TnO93anVMIN
8eq0skpwF0MCCB/pHFu3tGUHpbwuHztszlrR0A60FSjePBu4JWlCDWGYxJGWqzbW
9aliCeiF6iQ4I1FVqO12Fv2GPth6Bar3tLUhOSz/AnkgDkjpH0P3XAok6bEd0zpk
1nb7hYOo/elN8cE3J4f9ZyL8uKCj3iVpy/dOzGJL3fnd1YtalQ58YHYpF5rklerr
A00O/VujCSw6NM6tACxdliDjiVpYg3hUIjE4zEGLLlPQD8kwrCfnMIPf5q7EJp7G
Kn7a7JleUoqCq2VmVxv5Zu1qJIDH66EWfZFW4OFOoPpmNruFcdyXZBELynW0JWN1
WMhNbCMln9MUiEwZj7lM+WlyVwRVBQ6Yz4dnJyn2+dpudRbwI4MP89Dukfw2sQO8
fkeDIm+pTWuYNX0ljymbJuNlHZygK3Kwh5laGvryjVV9Ht1dq6fs7q1Ui0k1m8be
8K6n7XEzyYfNRXLYhh6BiJibcKVmm2+K2qBBVgIOk/It1hzJ25MjxpqSW9JIJJJI
9uDiKOGfetVyVY6My6gQW7YD/uqylcOKXvU/qvhDaaqzVAL0XaQkhXdJ105apB1q
C3ztbt1QLs/cDJHs40tQVahdxzI+WZngTu11nMdFk7tRxw/FnPdlPy51nYtQwMYM
mSBZNXUJaVwN3rKByJO8Jjj9CI2ty6L2WUXo+wBXYWhnXsCgtdc13kL3dSaFo5lP
Hp7oFAfOysqxlqPf3yZ7CK2NQmI2ABxW34h5PLYpuECBv29NqUYEV7LMNvIWlHAE
5Vb56Fhjiq8L2hCMkKF0hsTObaAbfpz3wD4yrfVFtWESlY8ovVbEiv4gRRfKCuNv
StrlhApA0r+PJZiWC6dbFq/N/AKnVJzReqAsh4y8xV305VMS1ZEqcWP7zNFRzRy1
QItB0CwX7F492shsLzg7t6rEOU8HKxZk70PHolEVEnmCxdPcG1msIOylEdUQzt62
ipmFEIavzTMgMDtJU4YMQfN2SSI1mdXD179TduYTvFT73rQwDpQ6VtJk2KwM2mMT
6a4/w3KvXASSm3ayEswxv0utGWd8REnUrvxNUNzT42m7cLa4PyhQPwRFUSvyMxip
yFKw5fhOD512LEfccHgraaqk19vlAMSpFz2zKoXnute4bCI1fittxnJ0jPsUFFIE
lJuD220L0UNhJXv243h4Nk3Do0STB335epsUcSENPwO9A22+5+8bFkvDSxqmq21p
gJ0hAXpFysqYRpXU2Wyd7KkAGLWUDadS4gHAu4fVz6/7XEUt9J0DNQnW9ePX4aMS
ohfaogyiq6Ss+WdVd07cvlebr2pm3G6d/YujK1LmyzBkn1iOOzH8MXV4+ek1HK1w
cUgouPSiZCjNEJ2n7xiw/Aq5+R0CPb7oi6A05jD2+htwQqIHkOkG0KEUUmTmzOuH
DUOxalLottS08NHW+yrso0AwXSUHy4zgLmyfFZsYVDeK3v5hR+4OK/jBaOOoD/rw
0lU+Ihw8AE9tQ+zFXnRHA8Fda23IJRffJBxmk0+M3k6a5P5JpSv3AETqBOZnkgcp
nzrpJZNJJMoLIrg6XL0y9JMVVOCtUP4WhSVdAWHodEkJn+SniQH5VdGln+o5ITmT
8s4xU2j9NfD61L0mD5NHmeIHsZglnoI9gudurdAtvmF7rF2+E8LjEq8etEhetNDM
gyuGHgLFpld+ytOplJhIx/yA/VD67VJX+k/pQ/LzVWxZlkiiVrguBHZD8uZsa+HZ
F0lXc2SjSbQb3zUbWjQH9lvWh/W6L37U8atMLjCNbKsnov5O59JhzPk22n6OWV2C
mBEQF1S1km//n57CEAjKFoA683kwH0HWTStnBehjvH5qiKTgclRkvnes7mSfQ/HA
g9HtbwK6oA8b3Xu50n/PKfYFn0IJ9BtubR7E/e7q4FB4DseCesJ7t6e3jBVGVSvl
tKJcQmB4zGd4G3Uh1m5VphKkSbt3ijIuekVP/h99Ou5ZuFn6JIoPk/aSSz4l9Dvz
7HWsOofEx+MAeUERk/cuTWWSrmL76DHqwSfiYDb1Vmqhdo0U+s+JpmezydCeC04v
VKdI+b95afmsrjPTTULd8glPNmjtg3Ur+dhX7eD9E806OqMptSEggmwHglrxgk8x
8ffpfapISC0HHF15EtTfzNH1EXxuBzkt/mJwVAPDWYUDJ2pbzE9SxGafd79ZcRB5
K8tuXq62Qy58QCy3sYvp52/wF1n7y+yU7Ls2pEPZjxn4YExbSeUDed137prf2APe
XEo6pKUpj99sPhu8PN9QvGD92VnQa53dfNdLZB666mr6VdgFB3ki0+0o1EXQpOr5
/MtcP1fOqg4IuWz5FFRA+zI85pp5jYuJlJVE14P6fdRd3KfvBEC6uaRIeCCkFNLH
Vjswo9pLNyrm7CM9MSfRnI5I0+EcxRwqXuqV8BFn7dKwyXK57CFMXEN6ScRUu9UE
R+8AirGAnceKjq4RLiadEfiidglS0iyVtR4mZ43XwpONw3qadnPty5UF/2KggTbK
BTi+JkKXILgmiGFf49EyO9IWBVrJq5KUkdO25jeev3Ac+5dEiMW9jKMzGMZHtwJI
qGYo1xScf6VULvXWualrw+eTAXogjc219NkWElJg1GmiQ8XUA3XH2aWb2Pe7L/nc
PE/WdzqgiYwjKN+P9G+NqPJpe238Iv9Atx96GwVSVm2nsTAt+gyYhoAoIje+N9tM
NXCE4eoHb0oP84AOtyMUuu68NNB0V1rSeqO0R9Lu+/9aLR6qXmg6X1ypoLzo1WjY
93AYxlOJUCSaRxY6yXTPXhrApZUtWUphYGiPagvmO+Ez+m/gdzMPcv3yKqp9et87
y1yIQYHpAroxJV2+hXBQuFQuwtDMrIXG4uFPLzzVneQM+auh7EI10xCCNwRs/+O1
9AzJS1EWc0mq6zMrkwmZr9P3xJWH+IUHARfGht/npg+aiCDtRw+G6obzcVYOzgER
0Ft/I3Qmo+zoLu44O1gtiMrqW1vtEtTE4ZAuYb8iXfM30ANHnLPlHwDyp+lMGcBg
1quLyspicii8hFX7Biz48Oi9j3Kw4gLn3v0JDWDZQ9B6n9H55CWoQGxwIugEbnNj
oGrIIMCs8qdvKHQ9+u18GgPMuGxrM5VsvYYJY6UYqBz5Lwd+fGR8OLmi00uSUOBI
rLJ8kJzxXlniUTBJ8cya8lFQGijGsSBO2cLKPnbrwt/BBb2fWnjGPt1E8O6gvRpE
9zb1y4vLWppc4MdqK6dmW0g01VEZolKRAS8Ns6dig2V/aEXZH2Ked+I//TLBgNsb
gq4bxNk2pq+o2IErxd1AGBkI8+yfqKSLJBMO5K7tWolosIiemOJ9uXnNzmEyx8dd
g+SsjPYB/LzP946o+YYM4chF2ZLV4GB0wnn53SubBQZg1Y36qfjuy3x5bejN/fpB
b8/QFCOr75E6YOY49sIdkAAU/E8zlZ1arSXkEvN7cfBN/VmPav784hpiRCZPy4aB
YUV10y8HxRxBlKAyt2HuAADuLB4Pykc+AsbCRZsgoGs8FNLhO1aJzVthzt2kZZAa
HlcbmM+oOo8mLub6eRRVRZ9lZzYVHnrjzB5BTZlPRu/DDBCMAB7jg0SnobMV+WSW
MKOMzqR/o33ewM75iLjRjubWz39hurS5uGaVxdLWBIRXUhg7oo4cucM/UY58wVZw
6KZRlPoyN40z7imTN97sR83mas+byOlPHwFoam5BMSwo41+4WXiOA791k01+qkzm
0msIbixXQ5EG7+xdd1IB/AUb+l/wx77p/ugAb3iNOhtsoniJ6Hp2z+bn6ozJx/GQ
wC/t3RX9dmE/tEe2nd4yYZ1bbwLe03Q6kAQxZbzDaWTCYMC9wscRLDheS7GMpqXd
kv/jCKcL8n7ya/Hn+cfhLUJjzzyiwgReCKIa7yug1ZxXjwt9xtk5RN9Rb0W6OnUp
lBqv6i5+2/Wd+3TgGwYMgQtK+FnUFDBS2LSWT56Uv3xKKmrFCRqIiCEzV79d7TGg
HbsbskAPimypmsJNRD9WvCLYxUS5DZnI3OBmO5+IM9GPnxVeHTDTUx8iqp5OwEkg
L1MpBMzmeDqpOmsoKaQ259/N+/qfekB7PHnoji3cbqiBSHvcvE429eAXouOHD8j6
EPkY42R2uBAg7NgYFqzF05wQ/RV8VS9QNNTQwVR8cdFLPake4AOCUA864d5OVYEo
O7/W1vaMMpcIwX5mK4wVEqP7IbobAk1R+55hEFIwQ1kGe6NWb0DDKSjLmxem7OSl
N8w+MH5bgIlNgOi2Qwd3EP46zMtQwZZgUXdkL4shmYZBGwuCjYaaz/JMJE+sIqCE
3/B/P9wIwmTen5d1ZIJutFz06QA0OAbXpt8jprmFIEi+rRNlVh6dT0MiWPS3uJaZ
NuMp11K9A3fkvrk2kyP/xLO6765IxfyglYPuryEUBfkO3TPvfIupfLlL2kpGzz6B
eU1fF192xzm3TX6nVrCWtzzHC+c5grZM/YfXdY7wAU27SD1u5UZg4XYx01W57HYF
VwkQlUaEW4rWSup20qrgb5olAhTczyboGlYZakgTU+QM/NXN+h6AP/QP5Lcr19+a
nxNqY4dcjX+UdH0xEA1Y99nrD+75W25a6vzI4hPs3kczSWqAzpihXOi/OcrEH0n0
nnis8DGNQNYwb27yGWaJ0JlUSxaEeOHO/neP9ZTYMyrDG7Wm1ri0iBNsy6muWLRI
u3YCqJPmd0UqMy2aDXosw7619wm+/58zpcmZ+RtgfvJh45+R23LNhrNFHu0eQMKq
as20NVZCeSHieJ8Vwu/1bZdE6LksPn4ZZJSU7hK1bWbiA629u6qi4fybl7PLp4e8
81qxmvub1UO7kYv4ClkLojG0Or6Ss3k+JqOk6ar+B3tEq8Eh3WXoP88qfx6tjx6k
HF41phr6ONnRs1UYKYsUS78zzyfAkFXd7pSo4Mh7K+XwIrmVhMzIrvDYT1BKtHUv
sW+eyDreKYjqlK3DA6RK59wt96NgASt3o//5wtBx+I//eABGG2VS+buwEZXO2Emb
uLStGWn+/yUWHPBCWFARL42N6IxBj3lVcV3ZSGYvfEHxrNeV2XwqsNh+Jogfbcce
4egEYG7yiBtObTiyp8JiRZjAPqCyvqOdwGW7N4nWUjYXzOmbrGSRvpc+VkbLto2f
iK1HEW5EyKnc8IDXKIuhaYOK+oNBl9UOLaxtrJxgzGYcX1L4NMxF/TZdhGrDS3+o
r9k0xBAGdXxt02VOLIyO0EAG7qQJqrpDEWToV9YZy7bjRLp940pMFv5TPE3dy5DL
iYzIcNrR4lasLup2VefwYxYFJe3ez3QFTz6kpS+h2l0u3Dnlq2mT7SJsGVeufnnE
Kuxm9pQCV9ZcTogr0BGXTIYdIEyGCNAM2FLnZlKRshp0Mbc9wmM7P623HCPkCRNx
vk+0mxaOfs1TbG1H0vxnx8+EIp5aAIeYj3uxGwDC3LcmPOta2UbLE4/Cs/iJOrXk
06gCnDy5Au7ApGWZadxvgEiovviMsvharNKRsopZN/Et2bPEOouGqFC27DTm2as/
rC1QZpUK3JM3EJHxac2d16In8QtvtVGCnguQWR25L3+JQ3z7vlwN/BcKNTTgVDUi
D7MefI3qpCY3VFe6dGi7t9dO5HamPpqOEK4GGnX7tx3QrirMU6dmZeuxRNiY/vDg
OrmTomtmnCF0/fw0AmAlKBQ47F/02paQGZMqJNscHSsX0BrSI23na0z+1s+Ks+it
YS9VIUOljkJSUjexFGxJHh8Zn5dj+67+DzfGyVJCbdomMO6iIYAnv/39xokw1q5m
s9Gy3TvWEMk0A5aNnjEmtW0b0uRTe7OmM7G8O/PCWMZM/R/uOlUFQIFtZKiRteRr
sPo6WZqoPOwF63gcSG6rO/iwi7NXgMYVus5urLTUYlAiuWCtvjK3AM2gtjoPAlE+
kgr1T01lGy/WYvkQnhpClCeKPUOox2YUm095A4uEWrz5KZ8Wd8BnjBiXeYBLV87s
gHHvrbGlW+o+zOP/suguzd+a8CeuUwQ2+W7nj4w5IzEs0eC0Q8tVwA/UOMxmsBXE
elOTsLU3zOgCWM4GnVN7khiUgA4UXClAfSu+YFALe4nFCMvCKjkh3Vr0lB73PKHq
qIS/ZRBvoRtbM+J3xB9fHD9sqn7UGEEuLLvoHASLrw6nnu2tZXGSJZGoEBMYqmSc
4BhqBqtWvUbOkIWr5Mp7yf6ysirbUsy5TSzgllumLRlaPTaUQ0a/MTPawSQwUk8G
/liUbhBB2AT+cKPgnxRioJw/+x/MzmBXIj7pBE44qPjhnBqLX9WeEjAI0pCYCphy
HFY5NnxcjfkeVCCEDlx9jXC2hJ+H6F6Jkjthu6FR4+bVwwBhsYbpIN0QgVknS+Jb
apz7tFsnXlLW8eUhP7dshA1oe3OSKOD2l8xsC+UlCsL24ET/aS3P0v+t0zat+M3s
RIgLTDP0krqpk4uIfCEpa7MOFzuxGPjuT+b+7Uf5pH6RhluHHJQno/0lEBvdFI9n
TFO83cKiXxVUZ+3fK0Q5zD3a84Vs+3WpedUznGj4ygRzoUR1rXZt6xlF9vxzgqHv
lg7nezT2ZFuDNgmE8MIpCtCUMx/DxXosBW69jI7PDpNhLN1q7vzjAtVnZmMvbFf3
U+nJDFYR5itiZKq1G/UuHMgcOirmM3IL7zI9yS0dU0sNdcF46CaPEtGZ27QcsCG4
bF0mJwNVw5V0lJMd/aVP1KNLURmDNAGwvepIGFO7XYZao2l5AHoinT4vgkMxvySP
AMZWvEyVMaqO930TsSwtoZmEQzgrv96giocpvPywEg+GiEJc7l/kXqVa1TVWeu+r
lobVmuhjQL7N/+mmwsB6RSj5GkJMWirN6+FHLXjurLmUxx5Z/GD08JLLfq+GGDJI
EGGbqtvGtuVBAIigwgLYx3q6B58NqFvZ+EmwxCz/n6WMMeMrrpcJ6Ap9fCZKgCga
WVI+tEXNTeMCpDiKalEkOq4izPBwocR5dbO065Rb3hVdtnxAxJsZKHNmDUXgoSIW
g9MyWXGrmI8ApoalC9xfiXQLFcP6rxXlTlufcxBUfmZAZavbUL2ouNwN4d3OM/fN
uqMjydEOIvzkPobf/dLwAiRNP9NF3bUrAK9V1Y8/rIIUaM7Q2ueRefM11JoZT+KU
Zl2LoDCLJiiQtqZLLhzc1Hl51DoissHZ6x2KBLHj30+gAuNSfqD9EeppOD40mOwm
8R0OtWtrKLO87JTMdpKS2DaA00wvoz5mOBm4NAk5ISs6B0GXEqQrNGiKiYtZ6CC+
Ye201PBQ+CrIj0JAoVptPh9K8yLGdTFe5cxurj4oLv6WCkRvqJfw7Aa9e4+Yv6LA
KBymCDYIm88l5rnO6leqTLZeexo/NUdgrtVj3XOKf02cck0DuAn2H/uouypoMfVJ
m6JtwgeYD3XfmF5gYYsAKemQ6Cc7KecYynbIia5wfBso9s1fJEeHQ/2U1uSYUUsq
dlmWaKRW3E7PBg9TFWkK86NVmbn1JJaY8ISYP53Vum6bH0Dy9reWqPRzVX9AT1ER
xF+0uxCkUBVCCrd5Rk9SwKGQH1zZp6UYgHhHdhkObF1M3CLDviVnjixrXFh2Y9Kg
l6Jb2J0aUgw4reJgFoiH2jDXhLpJrH7k4s2huRTG2YOcFhG+HFHMcc+TpeieokJ4
M3J5dcLtsQBP4rUXHJC3BSCQqKrW7eFnRW06/V6HsJrA8nPBJ+r/Y2cz1ygtkPg4
4A2Mi6ppUGu1wNX+lVvBnymlRKE3E5TzNHSaVLlPnhwNgSS9RGFbiD84sYXsxiNE
4T0Nd/D3yV69WbAH9bkAdMTOQBdFjc9Qnlul8VL+1r0grUiK9iuSNgennmXCPec7
5FTsQOfmQ3Z+sEvP4ox+Wx0z8HFlxHpoaSosDTlSNs0kL4Rdur/4Cm3+FSYsECop
nZem/299I4i0bxu803hh1vFerw4G9bVvJ31Lsi32iUmOzfcQttKET3YsVxHq63/c
z0bgiQUFXWMzGPLelSxn5kKTcSQNdYzekmXGxuDk1AtBheyZd1O16jXlECPt44jH
2K8krtvk9GblAFpsXYEBTXIRgtB5orXUpTy6fhck1wbc4Fde6GjugM2BifISXd/B
K8kcganeqpnYC6YI9g1Va2AObvI/vaJnLkGuiFTLBjPdob5AOmut6XBIgsWHyBs4
1AZQFeE6armVL3Zic7HFm8s+h/xOBMsZP8UUPIB9sp6Lu4RGisnRsmEWE2TZ9qyj
2JRCJByuFuBwAPLi0CiCD9KEYZ7C+ZnBr9SfRUJW4WfZw1aCs00drLHIQI+HRamv
IDumbc+6r8XEqBXZ8EGDcs4/C1zaN6IiISTvciClQbuWV2XAdKSd7O9A9zwMiW8W
4yUzQmUNd3Swi1Xpkakq2w9rtcmYsAfkAU4/n29ivX/3b2V209Z/Rb+LZN3zb6as
Vbw52Hw80kGugMIY28CHGpJsGx2+G0/u8fzaN+2TEGIadpEWwrd5Qj+poPI/Fm/U
X6DIJmWfm5aakP20m4bt7bfKGqQxXA+99HNNF27IrA28wg/oDypbBHiY6M85OupN
sdCP7QLFWTBc5rTxCxQxX8eD55Xcl1clrSN4CcF8xCxgR5kRKOnJJCPmFkRlaNpZ
74U8oLDCxkNCk/WGUJm81SUN/RPCJFFRTtcgelgtp9d3prdyDfrX9GDue2UoP7+l
Vb8qWorzPYei4Q0BBJm61N8OiXhX9AbE+8QSXZZ4iLk77ZbIVdTmhHCqUBCSpGpc
8dsX8Vb9xwvl4lz2AoDDBb/iAJFGAeQdzHG3jK5Gk45efSIo4KjuIQ9+6SiOzEzb
dQdGLBOjAx2EWI6dzAUBQWVG6kI/F+bxfMS1rP5uz+MFuX32LDqFd1M6j8C109di
InrVwGjmWCmgR1MINcpn+lUB2ja+746l/Kho//RVmeV980QYcn78hafD5+EqkWJf
4XOXYn3zE42i1VXC7NwBcANOjYpNjQhvKq+2nvd6Mk5aMMjwHjj1YiXi8RHQWZIZ
/BYrhL8xYamMP3miSWyrXdAiIWvSLi+UyIUbNzOABco0dA5i1+oKvMxDZliee1NE
EY8YUEXiWpqErvGUcMeRtvClVOFuj0v3CaDnh95MM/iYjVgUsn7gnyDkbYR1ruLh
CWTGjGVy+qQpy/7JZIb+pT8xYcYstDBv9qk3VtFbPFlsLGDQQvyNKferuDrZk+xC
hYJ/6Z4W+A2LfgdhEEZgq5qNMrUNycoMF7IYKU/GK0Om+nhIGJh+lxYQBPrNdWVL
lcDYkoAaOucXcgVUGUVuXOkVVgHuG5BXc/DnG5inRI3Axqu+r1xKRKNm86LRDJdC
DiKRuF9AqroyPzedLegyZvbqtGodpFKzp0ox+SEhqMGvFnGJujmtpQwPhs8MfWDD
fY1+fFyHLQxzxpvt325fIm3CSOWcm/NWpcpCMP++QXvn5GyAQ52Ba5KQdQcN98pz
wgBeUlloFnWb/lD0yFd9qiEuA+PxETH1XUolC7gN8C9j6yvUZlTCd+5wgjQACGbu
BZ7a2A0F3SZTttte//bkQHqdRFYP8UCFTlDACRzGTmSsYGrL3zSQuX1Jgr2r+7qH
aqoyTxVS0zBB8fbyITbaiEBZGMwzpGO3sur+FGDcUwrTzyMyw0BxyPwjRly5hUT2
+QedLj2MtCGN1dovjVkunZcVRmgHkVKuLUUnN9Y98DTSVt8Wy6yNz8TtzfMv6mNt
CflgYm2zdRI4+np1MiRfrjzs2UXdPpcCPC51F1HbjuFJ4pC61lr+ypkCjYkNhEZY
deeuiX7l2ePua5svBkww2KvZ1LCbwxo6Wz/fis851QZfQwZcIghG5QLcGc9vdfQG
+6OF9bhmR7wMacJEuriBreAUbZ70Ei6QXFcgAKxwxWWuOLKKRHBCeQYEv9tQXKRk
g3Rs1VE8Nf0ZWrty2orM8AU2veIVd/ZI80KWTrKWn51SyghToxeV0KH5baIm7u4c
Fx8/MOI8Uz7C01ay+flI/C+to5yp+OfZYhkOzkr/te+caONTZLEH1NuaHPBuwZLD
sjq3qIfabwelZUa/BQv0BYPLCvKA4vwUTCvKu7AGgWMDPzYG6/4X+Hlpfl0x2cee
UZYZuet6Q6gTS5lYN8T3CFcFo2+VRpGJqRIxlDFbl6Tm6oijcNuxqX5UvaNHQijo
cFsmxsYNWxEtA+FtuPyABI6zueOIIWWe1U8aML5s+zEKOuLa3SPHNTOaYR6r7MOl
4DX6z5pMVaqKEW2eeYMHGK7l/1C7PuF4vF+9mVU5KLuGPw0dk3cJS4YDTVCNPTew
cHhIXCdUnLOb13U6w2v7vUP4Me0oRHd7kLouoX5Mc2hyoZMpjnIyjM3GW7IqnnY0
3Ni8A27SRc/HmRofnLnyibzhXTmrm77/F5ehSP7vTy5rEjDxErJZnP06Yr98/Imt
+im1jCakRj3v1oHzRA4khUR45Q7I4jxPlGxHyNIT8XtrfxEUjUqJmW4UQPYWkOw/
obKyJZ2p+HX4iv7RpyBr7wLMX4igF9nelsjlzBFd2xN3tCauOI3kPoWKz8iAAn9s
n/KKn8zAGNrUTWmJF8s1tvl5uMYy0n8O2bR+hFVSZUKhsH47zQliLHHghPRxzGNt
ic+cy2lmAoltJ0/z4KamBuUqlKzNYSPN/GJ/ERxksLw7fDVdbEFHO4fQWojc2vcJ
v47DllUwv/AsdS8ROL3219z/0kZrb2ySmiysT3Ddp3UCL4sl/k39kG2+xHiCWKJs
oi4VxmQLTZQ+8Id+ILkTg1y7AJDfmVT5dexzTMVuWocDJmAaL5/Br9GEm6yJMYF7
zxwhzxEbqVjGhf2ZjlgZEbOR14+K5ekcMFyRgiFICpp46FTnDniYkc3gT3EtTA2L
ElrPqDs2/PEfz4h8m2UOcY3vtKU0pppu3+SkR7zKAQSFNHN3RTGdcp61S7aUMUTr
bFbFoXRFRVEt3iEN65R4a3SGAREMt3F+KXFbggkK7NxmZ8Hxjn0x7Gd5tBVxq1o8
psab3FfQbZMlwtPtU8zMokeIWcZvVX3C/6RziJt2YXj0XTg05/8hNlobO6RMVv6e
rfD5/Y5ogXDKmjDk3z0KzgEt99fC5kUneBxfjQlbOfRZEB2FdwHdGvUJwH6Tt6WK
FZScjEdRkDpH2opXwViGUSYGHmCxeaP4KisIFj6dJHUbq4WGxNk2Mz6j+xZg8x9r
nC9Gy3uDMKLanMp2G44E1MsBroCEzbWHxLSaplYPLI0M/9IU9rWL44S1UQJ2JHqo
bqaaFoXwO6hcZljlH48maORoAxSq2J6lx+TQhapgTpEy9nbFg4UKijb38HdctbxZ
0JVWchmd12GmahboPw70Ep6xHmpdVe6ek9Y31U0p/NJBfYsi9zN0O2c53x9pl6GV
xzjn+6SQ1mFe8qgEq0Q86XlAj2e4tMgChnaT6XeTT0iSbkSmek15ZmVrlaAvCGc9
DwwzUj0/Lyygr5QwIVQS9AJg/z5VlOi67uJQdD9IaqlMHTzGWmV591/Wj6mmoDYm
mjzXazMfqYxWhEAzCDsOs42bXV5V6n1GiF+44GOTkjc2DvQHICnS4IKGeOxArFak
+KChx9Cyj3n5x9bW6oHgrxzefHVLv/PTCBlhUhYmv/32BBMSU/MdKaJw4pOdRKyU
LjLyiw7Nu+9Yd+HWxbRgu5Dh9VVCs5vKCdxV6BqzKwCjeKyZduO8HTfSvCjWRecX
J4NgrhXRM8Zgf3azJkjn017fSiJFn70N8UMrHk+DCQOry/f7WXCLlvDNKbq9w4iE
BpBKY7Pw1Q81o+gHvTrQTu28oMsu+iP77nnBR9TTU/O1Gl3jZ75gCHaUUGKXKKM/
Qd50IOIwcQhZINCAK7F374xzkSNJ9Mu35EeeWe+f1y+lR3e1MN2t3JZQ7ek2YfQZ
jpxS1qUWCu/EHNpPqwz8fCZQUEYSMuNbQoPCcdDKU5ZdC/m6jePL4k43Np8RFPnm
oDeLr7QIjiFPqEUIxM+rQ/UHScPZtb2luBnpJnVMLxSSPkZzvHC6gitIAP4oe5V1
CDDV6kGmf3Ks/n5O2h4hRhJg8z53FYECPziTA/MO6fhkgOIfLIBwvmWNVzN1FjJU
RKXDjNGKfhC7uNV9WyEfFtBao4NYV8wbzfIdvWgUFzuCSPKRtNI/dGa67sa8Uuv0
5RfZC8Nm09ggtBL4MkVu2Iec0WhQQGcuMDzLvaVVCDu4IWF9SoeVPMRsG4INeyZP
Y4pa7Jg7PyduD6wJpTNGar45ayxGg/ISLc6uQ8vRQk5BfS1ixvoN07PydpJLDAUD
dxYL6IHEYCyItw3yRu7jJtOmI6yo55+17iqV7UjxCmKMNcHrfqehZMmE/NL1Spx3
5ZVfHWOsUazLWeDGbmGTI0hJv98uleEDqBNGfUitC7XMSm8JAghzg5ig4eldljEa
QOZmlPeAIuDwETJ6fPIZI+ydaMG94ZApVTlSU9xKp8WGFBh3ZUKKXCH/xP9Q9wrW
Kt8fBbB5jab4o8zQrvDvTZNDfxNrCOqUxuT/fD2lKbl0iDfRp2yUg5hO3xFAhbRv
DjLw2H/+ikrELvj9W6eQLiQuAACscrtQOzxhb2tFv/Txw8Gd4PwKhRpInm08k6TJ
S0JUbhed4ctivzfGFUyVx3aQNsWapbNKI7D9lXeyc6z2qUj4d0OPOuhUuOMV3GaT
Pgmw5tEKCng0aYpksqOil6kDMJsyNvNF7XcgqUBq39FUdOdAQTFrpotVnWHLkHe7
ad4VBGuhA5psCRr+A/HaPafxAUWNJOV6D7XM+1qUMeFEgLMvxf1UGkSYZrOKBEQh
Vn/CuPVAkUa1QTGofk1Bgt715R8LFQ1jNJFSPBj7g3Yg5y6dMU0SQtcTzmQojfPZ
LsYRRwPbDroOiMoUyPm8tadi1BU/mbif3MWYTW/XrodnMnHYQxAksEbLNSsp8t3k
b0JmFqHxVhxemmW1bCFC5aIdFiK489nDis2xsJZ8kxfF9DcZfCDsNvgX0prBapcH
ExzmJVZoOyAjD6+EEjfYhxFpMNbYcIF0kE6DtmgkbxDNSXiUeYBVMhLYbIVTTUxQ
2AK1dPx27QFWwyfP7P5eLLnXXgLUF/xv9Z/POggoBgDHhQYPmr7CvBpJB+szc2KX
0yfZdpwE702+gBrnPv8LgamTKaFVRwR3AKnqEladHR/vDXzEvtBniEq3yNpUWJQv
H18+WqeMk1CyYvGTS9O1hOnVTbkQbBAdyNHPrAlHSaJizqjj7L1pd257OUUbzg4N
5JEimidYfMXnutq3Q0TI/iouKMIaX55r70ZYNe5SXyKGYKoroJXyQzdGsUFRBysb
EEPPvVHYRXOFO+TmXUd1j1pwoOiEJVCutDK5/GnJuArwNfzlX/ZsGEyvbqqzlq11
01RuwvFq18rnNJppWEgN4IcJM8B7LxrD8fV2fgRlx4R+8YmWToJX6oQKRCcspguC
vdAvdtu11i12BgjXPlprWWzB4hLtTKGXKNBatz/edpBdFNqOXh52iT79BgTTnKdu
c7TG+eSRyocd2n3+28ea8tSG54MsS8RnjzzQZzmjQewyBVpIGuiY2v6dwjeXaF0v
xNu99egwOZP+Fmnta5LL5KropC4eP+t9zPpFtB2R9QF2zpY0Owj481ZVjmUBjrdt
fza7W5IznL6fO4OTtSBgvb7ByvSpLMiHoxghT93JkKcf6uGDOW13f4bBfLOnyBAf
6qX0lFfHPX5wKQaaSU9iVxdzpwVRtFJyoMaxGK9CSE9Q3TLyMM7QhQqlqyWkM3N4
gpS3x7H8uexTmG27HSx3gI3vbzYfBTeFGJypvMwhLFH65aoN5Q0FdUmuj+tdOzAY
5n4cDm1Ev7TdCZH1gh6OAv1LlwpyL10Qkg5nGvJSH3Inuu8jfvY/40zS16KhGJ5U
hybE0cOKOgj2u/ywHayNAFfCb8EsBvnVVK2kiBlcPCzwsg6cGLmo93epq5E6vfeD
OI2YS+tR3DkYag8VNOr+B+ekLxxpxEbBG509MbY47WzeT/oaKx9FChydnwrs+iR9
XjBJ7fW1ZAGcYAj/o6+4A4O0EJQCdPJkhDCiyR3Y+GzoelKhgflQvKP+jTFdeUtA
+Oh0f3b/I+Tx6RWXbyh1SQeevEwAR25WZ8EZNQKcSxWi+5dZMH/PACzNj5kCKqIs
Z61R9owjnyoS8m2T8lk/qS1Z7jZlX5USviR+uowZkBK5NDzg7fAZtUm58XMNflhc
2G6qdliltq8UrG53mIdjcMztRBvLS7ar0WPuZ3ftq4U3PxTEO0o9OxSiZBjPE2YM
9A3HthubH/LZbX4MCkxABVMvkWQXkLcjSGsV3ZrQ74e0n3akQpJhg7h/8/Vr7rHN
oFd6L7FpmL7NJKf4eH2TZAuHvctRhz01McKrj2qUovL2t0z7DFn6D1Fz5BSO/95G
v9HzQEPxGQgfvpU6+sk7UZhTvSS0dW4kBTP1S4GmWGHcJyEHFnoTSNurFw9Ct0K9
ULb3Wh1+aulPAH3p1sRAIq4IS9n6m69RKBtscUIL9SdFkm7gwpwN67LOeQFIFeUY
2NGd1cGuZLOep0/g6A/wv+BSFSeTSeiCgnK5CUBw9XZJBp3kd9OzSFL9CRQShWm9
C/p/OuzuaGr+5RU/MkVjGNcxjkldoqc3RPc/gi3cmHajTtZWn1qdSRDOn45RvrXu
B3J+TIPDxfPkP+sg1Y5AIv/tB+TEZgUDASW97DGwpGOIpc0DlEXtY2uZtokREP/I
OP+Go07tOeOhpPDxGqp0o1PDzOa3fHkrNh2ZfZ/XZeWM4qPHUJOzNGTePEU19KVL
YyRkz5FVBn34QHph+2yt6JtWa9z8sWC22x8A6MYzjHrXlxljIHZsmqIIWr4kPLcq
wF0d0MwHekaXWg5fbEXWWJE0aP8BzQPTvtqTPcWImRk3wFJrDCHM0FTCGWdkowDi
NdtuzAYRj51R2qj8lgcimIJ4z2owYj5ZrFNXlwhRL5hUZrIekVXhk6mMWZWVejH7
xdUieK0EzTz1fx9rCldwalUk45lSc7e6mvIQ5Dt4wW8AAQ/IOBA3Swcop1CSNz/9
htCBz5OG+t6NcMPWUeO2p5KoBafaCFjkHvqgi4Wvc7MxdxWjpUpDj0RgpKGEIKCU
9AJBf0R+Bp6NyBqxtwVGdvJhRpzKNm3q3HqBWKwtLrVyK2gE7s6CArBaWerMSBGx
NdBQkFboHBIAZGgUGBCvM6UK/PGa0JweHdKp8cReBxeUMMJ3AgMxSyLEdZ4q0LS+
85MgMKMOJHxuroGalpJ7t3P6o08wwtaGhM6JXPILAQaptO8vzakdM4x5N1iudbFc
8lPoZ0/sVqAUYPC+mzAeEpSSQ2Dl69PHNJQsu1ok52+HLrxtHDyIUUGfY2KmN0aW
CC4RBtVKD+cxgvSMQsSCDEp2+05j/PDOqP5IT/Iv+VfwXEYWvycxhL8hLOh60HBx
JB6jSpw18CisDskBaFd1pFIKYVnqBHp2RihQVgnI54/CS7z6FBGWQ/SClBVTiElB
4ElF7FANGjMOCbE89vtMdrhENgkAPceGiyp2abZFE+S2efPr/vtOTWtrlZLwfwwc
ZS14rmE8mw6xWLcme13A3OlzcHsdVUN3Vt0NbeZSc3jn6CV8FbZpji7zc08Ld4ST
EdW0D78HpeHYBGD+QZoc4eQ+bmj+Fs4LqYgcEnJrC0f4eEmnhKnyuJjsI3mqj6W0
FCcMWBWyXr30zvq5oYT0Cv0rwgAxpScnP1dTuYcUjibAw8dowyU++jmtwcMfbzdE
a+/DNkN1+RKcdKVKbgCiyc2d12K/kXnOpf5miIQJUbDzQ5NFJjpDApWO2K4Y2ply
Po6X3JHDB5cv5pQD5VXmIKcMTWYqQllHxuvxgrYz1s/w++wfM46pxCe6ZthkgUIR
YwjZ0SbLEsSywx/bk7oMxyMhXxhCpI9fsRsdzYoO7ls4iXBywXO3NVZx63qH3V9/
XWmJJV2k1TtC8hC8/PoOl/dA6d3XpWLwylMdy73mXI9kK+/5RsqbCYemJd3/CTml
bTBfK2039BxDTAyYnIiZj6P9TNiskzD6QDfzRz0mIe8Lx3TZgX4DqZ7CPb80km2f
EnLGPnturEBnOJNWcOtNNet+bxFRLlTub4L+fceIBdcFSIGKIoBuFGf7GvnsFv/N
yQdrpavYT0BHAgSDV6O06UmiKDHTvdICJb3v33lB90apNkLM3dOqzsggRq5JujV2
c2Hv2LDfX+aDXAKnJSXBWvsoBJ2jSvBm8srBSlaIK9XS3k45VID8LMO4awY1oaiw
VEgccyHcSXtdf409Nr0IF4Inl4QvOEwYBCuJl3MsrlqFCSFwJ4lKsod2OfBG2lu3
bhQpmXOL+0OrdnM3Fl7mOJa2jXadbUPQOEivTtQvPDROjc0j/MslpScNC0m4B9gW
gp24CEFj1TOHayIgYU0g30IhLM+c50hUzCL1Upqnow6jaHiCvbb3q3Ws1j9W8Ile
Wmv9iKEzOl+Qw+22t6bXVr0v7scOM9Hz5zwKpSuTa5ncoW/RBCQA9gIhEbxxNJtR
PxgA46pKse9sb7Im19Fdu9iZC6ZTGJVQohFszgXTnb38QbSRllJ9MdMztnt7cdO3
7mZf1lvZQ7daO3vc2lmihelyPKptC/X8tmgjBpQq73KYIB+lU6ipGx4VhTsozjM6
cA9+iXQ4uJRToGkUXr9EPQb3gidi6LIX4IA2JhKP1AXir7799xhz3BOfxayNSG3x
rIhO229d2kXNZ1iezlNKusmS395WtZn+HRsIos237XxV7dPI6x9mZkVpGe1qx9Yr
yogNLtVqHylsmJFu+RPxU+O95m6pulSQb9OvyGWdF7bhOFSDlFuvzmBgqGfehVaK
14kJqs2gaGCa5ZtsTBLncO46BK2joupc8YSYWuYVa6zol3GWazYu+AsKaZJz8xrW
/nyj0eoJ9BlU2FulL6c3N0mW9B23uhk68ijUcNxT4TCL0mQ7YvNndGoZNkud3tjJ
6BeBjrVETiNBH9j7+QKlsFhN4eZUL8rECl0XZlWTKJ/ZYZD+D6NOBwVaUBJG6zm8
0OEKjfxsRWe1c94M+EzPeCzaUPhAWL2ApPZ9vSHuR99d9Ov5ZkQM7+vXtbXRrhF2
NKVW5dJi8YGJ5Ko4ZezjOGr5bkljdDAhx8a1AOWUhaTI9FqnwsAWBGNcJwkOVE1g
HbhgwpLEdRSrH0si8TERdZTRk7QBMEKrKOFCJPbf4wisrT71HxlrxsttGAj0AS1+
bOXqZI9MQpv+/B/5HUDqw83wESOMoBkkJmTRI01eFRSKVmrgzOF9I8xwlu8zI77g
vqkEIW4Hv3MEWaVmF/sLZcdxiXqXaSpNxEhRObn1WEZ4akL4sbadWDZuDgO8jyhF
NYu2EslV/rFjvdNMTr24ofOyEW/uQvUb0IKmKcNfPCtU4W4fThTc64ajhMDcbQvy
JtNhvpfmz/Wf8db+XAzk9LeIbxkQb07LhGzmL3TTSMmGu6XkXqbaRbILkmcG0E0Q
h2x52kqPOiPoiZ6JqTGl0VcON7C9kTBg66t94MwCE36Q83ojLLpG6uHGLsqh+xwr
c21QHYMO5BFegtb2nq99YMdB5FpQTsXoD9mqcDQWzfs/o1BmIaNqrqnWXIm8AKV6
P5wjJbTi7HETe7wU/TmBF1e0fkNXL87YDdniy2vCMIOhJrRdcCpM4ZGclOC99DaU
RlVajKG1CZ48e0oz+f3vEgEKNvvfdbOxDVMnZd6uf1p9whGm6QSuGeBxuog65wIU
8iE/Z9nHLAKXVqYxDBDKAUfG2WLJTf60qo13BtIFV5SNdme6IZozPlQAeXb424H6
F/nFFkZrnla8L+GDNBnwWWCIXblebkmuTNa51FuZ+mfBwTT5OTVJOe8T3zuaJ6lq
lRGuC66xdntcIW5KEkjdnMKqn5lXY2NSeie/cfUNmG7AVXb2uPcgouFgr/F6x8N8
2E6A7HBN7Vi3J81JiVedH/YaU5jPc0Y5RmEqejaQNKiRJSlQhhtIz74KVU+GLuTN
7d0MqChuFfjpQKdNQzqJuPksgCaxokjXdlULqikUjLbAG7Bhh/ztsNnHmliBzOfO
doOok3dKDroL1BtkpBthgRqbKMMQryjZpaOGzSIY64TwlyPe5/dTcMzA/cRSOhnq
Gf0wQKB1Ye9Bre8vBvvlNzTrAyJ5xX4pYO4EwXZvrCTwGfKGFyOE7Noziv+IDTsN
KIhyQTbb58MJ/z+GS0cv7hB2bOuLZ6rmbgZj2z5Er5Ml4u1H9+UMIeoUbo+8nrKm
mVw81bhdLiVdP6kk0kSfMUTc/8Q4w7CLnYLRQgZPmd/SdzeCUgu4rsmnen8Jyr/V
+uEd4TVuDY14fZ5hQEnKfKBkJM0xGaLOfZQcyy1UyDutBBuc5eyT3IVbZJjRsN6h
cGsCqurh8BCLrAXR5wYo8IWqGeW1oK1m5veU2C6xQwDOPkaw6wsbPHC/ACvTQ3Id
XZoqxmycQ4RmgKmoGaRS6DD0PlwK9APDr9yGXyclBzAGhi1WYPXSUsI/jXbkfPmn
fbEKlHMYEO3WhH7V4aTFgpWHK3qJTj+4qK/TQYa/jEBlv4vp5d5icnFkSckj+mAe
km91Vne/51KFJdlrJ/qRej2hguQ9YrVXEXkDUYQ8hPpqkScz30BAn25KoCp/iYea
zZPxnrhExVR1ZfT061FkdZvT1g6ZLuaZvOpP6/I6qgJAFBzRXdshroP+CEQehW1O
O7en5DIQ+5dTZGw18VR+bSymqT36GR5CSuT9EC0e1A9Uwytj8U6Gz+Nm4KiTKKHF
Vkv4tHaW6rgS65nmQHCsm3SKrmquSZNDVAfDWou/paQmtWjy/IAwCWIKdEZfUdK+
atIRFKssoadHrosgnSqhGC7pWcTkBzgva9UvC3aEi0kSlJ1UbW+vT05TzcyGIeEI
TNrns22EsOOoEVxfAzr7/EHJ5L54V85+GsGIzsjLCcQo4E2h851khNAUxqS4HTWM
y6IH05EUGq0OkhzS17dr5bvQr9yL1Wq2kFIzuTB343+8MGCqDohoAHyJ66e1POn3
s8C9xyq5lt/hyHluEHu1P9Lc2O9lpuhTVZVSOG4CL5gljKd1SSNm/05THxbV1hUW
cNCSY8Qbej27wFA6pFjQS3W4pIDxtpe8mhxHKvn2leUO3IV19OJayixbVo996qz4
xYUy5T0lBr/M/Efi/z9sK3bgo0OcEviZbr9dyVpTTaTADQ7/gBVNZXvEzGG50iyK
Yne5gf0B++aQBr7N1Avw8DEORsdVltPGSeI/CfTjnIr+wbqAZyn5+fEhjLh/cSxq
H5YMNTNg+T8jSg0C1Y1CbSnY233bN4HaAvkyq1alvgEP/QOgH6n0go+ZffvKHDVf
rAXhevnz9dsjbda0UyTMA7lBL+tMHHgKs+M3QI/7o/Mocw+ziD0pPolVILvhiuZi
ToiRbbyUnlYyJ5a3v8GRbcZ0c1IDfDAlaKMOBHAAtCZIF+Fbrd86bxy0TJj7ppYJ
v5kTp6GGikLcqx9LOF3wfcTO1dRPgdLJNjXJLHB3wdnZTE1V3FV1h69MMeTSiZs3
TqgArjHfo8w9k6qzYir9ZXwohiHyaGT7PiFp3Yy5FMc1wLYEbkdn+kMmWePRYLji
Uw8lEc6hqd4gCFaUeyiaTTEX+0l1A8q1TToIOmqvE39zjPphxe3JcrH+KgJv6kPu
zAaUQ/DGpP09LrN8+LpXaaUg9iQEAKq0FrM/i2WXjGOyq8kFx549cIYpDGb/qdbO
sNi36SKoNEiitJRWNojy5P/+yFUck4n0o5vPtEmGHlGhxuFOa6LLtK4YdfJWMrzO
YJ9fDiUrmPiuM7zxk6I3WGOfhsD7CnomUF4eUq4kS871SFpLZqxxUS0kE4/1Tw91
nnkY5M8jvKj9hs5kbLYC17HjEkYti7Uyk/LZYECP/GPs6gzJxeBI8UCnpNDsi5W/
PeapiPR8syN1M97JnNiIb8tBUEm52cc07YGfi66H2lIQr9NUphOewH92JxdgACoY
zidMzmr0O652k8NGPIMhArLuJd5tqZb3hsq4FKtf077nnX9J4B4P4+6CNqN/FzQq
NhkYlpcNf4/3VLQD4y/xiMA9+aGVI0eqzd+qq7h2JM968cuB4m1NzOMlCt2kF6IH
crBbXraJ1dQaQz+1HrdJUfzW6qFLZHvX8/aCviZnRNeg5fXsZZglAZ2HQG+lXmQy
ncHi7n7iEcDCxNSFEsTI6RFOBKe0+yjRUxNqV0/brVX6SPSZYoC/jCnqOa7UmJk9
a5GRz+KjUGke+MRhISlwpTPlbBGoCdm/7A590/CxyEOyQRZxfgGXIYnSXERPCVgu
tYytb1V15uYxG3VvYWAaKnOSeBL+k3q7fHgbx3EKu8xum9IYexTfacWzVK8qUv08
1HvMIgAgYTK7Aqque7AYFRxzj3ZADoP0EAOMTCZ1MexxM1fdiHNwm3c7vXjz+c3L
pTzBCILZ50aUvWqfVOcbdAgnFSLwkPl0ON7QBgwrYu+nxIQTp9afym/fHIsaHma6
L6AfSqcPW20Z/l5DsKWhiyVJTKV0y6B7DDRQXtSCr5WEzDz65iJ0NeauqOE9RWJj
B4S1txKgyDos0B4NY1DRahuz8v41OI+Js7NDpvD28HeXoO2rM8mSScWuTF0Bg+bY
Ljpw6rZtoezxg6tH5FzP5vZ6ONMLRwJQ6zlMeLnV9wkaP+s/lnJOzZzUTKWOwl6s
AlX+0vy6LhaGN+F8+3lvvroIhKPr+/YpdswulgqPPqk171eBuy/nNF769CrOKCF6
2BYg5xCMNWlrjmdAngciiaeVahwmEk/PpFxhF+HEUQ37HbCJCb5xwmlC+U1PaNTF
7TlXWnAijEV98+l+IXr18D1CRdQgnUhHD392v8qcfbZFJUyexapkdyKdv/RKDG5u
lWyd3E7FL8wbUsfkbs0TcBUT9WrQovlbqIemmtCWLo//y4dqsr1dZQrs7d3KX31M
1ZtC3l+Dcz7/hML/DUhhKoG5ykUUYr5GvpRrcKfozRrYkpORzmVAkfqoYb6YeoKD
B+Q3+PfZdANltAC/znk5BHUDLMJaANycZKcwMtid/jKU0fxkVaM5e/klAChqBCuM
8qTA4vVHLh7BCG+Qv/jkKQVL42wbcwXwwJEFELb5VmhkJF5HnTHjruA2ad+Pb9pQ
4zw+Oo8aRsx5x1/Ul9PRGMhUcTIXXz8irybQWPPmAHN6H9wrY8/msLOCFAt38VYS
Oe3/VSaJqq2nKn/nBJraX32ctG2Q6JPGmV8UpFlBG0fk/gDRGFFFGV/pLXX23NP/
RTdf52KnGaOvuM42WoP4cRd2lHt+7zZqU1MTZbsdkXALLf2mNHvrDA7n07yZi3C7
10d5P2EMbOG41jPGaSoRdcyDf0UVQZ3s4JJxnfnbFuDvWFeFWDXtCnxGDlY8D+KG
JW+4j0wRBfBSYR9T2XKc2XpHU8liG0583gvBlP5efHDmoSEom5ryZC4AUwzZ0vGe
dLhdGH0NeVO19kh5/tXYsObKw5YyZt7x0Wz+mUwNz2dR3qmSvL3r+qPbkdIjkr7S
dGFclhbF3YsUPIkA6d2CEA==
`protect end_protected