`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
ddtXksX2+yylW5zu6QL2Lhnb2d1sD00763mmSITNX595NcHTEkwn0zB1Dry37fOW
FufOhVzEJp80NC5qZ/+F0Vk7Ik02dIR0elf3clrjeJRK85K4e3Hoo4xn7YbFUIms
l/8VZSb14+JVGURjfswrIyCUotIzlzVYZ6gzoZwDXIi5gQIBf/gI+KxNXPaKV+PQ
Ufys/12rjO6aI/pPlqSm0hCvftmBcnezN2hk1UeXgOIuKZnogjOsf0iJVX2aOOWE
6pD/psybjbnsNB6kH5uFTA5frkzIzkzl5d9+YDm9OyC+k84E83I/7/j+rk4L2dah
QJOvksSIzN867/4Qt8qYTQ==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="MvBXkzurAa5VTw+1JJ70nePUfoQXBvZOku/SMmg4TwQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
oRtzZL4VJ4iwysPsC8SXYCzXS8Fw2gtZTOskLcDV+1B9Nzn1zTyNtlo6lNICRmmK
ZRVu2BmCc2G+fmzynYlNTnSa7C0Cuel6FYpxCBlOuk3OF2tzAmLAuDyOH3Z1Yjzk
a0aHuoCdIRKv7BrZCdALt03JeUmXKPdOmIlkVGFl8yw=
`protect rights_digest_method = "sha256"
`protect end_toolblock="Jn9CQpRhJt4rnzZPRk+dOpzAubz7omckX1MrFd4p81o="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 2400 )
`protect data_block
gD6l00tciPUa6pDNTk/+tzLxvdHE2s3DQL3/JqqujQBC/Ei+vcAB8wM3doqg5vTg
mdfn9XB1bLOis2CVSfu295W2DNwHfMSTc/8BhCDRnTlLIX0UCJs9Za0+LoM0rMrV
T7EjVWppbP+Em6PkVKCwlmIQ7JKaifJ+Y+kjw9HCGboKYyicrgJPh4UIEYtmOThA
EgknCL0/iBtHXbfYsQJ/ksghc8kkC9qWfCRri9Nh6ymTMeDvAtn+pSYyoSbaOWXj
hvgT/WLNY9BvHOpqgB03epeiC8SpShZDUMWQZR6FJEPA45h7yeJyrgi9NOT2utnT
Qm5HhEN8IG9V3+sdLP8UskJCyhjPfBLcJo7ogrPqloniNa6/YocT6TXjHoQxMVAa
jCkyl2ghe/0rOVOqReqLKeC543O5NchPfRyWVYqO3dVmnAYWEJh1ROlEf/ZYHCOR
RMxry8FF7YRcgcEfqgn3HCkbMVODRKouI0iXjNvVf++noRGlWQPL25kyCj+DB1IV
SW0MoKgp1iRrpqe3CNB1V5yDWCaMvsjAPg8Ok8lFCI714A+vxXyIboPJwOz3sTMe
Zc3aWe+yZFcQaTpOAs+RMJVfqbBnnW/Zy7tV0rQqwFiA7tZX9EofiTzs18nHm/M0
3+4P6AEvvetmT7p/4xYx/l2V0LPqtp7mpTpZuImCYt9hna/6C6RDJCq6EVeEGffj
glR+nr1B28WwdfoSsodGCGi6zZmmdS7UCYwMgobuGru7tNMC87TUt1qqErE03jDz
NOuW0rapB20nfAkle2NmXZif8wmvzMxg/KwHXIajCe5xuwitCJ3Wo9Lf4Upq+Uue
wE8lww/lbVtcMAThv29BJ4XKoTjqZUsaguoJJdI4BKtMHk5kGMPMQicuC0qURlfz
2BhFOd8PuOxrsPwe3k7IhFLMeC0B3ac+GdZ/op+RJqHpyhjodLIrtMq75qaKx1j8
jIGvEvx4UOAlk/29+CZXaoM+0gHej6M3HiJlIxTGXiqTZEQMw3s1Nmu1anArmLeQ
q8j/fzukbZmnZ9O0iA0pE3+1AH63JB/L2hNe4Y9tKa39LQuZi9+Jwi51vwPc6lTm
Nruxj/rKEUez2fBUo3TVggY4pgscb1xGnBKwpdT2qnyF3yz0R16P3EAwgYSpTKp8
NQZ9haheOnLm+w/S49TeYBPSwNVLWys4dQCY38ddSF9IosZP6VtDePlEtRUWxYxu
tDJFYMANe+F7CMBsIvt9lksCqGH2aojZKynHtpNPQd8TWXH6W3wjxR3j+Q3MMVaV
D3LLu5AfKBhxwFZJcmytB50bloY3OXv7eDp+po8N16zMWJhCSEuvkxSNk5eDt8/n
8ICw7EvfaF5hVvjuT4l5EMnZ+fft1BiFTCL3/93HC/qsaBb3Yb7jnvzCIVwt+V3C
uCqj/6Ybps4dPWPUcIXs5pxFDzQPkyo10u696lk8ipTzSN+qHFR0wmHMWvXBgJMb
dW1yxnO6h034I3bdx2ULVlSjiCKSBwq3egex8SguSF2mvoRwvCboH/Xr7eUl5jVS
IOY4CDDONEN6HMhixMsQglO6u7Rgq9lPEqN04ekox51VwwpbalyRpUAdNlUHnayD
JLsZ7SYM/w2B61Q+hc9UEGDbvbdabA9tk+qVB81b0Y2Z8+j9oJwY6iHMAm/W0vKX
6dy2uaBVk6E0vV8bxJ3SYilI+nPEW/AadQXi2CwkIMTcoUta3luWePlgMTeszVJX
cdrD+qtDNwRZOS+nZHsqcew5tBvMnKnvhcW3O3Gjb1AdE7Fwqrh4ZeIUykKYuRn3
TsJJ3ryYHWVaUcMUmx8/oB0/8xo51SwihYEGflpzB5AkYiaQZnY+7Ky/nYJZYJhM
Vain+kHJVUr8lrd7/REwh0Jh5w79rgB0r/pNwQ4TFULjgDV7nYDAX3LNxuAjE+Cm
LCfiXUI5+4iISL2Um3alvBl2oLfZRKFbNwtX8xosjOUEKSvCiKPMdP1vDlgXumXx
jletad1rDQeQTNdzgpC+LWUaeh9exYAV/9eiQUseacFBmCNZSNO1IUdiza1XByS3
kKIx+Sn7eObGUrYcOXvMDYXMPgvz4qi3nXq7CEb/2H895pOeFQ1zpM8OoDS85WYJ
xpTa+r4enSsCdxopVcPwTNgmp7WpBjLd8Gmz9P2TlP2XGc+ya9Vg9iFV0DsTdFA5
iIP7rFO9dDf4h8iWG0XyiwmwtkUT+BlfDQkaWtFaoWxKLgLQs3Mj+qoyPEAc431I
8EQNZFfeXNzLQHIE+9/x0WD5hF5g6kb+120VoF2w2SDiFIgfIDWmnjS0ZkDkHS+B
TXlIY09DIIozUPjc9OuKB1Cgw+wrK+4GDQ+KzR+ATEjFuzj1wSl66MGIx/oTOJVE
RrUbmr6gO7T/ZKbj0Bz0WoAFu1dFE0r6vq7dj40aut0Ep1xYYLwDzDN23VbkSmVq
J2I5afwr5VPuzNuPvyxrg58v8Edw3uY/8jCaNur+S0cFXkqSPBw6UrGPpV8RZdmy
iws0i71vs7CZzXN/4ydX4x/7lkPItSZH+qw0t8sMQE4C2/r3yj7H+pfSJHTyBBBV
/Urc1e+94j95OUPaoybfjHfmZddklWM/fpoVXGVgV+OXM5BolUXF8/68A718nNa/
htalrRJ5CeIIwsNgZhpFPLrpssaygZYbyEfo5Wr5osGo1HqXv4Nchj7bxDcum9B6
Bo4MCtnl6WhN9yp4x/B0mtX/ZEqYjgrW5n8xCx+T8iXGsHRHGen2MUv1CHhz01fP
KG/C8ZhzEQmhEMC8+reOuhajSsqf54pm4tfxmOca9D1Ei5293TD/b9shTZL2u43U
TzVWOLP7u7YUrVlH/pDQlbp3cHvqgTJjRKHpVLVdUYBzYMz6MROTk+wikl+reW9+
a+RfYPpKCRi6e3EdWPAuGUOfKI0ev6nuv/IPmsoNZnbMWJTMPEw+jgtb058oUsG8
qBS43NTo0IKTmuqvK6oDkAOQKds5MEobma2mMQFPVdF/UYxqJn8+NvC1NoRuZu4V
D5E4DdyUhTSA9oB6p+blxtt/CZ2xy6wdO1UUMncVXNJBWiFfc0IW0d13Oc0vUdBW
5Po8eEFGFDgGxWMRTc9blwwFoJTpxatRUF3h7eh9oBBYnvs7t8Gps0Dz/KNQfcIQ
WR4ZmVj0jZieYNqQHh2h9bngZf0XO8eWImuGRB8AsVPr1A78EVF8P3sKDrGGog2B
`protect end_protected