`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
ddtXksX2+yylW5zu6QL2Lhnb2d1sD00763mmSITNX595NcHTEkwn0zB1Dry37fOW
FufOhVzEJp80NC5qZ/+F0Vk7Ik02dIR0elf3clrjeJRK85K4e3Hoo4xn7YbFUIms
l/8VZSb14+JVGURjfswrIyCUotIzlzVYZ6gzoZwDXIi5gQIBf/gI+KxNXPaKV+PQ
Ufys/12rjO6aI/pPlqSm0hCvftmBcnezN2hk1UeXgOIuKZnogjOsf0iJVX2aOOWE
6pD/psybjbnsNB6kH5uFTA5frkzIzkzl5d9+YDm9OyC+k84E83I/7/j+rk4L2dah
QJOvksSIzN867/4Qt8qYTQ==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="MvBXkzurAa5VTw+1JJ70nePUfoQXBvZOku/SMmg4TwQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
oRtzZL4VJ4iwysPsC8SXYCzXS8Fw2gtZTOskLcDV+1B9Nzn1zTyNtlo6lNICRmmK
ZRVu2BmCc2G+fmzynYlNTnSa7C0Cuel6FYpxCBlOuk3OF2tzAmLAuDyOH3Z1Yjzk
a0aHuoCdIRKv7BrZCdALt03JeUmXKPdOmIlkVGFl8yw=
`protect rights_digest_method = "sha256"
`protect end_toolblock="Jn9CQpRhJt4rnzZPRk+dOpzAubz7omckX1MrFd4p81o="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 10272 )
`protect data_block
gD6l00tciPUa6pDNTk/+t0OO0nC/UTtBwLB41d4inuAUA3i/ALrNyoJVcBnAmEQW
ptbcNp5fxEUJjnOxnedyZEuEBxWRieZFQnkRdF269oNqhn4BFXtpjb8m6VaK1aEu
0fVboXcLKjdKSrTx7foIyqARoQNAlfmqUY4KLKq3makXR4jhOVdZGloyqbJEKk3W
FbTQYOWekwPH9znidHem4z6MnhdYVH9b8BRSgARSLLB3S+UpFmdBM3jR9fNiu9AS
lLV9txbsZhwteW9Yk+5qZs2rA9kBgSRVVJ7doXyhzhi+TTTp68kf7iZkC5QjhiUi
QduknB/kE8D0A2r2W7GP7B08S3VgdglQlPKlFb8sS/9z7w57xAFIaM5OEYJwUgey
exZkbAsSux07Z721sFhYNJIpYIPLyyEtGV/1j8Ma+fXKstxmYhaAEDNrau/rsayH
PSBayvPiVf30aV/lH9wPm5adSwMUV+HpvyUuj3wqC4JN2K3OKorABPe4CqVty3+Y
rWdxwvlBIM5+C/mR8f2gTr+O8wzR1ZgPqr7owz710ymkjRlaKZhz6/MEv0Ce2c2W
4NiBCib3ZSnaB3LQi0ps1WlvV0mC+Tm7Q6iXX5tGVCWacnKu5pH30GPz+WIXi/Dg
hV7ud9qRoHDM64sv6cFaSPw2qzyFduhCNbUWfToXGctC8d3keMyrvKC3DAMvtFMn
8+I3vKvqOl193HTh6xJfjoR+tXA4EBOn6Vx9RloZ9Ufxb74wmS8QLpyhBk9bnDoY
2N9kQSLJT5rzJb4p6d6aeMWByS8kgRWBu35ZCgfZYRWbIrcZHpm3gAXREHIFUlSo
xq50Zx565YRyPELsIlEdWYbM9z5Uq8DMlclKilnVJl0jdpSMqhCEFu+LcNdZinPV
T+rY4umVvx01rrTCEhEYEYQGXw3snxh8c4UalG359dBXz3i0BFxAAvDTfaPypHEp
RerTfvy9Idh9jy+EZo1rCBA6/jWAvx6dQdJdHBWmsuJCH9j03uX+efhEUoGjvYB0
Y1/zYv4XoXmS8XRwnXff6dHkWIATSoLBMFiJPn697GFoybZaTrG8tGNHz5xgqfnj
w1sSLYZE2mTh9VQxdrdrYv8ss1nY7zn/SoWQcW7hIMV3I88N1hz5rHq3DAsIOZ5R
w9RnJD1+Mm/LnM5pa3TyxjN0VoZ+cMd8u9RL2gobzwfkB1WAzOiNVH1h/Q5B2MY0
Qex/aKhp+uK7bOpfRRvviB/eLMX2MDbgqN8+RPUeVQV/waNl/q7miiIF1KjkhcIw
J4K6Wpk4sSkSmtpILjkpRQn25NDAXm5u2A3Ot0Nr2ov1ue/nQDYd1MorbQCHCSSP
jvHTX+fe3s0LqhqC1oqRtEDZQIeQW1tHG8Oywu10Htg052J7A6GUDUu6/JIdvn9S
ntnfMX1lbr1u1Da9nLi5r+bKmBqWvTzOSvpzNLuEathns1pXA4DJov4lWSjfdgUG
Ut1z7b/mFS5iYy27cycDOK9Tw69HglmVMsjw0njFq6PBxq8KL65UQYdJ8/JF4WpL
IxFe5JpXHeKa5E8vzC7BjoJ/w4suGABlcOfezeUxuxubAxbwXVm5eLiLt8fUkURF
56d0FDrIt3+CSBAVX4aVrXMXsENd+WJBH42u48j8VzCMpi4eBmeWfbAgyhlBC+uG
QJxd56NAa7Y4VFam+Wk9SDBetpSqRReRTeJJUYVp9afHKYd6acJbg4xOI1NtdRnG
bC8wqkNOZy6gDOqZIbdV7TKpXkTidvr4GMjZScRu0UwpS9OtfBrJ/Wq6NoY5Zeav
Y49VPcr4HxBGD1IhbStpQaLSbNaOF1j4amKJWSkefpyBexefhGKEm08+TeJaMRkN
2TpvyId3p5JZI6fxERcoyeJYEOauYTrw0LiKA2RUpJZsb6gPlUnyHGS6pFhXlj66
7L8JJKtGIKYSgplJfKOFYGL9h3dVxrQIpbx+aEoKHOU88oxVotezzQicPaZ2dKMQ
eShQeJ9YB1JrMgfmHAQwGwKlGVPegp95O83V1BlikeXhGrt2jLIwCsf76Ju6iZLU
4iVxbzM2eNH+5o1CGjbJ1cbXyKllgNcKR5S9OEXOfe2/nPwbMt4ORLRT6W7lLYfp
+hqQwaIZSKtkO+qNaeCjKjXU9syabOT2m0xfA1jwVg0sSGiliuyRdjpKQdSh7WvA
IMFiSPJpySmlV3qREyayLi2ytYIK55hTpPJx0iKxHCGg9R24fXbf1jjuw4sfSG8t
DhnO0g9VR9IqnN5nGnXqJyNEqydsxBp7DpLPNF93ITBMDDbRfOYCrUEj+XEpqFkc
T71AMSHhQLKVAvQHYpGwiYj+f3EIsssTRLHDnacs8Fg88+TZjHkNE28+sqmZzOjZ
whGK/1Q08nzAJ8J/O6aLN6NHE25K2KHeHnhCdRraEOkzbWxzeN9fqrNgefOvRj6+
hhsU7oWXn+SuVMOnbSLRfq1izk0WX7zV8WXTPWxC4NZs9Sufv/Gx+GYJ+jH3j/Am
gj2kCwp2ZC3slj39LTNwcp1YbAgxI6YskxIdym/BEeqQH+z1dj/gqRJLOlxMfRsw
3uJzuPLDj6IHu/S+CwHVNI5kGtJOM6HYieck5fOWfd0LTC2OWnHzo9Q8v2ik21Zr
riA/3XXLqfVOo9DY7HgLFHq+DRJVlpkkrCprL6XATb4tyVhVMTdARv0vkhJl6YAj
6B8C7L1SAGnfsOI8Qf0xmjzG4LYrrb1p/g2jRR7FZ4ubhkDLzE7hWtzzlQyNWeM/
WXvPtVw7wk8qfJUcStQzqONRrl5foNlZbEZMXbQqvZx++z/GqnK8e2x4hXANUAI3
is5rIB+v8fBrL5kgvROzlRSFlrq2VzxKoLuqUmjGBW0GJEKvx/KtalWmoxFx4mQQ
Wb4l0yH0xogq3HIqHn2vdoUg2dgC0/5BfAou4xdbhrshmQkQiIKd+Q7MCNxDO5Z/
NTFHmWiKwQ+LfiiwrlKZRLVy3PDdFXqsHtD/AmEh8qcCe3gPncOl8HYVJYaBE4ly
AnofLHbNgXaasbDsazqYuwBotGHvSApd2rg9/Gqh2Hg6IMIH8i9NQ+WKKp9WItCo
jalLoFtvO3lTPDGDu4L1gz8WjX9kpyRvI+J9PXcAoeivktOfPfpbpJW5qXh4VZl8
eJr3JbdtsM3FZEhl+b2ufieD3WZEGWn7Sjn+56ZgsS1+T564Pqw/DlF4o+eFKTO2
dhjZHxAja1icwutpwoHrq1EHABuSg2+iONxUrkc86pwiCLRO87SlLZdGnBvLTMli
TJpOW3s7dME/TdQhAx2qOZ8qolvOlWvKX5m8wYr3q8ulbMESmqyI+iPEdqtLo/TB
FAhImfuBwE1soNZ2o0rRn+MDp0H7N3/KNYk8w893SwSAoxH/sUFuKpR5CbhwhR0w
HGaB63Wx4+EVNYgQPn8YLzzVJ3OJTzk/V7OjWL3mptqUvTvAHWvmIzKxUR1T0uMf
LnJet4Fk5CLco3+CTXhnrzr6zREOksiehbqzspdTMQQOSfRqOCEOIkGWk7mzWTux
DJsrzclK6EEG2ijUv7TGl2SK1JaP+mWwKl+Dg5j3/m4Dxo7AbIToUKb5JvRvAWju
VPWcP3vWCkCQ+BBkK/rJ+SksugmvEuV0KjQg8I822ai6c1eCDOtgRYVY8++UdI6r
SgGJQQK1cf9TeefKT8FRWzUzvlPNMdIgqOAuP7nIKac6k4teD3XwFMuKSGmdyq0+
aseHxOKTrk6OI/6qtLXkuAX91d+uSU8SN+MyI2bqCZ9bUcFSeZNjJWfKj5zroHar
cyupVkPZuZmiM7ezcfTnmplpDSOfOUczdQyVG8yqgcX2AoJUJV5y7HJhH+AK18pj
j4LP6+aMeqUHbZCmTcCIs3DRFqPKMKA7s2BaIN84uFsQh1hPvlVos8n+8mmF7TkQ
1DhZSr9GeHIZ1rNjt1oC8xh7wFuaRIjtVFxq1PmpI3Pnp3JjOcECYwTAzStmwzlf
aZljR2fNZdib9KFtgy5jubcuxK2zet4h9SEHCQ9Un+JrvPo/06nf4vhUKwxTmyFw
vDp1BSyHcSzIZdvjCwJImp2SeU2U+iuc343EPPYI7vmKBa6ACHN9YSgWK2V4gBpa
1Z/rmayG+tXRDc5GBX/f91tKq0xJ7LVXbufxCGqfEbJg9S22RF4byxSUSE6zG7pC
Nlg79PW5+UsUf95Zr3pxgoFdQhwkIG2MMRt4ol1h0+Vx2LSGJr65T7J80rWDmvlg
g4LJxgCft5+UOayfhPMwaYNwFj3AiXjDiJ2urlCdNviyMYplRY6GAOP9naLeCCba
0UBq4Jtkv1hdHVnbG4Mf/OQdrzmJcTWjZapbcsLjRlmEAm94KL7QmySqNUB84lQV
wrIez96MeiHh6YM9UmAjoYRfT12Oj8RqHZ6AYAP9cE8aiEgOynN3jqu3mYRvubEU
/EnUSUIIMf1B8QgqghbOayqfbsIS4WwjnKKlQlZtDAB4N3w8zmdT18LUIu+jIBob
9AsjsW5OTPsOAeVCCWwbNGeGhXpPYTQgZ3fcNG9yxirDwwUiKXJ07ChPUpmYeGxT
icugflxpB7HT738KdW8zzgeMW3QEHPW7qF/S8Ggr0MhzzdYHoQ7UYaOs6doJ01xG
DTd9S0V0HUc7sM0wdFNyzFogYU7a5/NOI1refXaBy4wK+z2vCMG43xQ3xfsB7vgM
ZXRuIaVjBlpgkZVyRbswqk1INXRhg8avE+BDqam883Uz070A++5mizp1MAkP7QPX
BZ7PO4Eh1Aox52TBMMoGzP12pX7ncmeRqqUcKkJDVd+6+tndbPPr5m2bi0vfe8I3
I4FlvFMQu48t8Os4Cn0b8yNSqcb3oMFcX1nw2OgnOeUObkEcWDc0LKFEFRDD98Dt
keeLxctII207foF3Has2M376nctBj1S6HqEigXJVetQqnx63JIp2v402PvpMi2PW
BKkohTIeg9FdOLaEhtPsO/6O3etd8wbsMlF9o9SdIgDfjsHfrD4Rpzk/Avhqpvmb
7FBkbbK+uKzSBr8KtuXKkAU/5rj/l+xRxlO6RpkchvX0Hi8Ll0dL9NceDk3PpZ4v
7z3jcydN9PnI7aAtRjQjt+RpKc300t6CG8fDV2zju/0it/rJj4h5vQf4EveSK8jS
0EOyhnhSjPkgoWsGZcygUFn73J+cbGu1d4VZElhKHx3JOZo7mKqy+A1DVbq+eZ2j
KENa4N7LVFD+oirAUoSYwqe9ZrGwhVeSmH/mKhZ4ZVk4viYso5u6xLWMh/uqiulP
8zG5Xf3YitP1H6CYcg+NHoauIizIPNAcyyDsgEs0/APTp3ujFuFMuPIZOUiObVmK
MwA7nJUc8tJoq01X8d91wMbd9KpKId71SErZj9+lmDn7E4gnrJGfbGirt4Jptocz
hbf1mdGjGX2Mxm1V43nzD3VgEdzvVMtb+BOIGyujmgRju9Kf2fcYGr9lf+OYuIHB
U7DMmOE89P1n+62h8KnRXziijbcevn5J/BIjX+B+/zDV49ieQ1sddPJ/Nxw0QMgk
i34p6ozKgUPYbcktd0+6Ib6cLuT/qqB5a6CySErsKrDhydYrIigB3145m/yz4B7p
3/wgpBz7YQ1ir4Fw9JqG8sgyPl9FLkcUCCLhYu/T2oRHNcC/PJtUgtokY+/yVM/4
pg52cEupgcLcr2p4tImVOZg0DYui0A5ImDBoHqbbDIkdKvzaOxKpTV2fc9PPz2nh
PP3pt50/mhEfc1DmOgDYI1N+ramKq7F6E9oEZmKtn+odKSiFrMafEKS55oia/9FV
psfYco0eLpFb8expTxLeVRbpoQ2gn6pbnknWCWxMrm1/E1GFUZ2RDtE3G4j7JM1V
xJjumnqmriiSBNx5XcZ3pLF0ADSMh+0dDfTS710s9wbh9yhEKt7lxXMjbLOvFgJK
4oDDaRbuJdlFm2UCwDcPEybd5fxM8fARKNBxy+EbbMYL/Jg/OOh/nbKfxtrMASNm
GbDslYRG3OhLKZOeQ6ruqr7mW0am/WB47j646YVtywsm0Ymdjvjq1YnrgIzOgnVP
SxIr9Dsb4coCu4I7KHN/DRd52QI43M2l8s6U3Ri7Kv3Mdaw/QWM+b5nL+fSDFni9
/nuIx+lgBiacD5EgNFOiMxvTBBhP6ZcuS6sOUU+M2CfUMwOULeA1Jn2XxM3Ve+DH
OYmGqR6gJGjadnnH1UXmAepoEv7jKnbIHmOw2v3pdxnbYZ46b3016MrUC/TdAQd7
6QJj7Vjy7GwaGaV6HddKRnXLTVRfAFC+GeEtYpYjRG41UqJcz8p7SMNvX8p4EUuY
Ee4NO+gobXi1hvYHRhnFdt48p5jbqmI8nAlxUglU+SRcaOnMHOoFR8saYBq8sZYj
dtYsCs2Mru5pjKATLUtzwsCgyRpaTD8LrAKkfX2blAAfSt+aXw8nEraQmY3Yxxm1
DD8VbvYE5UzVDjnmxkisJVx2E1JpN/v8b6vVAJQPN2AeEpF608nECPgJ3EKAU1vv
34FWZvbbGfWDvIGoKXG6VneJUC13qAWa2uDT/lDh4S4UrO+GtGhk/9ZZcdYZdJzJ
TgwYWb8wD7eFdg76/eHGx67as5XNk1sP8VrjMWbWsC1PM0Sycd61zymV9CWT10eZ
6tDqux27jQNgZxkBbj7jZk7gVJ3yhastUK2pLCk+3exshYsUlEZrnYBrMJ0d7SVV
NcIEqfBTClpnmv7gwoP9RG70E+zw6lT+r9Cxzhd6F+MK9Rc0xjjr2zftWKLhtZ7P
MxMmDfFDrho/ReCI3ijfEi1f50OzwYDSDbMyoZsT7gszZv045eRxCX0KD7FGWxqn
dXtsj8xgjMZODUaS2VxfwQtxZ/NcBrykYVN33/D59s7gttetnPzA+AlF/TFif6Gm
ZlCvMxS7c2+VrylEXRCNp/722qwFur+5No4PkjQ8gX+zKrzBUnQhX/9apEFcuyFi
GnV3NiBdw+4s1SJo+3hpwSl7TkDW0sF3BE+K2pAnlIu/Rcl42qnkcFrUkr4h7lk/
1f2+E9kF95m6HG0Mgzm+tB2P8LzvlricoAV8rmPcU6usBuLmSQqIS17tXQam5Uik
UmncqGQN4s/WSpr3YIsYasgzOi6BMwFPRYi6jAjG1N4KmJx6jSDRYnnVUmB/n0y8
TLZxdWdxeH1jnX8JnISKrDRXij+SyERtGiWYVnm/ZPVCeofpP0SZLI90SFafdTcY
wdVkxf0C6tjCCI1sbPUm7HOz9eZ9oeq2N/xpwtf40H1IQGpfV0w8cEhA0ebcoyO/
xMJcPbz7OL7qUt48FYKOrmZsd82ypB3MahmR3ouuB1gvJNA+m3GhmMjUSvC717YT
cNT9KSxL2qTEnhumfyj7S0vuVLx0Gu0y5JXMfhHHefSZAs9Bpyl2MeKf0Zid7kcP
hyQcvTJaWqJvRdG8jKiRRjNFEdz+LwBaA/HB/KJmruAV3vQ2XWJBCcd6WvHbaCw6
HtEUdK3Q9bjKpuL326FbASjuSXWBKRTHjiLTq4hMoRDQGd2hQIwpLP1GXgRJJtyh
yf9B3sbG4Vd6l+CL0e2CN6KAMGxpdvd0MaPnET1E4EJL22M7K27TLjavrrokEBy1
aw/8iBLGxWK1YUDk/YKSFheWGMdOKjlQqSU0UkWFixP/dbWY5vvytdE1JKwzwwpu
rLCinyt7KBeZqOnbKNZkVUowXfXKasT3pvnhCGKSnIA/Ukvjmu3IXf7VEoyCXaJL
IMLSduC7EJbOtha7rgSGmnpxio6G6tDmd/Xa4uYhIDzQw4Roe/62oep6Zvlcdvr1
WlzWY2X7JV0YUL6u1ktrycys52OP/7GZ//turv3RKhE/JVdLnu/zu5RwdeiB9eX2
SbyC1FbBZ4ygATU46PH8gGVkFX402qr3m8EAkjgAuw41N3wU3KnoFi0MPoCkJQZK
Kk/5drL6CnEtTwGkm/ZN9lzBrkXCsISfHMEtXdOsc8TjW0bUk6J+CTYDBmiVGUuP
RGWWqvjDjosMxrDf87JM0zW9GGxBocDzrDfVP5xzq0aSBGZQRF2tpGyPtEQdOlCW
dZngZCv9+NjlwqFsA3u0rlDskDLHoHOMdy/ps71xnhm0XYC7YpJC9TPFAawSvlt6
MLKrdBNS8CM7VB7uBr3blTVYG7SYh/IN5GyUSF3Q5maGT3crCwuD3wTLttj5uC52
eBgzfzEyqwQTgSR4mM2JxJQ278nc8Kug/pH/OCUTNyq0d/9gz/Jf9VaKMiVfXpu7
DJ8JNeVm4fgJfhBXkzqyXT8iOgkUDzjLh/CwxlvAD6EDSDgbUaLHCwf0Ioi9hk29
s52z8NGDN6js885TFlKs5HqtTtTnuiBeQEbPCCaAdT7SUSPKa6wLA/OXo0z+qdIZ
JOl2XWvvdEGD6xAh8Kcwr4wnRDUl6ljhRtYjLibI0E+IKH5jbL4r+t3QD6zG3G8b
zWMlaJvH9KIMKdXvgJFI21HcDviSMRH8JuKRyAEylYdA1mtEQpZoxnLYtnUSvQxW
T6/DoVvCgB16MIqMh/eIId8m1REtL5CQRiRxkAyMj0o/BjMINb57g9lmUdnT1oK9
sxM4LuPJfj/+VuECexXak8S2Ykt8wVoW2TzYd/R5BHty+xD6G691Ygd32DXSUeHM
WomC8HCfTg4odmbCfaY8E7yBopOYr1FuUmMpjhcZMYCrLi1d1k2jVxO32dL2fNEa
WP8mf5mJP6rQPPr/z7FIAZZOEQEsEJzFTE8MjNqzmNbxi2XhULDcmCNmHQe2XgQD
/JqpESaIwM7DOQyiRc+PvqMY9sfSoc/qUtyHMlamb/E96z/6vw7Q6hOxzCEdS4SP
VSIneZrekFVFgbp+l926l2svc2pch1PNW5yq66WWuSCkIlgVkSLoBYYyduEBEpE0
lqPcMGo3/9QzbrqLXKsTWpoRYRjTvR5aWrqKMoVtrwVy3+4yMBQapzf/J4AJ6aKa
38qB4TzwC5BRuFaqMhIE1Jl3J1PaB50dSlCzrgWU0maU28wvt6mrTRdxF0fINEQO
HQuIBPCNmZCO8jeqzeHRf/ZyjWTGgxiQfP1/KeIZktS2OM54KViOET9ScyLui7pv
0NZa4OtQtEwIJhM3+g1oaxvUb9S5jGm99k6lGklupqzGcxEb5tdir7uOpB0b2nYv
aNKaWSKHlQN33oYTHa3FCDEemf71MCf+/2eQ/3hAppxyJcTqpApi9r+egD/2NDUf
Y6kt0ME5cg5VuJa0Xh36bWcr+03+qs5WjU8iNC953nfBhWtZwiPibpbnCBIzVbBv
D0+CrOvio9fxfo9fyLlSXyBERm5S668GXqBVxqXxybybpEj8HQMJAm4RsOqcBglQ
pmVN+VHEEomtgALHOqbHeeuUiF8WIx8r5f0VDkhr7HH5Fi1RF9hFLDGztUHk2dAo
ZvVWQfI186bG42kVrrFedLLWSWBMnOO1f/iRPG0y0lcQV4or3g6MmMSsJglJfLg5
zKjCgvrkDEk1ieXbvifu24kMDwCPs9xxvX//iNtnfiMyKw0NcGSKW+gYrduLFUG8
yYIItpN1ZyasOk6AOMVI7KOJPGF/KUUra5kV/FtwnuQky9tOs8svQaybNLNv2Q66
suOS4OKzlj7CbfNafDUvakOxamPgaJLtRtekG4V35tJGtNro6Ybc2527+HRX+fWa
y3ShilY107PEL+MNa2oCc/ovUf2h4Z8fo1/OOU8NgoVVqut3gqTVFj96PNao10J/
I5UlQejjd40DnWJwyEMyAxlJozDovX3m0VSxtRoWjKD6ZBIAjdoz9+kiSVsCntcw
Fo9V9Is9ZP7ssEja/aaQuD3mACRNYUiJVaSob919butEFfd7iZZppHHKUVvgk+0U
w3eiFpgd73pQRbl0UQuaTwcZ8mHnWmYMWze4OHGoSkqkFzS1Kq50RenuUshpuSMm
Cr0egv1iET4W2FdulvMEM/cfTzf29cCITmQAGtPEvIM7la1vbhavj1bzKfLULsRD
MVv6xpejWLwiCk7ej/uzR/y6uTAWjNuMYvdDwt3xp0C1ZSjS86rL+2V0raTeKLc6
hCGFUUXqyezIgkA1rdB967M+yaldWK52yY/6o8CRDOUoGofoM1ACPWejxhxwZRP9
knde9j7q+K7wUZNXGgmm+pVbsGlnigOtoAF1LRsMwZuI0k/g+JwZsdCU995ilhJ6
5i9hyn5uJjkdV6Xsu6rk/6Aah93Yru9xi+fNXE2FjwPt5/ZcqjCaQxXL8Wu1C/Pz
vXg10o7bgcOCunANgZV8keEYeU90BeKDVofB4+WceX73JYdHyPl4wAwgMNBZBCPr
uvQO4uNnfYBNaUNaWA421lsJiKsxMicwP2t0fF0EfAo6VjQjumM/9R7AOjqwkDkW
SbpK6zATDDVDPjgNUZk3sI7xSyEYBkYP2KrPJIK+76c84NGdxpyambwXJ+wDSFZp
k5IfJ0n6x19zjnzz6PtdSoj/1EjlJfGP8T+/lnhH+1MXepXZVTBJPKTPbGVgyw9+
7KVM0U2KptmjZRPzLuSo47Y3cxOEGzslkZvUYR6dK+Uzh0tFsCWQfcagxtKKGtI2
HAZ+LdAppQF6zqXw0mSggsSjJgvtnM57sSBbAYu9UQhXkVOhZBe/bftPlmNI55aQ
9O8mznsHAi3QaoTdM2jJv8d+6Vjfro9ipiMamdeG90zB9w6wn/ppF9bevcYrHptt
kt5Bey8bIUe61sJbbf6dSr2YXg/qX71kq417KaKoD9VzeOMNaIh6h5cXfGltJk8H
UQ96zkiLmwKPaL081rrPazSmOTws9goz/CwLVueYWNUSxEql6O2HV2hAIitQeM1a
uHLI0vWXIhWQohJ9u2ajTq/dyCNlkEpyvEXP8wS+wZoYaiRUzK4Iib+Ez44u8EXB
rHDJYKpX6BoRwIr//MrR7aiA9OBxJyvSb3xltcoKDCP39JR3aiczGXcIIebz4upx
Ks3otAS2rcLNJxEZDGd5ajCc1lZdck6Zt0zEAVRlx8pqexW1Jk9908gBYT38TxmW
2omYlA8DLp0HfXkeP/F+inmi/oi5hu6YPh/Z6KKO2PmbtxiCYfJm8+inxmrLP0DB
JCQ9RTi5wXqbDFi62g6jmEssz01ffghz6t94eCyv1kGtSbUHYpSCiw1j15ijsq05
aCuBA1nT8IJ8BVnC8eJtkRlD7lhhtXmslZczAVPUjGtXBE4MWVVy+OBe/65Uvu1D
6k8Vs11PSX4GLZjp7xKoSWRDySESLlCQaD5ocPMlCmyRyERWuIm9L1ArC32Gn0/q
nVIvcJ/kfu3rgpT8is9TswqW2GI0HZNsE1azgCuxcxNIgocgHheJcjro7j8bhhlT
QMg9TVuPedrjX4g2F5/b95VZJeIyzNmOJZUEM1/DHc8uH0idILoNXQq8j/3kmcB8
7uayDNUjnbqqA4juz5sfewqPO+IfWW1BUO9k5VAtUaExEK8XGEyFPT2hqxWqFDFJ
m6MZ4vT8Sg1z0ciDVWHOSrPfwe8WFnM5QmVPgcMNoRhZ0aiKEcDmUYzdDeypp1r5
h/dRGiEwcxOmR+FDlzgKa40R7mIhm6oDgOTPV0UdXZMw7Vi/uhPyySJWkOZaUq3N
+8Hr659UGfEFnoq+2/m0kxCzuFcosw+l2kTid4i2wDzeY8h2XAmNMuu/dy69hw07
MjJGmNOHv1sbEn6Q9ir/FzKmFfsEeB/ndXomWwjWhkYt2ZHWK+KGY2fW0p41QUaV
u3685mAoWd3JiDKHWfLR535/YaPl7E9KnnQpBpnDOrewcoJyy2uvVhVxuyJI9R3X
kxfG9fue8OlFkiEw0R9JCnXIWgO776Jbjjrp4vHEQExCM5XavhTiwMSqLvblZreV
TDiGvFUscHeIDRF7JSOynBGeKO964qfSonAxvbNqnUBNYA+mshreCkobiJUbYc+3
0yC1d252I2FGXUq86koZKQ3+Gm2MysQUy3SxjFIWgyNulSfiMq+4/S+g8H4ZWtjH
QTd5PjT/K97sqrcYM2zJ2ypQEE+0OR/l8spOZ1BJfXMAtHGzhUENBrk26RmgrgCc
991SX3gnFa4z0OsoDNDsQXa471g1EaRhPBwRTz9nQCqzDUxd46EZ0OofrqK5GGXR
00R47wWjSol0Q4/wDU9IRJQsdldhyZdV2LRvZATR4xIcisLb0rynYlf7sYYWthuK
XrjQGFQwPpcvy4auv/yrM3htnblAVRWbNvPYSbP5jGtpppJsWChcX3KGSmFsK5xk
dpfTjXymACg87NBhwiNEX7FrkayQbEF0TWNSTM3RT9jrfpspkON8IogfrITcNaAj
j3Kp1HRdo00gVVpX1W/1xDacE6RWNe9OhlborHJu7Z4+VIgVB4hW0JISsKHnyx2H
kvq+pDOurIgjS+akjAGDd9OMVAJm75slVJqXnO2nROM79hUun5fveTTnGk6gO5o7
7BrkzTvSe6Qoz926qGf7SjWGbDOEs1shB0HodyuqJsag8nrlzfhygYTu4jENHCZx
rabA/tD2WdsYI+tAgoZHEi5affPLMVTaclE/p/EOhz3vb9e7nAQlrHL51sz+v8PB
kjCXVqHQYdsvDRr5dyXNYOpexFFyW3ncQRwCZvgnP+v1wGoFo81OZL+yrKsTFXTm
FdLUF9rgpHQqTXo4Rc56Kjvb4E+1Ez6dO61lHKshb9fh7WDRFWtfJIvCKuMMPIjo
882xHpzYV3UqEZ0Ew5EcP6CwPEFghohUXF2xdA/GYhTSwSkhNgUf4AwuXaVZWDWo
YL4OIB0iBBjLTIat5zSGj0gMKxvYmnbPitWY7Upjr73sUhO35WCmf5Oqilx7wc7I
Cexmb+3Pxjcyq//PjyB7UPGq/BpsS9d970qUvbO78z/Q2xRkKwnN0YdGRfG9NbIM
CeI1uaNDM8HwgZzux38/iIyjoaBGeGu5HtyIuD88e+r2vwfp2sKkl8DlZTFRDySR
rPlh/0uS7JMVCmXzIue6o8nF3YJ1GLzGfrBNqlPI583FQr0/1oG9zAOvsma0fd+f
IOFneDmBvH9edHKK6pZDY5pSB4UkzUpWfiLRYH+LKQW/818WQbHH8Lm9lQLtcKSF
LSOZgCasLrQGJ45Lopi+9eZuIKTWP729eQs4OG53u0im2m9mdk+mIpoWAQyVACLp
v4+IktuE6UNZNjgre9F9wReWFhgNqp5kckKYbBtwoO9IarecoivkjxvwuOFnVJAV
YLqCnFdtZL3b9E33riS7VibZSlzHKR5tovijUoYGHc8LroFDeyFZcni9vTdgie6v
OIkMOunIkDJzszIHF7W0lrvQ4l9mAKhkVdCLIqX2DfL6KIco914R7fUVy5bB6xa2
qyOe85IxZE0N7CMLWMAJOyhtMeY5DyddKzcltCJHMAiMEQiZHeCoi9guM/b+wrlu
s99yxpFnbk8s4N9JlI1LQWlGRbA2gyLnDhCuuMdKFQGflgc3leFOUDINbRC9GgUq
p1rFUWXELuPKtkGeZRgKpqKTVmE+YBvyrWZ+ffuZkD5K9faKaN3QOVyS2FjRahow
A2o06kM8c8MqmkysrS1uujHENR8cs2y1mGHP5zNj8I46b3PH/Jz3IPD2iiWcpcOl
PYLKa4GBM1ghzqK7dGBiwnCgMIGASIPWPyJUBnyOwkCAGPf3r/GIZWqlwJNQ+B1u
YuCiO2Hl08BOhdbS0Wg7CHJrcjlsx00jddq3l7Wqqs3Z6YjWoVHZEtxrc+/AMiiq
ZdxlXBgpmvanRx7gXO98GSLLb24hfg1PdHrGHHSyopQcY04398KB2/xzuqlYoag4
`protect end_protected