`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
ddtXksX2+yylW5zu6QL2Lhnb2d1sD00763mmSITNX595NcHTEkwn0zB1Dry37fOW
FufOhVzEJp80NC5qZ/+F0Vk7Ik02dIR0elf3clrjeJRK85K4e3Hoo4xn7YbFUIms
l/8VZSb14+JVGURjfswrIyCUotIzlzVYZ6gzoZwDXIi5gQIBf/gI+KxNXPaKV+PQ
Ufys/12rjO6aI/pPlqSm0hCvftmBcnezN2hk1UeXgOIuKZnogjOsf0iJVX2aOOWE
6pD/psybjbnsNB6kH5uFTA5frkzIzkzl5d9+YDm9OyC+k84E83I/7/j+rk4L2dah
QJOvksSIzN867/4Qt8qYTQ==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="MvBXkzurAa5VTw+1JJ70nePUfoQXBvZOku/SMmg4TwQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
oRtzZL4VJ4iwysPsC8SXYCzXS8Fw2gtZTOskLcDV+1B9Nzn1zTyNtlo6lNICRmmK
ZRVu2BmCc2G+fmzynYlNTnSa7C0Cuel6FYpxCBlOuk3OF2tzAmLAuDyOH3Z1Yjzk
a0aHuoCdIRKv7BrZCdALt03JeUmXKPdOmIlkVGFl8yw=
`protect rights_digest_method = "sha256"
`protect end_toolblock="Jn9CQpRhJt4rnzZPRk+dOpzAubz7omckX1MrFd4p81o="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 11456 )
`protect data_block
gD6l00tciPUa6pDNTk/+t0OO0nC/UTtBwLB41d4inuAUA3i/ALrNyoJVcBnAmEQW
ptbcNp5fxEUJjnOxnedyZEuEBxWRieZFQnkRdF269oOMJeL3B2AVvPhknnkKxpY4
DOJ1gLYgVRZPdSsuUIhPN8UEdeUmqmdDovuJP16+qt7/w2qrfiTfSuDGYPGW82zh
3J4SabL2+4ePDzDTMUyqx5dkJEoW1jOqj2QqsNuxnEmtsApaD/odQLOD1U11Lw+q
tqo23mJS5ldvAWMuax8sYOzEqnsW6oW7fa8ZmVyJ3at5ZL+QgLp8H3vgJnuqScGB
rGg4VN8O2ybGYJRAjogUtf02q9wBMcTlVF4XLiajaN25lCis6C0js2wtvUMH1Ln6
tFUxEdlzf7jQstgz+x0SfuZuDuJwQKcQm97DnMlZCbMGzAwikRsyMg3tJNPmnHcA
azSNNGewMRHh6yK9FFAWQz96929C38L7k6LWh4tbK+XGDvh5UdOtpifUkb9igGaJ
n8sEVyqcrPvKH9hNtfN7FVMSv4VYVV6mY5dT3JCBeGGgx26F39SLgvkYuIWPPub8
eqnOrPDKxYcmLL89Uq/mVuAXKqpOmuVUP6uA9k+1a0fVHnOBBnjZj1QrRkuE7V1s
AjfoSdSinZs77VXLUiq8SjchMW4JCtdVP5+Cv+giZRfKXbw/xjl7JCBWe07EmWRF
pg4vMnLzjPMVsakF3YPwXyct+iCLf3fYyfd42NBEZkntxwL1i9v+Dw1mqv275gD0
8QMJkmHPRl+YzpmHLk8x9lGx/3Dg+dAmbJdNSoiXb8fd7ESxsOOGnWtDxCvhbAPM
Ye9lDUo+W2J5Yt4qRO1PjYklMm9h9b6z2s11o7U0QDNEbh8QeK9YaaS27MBAO8CF
zShRIizGYemIz9A9We/hAq9spyrbXu3BI2S3aiQodV4sDLy3jTOFlN18exHREmZF
o1jQJACXmDNGZvNk7Spn9TjchZrnsS3JiE4m2NBmdGMqLYjGdzGs/I2P4togpl31
9a77HqLU8ER0IBBqrkXsvBI6zg/oHBYSWa+1HFvbAo8ePlmh8NpwygEV5t1vZ2CT
3nMQr6B2mATMyDQ7Qv+ZmlxMBaFJZfH/XDgqtnwLGc6X30oM72nu7vVVBeNVZVY5
99q94p9GFfDjhv4jeEvng5uEAi70aEh9a093Y4w2UzdfTuCI91pZidH623ELJB8Q
OxZCb/iOueHKOQ0aDR3hFJP249Q+6oZQWhLzTm5TfAnnyDjILLQn52ki+8xfLtp1
bbEFhFNKiXWpuLHwOzRsOmQW0Rg27lNtnLLyJsTYI1EH2dm3eDNjB9dgBbG7oicY
Sf/3uKTtEwzfJ3Ky9+aZFsLfyspp19+aX7wdWP0BCV+O3vRByQg5ROzZtcjTcrxG
jVwMfgxo/nabMjNTxEVKYBqMxFottWqUUtmh5bSQ4q/IzpAl6g3uUXeN+536DY/Q
5cR+ehYIcbXFVqbmOjqxFrbWetJ97wRkgXHA3pe7ZgcRK8rv6rRwADaDaOV6duIg
ZEx7C3VJvXQVuWoj8DC48BvmBnKbnLNRs6HxtS+UgskEj5sStbuw3nfERc1Mq14C
fynvk1mHAmFzdrPrdacFPtkHlptVteWGJBl6w3EzTc0jq/p6DuZLMSUagPKFTEts
XHQv2kc5DfqwP5sBMwQV4hW51pZ8A14eR2VJkL8WKc01+PfE6/0rDRDTvqwf+bjq
az7vYkBRyjqOw0SRUL+h0CxSsOQ6ccWUCerzyyKZDYY8wq8BHlg8L+F5AYlNOy//
oOEzZInRFAEH632jAFOQwFslsjDGysS0lRT1R+l5scQ2SYKMXMhBXPdairiN2Y36
dv/6p52SE9Zoi1OBBnMd+FP8VCJokEMcKIqpbGJdS3cUVIO7v+MoXp+dmT0pKguX
dPwhoUEja1TRFeNUEHv8B9cRyxicfxUJtLplEzVpW44GGv7FJPIRzL55A+iLigi5
xvirnzIHJyTb1KH1rYHr/jiqPNkwgceOMxL/4MDgDiVKMqlpZH5cbDQXnCwwWZuF
mYII3dakgtXiNP9GXL8tMe7iUrjlFow8t4Hv8E8+gARD87cpDrCHjKhh8xORCmjc
ZI+WQAFz2KFCYSJTPBjgrmR2tAwy/fWzPxmfpnbqQESV2uICuK7H8VNUziK/gmLa
Zo+lnOMn9WztSDQT4MA6Hm3Eb5vWs34kAy461hs4v+oQC/piOmjx5XExRCwHSr2h
ILpCQNT11SP2xDB1pF392mlRoiU0Rc69c3DpEiVGKGAlafmhwqb0z+kWQVdkZkMc
DZLkc7VMUJL3wiowr0hp9b42nIXPPrBIy3a0/WDtwbXCdm0q/7q1Xl3nU/X601FT
F0QWR97ZppdboA34wBHbGamKhcLeofJJEzT+D3KnwMtygM3K6+dHUpVNNEDa6umn
SnhhmU3ibyBtTHTg5L8OkAy0ZQRFpCc4pvbbqYw8/yS+FbB7pY+WWhvGORjASXSJ
oi605YglkMAKITbO3DUQvaO95R9NV0nXmYBBFqRDy3uQWKDsDINWZ4jT6gPTrehS
qJrY5xFw2x0n9Cip66rVkSU+lrTzusNpw1VbTajCGgleFoxMaij2VLrCt+pL8E3g
WT1GC7pial6wE5NMGSh1uwIafnrEMXqK1mnznwF9a8VX36bnpzLN0dWHIGEW/RkD
2rCh8Z0K7knpAJCz8p4rgNuMDI9U4IclvHzixwN+ls0otO1DyhkN5xEZqJsEveGO
VK9/X71JrZc7w1TYoOtV/wJ1W3bsx7lsb4/mVYrZtyXBpRpoAUBAdMaAb5wfggEZ
rPwB8dISkMNf5Sc7SQccRZE02oG2mxtPBIvrGUzugfBPOusTu8KptgR9iEzN7Bsr
jGdmd/L/WMb+Lm35GLtHpUD3QTkQGisLFGZhCyyv9lmIJXM42GBAnMljDsJS2y1r
IUnbvaG2leXKjCMovQqx6/9dDM+oHhuNxxg4kSy7NQoCBc91Q2yXspCBSAZCcROB
72ReSoJruzoDgolcUeErwqlfOr+Z7vFWT1hvSFKfSlt+kvwmEZpL1NB4RzKQtYrI
Uye2/yApwfPF3p5tngNMEFZPRkGj9QEsqvfV1ghFq4o6j8/asLAUpKXnb+FB56ly
snsnG6Adt8ajk7lifiPSZDMj5TGTvRoWTs4Q3wpUusbvfPw8lTOQQfRnBymEAyIf
dbks9i7d/SWMjNOLmaP22Ex/dZ2T3ZjQQjIg8nVm6nRL2omwfKSJ9y4acPvnwl2K
NR7Srdk5qw2JEYL/OW6t1qBYtgpXoPoDPypQTUAt37DcBCNN/KWrHH/vSUirDHEo
5XVOxxtIRLbNLFEmY0RsuzQ8A+4ns4YzHUCUmnqoXZ+20up61+pMI5H06mDqXj08
npmrcEb/cIW7PHNT8zv/9ZnCyy/NnBnbuj5PGvLiWo39FmI5Z15Ta6cBXV2xmuqo
erI0jvbVvIltcDE2EwfmBrh9KaNs9lo5OP1P7qrt5OIKRn9rTEUgqUFHjx92b9Mz
VOqlDi7dPFCyr5eSWlQfv98Zjku/VXCCyZ5uBH4Yypvv2Xb3+8h3kMjp+WHaWIl4
wRkDIkoumkabph+bGvOn6JqNCACgxhiGYtD5E5LbLW6/yrMkqbvGRqQ4eEM2IpWS
LuWJxZo7i8h6GZ2L7Rzr3GpWrJVj4D59G0yFRpVwGG2OQOy+j+9M3Jlu1EFcKM9p
wn2B1Wo2wVcf/tvgmrP4YEIR766DoshXU1vs4BT1TaelJkFMOWp3JUANx19qxz/C
Y2j5pS38QOmWCHv01PB7uplxURuME35uVPNlK/sHZj/tvNsJ8ZY4my+bZ6DTNTUn
v369LCWSezyyw/3922kZz7xSNz7PXu/vwJI2Mj3DLLzl4q4yAN27fMlX/HvO9lI5
aUGBQw9nZA1NXq2WXLnGMUXOyJfK82c52KdZMvOc0B7+GNMeaz0BisgZ7v8Eaqn0
58K42aOQf6uPEc9OD6J81prrt7adEN7r5qDZlIt4vMeSpQLtsIjVLMSh/K5K0BfY
WeP3pJ57ArbUzb4WugYaTNC0aOkV6GNYXUtPXrVJGtdiiafQwUhM0r4FYTBx721E
kCFWqXht8nFVOkBKG+AAQMlFYCXFqjpoVcV4oOnl1Y0er2AzLAuOWSoXCCTBM8Xi
SeSQ/dt7YH+sgaS7HdhK+0687cuW6GUJDp8/2FZ0bthHDIfKDt5JsLiPrpn2WJJg
92/nitojG1Ac0Uh7AKKYsooN/m/IDI8eDS4zxtdy9b/8RN2+y7UMhapfXhF2jnOr
+SZLkxT93+38EFYE8uOaM9fs7BsUhmeZtZ18tjRqfmYU0JogWAPvdB/icfHwEKgq
hfnPkiRUfXmRbUJwtUcAwqBGO8zmTfRVghF0yeg0BNEIap6UHXUEghlYFgVqbDpV
Apk5xoeCufOYcrZOx3da3zT6MGybocpJWDdZbe+Sv9G7Wqg33hFiF8SHs/AsW/iI
hJl6fvrM3DJf0/toiB4Jv/BWlFztTQeUh1y3vlJ2dElh5jzxm2lQubKmqvZEPDdV
awf5a7B8RbPg+Oa8c0nCimt6vZLs2cKuYOkWy593n9lMtDCbYir+pGIbTpPYwzWD
zPsooOHa3iksZD7DrgxYjHTDnnvxlU1OZSRM66iuz5l9pnhyDruq7FkdredMzBKO
CeYRR+/hCU87/OvXoyGyq6SWDxsDC2Svg6Nlckjrcw0xq1XsoLqg5PKqScERgQoW
JnV3WKD4VAa8gPWqPxIT9PUPPuIAGCeqbqW9RmGTwd0WVgKf4sITha7HQpK6H2jD
TZh4OfIo9aM47VCFL3wrpVemx4/tmxnzVzsL3lDLdAn7lB5NwQVvjte+5im/rcYD
BBzsCDQ3SNtJTxlf2gKtDHe+WcAUmG8D5ajRUGQJzo8BfrMCYv6edINVLa9Ftvdw
bDZPiDDJj/ktp+45PjlgWI0U1Or3+8l8EKSMge6PE8419117rxnJxDMU8Ta9YE8y
PeJC5PrcuCvvrPEUyjWkuobsuKSjhJAJHTUsSmfWEEpYyeO79Hl5Gt1UnGuiSBEZ
/OpiswNNKWp7YARP3KVOPXehbx3/NGHb7kTJLAR2tmM2K1Vf/c0Lm4XGh/IJW8B9
gBLMgcLNbvSk8hdxBcElNvaya3Peye1+evABPi/ptg9KacnyS+xmS28J+7LaKIgm
8uzTwOCHGJ0NPnWnzaWfWUWs6wVj6Urv8azgGQXbldGGCzyS9ktJgiCrn6mQbofv
s/H8pR1NQmUsG5IaMe1jn1pCQJAAOjIYBSoKWp6/2lkzEw8a2K1PbS9ns5WuKo6F
I/kI4N6usrNTd2aSjkGcC8Dg4jHt+PYaO8Eq/xdD4NiBXn3xM3j3uclPjExxHFY5
0hG/SQd8GuyjFTeSEGFSMTBc3kg+z2pBUuVnck7r2A79l5yIgpRwB9YNCMfPm6bw
XVJ5ki0mfkA3pZz++UolHEDaJV9Stfu9iNbDkMXydJ9Tjg9gnJoTprSlr4Yi02QH
iXCxQ+bJC3ayUexGfCpAt05qrp8BKk5+yAcAadmCr7tRJ05LGw2LlVfUkqCij7ly
P8Cn6ySl1O/s/b4REIAorG8SNpU2qYNyiQaX2eT8JQggmunCMT7vAiYD+85S8XQ/
mIAi+3G80cZcAEc/+EctU7L+ecCcyKQFDJoXZjXAvADt8cWnSaPBTm2+HOR8riIT
XHNlkpAsUPn3pAn+nLnxTEb2ZxLYiBDiOrF+z82+5ClS9C77jJoWI1NRI0RMISfW
DnYfiOYW0+j67sXPQAcQXWOiVOKGquVX7plWQ4d7fnsvwHGosTsxRWVu07NV2WEw
Pd+oRki8bTboCJ0GDTk+tViZvq6pJc/p28n6LJaO85VN/ujtaTeqi7Ir6zFNdEiL
dDhHMej96qPsHocURsDO3zBimSqBLZyrRpAjKLpGoY6XE5P4t0r+OYWZDqlRkPec
Ktv++ZFi6awzrcD0F4bbAEWRtvDbCygzIi1fXHojLAsA53c5GABGLrk6Aq6CPcUy
9atYDNfY57QiKbr2e3+QkpAlYT7Bs0Xhd4X1geWY4sqNX3geK3n+26mccVNXN7C9
7MExpYQER9N7fkXwKXRgdw3Wa6LlBYTrGlEoPmGFDQdmOq2FW4sGtasJBd3HiWVJ
YLwRaVtfxKzoIvlZ3dJIeE8r2g8vddz6dLZVeF2FXRuyEFpr6P6wZy8NZk2mfA8K
tOFCCgt3dGa80ejxJabKpxA7mnz/414L/uPBNErtD/kSvoyvzaE9OTffd3Of4rUy
xCspXwbpzZvZ0oac19Hm+aSBaDYTsDFpCBttQm1/KGJD0Uu9ToVf7WZHEgP8LOfR
gZAxrwZSxcnHV6JtArlc2aXBqv6/11tTv2jD5z4yVenQIB9Q4RvN/3jDlYPZPX9n
mty+h8j49grMKe1Jv7svULJdgCnwXRJeCB8ydues37b7AyH09OvQW4hachHIeQ4l
CmduZ/MjjPZzPla7LmpM5S5OsIeVR6L2aeR4liTfm9QeM3j973PendxDnZEgL2Cq
uOmeZafZLTNpvKO5PjuZ0WUv3RQ1XvTOpS9zVnMEQaoqx605WG1PXHY4JOV7826D
lCrnlwfpWFzQaP5zkzVkzsJWgdEu39ictaUDCmO9Q5Ewfn9kb4d7pMUMHQP8Twr/
THRFGfC1LK449+7AatpUzrXVHEdYhVAN5G2L4Jqa401Xr6j5moynP+7N3aLzb39r
zZYo/J79CNoI3HH5mq+ZZ9erNPRUHiTerv/7uEQLBze/4e3IlxQq8GJDyOGVhqfD
2k5Ix3qQKeNRoyBhHFaA5f5LnVlHI64QCjS2pTp4jCxRj2WGMwE2JRMBB7KMV0sP
G/7XBxOOD3goQRfK1/hNvOXp87Y/O+N/Y+lsq6xJnm6XA/rZWwq0LG/baSoRXq4A
W5NskGrNx8gFvijp1BenAH8TgYMYcuN6iVfllOvYXgAwuMU3+SpB1mGm1/myyGtx
pvE24oPgVgKzEl5H9d/VQTo2iFSu+Bj6PxtDzTg5DLjq7ucbc8q3gTIP/dh2nqpp
qxk70PYgJKz5/GJ2NCiXslT0kzusz40rSLgS2dI1u8gcPb0tMbtM+cnjbXM8sLzk
9g8VoNiwHHYPXk75SL5MuIqca1uSY2Wf9Oc6xXHkURhAzxJVL3tXeuzOwRlmqShI
a973GBaSdlX1hMuV0cbrT73p7euc+P1XeUksDD3fS/ekTaiJueC6DKHdPAkJ5M3g
9NDpyTaOFsQu0PFRihqvAOYEn1T4WZSaLcQF/nuDjliMcroT+qdiqLai+IuxrQBK
cVg6qK1xJ/AfqbeVXMffKNkmWensQWlieB8oO1ka3f2EwMvR0HPVAZdZqCrKHDf/
lxJ/l0eU5t0j7NFH8T8y9UDLVvMuSPqhys2h2vo4mgxypMBGA9Xn0O5J9FhGm4eD
fz4/nQEDN837qsu3u1PzVGQMAzvQfn/m0Ec+bAlcrFWZKqic+PRWt+2n83eD2lm/
IkbBFOO4Ier5G10WNhnhHx5QRaGT2DLZqwQ5m3nsNpUwsZN6MuKoM2cPvO88izxu
Gdb3KdOtctz6qquuxKoefHgLHajsHOu/DDeKsDwrniBrvBel5agsL9ftLDVgnhsF
SHGWDD6ymqloyhqpXSZ42v1dtGyskJeQoPePhRr8PR4EhrbVaanQk3fbWErqLS+/
LLO+CJLOWIfk6ebiqdiCajXcWxVb+gZdZPZR6s0PzzCnDzBO/ibdFxBc6KmlHuPS
+blgRsDhWUdiHr3hzuPFLqusUGJjXZld1Run2B4zFLfZ63SNzITK1rlvlQ2v7a1t
aTaTZn7szfRunflQJtRRB4ndxpTHP0I/MGsU90Cs8DiT6ZRw9iGMyk+6U3wSCm+S
7yr2lkLWy/FMSZlTOjBqLfBY9+x7lRBCVEdio7lSK3Y4ETsfvc+FAZYEJW+EEeyV
evt7eaDfnDMTdb9V3GoFUuL7Axu9imKJ3DVTGJR3uCgPYp5Ha6GelmZFZqoaSuN7
lj1PQyBwlbOCXFZej1gU8ueyCTCXD4Zsn0Lf7cG/F80FKhgX+wsj2cDCCCa7nN9d
P6TEsQWfXcESwbc3gK0Z3gAbUl+ZQ+BCHSAvb9kVHwlWntv9Kmqk4igw80DeDEoz
aQutcafM82acjcD1qLnP9T391MBxUw5MFyBMxabwzoH+rqbgBqT0jROyPK1PtuUg
rPCxU1VWKSpyhMCNfQyQHyuchojjgXjx06hFMakRQzN6auRgONi+5LNeEVWM2EIk
cddIeZQnO2dCzjgDKO9EC0tOqQj3QPy2Q/cB4uBlkS2mcaks2AGBxn28ba8J8U5U
nlAKz8leH6VfVHfcLuuI/f/a5XlKuC5PWYaQjLLg6NTNSEM4wQkPK2UeFq0cP/Yb
ZdM6rA0xK+NfD2OL4hpCyyMKKRwBpXjLCfArUa9gEk+f/BmuFf66OYC8HEHqYo3V
W9mmFSepTWoaICIUyJoARQHAkzbfUCwj0z+CJLYUORRRzi21Bi7leJf+15aHaJbs
rXrHt3ZYpYaTpKg5j5On5lKL7GTrMe2kW27RVbLZKhXnGPr239cKVL0HPsKsIFT9
vNMgO0ezlbacaYBZos80QVyxZhlqVrYdvLoROj+Dy+LQxS1Eamxpms8DqZsXLaDv
mosf0BQFoxedJWaDGQ+rPz2JnizL+qbfa0jIUBxEQKaGMiWDpuof2q7qhw04/inS
peZnY8pmHU0bGzHD1sxq4vvW2fgJd0UgBBglVUQjfHu3fnf+Heia67uteGgasUVR
osNHxUI2+ZPciBv81GFP0nTjr326m81tlxuhdT4N78LiMARg/JLlC9XuqfnsYOp+
DRTKGUDNvbZH7Ox+sh40DlGo6L9yB9ajWMWTB5G6j6sbn02CgBoQDYNbS49cJspX
2LvxNxQ2lS0uaNND0py2P+N1Icu/uKNfg8dl7fE+IHKzYqR4HqL8k7G8bS8NQdGc
HqcAJqZWG9uzHJvrP/JmjQGIV28if46ASdMxPDczp8G1jUiD8jdyVhY50ubLGaot
cLo7bo32iiseCuHodvEAyeWWdqv8mmZEaYVZGCzz87E+yy0CpSPwici0GPVc+PuR
Pch4dcfhp+r7Lhu9lkRiGpuxmuMDVvQsJXsiWLE18PYbc8uNHAKJjhP63MeHtVA3
Zv3Voie/we1loLTK2qKu4x4hMTLKg3KEk+VvPivhbsWM0IsZAq/uwy5jPOtrbKpz
b4ZqC/egdEnW3wOmuPj6LZrpS8ojACUypYtatE/Fz2wmwi59j8gyGdAA/iWj6EWy
aAT1CsruWUetHzahx6fMUjvLcxUl05k3OKSOZQPOLJCimaso1ek/Ty7PbxwCkC/v
8K/osjvd4zrFahaQLUHfE3dFSlTXgau/0oM1AUS3nSr+ZcXVmV+aidpKOwlMqf20
YhltAMEDGYGVoEG90BLWm6O+aMSNFJUCFb+kAsXzzNVGZD+esKm1Nbuw5RJkodpk
vTuvGA6YSbEZ0wwnwvDIhWr0NDeoEOEzu3+Adk6k6VqkzY9qW1dKxjPpx07UEmZF
e+p13/snBdpT35sKWJildMf02NtHhbK/FLO4MlrrBqT3DqIL7ZJYmKB2c15DZ6H/
T7/EkNVtuzLhtrvXlKBooeOla8x/TIp96hhwxU8CmL5ye322wY+RLZlUylDjcgFH
5WuBJtdblvr+tA1KIFtsDJTIeoAVEvBGErcS8G8uKMg1C+iMUGMdb5GNgTTpe80f
aOrLLHU131drMoUAuSCIeVQCbocMWSMefzvrlKSWLcuQyM5u7W3jIVb25H4q56yQ
fl1CW9jSY27K6tThCHw22S57k18ji6vTcmzk8EoOuIpFC/rTwqGvT3BOHGRPrNTT
xiUBvV4u789dVBVswv98yA/szV9e1JzgqzeIhyzRFyEF/NVHlCaNubTP/TozXuAV
TTO4S872Wpib5tbMgJ4o6rllm1VEQDQR1eQJ6sqArOU8hCHIoh6RN8zACx0TkvGO
gTz4C77irDMlgSIETSIAXsDWA1g8NvT2ZOFQiFyp6Ko+xfTZlhyZ1R/QFtzyh7MN
gfCCy4ABAt5VWVOz8ftwYO5xdgFu/pW6Nso5WbsEYXG0O2rxiXT/t4m/HWnNLBKx
/v5mnDztC3pvTd1aG3MQrt15wrMvdUR5SAmg9h/j9r8ct/N3xKwrHFzC1ZvYjYsD
PMV1yYJioRrN11d0WAGkpazLZEJF30vzlXdtq+C/ksQ3KLAVCiqtucbFFUgYUx3/
D1Npds2+D8AWUbirnrRKCbL6G9G/wxC5BSuZYqD79wgn6gtL9UOdfrn9Mz6HtvFG
g/7xJKPdTRrS/4Wl+8KZl+qeQ3y3znR1HCqX1qdVUEF84MIMyU+kt2wNa9ROpfId
Z4HVKv7lRag89eo9+RnnMlej+WqJz7QO8W6BmexmPLShHaqNd6/+7TnX82JJ4Kr+
CnvT6e8V1SQmIQyc2oLm9pzWo650/44tlhYPlzDgIa/GCHPviRUlc+o2DLKfk6aK
vwKtjOQb3EktBR+1LwHdVbfkjguXdlJmR6PpPKHYgT78VE482tjJF90DUX98BR0b
6aG9FamksEPOjGo3874B/whx9XWrCMJwnK+yL543Kqrv31Pj+k0lnytXLCvKpjUD
xUnu5Lz22JxCLPa/IHlo8O+tReTzKj7JlKSClwiYaZXIl3KTl/tmJpn2kgeZmntW
OJLpi5gWTdInrbb9RKJBOnOwR3b0Sd7rUa7R/PBS+kaYd27HAuSpTyFuEMViKSlI
uRHF2DsBnyWrwsU18uHRvLGNPSF9tPN2+OBAbB2x/aazEf9JB7qkNSQOFnKcr5PB
2lsd69fS1VUztNOePBQ38cl6xIWr5XTvmm1ciSM+0LQUiyqixzQZFxoaEYxByJku
6fE1VUN5tkukiZXR08mNkDvAN1tuzS1jR9E+VIBACZsccB+4JLzBjVUxBKeLG7ki
diIGSjbI1UzwJiu+jLKZWCq1j6OQAxizo8C3q0Vd3qmmy0BGkPfESr7+b4k+qM2M
d2RZhMOyjezZjJ+vG+CbRij1wZrFUZONFvPxRIux6LZjm2RZzWMwOhCaR5WwDind
QwW2f4SLvKgZOvzpdLzNOnxR0juZhpyG5M3rBHygFkmlxdGrpP0+bR8OBCJ8mhOH
K18ZQPkEcJ50RMp5fybk0RNWpjDRCObIdITm4ZA8g9WyuEtPTdTN8E+e4ZOkLUX5
vcXt06R8rjP/Bddaxo0q660/MNu3Fu2k0/VmbyYApv7gGt1MFkIABUHSde8KUazx
Z+/fG93tQ9kz3rge4qM16HVdjlZztlQX/XosVHCFNrC4UKvEkCGaeHGy3s4jGcxS
5uPjDEKNAKKVQ+CjjdAtN2vxcwbctpt///Po5glie6aSqRDQzCgVZJhu+5EXoCOy
vBxRIJuLKSEYZbk8MMnY0fnMBX1IQA/NAX0vWkjdXgTp5fcb3H/BHjr2nmSo+o/i
r1a2EjPtXcmBAAzmlYpJyL4DQdLapCepDxgW9eeHqlXFGTMvV+4YkXLf4iZPqXIs
6NyqPkq14FzPlrZpOI8O2mwhfOlWchkXCwH/bCTZo4RzIBZXlvz2v5cdgA9JOt87
c3P5HHRGk4zOYegvjctcNOyqLWE8Fl7QWTvoHk77gy5cSTP7nLWA50+8G9WxBizy
QC1ztVqLwFw5TBMyN5Yb0+EIg98SR6sqtla8x9CjMQWs3UzHTEw/RYxX0mfbly7V
KMLrQ17AOqi/6ZiVAtj/ZBGuGRcOXQ1WnRYScjyelX13mdBqlquDeXjIexi2FpjD
XIgXn22NqE/Ym5k4kMMEpISMPr9p2ILSRJ4eCmzlgCdc2FlYByuoLTkZU97Ta8vC
zW743f7DNVQsC3wjVzOotM9OSVmjqhZnAPnmr5Lq82RimaLEpurCul49a0jwYGh/
1ynEP4KYQMkhB9tnDFo2Wuzpcyd9JhgJl/4btl7IVuVKbOEtorvCVBx97N7xUnRq
zm6n8C3/cT5S041080p9gbld9yGpjzqQSdV9U/tLx6CPVqzeVKow9rjgS1DF9ikl
1XFgkp5hVep+TZaUpnQeBWrxs/4+HPkzgUWNqkaS0ngYmVt3t/78GgHp/74Q9R0k
1qYRiJezMyI5jTjCl2PLtY7aDjyMnEcISC923D56xfiJSpblYdwiP+bgITxnumuU
OuiNse8zBiWaKNyI0/KgNwd3VswJEi7Quz4fz1xDaKIKRxTeSoWCgumJFdb2tvu2
XPBqCyvg6M9GqqReMMPr4jEqjQEFAXRi2HUDPoTpI6CsU83975CRznjus8nhkCaG
6xRLLaYcszaojQqjUuqalukZoDeDd3mS6wgDe/g6un4mOXRIFiBJtHbR5B8y7wp6
/nvrF0vUqcMghdbzGYsHRYN8wjXV1GTcluv6lDAYmXbHot/uxArmFCDChP89I80k
ckVzk36Qx2nVmXxjDJa7uph6pUjiGsc0xhL+JWLgnCKvZ2UcD+14sQ/6/idLGzGq
DAYdtMDX7DV4hgjUqGKLx/pOi+yXHzac3cx4qAhuBv7SaqaskYsx1DU0jm/4Zp6I
z82jaHwahrS0g89iGt3W6tm+8gYbjCDvIQO7QUoVNoNWGEP6+PuPjKTc9z7x+z7b
JxWPR92vwLAPSJQI8yrixDdaFWnWVYHPe7MLsYw99WKBSXiyUCgrS2UOEv1QE0A8
pmGTtKZF+LxxXo1Q3jsuqQ+uIjeT5lWIlttocmRHg3eIZqRoDLCK6ZQCvnvo96Bz
X+xOqNMkKZdIVnqSd6GcM0SorSVT3srVFuclSW95zuuNbNsG+zf4MuSpqegzb95P
Bn53ljxDAd5TWIqU0/P1bCoXB+w/Fm9/5lmY5Za6f8Szrthm+0gL/Ivcco7vxxOZ
+vCirDVg0sQIFIDxtRFZKaWFuQKjl31MFLkmbIaTcnqXGwD9qfn1eQblEHHlX2AJ
CLBqULBzx+RqCb8un6uyq+QMraXdAUa+vkQJEn3+vepVThK0GBroTJ03osQEKFYm
DVEkTgiszkUDk5TRou20h7r9dgwQE3e8lCtdXJqrqi29v9KgYTfbYHIQTDhvncmp
1vGLyACn/vl3tlUYZKo3ut7bb4IvfGES4SAKKxwDV56mUkbN8a2dczgdVTKK8MNz
QY7SsPjDrTWf94GhhV3SK/1o91znt0H/U1VnQXhXerZgzXmeRE7SM5wVXejpjBQ2
Cw+3jocV19NQizQa4rZXJRkDX4K3rgUklc02PNK/BZbXeJysoe2aNPgwu9zIu1bG
VRVILgvE1AMD+nro8vGZ/Yz3eQ8onOdihC1FQS9cdCTWGJTa6BmjNtjZ7UIefL8j
tgDBqMOIQqzrm6JNtDqv++Rh7kon//rc34PUwf0iO5b5mV9xrTqCLcNEPt7ZHeyh
CgAOOq1RSZsRfcvUJUcqbUyjZUzVXLfqXtDMWGXwpsoxSO1ptbkctYs8yyOzZ7Eh
GWS0Xxsc9Xv6evBnQOfAuv/ct5pN90y+iYz6m7CPoCLYvmq54EAmgtMnmsKXRF+m
hf5niki/7XP49mwmYmOfd9DnQFasWdwELF3ulwIZ6Zx/sPa0mF/9zUEooBX0qDQ3
uDck6NtL8O0wVxO0njAqjy+vOpY18xlzgD8cnY7wRnaqwZAZ26Y2wAA31diPNSBq
7q/s3BFqCDiSPU8SviSkspftzpZEdF3mfnsAjvIS4CN8P2PkxHdSKhLue/YPRWKh
GaMvCnVJ9gjRhnDTQjpTXmKvoi4vKOEXUvclBlDi112610CCQpgs93JfYMs4oo1v
eddbBt0N7tOmmkMtMj5qUp4W78yQJ3UICCYdaaAF/bj224vQgg30zbrveBdn1Ebc
NimqJ2jCliEbjGyXo839yru2+sDKdsbajF5dQXqNQTtM4RUlW+lI6EpoiFJ51QWr
gfzF92AqOXtXRTul6w6qrN5TRebP0w6zGKLQ5M+o3gS8OisDRLOeRw9sWcUi/7hs
L/apRSczcw8FN/0DEyippN5iHghr/lfQ3tomQKv+xuL8isFQtYdrfaYXJOu6YFQN
wguC8mBnAQtPM5lLaKoUoVNyaNyMb8y0n/h9vdLcQn5Xoa5eTxfMqS0vRKlaIDkj
NLPPTJI39anFdnr/epv5I499Mz+pFljfZk2huwHnUnT7V8YeVwp0t3/cXH0uJ526
Rp1YaE4h1VW8wKnmCT5kJFbAsClFlo+4WWv0osYW4G1ohCm8cgOFP4ZXg5YoZ/CL
qcTYEwp3NxwjvH2VXNSHCqf1ZBmz+vWVyIw3DPRPsMGKuc7zyy3T6gE8Cg2OkDts
l2N3xbjqCyAOyGXr8UE3CneceiwOVCzXLEaVsK0gPGnPVqE8xPE6y2MQ8gaP/2mZ
Ux2qz4Bs3bggzkTsxyC+kLYQUvbqVZJimezRqzm9Ct9/yM0hv22JW9foO76EAabz
jPfhSn/A3xo9MYoExO/KuSRe+UK48lLT4QLq9wK9mEi3ABQMoborBnZsqnIJtQ4g
kEpctx6f6VFKcQt6ZNlSSiNbV8LU1V9qn9UdNiYkMqBJKbXOFlhF20HH5CP3ODo5
AKmEgRgVITYUWdMd02K7ql/KH008tQ9nsZrwULznIPbhw35x+36M2q7UggmbvEHF
/tHJ7idyzZwuqiplTS3WCr4YMsStQfp440mhcqMClx44AfdKtqDwj23ocdunNSxQ
sINkxw9+4bzumFInNn4tk0xoISx0DOtV9uqUW3Ge3KVWR3MciAWaYJGbi1RzpYJi
d5NG4sK0W09I8WECgUUiz4iqo8DORT2zSP2IIcW15CSQVQUQCWqcJrnDaPUeGliQ
hTyi9GE5XV76ZObhzSRrTZuvialQXhUf6suJstmWnlOLaD8YGza8nB6UJCjE4F8D
6a6sLI7AEdWiBn7w+t2+92AY3IyjKJcTN3CMvWrHS99nRdqAKDY6XxBrH3LiF8Ha
cIWN+/ZZ3m6P3MCmDsy92tHFmp4AOzexPBhdHtkOaxAiaKgL29NB4lWM2kJggp38
2eEuy+xds1oFta2RypbWwbxTgQ1BskUDuZ0SztNIbNe5b1uA9G73NuagAr9LhzF/
AvigIpNTk1+F+/HAShQr8Pa/reYeyr9YlzJAo/0taFQ5abRorMDxjPx2jLvFAln9
VfA4VEfnMgVVRtvU4yEN/6hBs0i/LeTExtf+ORGwhDr0ZsJ9S4JV94x5PPv7/KmX
QVfzStNxpwcQV52IeeaYnO7duNHWJAGSQ2WdrmrKiMkUWGpH9hQWomwD0ksoTlJT
sAdTm2vmuVHdvdhMYdL7MlBGfr+nR7chXlBH28z29CY=
`protect end_protected