`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
ddtXksX2+yylW5zu6QL2Lhnb2d1sD00763mmSITNX595NcHTEkwn0zB1Dry37fOW
FufOhVzEJp80NC5qZ/+F0Vk7Ik02dIR0elf3clrjeJRK85K4e3Hoo4xn7YbFUIms
l/8VZSb14+JVGURjfswrIyCUotIzlzVYZ6gzoZwDXIi5gQIBf/gI+KxNXPaKV+PQ
Ufys/12rjO6aI/pPlqSm0hCvftmBcnezN2hk1UeXgOIuKZnogjOsf0iJVX2aOOWE
6pD/psybjbnsNB6kH5uFTA5frkzIzkzl5d9+YDm9OyC+k84E83I/7/j+rk4L2dah
QJOvksSIzN867/4Qt8qYTQ==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="MvBXkzurAa5VTw+1JJ70nePUfoQXBvZOku/SMmg4TwQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
oRtzZL4VJ4iwysPsC8SXYCzXS8Fw2gtZTOskLcDV+1B9Nzn1zTyNtlo6lNICRmmK
ZRVu2BmCc2G+fmzynYlNTnSa7C0Cuel6FYpxCBlOuk3OF2tzAmLAuDyOH3Z1Yjzk
a0aHuoCdIRKv7BrZCdALt03JeUmXKPdOmIlkVGFl8yw=
`protect rights_digest_method = "sha256"
`protect end_toolblock="Jn9CQpRhJt4rnzZPRk+dOpzAubz7omckX1MrFd4p81o="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 12064 )
`protect data_block
gD6l00tciPUa6pDNTk/+tzLxvdHE2s3DQL3/JqqujQBC/Ei+vcAB8wM3doqg5vTg
mdfn9XB1bLOis2CVSfu295W2DNwHfMSTc/8BhCDRnTlLIX0UCJs9Za0+LoM0rMrV
T7EjVWppbP+Em6PkVKCwlmIQ7JKaifJ+Y+kjw9HCGboYo5074hY+K/CBbfsBQY86
NbkSLCO87IQEY+0Q2aP6t3HaLEE316UVfxLWDIkUXZ3xXfjlJEi8rByLy++RZit6
HXeX0O+Px9CZZ3nB7waHW2uEkzFnnAGCxfnL0BOTvri0Kg9YIhMEBztHIZ/JKDks
vW/+D1DDVzTXvxqGEnjT0eZZ7nrjz/j7IaZYk+cOw/aejNM9X/7ieNYqKR+7cPcX
oegpIo1gFKX99fqiZsQFC3WRfWWt3CpJvNp2poPsG/trHtHLpXoM++4/0+HlXR6O
640AhY/sHyISaMPfDbXMTwYx/u8tmaD0zfPgg/394xPV06TTRT7IMsg/HvunLmOj
RMTECziCBZmeYVS+eenriPZ+1Tnwa0SJQcefHnXD6AivFvtGqUc8ahCKwrLC63Xl
rMDG84vKGvxDc9kgsyXnSxfNN3r1UlqacptxAgGjtyJLPiuvShlmci/mMMhVo5De
SmE/Ws22x3BiJZBkKr/TCUrA+tD8FAO/K1mWBLavDXT6xSBb4xQg6ZxlmwcsjfNY
xR8EZ7QsGjI7zUNPT0QJPB8BsFGUJ1RgrWhFzKU410lIJNiZoctno6KYKu/kXNG/
ZHZE4+pwYHr/ZO5fB16fEMv64mJmrmTAWghzZDZZ4S5G/uv7kXayPL+AhkDd44T1
3MDQRMs/o4+r5sV5vaDo8FTgJ8BGvrC7PFUD0dxm9CX8/8cF2jre5vZRH8XxkmO8
MhvaZbdZyXSwyzW4+UnH0nspMl6RnF2XgBrgXIe9Ff6ql4N4QSWvT1NnYYHAxAJ+
CKs5B/SC6ifcoHtl+xKpByUm67a7Zyp7r1T2jA9b/+8XHOmQEjP0UW+Voxbmceao
XdOmMgdPEIs+2IzjHYNACDCVadUA2Q3feJART59bSF7YCJrwBWl6A8z2yhczYNGv
Fu0xeFYap77+CfyzbdeI7p0WO/3VqrMV24/C3PCvwgKgSDAVH9habQIYNovf9zFm
r1JDfZQN+5hiZ3pUXJ/2tBwlaHtVteCZaqMN/xNcbcRt548xK0z1TZm0K4w8O0Br
Cjj93ZRQkGW+iXUjYiSIGHaXWXkiHlAwzBc42R5tDFhTRRpCSP5cnfS/UQUhHRyy
i6fchXtBxFOkHmlLoD/ckROnZ0lqiw1MJ6y3Is2jf5NDTIBRZgw4bzB8yXI85a/3
YuYv0iVr1d5o/skGhRHTkBx9BIy4fhIYAXHLCo5KAWEEfczgOAH1s/FoPex8k+8Y
+7vhfBI5r6iWHorqH2Toyp1sxwwQZHXgBkyuUt+ah4PyoAz1lY/ahc/75Wb2g7NI
E7TFjNLi9+pvqC0s/wxT9yRigD2QmDfmb6mwyrkpkJL0y7lBmO/u1LWQFPYKuNPS
EHcVKKzMMiN1y8s0NWvRXesIwkyVTb/UzZ7/zu1IdC0YYRRzXLP0FDaiB4BWIZYN
2UUdBbW18nMWW3g2AvWlooBZn4mhSHH0LRHGej/GtRjYAiKRTEikb171VuE1Cxmj
ZB4P4mM7UBNTvRhaBOae8Iv40W13TnBS1TFcgZSPiiLFgjC7dVSlTW5M8P7LCrck
U8yiR7m5NR9UfTYT4IcwIzDpbW+HKg3VR3+WXpPFlliuUdQaafNnq1+Du7Vsnup4
rYvUmmw2ZEAJ0VHbcDqsl896KA5xz6fR0x/H8nz54TtO/MHqEHKTFi8udMAjRPUI
nwwEwYARNnKp5gPmyVbGx2ZJ6skHNqmKwOuuCYvQ8/iIQUVUUJ5WomNKlqc25nA4
8mcP/I6G+IazsAqBfc5Yd8kjkOGo/fd5CHSw7ZeqCr8yNkzFNJKW0tvp8LsggSHA
77eMNhL4FKIFrQOOCyHqdULf7miuErdU+uG96Kc6kBI6Kccrttv+2QUNl0ZHOa6d
y28yAjx+73I5k29wifmLRrQotQFyS9/7PcqE22ybhEk2epCjzZsT2d1u4+TZM5vd
K6EX+mQKXyM1t3FbLX1yyapiDjTlTMDD7Yb1heFjzpidHloAcbxfUhA9P5YErrf/
cL3VJuL50Hdl9mg9CJkjOrVvJNnWthdvIXYAM90bU7gNXCMoqHUPmBm15ZbTYOG9
lmmHG94fvPYOJ0f9H0C6hTFwDWC0DHOcRrIwyjHgDAYofOO4VmsTA54+eFxm4HnV
bFd2JoxYO5CEUkX2R6womqd/4u+rL3Pc7Xx3DqS2OkS4g0b0lZlGvyWnIRVWQOnm
133udEqpXKTuc5xwgS7XAjnCbYndYFECRxChV6osB1OYMjza6B/5RZXJX9dJxOKb
vGizucgE/2Mw7Q/xAJ2xEBc/KDYWRISLTxSRx64jAbqRIcVoLek8oOnQN8YGV8JI
Bqa0obBHAIoOxLNQpTWSs0mM15kzX1TuQf6QLiSjJaH66lOh3F+8tk0xcZLOYUSb
Lv1X5EYJucK5qzEL3qFEa0+NNNAnLkZx/HAwllq86jldAnLP8OSXFDd6wu1sS+NH
Y37sdZMbGrsnA9NXGA52xt/HWMNINKbpg/jfx7huWkIhwSNbDcfjat0WYzpafNSA
g225imMaz9zUy70ZK2y0Th+sripRKrU/QUfOhVLuhm71ZkUMc0T8nr6+yRWCkkWC
4TYz7gua9yFONaiSqgQBhoo/P6FzhZizovGPvIy3fXZCHZNLfn9FrXhdsZbJSDAO
wdHejG91DDVj1WNAN8N6Cx7H0I1Vo0fLwteukY3xbfv4JqIWDKY3WRDar2SW8EMd
EAv/re59KfWP1857HLEvxGApKxbNwxkqWMxLDGcGUH0iCxPT1mBJt7aeSRNxSQgs
nQvDsqwOBj7ZPQ4KY2+LT6NQTSRS1M0r4qJn9IgATMRjr80McrclXTjyPtzv3Ub8
dtwBalL9875x3j7JuU1/ESND5+vbpgbERvLJFKKVNi+SHqxpWFLoo/fjwKk8AEqi
YsS3Ydn9nr5CuLo7ueuyQ5RR9lxDvB+k0dt8+uAs9ZRw7XCB0Yv2loL30ow9Fxpl
0lnFJ4qSzRdd6nCTsrC1Y2zCqBMJYlYzDXJupCoYSQaBh7ns2eAKxjrHSH4oNvo0
W8o1Ek+SkVArjVJJTKGBMwJ3Ld1w1siShez12qFqz3zdhMUGMOYSOeqfsWCX9QCo
B6heSwlGBWII08mLsL+fqRhPPGsWgaKPVU7ugMqCq6bKTPco2ozKDuFF+eq8IpeV
dCZLRFTZqB9YOkFa7scIK/S07SOi133V4OSAPjZcEv/DNdfFp3nEETFlEJhrY5VC
eumO5iGu5vWhBs6sGHN5Lmsn1bFIyj8ldg+41d4tJ0xk9zof2gywRfM2XnzvgWNe
BIFPi9NN3sVB/SNCeaYWZll4sCwuributcJiAAYyvgO6pfZXPqZh2vZpxqCMQk7B
HUdyZk13mMcRh6nx+zo21nLUQ+2dZ4VYOVddOWbb4J+uvvYXgt2y9x+VjbYgQCUZ
I3yryVw4i8jZ+aOR8NcqsVEb+EDbQf2OXOa77O5W2eo6tShZWEEEil4xHYPuhxDc
cPciUw31SUPRJjQb8/0a2QLt+i8+x2Pdhg1BPnlo0FqP6AMwjRntdAZF7SFAKVc2
P+6JHUjsF80fyrYopgnLQ2JDabRiEpHCS7i6tPEhuX93dMRUsmX7MMgLa/ypM+IU
PDe4kFiV/A23kKApgPl/miCWoegRx8LSfWtbmMIOtJMkkoJhJP3yRjGv4sl7CK1Y
Hba0aI8i/QejArZvHTECKtnNI5cX4ucll+QUHbNOaxl3GcebXwPTSm3O6aGO3RUA
dvhFdUl4whge7F6tjy7Mw48V1j5/Ff4dS64jUCuWhLweetWXGbCBIRnb96UFhEVD
btV4Vwawkt2IvHp/4qT0zv+sMZlnritHD2lUmbiirZfcQUQPITS/D6CMbH/ZoR53
JiaVzKE7pQmh1jGe6tbg5QPUEK8Uha86vkGJ+oeeivFLNjUlbCT+mzK7mIS9Vkgy
fqgWEQaOykvdZIDEpEWkwHi9Pl3sSFQAB+EH26tPdNDZb3lzc5n3fS8E626k4oh2
Cx/VcmaUix6ZZJHONIf6JEp5NFsRFRQDbyiRY8RC8NqcYbHUFNEYg5ZXnzliwWo3
7Z3l5HLm4oJws5C0TMfJh21pVMIklyUqJuy6SKCn4A6ckrI6MPWgTb5HwSx/jbwc
RIbaXO/9GJzjy4xTGt9N4BTXrLfDifhWdCrV0PJhD/VtHUGcVW+cc5DH6gwpcduR
SMGdKyZOcoILMvzlSth0UDpDbY2IBvDb3hInfgVvzJmK04WwM/PH6byR0V1gN9Gg
qYiBUjGV16XCYqN760ZQnuxyXda8IDv55BYurZniI+3uWTfrpiDw1QolSZXsS4SZ
Rv9VMPG/trNE0Y5THQeNe06NSlY5YIIMR6k2ByDlYCM1eDqY8VhSukKucPfcipWG
xdvFAnV98YncZuOl4WX0aLpmiXPxX0udu8UfW6Eoh6xntDCmOWA8gvkQ/a6/vR45
CY23R2Oxew0xJab1HvCTwRSdd/WJ1goxFfT9zreYvMXSBmuil7Mrj20JxSWK76fG
0VBCkbS/RjA7tkpeqFefsIuiT3R89bP/22cxzWnL2LGV7QbBtJgAo3HXvDhfs2z0
GGv/sJro3Jlx7aUVzMvQQvRq9bju4sPvTs4lVMsJ/YfZ3Xl2O2uOkumCPe+LDdJa
yR0kl62R8u99LbnAdirdIO1zKq786zv5C09Vrr9wndkMU80MQM72nj7Hu7v4tMJW
behTk3BSVASJUCsqwiJgt8QfEqLKeoRbzna78m1MKpI3xX4kNl3TbvyB46X0SotS
UvTMJTbUyxp7PMXI3matwbEHXMP9rjRT8jiaBJY5cofcXTDbfln4Ci9M8hGGrVO/
edcnad1ev4mBaeQg+Kg7rwdeXzYv+qKg+rm5QPQPA7TuEAh5TLrFhMadPNN6CpK1
/WlXZ/6d5394TkslgIsRtz5HmHmKpWrEXByD8+av039er+kNs6rJVR+IXu6igweG
Ue838o5H0A3Zc0cjXWrtG7vm6L7+FMRIpsfZ+MyRaFEOVc15yQadYxCiMhfHiJry
uxFu1QeDYwnlxfK5nBRYgNkPRPewFuIQEbWBcQlFMfq3a7pZJp0UjqBpJKRKeha/
RSXFXnAkDrM8al0Nz3TTC7LpKsmYtQSrR0iJKaBkyCwITWqJinS+3bK4mdGKL5MP
fpFtyDURXOMEFt62/gXwxtFjsuJgfSws+vwq1vp3wkuETkDaXnW27/JBAKNxO3rp
5htj9ENg3wh/9Dswsq67qMJ160V2AUTGsbQUdPko4jruMgXSllO9Y3wd4f7mcZq/
6KpXU6HuRGR3i8Cb42SXZUrqKiPCDfSlNX2Ghg9fAuufwy5g52YZZzJlOG/541Uq
pXP4dn7AJdH8IL/nN6KZ4iM417kaZ5JaMBByBtcQZJ+2nR3Y+5Xb3QzQB6MREB4A
VB3bogZQb7Xqw5QLHBqUZ+rgugifsAmc/K1RtQbG6s+l6nywFx/k+O3FigReWVVr
7LsYKnC3lSCjnGQjnFnUGMu/y336Aew/JbJFWEv3bQEXukkLrB/utb0ppXIgROVy
jWUnESDjqmRy7Bmyrs8WEgzl2kidp0rkU4i7b9uHn5S5sqcHZTa6pvrwDjTovWaR
VhgM2/ydFFpqIzVVZkkhTxVI9/D92TZxdXxqTQ+lVREOQr6Hg7rUOa+OKP7NnHnX
8wZxfC1rgkQca8jXElmOcoZ8b24ORHg/i3swhZj9Hay7uC0k1P4r8y3+hZ2I7Aln
MfAfE9T61tOuuZO7ot640f8yWn6aSMSXj6nrM1K0jbtOQYzR1tDV2YHaXELhRmAV
P8juPtgKm8mUVuXHg9knXLSF929Th4Cw657+zJ7TjRoBdzw8DSMlYJ31ds8WOzV+
B66BMYng6hS9RRaDhet0bUGgLVDt1unL1I2GHSBzfRbKfefmQW2M+X4gVJUU1Gfn
NHXH+E8mOoCtWyPFvcaOnbxiPpTPZU8XB8G+3B4y3K0SWU44n/3ULFnEuvGCIm1w
AKtdJEpyn1b/t3XNcusK24i/BuG9ZWD44nJvazdvuKn7tQO7WHcJBsY0RQNIEmZS
6KBmh+Ywec8OE+PpxBiBVgKjQmLTG09qCc3AzFTR10ta9ABfDSKMpVsTI3gYJgVL
VWNlVLLEpGn7sF8dmmpX9t1G/hBP1k80mkV9iXMlgYO0J5CVz7UgeVKuLGxRdwCt
IwQMxrH/7N2sfKjwIwDUzLJmO/0kd1IyGQ9Otv0+ocYmLNe6dYPJkEm2gHZv5z/A
BCGlB+eSNhkyUJEzwQDvLBknjNNCKHfCzgyzyCgpIftevOxeiiAimq3AMxW9eWSj
2H4hOfei8iI0vHh/K0NxpNXioNPJSo/NdXSthzihmOydq7FnM5oBA7H5ng8aLkEZ
fZ6GRYGrPXCFbfOEGhCM99HkGVsrAYGlPMrbcs7FjmV9GbxWVp2V6Eu4gAiAXamO
5WA3PBD7nSfLVDFdH0yv2OPl4Dy6SXRS77roUw4W0XKHaf7CPirEMbEjOBOKhQO6
ecFwIM/yMnsr8/fqW9WZq2Mz1wIPvZh6dpvQ707ZUIkvnFp9gBrfJvVdBgVWQRw4
Qe0aMB/Aa9EfB73jvvazZRk4yb5kokX6e+z/QS+kTwoY8ixDNcR1To6994M3hCPC
svwz+72sg4eR+wH0hj7OOUe2zd34O3muQHvif1RBRj0+BZBsXEuZgBkCc7W9DZ2S
M+E8FAQ6mgFUF8z4u3j7OwuaFRlWxksAZMfUoRG+p7iKXFNby1cnYRTNCUsgOwPn
W/ad+CvVEqKd93TuHfhT7/aAOWlxLVygw1N8zf1A3BiOeDYp1yOKVQCPAHfNohVR
8Q4M7tNRpur1lnmbQrj+jWnfbQT6T1sawep4BV6c2PR9lsR1L+TvIpJfg7GSoR8X
3HEEZIlfdXh6+k7LFIbl4YRmoCMDcudLq8SKn3A1EPfh6jtEG2OBLcZkPoKxPHUE
M8QGFDodTBo25KkfxMCkRdf4xQ+VN4vL3k5FuhUuhaTeM5YwmIdGjOeZZuEc1RVc
h4Bl/uTAIDMYvWppefEQ/vteWo+AIRrG/GHkvzhVkidpiyq+/zSlrptkm7wksP2A
8OF7/IRj08ItLc0nQxEcLkyYGc4ylUFfvKX4310U2V3JiuPMRpfIySz+Y7+rxsxe
pQI+GY2HdvM+Z/KBKfRduw1gTNa/s5WJQG+IEeXRUehs2JQ7i9PFzc7VWsqV9L0j
y6/ggvXR3KM0psfTZvmFkCj0ITgrJMj05T1gVho5BV2pL6mGqbPz/NLSwtFbdwH7
ZVTfgSkQGJWQuiVcr51WVfGujiBnTF9PMBX9MLrZsHv+w8BZuKZShuPUv78mcb9v
mAEWTlTIgf+4xMX11odPVoVXrnKrYqbq0SZ4NOjHMVkqkIfA2W/GbKKl2cVLTCF4
0BFiv4V9ygOWjhAXU6zrFavuQpLpwfZNe87rfqabmKOLt5hUHt1/OBj8BuM8CkB9
ova6K9Gv5r0E4rsrCCTCYtH8zz1q7DJ8lL5f94XRxdYzAmqqIiGfZPzvEDMFWevv
5tO4+0ijOrEQMwdE/aXHZh7C4pcUhZ8Xy00H0kQoKzhNVtPqxOr8LuZH5YKutlZ3
c40de7Z8LqUHoqYDv/dDhooQCo38JrAGxSQNYIqogfOI9/nnUpRZciv7XNTnX1W+
x4YOst/Tgj6HeHggnY7mSRjlAsa52ueS2XsnM/SLde5+mHAGCQ9yqEqmZjYay5k4
BsW0i37+GS336Y5TTR0lKhrBLqDdV+LGsOc9oPiprxHm0RiyQghD3EmJmg+gbm5T
EOFMikFj2bLYRODCrGJOfmL4pKYXJV20Nis5XmRSluYfFhv6ApCCmNjsXv454/Hj
QffB61qnCy5dYiLYNuTH3WXDCRNBpFkF5EMwS2JejrEESnvovbNBrTQm1wimfHZZ
dX1Hu+ZhyzFrUALG+sNusQugfPI0n5vEtgEdsL7hbjunmn6HeI33DbmONH4PzEPQ
AlzuywXXNNCn4onBb6iEYAMD6W4UZiuvQo2WjcGLehujze9aOy4Pn1dtOVtR53vc
ypAKUvdpHd9TMhRqv0hWSxUBa7HJyJ3HGjVr03PiQEpLnTTFTiP0aYiA4uFJjlds
hoszPfyCu30H+wEKy18jTX+Ba0yCaK6Yrgbp8zOUveY9R1CRWSNal3zRTK1EXiDz
l2XLHqzRnTC0DYaqdWiJBpb5Ebv+0jgr73gnb4Hibf6RV0mRHdNWB7xJlQI9NGeC
In9pRmOLxkGNXW5FssUZYidvzEjcyDRi3XWHV0LNOEHzzZA4dLTHxSi+sHAP4hZg
hCZv9YbuwE4JNcr+PLwxCrsSg3qqI68Ki1+trGQ6hLw5zeBUEfE9kP1G9qlg+oVF
x9pyLd+CBZfsI7FRHlJMg4Upglt+fddiaFAUjuv4pbC+nXkbnjgHebDyMw4JtSus
PGsEKxkR5ueA8bWlSx/BRe+ShUhQEJ3kHKg6pSy2+e0I1qFmEM2Gjdu725U+kfZV
FRNReZx9E0pFov4HAHEkB6K2oKf0JSc6VHDNeWyOENhfCWtdWkDKc37jlksQ9jxk
FlYrSaYKIjYDyKvqoIr7uzJZTHb9ReyNPZUAcOvDPcPkGF0rrOlfOnWpE1GdMr08
4KvsxGiLwYjJHqpoK37YiJeYVoJGU/U4SsLjhfevb61DiCUAMpUm4ttL291HAqQN
cqbuaz9EGX6nhqz1PKX2ywhoNmiUpIW2qfFhnC8Z3R6xwnF3SU2695HZAJziYZRq
YDlkkTXnmC9Q1D6oGjNjc3XnRCcQeFn7JDw5XTxtO17W+GXdErsi0/SvNL0+cQAh
8AZ+Q8YlS3CBfu4Ls93rn7sNcipM3kPSJN81i2xBg+4sV+9y0+4w3LEETQbmMkJ8
vXyvjzvi4f1DlfbJqNQrMiRjFv2Z//b/VKcq93IBi43R3bZfphLuoptQjbGYXWrC
ykhQ/+UZJ7WPOVCMJKsPn32+W7z4A1uNrYzfAzLJMUAk9pu7cNNhEsU5/g9p4iSw
7YbSNN9+P+oEYSAojuxXe6M12XDymRJSUHx0unXBKdfxGkTVoF7W+gQJlj3NV8IA
4fY1Yb8SoTpzR8gxbIbaKLvR7fR8ww+G72GvM91RFDs2y7f1SvIaDh3Fenp54y2E
bO2KFtWALyZPOwLaZ/3KJiSrfeiNru/uz1AxdGSqXYzhknf3e2hHvfzIdVbqdjP1
A/Yj92ogwGwYUvOxKucfmF7DbyH3hXQVCYOzrlHJ7MUiCYWdwr+ONzUU+hMPSFuR
pFJrOkahc5gX6zNjHQw/3jNRM030Hpo3uS6oMXIaoGRP+i9DJ9A5DIw43u/lQZva
fRjStqVnhNVJ6ppYLZqhbbTsotaqRuoemObrtyUO431X6VwO495DBc+czUbE36fu
MjZpJAub2A7vdJeKqDIOLsqMeflOOb+6lesDYvOdfGq7RxVnL7p1jkBsjXsVXK2r
/eG421KUbdCu129ilce+BJyNJCak6R3sqEsEQzYnFSSKdy1MYkLXZ/4xsVOKCFyw
SJ3xt8jga7u1H9z19xpyYtY0sJzb7njnP4CowAznf5f79B7NKxlkPqHtIsineSHi
j/2GM7gfljgJcwAqxAwzqfq51YW155K58O88hamwmLTNFYOmRMrn0R8Mg5ACaF5l
HTWj6yhkMjH9/35IX0SqH6xmzVNN86wJsa3T16Q7/I0XnYD1Q6bSEQVh2qo4snF1
J6bla/1l08HHzYoInpeVFjEDNef9qJn92gK7daH+K9zDm1wFTTY1hVIUmVNg//Df
ZZUynZr6U8A3qysMfVy3d1BwEj7F4A1h8HDh5ETmn+U6cohBXd7aFI260LMxfQT2
O+Uj1Hk3dA/EmLUsyMcZbGkZ0rE1xriAeRod07j0VII4mbdGdR1P2m8Me2sjIuh7
eXYPOYCyRVQ6CIxtBnsXkROUxTgdbZvvUfw+0NUCfEoCI20ZWJYqPD2pVF0tS4eX
UCPmPWvE5nt8ud2tsuvpJ7epxUsf20HuMdPW8AXfbalZb3sLjcZi3HyUq1+RLUX2
q8UAg4bEdFqbiyFHgn8xWwsJDT4ycwO5tWfM9/UEYZnhK1+ZtI2sLkAnVMswwIHu
TOtMob+rsL83vAZBKgfn2fVPfiUeRCziWT2WOOsCTTgqMUmr9x1CXGLnQBkJzP9f
NLq5SCjFTxCe//8/jSW16Pxz3o34TmvdvpANMfZzhAWLforbDEhE0H/TD+Y8Ep93
HZ7rBR5iFkEv/c1+Xu5IC7B5h0jEhrkNhN2jk7pxwv497dY6ZP68OdgRMLiLL1Gx
jxnTRIVNdgW5H9Vcyp+Z51v1wkK1Y7peaQbXT2ki9Shoj+qPVkmIHIrv0X6oCLfl
HizV+qD+1AKDJ/umX9AJ+q7AiFvM8uID0ne1oFQU6FX3AZeekxY0KnuD6X8TD8+N
hUOFh4qJHLhuftfEotjIHhhHhz2gUx57Sj6FRGcLAiqVXXAPP502+gX0wYPalz6b
G7cPzhIABSAdzRVpb0GQOo2uGfkum1lm/QZxKiVky4grCvA5CHIsoEA5njc6lYk4
viTVqa0+DYenw9CY8HX/i1fkRb07yijewGRtJPDJgNf1lUvVyhKbR+WoGzo+Jx33
kaLqF8ZhwVl98mbk3REhYn9HKkGlyTAjsInSnRu8h8t2KEZ3YoOhJCn5sPU3qE5s
gJ7ce5clp+zAkhZQalgvfrPyR+vh6r4ArMGOF81mCFc/lsxAB/Ltl+mzRC6vpSf9
2/XveSVGiuDLCXNqUbBkYmqxo0iUTu1hg3kFFBKs2Ra/gcNTuJCNSGEtq1PLagOX
o5qAK7MTCTxVkIYI6JAbAk/SCzRN2MUlz+kNPpGcTl3vk5gsEKskJOqP5sR+WYLM
uJQWZrJwODFzRQeArliU0d3MafjGqy5cqgtQeDFQ4bIVfx/RN3MoqHTLM1BKom6w
f3d1sk6yvhqUBrXGPXnVzya5c/8XuLG1vNtvKMm/Iy4i17gTfzxr3X/U1PUN9q9/
cXipeeNPhDFNo3+4WvEsnBXY2ESmKYiKq/oMTlvUMMZdpxFG48xbX1WZECYFXnpl
rwM97M1omT4flxFLWUbqh/GpbyDkuGr+9Gdl1OOLEk1XP3/qkRfoCPTyjxyGagSw
eumNXvnP6oSStLhNAu66jT6g3bXJL6BBZ8WpZ999syDczXS0pdZlXkM9M/yogDgk
QKZD9XNu5sl699Iih5cYZ15lyJfNh+W99DCpko2PEUtMLzfoji31Desxw+Hbsqf+
MqPV5hH8qUNnAOWgflv8vsjd5xcyemuQyy2bPI3DI0Zw/+mrbjWbf47/vMgD/lB5
tQqMAjoVouEgXCkhRzXOxSZ3OEW3cRGQ5Y2zOt8pFim2j+cp8rqKF5kCv4zyhFyu
6Z9SGUTmGh4Jcqg01kKbufzltdSqSPpvasH/jfTmsF7ZjWB3anktbbnD1w67LMdS
jEytrntxgh7etijS1Ce/BBq/kbjTIVr0yMhyCN4ITWHB894rhWFQ19NDS7MSEv2C
TAXdxhMV2AaxYhFuiSyHxtTJjl8p2q8pcK9Vj5SB4Qnu3vrDPslMWN6BcjMuVlCF
ZFwfN965lZ3p3/+LKb86Emom890b5+PEBJaWRbc94Ouja3vEVdJ1WlCwY9HYR6tl
J2/dLzWciVqqCR5BNyvVAVKCzalugFLRT1xbyHqL2NZe8OSeQkKh8wyXzhR2+ZQZ
cyoXuMecMzvQEy5O+ObovbD4jDo8pMn/LcGhFmIaVMgB0mLZWtHrCvvzb3gjjE7Z
IOD2UEDsZzcIyC73cQ0HO1r4vwRAQuCzRO3mpHGUrCRP34MKZZDKH1x0Niv8YjpC
1NGANUU1lc00/nd9bzGTlj44o5dHT5yTnCh4ZADCS1QgNzJ8jCUWN+i4jyH1BwqJ
N6ufRy3XIpTeNBK/mgqr3VjiWGFjstz/oGJuwapofTs32ndpd4Aqb3XgUDe/rU1S
MKjzE/yXK70IYNnuIih7LL5+bG2ejFHRiL7Bs/fFrj9dr1+uVuP+3K7dyV4z49g+
4zE26ltyfVOOXsqonTXl8ZtAjUVKJkRQm4wDf6fz5LIvjMieto0IRwANFVlZBRdJ
pgJWHkYLrwnGiZxt+fhLNToATeRsA/aEm0glg+LIiDd7DBmFwkFWH6dTI0RLEknd
5q0ysXCILd9Al4lrtL1V4jN5eLDdNFeohdNFUgamkhxbr9o/fhL5ndpLa45Dryp+
gi1RQgIUBVrufj662iqOTvDwdjLEjvCKcefuiuoeiaukBK1pEeld6bFcxaIoJa6+
DE1bD50XLpNt9iiiCgCgX3mcBxraMIgpuWI03Nt/JL7NiqM9zHv+aFVwri3UZbug
ZOxAiLZ8/KL22VryoFBSvf9yo5o7gO3Z7z5QiKkbxZrvOYO2imRAIKqbpqRI2WTo
5O4ujxxvEZtMr+N3+JUUvyGhKDt236O0rl8WedSjWRBCZIb1uG+SZBLPkFSYS0Rz
8l2HwN6luWhuGcKdaSCghA0vJPd7ELh5nSUW8ru2gZHcAL9D7sHSUl2Aa5cWz1r1
QSVubT9JZc4DbHEjC3XqMfCTeQuotzgXz2XJkT+vMTUyx/yL6h42Xp+1pHbItxqN
sQs2m12Ut00ci0xjgwkgap9takVKUwJOV3mMdnhl/dpkV5uAY4mf6UafKPxdcoIW
1oav8s1VW2I+aXTbhCpowR2xmIlYEOU9hp1XlBURs4jAA1oCi5JtDRejDOl0JYRr
L41gMYPdunp94Ne6ssU4RgXEMeuugkjw+WiWe+nu4H/AZ4Vvd1ZA4wb4BIAOgxna
bSRTSxD8NHZTronOOuf9YBXuPup3lc3O+jRPU6vHpklcbc1ZURAzJ6K+bJi3k5gd
aXVqv+ijAYvAD3/7jEg5YRVHoXC4vCGvGg5QEfA+u+pXWyyFmnVGUaTeBXzzXRGi
a3Fjn/Jv5RioiP9Mrc37KZGVufj1iHy7GVvfCW13Sby6yBmo7QAANwXQ4AP3SNNC
MQLjDFdbWQ7X4NtLPQ9Nq/9JtWeWIlFHuCTMGtIT/kQUak6cvU34ugzMmO2iwoMW
dLib1oNvLX8WQ1GK4F7jsHEwPpE6NQGJyvsZAlPIzSWBCTz6ru0BHyHGiWVieY1g
pz7UMZZnUWkXE8sG6bjeiJ7h0BVX3iunRWiZmdfKk5PwJrvgU5xckS1mRL4i6Wgj
ozVU4+VHrcam9CUL2eig+WAGLw1aghNWAYDT2QMTmNy3n6czUAvrui3Fr5syWpds
kGRiv+Ezf5SadAVBqo9Vla4lDhN2I0bvRRfN/JkGGTKOd+lFuGEoGhH1cIogM0CP
uWRNSHEiSDNmI5AGX3S54YtPe2A8GuVd5HMP9AtV9yPXqOJ+gYLBDqa+pE1TOGtZ
vdt1uSflpOavoFRdOiBWhDJqFGmRNMAzddf8Ww4TJpo/VsSRqFDjv33reJRFkwMv
fllyt5sdOs+3WQ3/ynDwrXJVOhdY6pgL1PElMd1TQFg01u2mfsUIOzAt2IEY6d7N
EiUHu3zob0bu7kj9SWynsnKXx0YhiA4hy9ZJ6Wn14j8TXtVHHJyOw7iRlxhIJH5+
cD8si+ThF3Rolu/svNYs3kHC/oA6z7sovdceKGqHfCksXJ+pNBuYtCkDOhqOcr3r
pG3bI5+d6qBdiE4S1rjvRWHEdTaB3aqio9HeUWC6hWwSQeUubc+tH6TW1HNyeC39
T/Z1I3yjDefMfLMCN/8u2/s/s/Y5m3bP3gU13W/RFhgRFQ/6qsRzw3s6ZLeSUJ6P
VXgD75TBRbmWv7FAOnwgbVwIfYvMTfAbJoNaTYqcybW3ewFwPuTsp5t4mkpokIqV
61emRHkOQnc7vUAJR5cBt2Qp2qC96S+J3OSpy5dpawxmMXbRwCy0UGgAiC8lfcC4
Aa56sYQeXkpXt5tFFs/xqSxiFFSOvRBMmYqv52Mdylt/oNJmX0Ok5YaYOcFKC3iL
CAvMleXQm75Y8iKKl/MvxXjAwuJ5TIuVkpFUJq3TO5Jng+7TwbQtwKQZrEmTypaT
1r5psnQCBuPFBhomTAckyoDdVcKpPkUMkmjCX7NX00TArRZLFANl40FwexAAeKfG
hjBoPoVDONNsaGWAHGKg1FLOCVJXr3yOSehbyONrxZYmxsNn9B1NhrQIzH/701+j
JjCjpNJdNOloNmj9WsfyOwcSbm+VCFrAYh7bSEdaDpK1GvAGjDfzpgdUmaTJmcH1
70haZ7MVIyntHm32s/cyHR4k74esPKAgdkThkaF8w05s+Ww0QulJBcx7zVWKM5T4
LpKqzecCl93zIeBb+vyQzXuTeJE+CdJJfLtUBWBzIkTKYeeGB9TtlOi1iDZ3flGb
ZBxzO28vKYaYIKVb/QczIcruUFqmscI+1zGyqvF61RlKaWejV7bJhFq/NJ67kSof
cjOO+rJ9ixhdN4jtMn+K5n6amroSSpfCK9z9OFK2FxemshQKppFuBXtdKFHJQdZR
OJEtvaHX7UCHWsCDSEu5eqXJcY5UZZWnxW4EZjfB6vWl9C2MImdjawELC+YOKx6F
VbKKf7yzAopFTei19Ajkq+XaNf0fUR3rstdsMBNiTC8TtiPuiOUIqVvlaaO7JZ7d
1oId9z+9epetjwdjR4c6qcFvMsdquWw56GBtbc4S8+2MHchZy3JRMl3R97I76c/T
h6oQUgqSuzlwpRsyFk079GqVMESvhf7jmLrFAizvZvfMKC6iOuQkoDLSExiLuUD2
vBCOOARQPw2yFwbvIJaAgq31YDZxktxULFLEjsarDnCswZhqJi0D0iUxVqhuUHzw
CT7TB+TwAxFo3QSvml9i7E2KH7s96TFj5Wt/C39A4hWl+4TkG5jPbpZfWEowP6B/
28t40YknIYxvakfmZdn8XTq0PhCS6qcttxI9M97xym/CanYoH+QHut1/s0ErHidr
h2jHFRlDNPDFvGlfad1d57ts+XGVP36Y9bDtx+X5FIYb1NIB2SjT4TASz+TDZtif
cfebbRsS7L/MCA6iGXzC7sviNQsv/ZUcJXMEAeyn6tzDwe42dBSkCqMjfl8zZTrs
AN/Qa2ooFXBMpeM7UxXHijtxgbNtKMuYo8QLFE8tXZOkqyaDtNab1WR7GkrRKI67
ZxR02WIz5nsAF8GAKaYWyv0Hc0OvJjMvCCERBGo0GosbdEagnfJgmLzlps4z+12L
/YFxrGf2eqV/4PHU2IobEa3RX/u5Tg/+SvkLD/DAqpi+PyXef52bt/geV51yeT9R
2hxt7QgMGb0oghenZa8KFVBXhFC01yr9oS9FshmXwuSbGSn1Nu3GP4ZbpcVlI0iH
K7DTWXEz7NYVQehtnkDmPRe0eKmqsLTWX4PorpeUCtc6LLkZJ9wpd3r72nTdh4qf
LE3/vCVitLDGISYVn0/SywyKtFQopjdOBdb7J6PAx9rZBqPgNiwD6gCoKY/gTETm
gzSUPu1vvkmy8JPp4QwjYjvmLKZH4zABHT6vKe8lXmTDYOd5AnJAEkA5TevnOMlg
rB7kXRpWVBmQhyF8sESo18zTMf1yFdinYao3RhSicM31oNnftuvVbSOYMcSiqG5j
PbEJ4F6A9JRdc3qieEACgOky6704JzUvtqp82zdhlw4kkTTqu2KTP8ZQNLgqG5Oz
2oTdfoLDsrYp6PqCyQafluJEFTyp8zOGuhylGR43AJlWf1NPyfoq00MthJG2ehXN
l+TOd7NRsNNRdhTCgxJ0BjSaZYhoSZTNeiY/SslmChwg9VFX852fIU0T2eDTXmoG
d08mGtCQRgWYN/U+A9nG4IDvERCn6PxbvCG8v/ohP5Q1Aq5+P0ujZvPM6ppPxNgI
Dz0sAVc0z3Rcl//SDjGndtxQ5fL97/hZDl+YDvfcN9xICgkVX6SA8BAPZb4pTO/T
KbKWyI1Ujhof2sj7yTCIn7SvnIwQG1Ax2Ha9JUlxb1PoYEu6+wB8+8gGPJ5rCbls
q2X3x0sgs1nxcRQFnYMK1g==
`protect end_protected