`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
ddtXksX2+yylW5zu6QL2Lhnb2d1sD00763mmSITNX595NcHTEkwn0zB1Dry37fOW
FufOhVzEJp80NC5qZ/+F0Vk7Ik02dIR0elf3clrjeJRK85K4e3Hoo4xn7YbFUIms
l/8VZSb14+JVGURjfswrIyCUotIzlzVYZ6gzoZwDXIi5gQIBf/gI+KxNXPaKV+PQ
Ufys/12rjO6aI/pPlqSm0hCvftmBcnezN2hk1UeXgOIuKZnogjOsf0iJVX2aOOWE
6pD/psybjbnsNB6kH5uFTA5frkzIzkzl5d9+YDm9OyC+k84E83I/7/j+rk4L2dah
QJOvksSIzN867/4Qt8qYTQ==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="MvBXkzurAa5VTw+1JJ70nePUfoQXBvZOku/SMmg4TwQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
oRtzZL4VJ4iwysPsC8SXYCzXS8Fw2gtZTOskLcDV+1B9Nzn1zTyNtlo6lNICRmmK
ZRVu2BmCc2G+fmzynYlNTnSa7C0Cuel6FYpxCBlOuk3OF2tzAmLAuDyOH3Z1Yjzk
a0aHuoCdIRKv7BrZCdALt03JeUmXKPdOmIlkVGFl8yw=
`protect rights_digest_method = "sha256"
`protect end_toolblock="Jn9CQpRhJt4rnzZPRk+dOpzAubz7omckX1MrFd4p81o="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 50224 )
`protect data_block
gD6l00tciPUa6pDNTk/+t0OO0nC/UTtBwLB41d4inuAUA3i/ALrNyoJVcBnAmEQW
ptbcNp5fxEUJjnOxnedyZEuEBxWRieZFQnkRdF269oNvAQza0TqYmp2uOv7pIEDD
pnCQAZbLD5fnGZSVWQFTkgbhHHezajiHAsX80PJJKlq8WGEG2MfFP2dcZYRPtW6D
O2WrBul9L/SVMe4lYpOPZ+zUZyP1scHD9VnNyd01dxH2PeC4U6Bg6b8IlDxERYF7
fWxbrljNogAfOU3ZtNZz/FXdniL3mGj9dHmLSw81ZKRFjlMLhK7Bpz4FtdMjf51R
Sp/VED0vyppzLsoy+BxmM9BriyDcT2PCTGzWGVGjYa+Tbtx03xgi9AHBthomUful
vaWx11ZOHelP18rTs3bLjFPi9zDKUHYE8m0K82JOtTBdUs/XR3x133WecT/ZZjCL
oGolbWWbjyOJBt9M7jRTcMArONrUVWucLXK0AC2Zw5xH+PLmJIlmcW7tdYoGeQzO
qOKWSLHwOPQY00ATJruta1Lm6OogMUMvJG/8+3um9/eU79rTyHS8rd7AYttn2Mpl
H4/0fkQz+LHTZY3WiOOI7nUkR+xMTQQ8bPpb9mnzwPcatR7SWDWve+rqgAg6rn33
hA2R6lzh/XBljVgKqtajYj/NKHHzB8QEyaUZdw0DYIGgp28rpErnjx+UP1SXKWsT
lPVaVUX5jp6jQA0OedVDP5jyraweCaOvrdKSrf0YD1a4bEJQev9FCtVNINmnK3SL
PGaPDI7SpW0qZSk3WS5ijq7UJC0wlCwb4VLrx227cif57WQoX3hXc1ShO36l/mO9
V9m3WoddZyhHH9BPidgnZujC+aVCmRC8tdECO72d6wKVXRPC0mtBi3V66QOUh4Gp
10G9OuB03uuYWtfaBLkfQbnCd4N8gBrKP06X0khUUGCL7qGiSOQvTGdVDdQ3rUBx
zQBHz4RupuzYBF+4aIRmQKuTFYdFyIRQZFyWu1GAaZBKMWbIAMzscfWr4TgYfXEs
9xooNJCMGSp7vPpHF/rHez5ol+KDXVCispcF8Q12jIMudT4QNSqO8oD9JQE2tKwh
5zi13KjvYeW1yDRPq5ul0pn3eAq1pULqYf932kuFcoB1Hz6MsKzobguJ8E+SS/a8
2Vm5gO3RXaXbvRrGKoBkrXL2jrgwvzm4GLS83dfa3c9ssWVVvwUcGsiMG/Kd7RFB
yZhrZPVFo5cS2Cx4j15+rAsQ8zXOLPbY9mS80/LMp2lv4eg9Zg7BZxLvwXR7pCWQ
51Qfler3yXs8kfpp/TEKAu6VRc6OnQtQj3oUYItBK4BYENTxB5t8PvvLjV58uERZ
iqqhPhfoyxJGO/T6lfpsRZQofHw0lpZ5gQWub3e09BYu8lJVCTT5G85uvTXKlMbU
1xnLu+zuT9jvCMn55R/fzlPH0nRFm+zTmkb5xNDlCwVsbFZkHHJSUbHGv4LUKlj4
otwot0iAOfo4EwzCzZswfbJqoGp+Kb/IAL3y5SFim02zxPOz0gFQkO7+o/1SfLIq
jQkUMHlGnitoFjkUMgGN0lgkJZZWT8y04m7ztk5XSTMt3xp9dQGviIcCjSh7KMax
EGUjYW/XshIB6lVW6bL5eccsXBl21eJhyDZY1lUaqzd46C29fR3qiYPDC5ZEFYrl
2JB45ETcI4Z74yx0GfPPGNxKdLT6VpvVtd5nfyqDZIT+JNp9YgltHhW8wRuxZouW
ulARGOaDfnC3qNfbb1OaM2Fc8ZaW3devPOc1UWU02I13KA+hOCYGh03N4DWTQw3k
Lf3zlGyW7AlyFAlY17dy+oZ06+ExARyMxNQeUxqFpMoleyv4Av8pOWnG5jDtBd8/
IN+V/5ZoZ3Xqr1M3Kg5YGXgX06M7tG+IqyunME5LtRRjqb1Epmuwg/lJ7Pk9DqDD
6FgWgTiALYjDuaGMvmb+OJSpuZmKD0z55BIHx4HVWM9FyvoHLV5hI/H4WTayFdxG
ultaKlnzf8mEXxvGY7PNtRsWYDIgaS/58dAqLMjY+Xts5q1sUliKuM7GnqSufria
6yszmrCorSVcezmYRUPZkVgkOl58cs/6lFboGi9GUN42vu+qdgt6IAAqC0Zy02uu
5pUVVso36Os183963HibPHnPMAH1cWYIowQCcScRt3/GtasI65HmLbFvucZgKtnb
HaoD1fY2MsQqi4QfPzsEvRVsGoaZRbD8nVJ9d6NtTINlX5teAw62N5uRMFkNvjT/
S25mw80WXEBj8je8H6qcDXWNrr1tRARBJ8q6J8i0raNoL5wX7f4f7ublKsqyyHrv
Vf2TROABRX/6Nq8CAxSeDr/C5vQDGmZsw845qZpRKZhKVp7dY9HY+qSwi70m9+s0
B6ozPjY8k90g2aVJC+/yOZeH/OXsGbp+UYRaAHIh7gWqedbkQapz50RxWyO4UlIj
zvcU3axmR0DYNtMp8Y1/506UkBUtGNVwO4s7jacjfxXYxeSVypU9IejLKArGFiHM
XW8ciDUdg7ETl3psdghd+AdU5LZMoDTWSnppagKjnWCxSF0CRfyJOdMcDf2aS8Yb
uy9WlR0FBf6nAAKC7JtQmc7AyyiIOmAJda1zX/0k836IKcX+jgtjnHoTlRfW5wMw
rN+pVluZSyiH2oVoJ/ZKcvckTCI5SFekrVdWyRci86ah7C9HAbYZLMQJ4R7OMEvh
IyG/2H9iHijSv669NO6VvM2SaSGYJpvHBV7n5bb6EtRGY+szwdF4cj8jZN6wZGtY
uRwQOkxI2jY5MKXRpmBu/VUop1iJWn9AuglRdhoDMxfmaFcFLGIOxYqc29DmIP2i
WnlH98bYZ1Cljt9ASz5taJopelL1/RqzKZxs2ruAhgQjwmU4bcAUU4lLzSBMA+KN
hSzfZl9Idi5MO4nUGZJuwWKKtT9mYB662FFkp2Tpw4camwwBy0AHySPps/WnIB4u
e1uZEzTz35Cg2h3EFYE9ChbUkb5R8YN8ll4fjVNEW55uxEUbBb1tzyz5VFiBZWId
6N9l7nJuM9coYG2+WGWXaKdbY8fip4+lqrpl1o/J+S6WLPLrAvhWsQY4Edns4Z1K
GIScBqn98uUjJYEis86e5FDaVKv6K4KTstj9J8SyIUwXDVNJPwCTSH/uVSEenJPv
ly16GtjkjjhnohZqX/gHfsahH2pJJcH7nbFMgt/Mk2FMH7igq0CHCnypTWWNDxf8
0uaKumXyh121fcOceCpgA6KCvkTYGPi7jAcHjwGJQrJFjcj3eSHASIuoCCpTeJ8f
66ZwbD74bZDjcZ+HLQQgIpTZRS5a7M8kfg3Oo8makUADL57sZwUY+SipS77o+qTZ
2lRXyyKG1k/VQM8pcb+5zNHsWsI+n1NkU0oY4vziYQzcFst9U1xKV4r6PFXKkl6r
3IAg7GwhXqFEY+6ffvAsYd6agUaTYAEiqrnn044jkwSG9Kk1uuq1V3poLcUuzHjW
eVQFjBCLG/dGb/VRYPpbIU2GA9vSECP81VbzxyVVT45OqYCag5HaML6+YaKskOaS
oM99qlwUzDamxAbXsNGnpLepVD0P3pjXYAGy5Cj721ix7IoL5t5pDOYbm9xwNu51
BHrYoSHvfxH2e8nJrSfbz1/Gx6WGfbm/5szYQauCVfUoSH/9A+tMra/BqPStnlQa
48cg6wDhpvHvPG+syB5nf/esu2jagiAhQ4CSkQpmDRFd33a7+AU9pI/yuhERphjv
OY6jcSzK5VntnKCQ3Vsigbu8+vwKXuB7WIwvPssSO71vHqjDKFDpzqypWTtWokae
5xR0ioXLJc6mU7pS6rDjsiM+JBbjPr/73G6kqtcbsYTXM6Eex8U81X4oWYIY5Q4C
dSwgZYBIRjZRemUKBUnFzqzonG1XnAGtxe0fPnjQuWg8jdupolfQbLgt8DZe03q2
BQICQe9bflQ6Xsvay1LahK2MtmaJdIhWUoATNOpHgntuHDJA45siIhxXCUZbMoU9
ST+fHOxZ6tSZi2iQQZLeIMGIIR8NBVDtYgU4im0EhXhiD8e2guNO1pzDDeXkPR84
2Q6guLKi89Y4pxZaAsc1Scq8nv7dFOVbdpAl36to/4cMhjY5MXox3zEfTjCSdK6I
thpgEpHZ2bu8KRC/0x611Yp4oQU95kaISquJF/BHXMdfduR+NPt+JO5bv610JaNU
OrPfpzdCmt3Q0iA5YZ44AwrLDOathgEKSHSYFtP8QhXpxYQRcqFZMnS293B0w67b
wO61UVxfMiQNe1xPfsFmYQ8Asid5pWtYTPNIVGAHedSvRfBfrhpdeGu4ViQH3gzD
/eGwCxJh6tTTwQuhz6xm7+m1j06Eqd1AnsaY+0rjcNlw7koFtyxoJMRLt7E/i8Zf
0b5TeTYAdVKXSv9w2maZbOn8lzBofn3ABVpD3h/9i1MdGbY3JZ/oV8GhHs3576yk
DrIC3QPvl749NgClLRDZEI5beAY8XimWqMzaXW1H5KJNn2BNUydajPtABmCLeOLx
odBJvYlIcuQwcxPFlRseG9qLAN+tm9R0gFfRfQNTM9EniFAzSvAqGPnP53mNIK1X
awLkuw4jiPGNALvstlZNbEw1dDC3uYl7frg9wE9iSktJkcmX7Dq9K47qEku1hGvZ
pDexD1pxzAGN170LGPFY5nDmJlzVJnwB3Z1ep3aWcd+3+X/hhrB1hre09hfC090Q
MCvqyt2IG9Ibq9QxiQlwIl9GwoaWWJ/X6zFGfz+m0gd6EztscSgfRILUsRaBmfCa
Xf4uteleA4hwDlMT6sk1K50lF/0jmE9U8YMlxnFjtP694T6YsbQM3sm1iGxJccRz
ftB5vKhZO2O9frJWiTnLsK1YjZeZpezDAKCvyN0ecY2ZY/QNZlIVi/sEm2kFn5gB
dhb8teWVi6COdWBPFGzK6v3fRnq/TyXpRqVdrAeGRqp/1up52z+17XsYnwR+cRow
VQ4uT3Qa+irbuL8Zgip7PAR9oJC8z25rlGpkV1l+evBKBTOyRq/1QhUFdtr0Qol1
aHDRRfIIZTwX7ryYcNaP6wj62zlY5Mdzlqz4tOdIqwIOEQPM3fuGCtajDGnoAKur
+SibYsFAlVtMESbBgYqu+wvIdQOTDu0kn2kp7wgtwF1VQpO0jZ9p0WmsFa96jn0y
skXEP/kbZLmbUUBeas1d0gLFmLP/f9wgCu6MtSKgQf2G4RvqjpLNoB4os0NENw15
E2mZb1vNdSWvUpnhs+QShXV4Skt+0yzRPwh9vi/56zcHTF52kEYlSqomSzTo5ORM
nlromHZZWZyXQteXQYkKEhpITAAPte1y2AETPISBXMODcdWV8C0cV6EmI58xoTzP
//0SKaXXBQzL93WgNIyMUBoI2otphzz5cELpNVx277gwpWJM3c89BeYinjAl+PDk
7ae/AR14ZYLyxd3s67Z/zVZ17WONijhIteEGUS5S5xlWOQjhW7cbxpSZ8MOq/cHr
bnFBrpPSQ7q4l56R//nVfe7t54INQP81qf8z+AmqvaVwbvxlprPTFkFcOhv3pUYv
SVndNnUyLTP/begNx9Z18xIdTFoPdfnMxjkjx4fAyUmmq5DueZ7JnsYnFQHwQF0P
MwqPBhaWqX63xYmjNCD+Hn/lvhL702IhcgPkVd8rk09YjK3GRAzfkUU4/FikmgMM
CfIehASl5UzTHomDCy4uy51Y9mnWUQkKePl85AAAGk6EtOHxZxWn+QEbRJUjW1Ki
Kac+YFlKMqjPgngZb3Gxcd5Ri4XTkpndcOYIfJgSTC0hWHj3aEzrKkgza+6BjEwP
3hWanemqZRYlvZrI72cbAimhs+30I3HbTuwpe1xlSL00pW4mm1lymeeuPvCbai6W
FATP5TJuoQkIN2t2ZADkAp5gxKhHPH3G0eUN153/QkjRGHTxwYkqWSKcTFeM3MU+
HfLNVbDGuFU6DFuAH2IsGwoARqRTqGybHkWgQbYgbUUo+A15M+FKRipbQJpA+TR0
/HiN0mLygkknilAZ9mg8zjz/maIksano/nW1ENkBDM6H31DZjrTOa2xHhslZVg8Y
nbfo7NLvIem+sLeMri7mVYOLDYkp6aGyTjWfE1uZQ04wyojygCuLujQuL4xHsMSR
QAnwjR6j+FUVAgG3cueItAdyaNYXJLJ6t8GgjmDDMXeiXragROwJCcFdRq1zhJTk
bxOmUXwOJyZxVVgHLKNATYT+laOPPQf77fZx89PozN1iDlxywJVPfbqk82pyPyY1
GE8EEOna1xLb5npu3uQaPF08AkbGWjxrk8kpc2SZn9kMQlQnGasYRCkX5BfRORpG
LfS69SBQLouU3xMC/aMVyKsd4KjVJAmtUm7yeb2Sau2zsEzRbr019U8rI6ic7s2s
v63RHrx/mg4UONpkwbqEnuB426Akg0Bm9FRByhQdCyOiL4I0/MXa19ecPlt1JzbE
PByojVvDkutsRgmlLweXydh4CHtWOqhyKlWCBiiVPNfPvXWo90teAbydZ0dstte/
gcFEUHSGmsTHffCEbRY8+EL66jrZDQfj7z4ZRtMTGMNWYf7uuY8IjeLzWxmY4j4J
NLNi6Q+8pfN1lz6xvhvzeZCWrRoHKhIUACld/5dnYQ7wJbAtaqYmt61xbXJU73R6
EO6JsPyMi4ftk8AoxZAlJD83clrUcTC077t0e3DqwW2+yf/Y/SwYR5Tja7bHSdfm
agq+gcpuND94jhV5WS6f+iEdkDirk5U1JIadyVprK/iA5HPlzdE6fbwFM953kVP6
bAG2LyDhYywJnksL1AJ1UbIdrslZFHyrL4t5rtuOljD/n0vvVFWnI3eyEdnzTT7U
5dBVPuFg7OXwk/eDwfAzW8ey+zXU1CkCQF6Dxb+NYHvp+arxGTgRnnhHyhVADAwk
vtOhs6xdy6BD6qA3dDCT0ENM1JabGvZv4DQtslwnATubISI2NG1cxD4ZAA6Hfmig
0P/8Uu3DMu/Fsr1NS4Uk88eYsthVVJ/NVNydgvMlZdJXFsbPO+p8dPGJyxCy7PL+
nD1kPrw+b4Wp5Z6oRAimCxiHiFi7qiKOowh1OfjX83jOuBjmQDKnlqoBGV7ZwkLC
zgcDHhZFxQxkZGNxOCAo8r4D7s987/XSmT3cNJcESpBpvqjxmqx61En5Gac1xn3c
Ae0lwaRIi/j5J1F4Jm0HZ5osPGGhlkCc5M+YxvOyXPIgkzPr/v8KNaKG9svc9eCm
D3I1oTHKXDvVPqLoLuKygtmVh2RRcLm3KaFNn60ZVesMc6MZaMyIB5XZr59j8tqz
kSktsr5JH+y06IhyqJ9aXTZjIg1bK3m8mMXrYgSkBZfaO9Ojj/7k4RqJnPh5VreZ
6uWPwI+JOXopElkBvdZMeReZ+rqX8TGCqpnTNHQRNSPUjjyD79RNLOEoNyw1AEPj
jmUQUBhM8hcdGOJfdIHc4AEzj6S+PM6KgN9gvP45odrHCjnc0yEdenysm4HEehXU
vHMihQ8WPRXlvC4gtW78/izCmG5ZnQTKMXf386xP8oE6cTsLIsej6cjaJwRUT8I2
F63XEQq41JAC0BW/EdO2A+7L++XUKmwaKKBQ/323XYhdBBMYKor4uTuWSY/jDEgq
bFWZJiHSiondRVId34avekCmy6xsBJJqn60wQbHGGVr0TtcnnYhy7n2ECKuFGT2w
tH9HEoj/IgmqbX68mkLn3ZCXE34ncKnBHyVpXGwPmG2iIUISWmC3nQ+aQNCgp2Za
/PAoqt06WVAGlxdKUPNVrI6NKifF7d/KWAt76HwHSpjG+JzFdAQx/p/USzdOzLnB
ZMi4fE7kd+cmo2HVf6Iylnqyi9cgcQJwcEyJlDeGgGjc6mrCg5EGo3AgHIdN31FS
BTSOEEtKhvTGwT4+hdrGfTWQJ/s5TvM+UKkxxDmcMvQpd6hBVtoGF0Hwju8n1cS2
gyYpQ5xqxrdH0sd/KA2DjC88Kg/mIp/CiGe05J/pndayjEQm7aaFHdF/zyh0QAfn
h30qXhatMK4bZ3b7bz38TsgSz2K9TIn6te8cnz6N4rHgyO8aVoze0zZrguSZh0lb
yGB9r/wzwL9WPhvkRd+VuEhPo+z6kQq8ILpiYdsshR3TifjbIx7JGNb5y7N9Io5G
tZGja1PT156ehQgQIAoL5DxPUZLRbg4qyouXMYxerncV7/6SRynJwWWW/Qq8CRqG
L8JoR889oezaWVaXc2fd0M5CxeDdeBEJZnjE1QzNLG0ZUQD8O7yo3UXWZniscQLr
aeC2yHqFLM7Lvs82dlWrTP/RwFlGVMBBeSrZd9xavtNNSKVhcstOiIh0pRnBLE+n
4VccRv2A0/2FvtGP7FRf5HjaRvj7cxkdJ7eErix4u5QPqoagdQTwKIDAoDeZO4Vf
/oPlnnOpumOOD5yLbunhY6gmt+YuAuMFgYBnOnYJy91MmAoPMPdY6wIfUBir3WJw
NYxhrBxC/ow5aB96CM0w1E06RCxD8+VOc6cRyAtOPeOY+yXPktY1bOmZ+7srcOty
AMl1PFh41VS+9SFq2Ex/+BD/eyBsJ7SScI+yJQ+rDyP9JBPTlAOzETTMSlWBMUh6
w1+sPXB3+w3eAjRGyQfZBDcPFljiufgMxHBJmhbmD1Abue30h6ZYi1lV1AcFaGJ/
XhvLb8biwRbHJdqOLstuqhZ3qhGCqeLqDsZL2d5jWsuROOpgTSz8lQRXWpUBBAh2
l8nvnbfs3cA+5AwdFmSL4xpZ8vOCbjo/ew1UJwHpz5dPtFZ3iiz/rJ7EulmuvoL2
nFAyOYBFphYxyECzeRklP0l4cS+HegQQzY0OkxlLUbY4LKFV5njAftYMQG9mP8KD
xdHAHJPM5j8PqDIksJ29ip3rJBBKW9XFVGumeIPe0147ME+6JNK+tTKnQ1fq9XT9
pE0K2LMCAGZYWWilfbBBLThCmkAqJj9yuSLIm2O+xJRBb4kAjmp26WZLFFtJBX3O
6he2XSt2HJ1ENPyr8CRLiFtylUmFWxehFvsrjtA0buZ/gic6nI2sJsfPX8WI58C4
TEgGlBckV3qE7C3K69UmTilGC2z+aW0dLqDXkWWZpJznwfFaYiAX5YkvXT7nNkX7
D+LBGTFbqvk0cVvI0bJVNswbWWMjVpcyr/m58+MZuuS9MUCBRyTXRCyBVBNkUo+8
8R5HCvpWTdaZb55NqM/v/iDR9ShorqHm/4y2ezu0+BggJYK+dGXOlxB9UhcU1vUM
4BAurccZZNY1tndBPUXK+wQuQZiGWeNAvSJDE0UdooCQ8MnkzY1d/OaWxsoUwnXy
eEt4G0uTFyiZGkP9V4KM8/vyMmP+lMAY0XiIrDN39wGjaGuLOlFQZc18NGlt2Pj1
5z80XNArBOnQIrdXyosUchHi7soSAbGFHPJqKDRgnQzKTc/Ey/2eOZOQ2e8pBc+0
/yyLd6OkDLILqEzrOpDZ6/NJ+Z+T1Ez4isE4y/nfopLDXol2Bbfq8fsxurPoklnh
H1s9pMjRBtYn0zBwRJJUwKK8oOybFMKSXa8G0mip/O12kjnXA+O0r5+TQ5WqfH4Z
E+GzVDRts1rfxs3DGPC1b7BZR9vonkvW2b8pyhVwR5jCmbDk25V8oPHF/fNQSDTN
Ep6HG2y6FYdOJ2J+mj7N8CvkEZmT2rauitM+YJvRM+9aSD7ID/7T9NhzWQWApc6k
xChjH1qbfl8PKlovKQm7rL5BFXAV18OD3DT3mOe/eHQMaiq8pjld3Ee+QpTK0VvD
PzwAwyyFdL9uV3CSYgeviDXBOqBmwbDm/DJk1KXnJYOl2ocRMiWlnJucR+LF4CVY
HTKhUTgSKVIAt1+R+7PRf9mRxtV7MLyG/wbxaLBT9mJNy2Sk2xpyg98UbQwgn1ue
v+Z17X2c9DtyexcJzwrZr4Ef1WsrTQNpiB6zEe0LuSIfKJiZ5DxI0tW7q2XP4PDL
Dh8VtXpHtzieueB74NjJIdW78OvyLcAhuv2rA+2J65y1cIf34PThHAYMYcKxUG4q
KnEJsVkgk56xTl4Nyz0D0l0zlJ/NGX6K1wWWj7m280hOHZrMjZlIhVBX2O7/QMCX
qGVLrYKw4oXxLeMznRB4hej3pEOhLIQXULB2qIuXSdypL3mpB92KaTaw9Y3P/w3s
vXKKjdmo3b8NWt1AExN2B3++y5xoZOcHgG7Zu0BI4S7WZzEbJRmkvJBvYFulw2Ai
wz1fpdNuqkMEH3L91fwV8nJse7yEcLGqxVyz3KSAwN629FG/NQtFb54QoYEs2Kf/
ncEmNWc/NTCwCgEPrq1HdoKfxmdYQZDe4jKgCvxOq1Dsy6eeGv6kr4OmQNJTcLvd
VVv7r/XjqriDj3d6kVmMHikdPnANwvaQy/RFr7ywl5Cg9htUbe4zlsKgYpmdRDf3
5KpoUo4t/UsxIhgNuRPKO5r9J7Lmm3H8QNgo8hMZlLczP8q3C+lQ/7Zg33+ZJJGu
+r1c3/bcFHYPBH+IXntbLacdvl4NTFoJN14Ec707azJBcyuxhlpNIp3xflMRa6oc
2ji+JZIBKDDDeT1+VPEKz028KlzlKi0XUfm6cHrwOLGF2obYL6vm5vxo67XCJ3wo
ekO29YP6rclK7H37ffR57dUrQtrNCtJQG+KLCvmxsrbaDRxWlvBX4QoB89HE4P3p
CHr0a/R/kjpt+TUfVO85CAFufhFjBJb/uYQVI3rrDtFIJXIwGAyLw2bvaBX3KTmC
xide0fv0yWVYlWsYcs35kKE2eGdvEKq7J+Ui0kNQtsiUdc8r0IXbug20FzwnRFEs
TkTlLM9E4ZLUje5g5tphGauNn8t8x+w4pId0Pp0a/Gk4Plu0SKGPlrhZ6Le0p+Xn
ua8vDCEDygPDIp/E8yN4Lb8r+u8ILbz/vSHqBS48cGRg3ugZJ4pzGUoYYQiVGzZ/
68iLxXCsEly11u5gRiTwCPsFLxr6XiSIsuwKc8RBEE221UsyTQcx5wh5syXzpLY8
3/yovzHWizmjPXQ9AnyKBmlnGLvZazud/0bygHXWHZrImN45EUqDi2nZKJZrC9OV
4XriV64A/PDbjKPJ0YLtyCdVaJRHIugTt2bkhTboKVHRsPTLXwB5/SRxLlXO+LVN
2rMz0WJKihxlq267MatWDzPqj5HHBk15M/k28FtJ3opremzpzPYPiN59xbzjhpTn
03ZJfWZ76Z4e2/4VTGdEunmvDA0IOknJLnsqGLCA1YEE4rkbzGaqggKq0+0Ma0yD
WzmTMQNbHvK1pGHWrfE14Uv++I1nuq7IoWkWy2OfYTLueH3wKsMTrYuZqSlv2Fzk
kgeC/8wic3i8EYFVQHhqMe0XV15itDNHhKK1uQIWsR2UNURgN2fhxjb6ZQxH9mOY
iwcoXoppXSQlQIFIzrF5cCxy9vjDu4BhvV5AwlDwxm2Xrg/zaYO6JGzJJNIxug0v
Lqrqg8nIX19hc5on6WoLzcNalMJCjmQp4+TosfYNh48q8TfLDZZ5FSMW9YPZghrs
JDXj2l308vEMYqD1DBbrVKqINeKnpCKVCwCaIq6bGJuk6BzINg2cp+KlmyiXNWs4
vFeW5Rubk02Wf11gkHfQ+uuuYhfMYeh9wm8O3ZpuPlQeaQfwqjFbXLZwpfHY/lIr
Z2A3E6pHrpZRv2hNSRA5lg3YB6udecMp17+W6n17hezlmYR2/I+6FTU4NJzxPMM9
7SB04pjZPmdk6ublaKJY13yv3oLH+7Xxs2aZ69cDbxze7HbsxjOR9bpOsJq41EH4
EfrX4RggYTOmFL9BXEvLtPobrAZM8GJj0tAuAd0ILKt+VtCghUb2Ne7Fdz+FuQ9M
6bOjjJhCdAqhfmvKpI/fPVX9/PaOfgU57Qf/7EBjyLQjA5vemoKNjPEALw07t925
HZ4Fgev10vRMSctVonZUCZg/iEs8QdomHP7C90fOdlP7iQhFZJ1ON0X0gQV3Y0i5
JY5s7nkb/krMa0a5gttXreadWZbp0xOgPQyQSqxg7xZrgW36ME1aVU5atwJ26bf1
n2+XY9DrBiDuMnrR9u7xG9+ElYP8MB99Ygsxc6dCPcTvOlt2J914i2kvQPm/DZ3T
FsQ1pmRc6cWkXoZTPNfFT81Irl4PtIGE7HPg8s7LztbuQ8izlczGmAtdwSPv9M1L
FimRtsfi3oumxF1ugraXH377LKeDcN56OWcPrpwVzT9tywrOoJp14Xr4Vy3rW4gl
oQp6YkKnOYISvO7EaZC9JHZuCJJabAkR1ezkIbiZvPLd2H+wGGs+CmPbJogdQtsF
zKSN2t8eFN6vp+HTqaOnP8+LIyH7XB6UYMqi8CSCAlvbsRhMLpIw5N/byQdBPM5/
61HBajpd3dU0TxqhoiLNs+N6D6ceBEnrNRGVuhwtqWc3J0NxG+Ffc3OhPOg1crAj
funlimFQ6NPemYpvvUZAyZKCAMN+epTOm4v91j0y2qJYku95PlN//WJ6E6sYVGqx
0Xpf5RVH23PghHKp1EVW/3Kr44GYalasSU0WU3TD2MUiCXZ3LOerlGp0ytWK+gYm
4suBNWAGmcNpqh35RFURq3l/enF9AKUtgD2xSrMwtVMJPyKR/21cf71tLfcqPcgh
G/N3Y9vFFOaKTCpOCh2/Mx02p4Ywk1p5jKIJ++kXRxil5PuVUdwRXIUcwaNmy6jn
SYq5N3/COZMESD1GbcFytC8mDcf1w0k7iDS8SUNHiaeUtVCYCoIPcdJM374yoO4A
saTuXhrSWPPboZ2rahW59zRa6TDFEZSelLrjZkT4ixU2DaFU+kIZVOlXSlUsN6EH
ap5gO8ctv719VTt8iV6o5xlEUmXgh2a27666wwl3u2Yvuv6YCYTukBRqaT8sDpfX
U1OW4dmiwhq7obsLVFp3nZXG49BTZr8hVZ7wnjIpoAXPzkNVA1z6kHytVNuNjVFM
O6XFWPAXnsu1P6JM05ath16wuBtqlaRkrN7O0Bw0W8lSsGSfRzYa9F26mDmFcQqj
t/bw2MdBGEqHsATt5gKiovOq5ervbhPSWQZB9x3i5umTF1WSkY+++zXP2G8UYvP3
ChpTR/MND8Q7YCaFQVD1hb9m6KUSx75Oof4QXSuddQoji1/AD//5AkeI2rf8EhaP
C6xFkVPwGrncaiFMl1i1ohN8328PwoOqZyIIpZ8Cc1QMkh0mP7Hb5v8FeQI/Nrw+
B6R+atenVVQYkkP50z2W0/muKwVYpNK9hIOmMpEU/AtY38aH/lWHTHe35rFeLS0R
krHZj212vCVPy0Wa1NmetEaRDkhLYfQf/NWdAagY44V7IiiNu0Crwvr7MF4Czi8V
goDWLXvKvIoLQRGYOmRiItAG9wZ/rizX2ySheBp+d2NqE2vTk60AyCU7w855vmic
QElLwQL+KpNR3TtC+jQovib0V7kekRuoPlRi0myNmP9EZ+mzh67/M+KERPvENHjX
wEX+jDzbXwOcuzcbEhlERuxxgFkNTiFxzlvVQ4WGP014/afvvxyBzPExJV8Cxy9Y
lZWWLZhZK3FWPNK85lmGgeRdwKDoax4u2phdIytPP/xScSCAMlG5HPn29TFGSLXJ
mrxCG9+QE8yxl8fKxXIqb2DvzUkT1FcM0xnCKHR3mWJJbu0cVGokLPhdxZFhuf6g
0/5NRC7ptSvf1cP0eYyyATRSL/yjIKdu6wesM/knCZE6j0uatPz63BAADYXZ++8C
jYoGbXhnW4PEy6I+L9gERJmuefnH9hc/FXj8l7/V5ldUHpzHtMbPDsd/nHV0UbKQ
iDaDgYzCezvem22iwWE9wi1tKP3z/+F3t0slMObwYSgwFXTlyFZqBFGh/OQ4MiWk
3sZfQTOMM8XMB8JldcFMgi81iGLmRZcMbEM6Q3xGC/9CYMoDmYqeKtwFG23nnrJW
YaNycAiyYPTev3t1Tn7TiBta3hsHrM4T+XzCqHCSAEjK9R+d+JqByiHnXEZYTLOT
b8r6SJNPJjJIwW+0KBOgrFTuNQBveNxT7dyFovekv8zWLsZjJclx/+H1q85L4aww
W1JMto215J+BKDspdbmh7ssiNfP5ZMVpPgiMO8Cl60WADZGm9EBHrbU9tD0oxfoy
dAOSqF7wJKVoe1F5qo0mFYBO0or43XXcg8x+gdeZATSCmXXB/MQr8uR6jI4O+OoL
ZdlWIn74rVXI4wkEKiaSD3byQZWZQZsI6yLzDkJjEgkGwXN30tFvSmPtLhoy8ps3
tyVwoQ+UE+yKpu0WTmFC+n5GRQmD9Hikez3GoJICe40MhUnGx1/Hl1d1nuB57Vkv
308dL8RL9t+SZBnrtVLDZipm0T4rcCjTZIGtS4BuuV4FSTOLsSpbLkKAAOTC/uvR
7mBrjzVXGqsV/o3q/yETbk6hq/u9yrpg8Z8AnZCc4YzYAaBaRodxDomAwGbTn/AO
E8dQ9HHwTOrq/5dxUnv/kVvNh72lWpO2IjqTzpXbdqeZLhO4CzI2NIVCZIoEhNpx
5ZoSiAivcca9DVgRWxlfk6q8YLaDaLxcjtxwSTF1fZSajjZi5W/ThEXN7Mxhu7ci
q/sxEtzbuNk6Q8o9xkHR6EvZVUJ4k7302+geT6datuWkG3im/bb5evkILIoFZtDN
kmb/prpB3MGBOtUrE3h1X5HHWVKmK06C2QirbUj13bluk/LW72UaC3UIt1bJiIKR
83kaxODsIDOKhVfS92wVAr8s0L/2FKv966swKUj8kTmYvQmUUjJxLxRTgsTmgxvP
jwvCNGJsxLrKw0TNONs48juggzNN25GFmbBvjOSjap8CpIlmFfjyYi2K6AYe9cmC
iuVubMlH9B/8v4PzE/gGX+PcZ7tLO7lmDNiILUs9vfMlitWj5XF+ec6p8BB1jcyt
znvH/RAJSmiIyomvPEyRf6nWLftyhSUcQtYqcGgdwZEsIMllG5DAGBjALuD541IA
g+ar5zOhAAfo2OfrnMjzKEGyGPvxtTKLpBHoTL+tcuZ6hmi1r/o9P0Nb7umvkX20
zB/1fdYl/28MOK909Q4i3DQBBMN7vDTpl9UBAcJUPziFyLUQG2QSXJsm+P2NWz9b
vmSvi5LThr0sDeXH4ZqPzdsE7KB4lhFSFmc3VFPqgwtI2LJ6fizc0IlYyoZ9q69o
O74y2RnOFvw7HRYEXm0ehPVBaLvk7zDrKjoaSSk1bXRexQsMLyqYV75K903yFA5f
rnTfezF2uHTkTscHOy68JxEiIRTCpB4W9dKuuM5+XtQXF5tw2c+iWy2QbiAkE3WU
SahRdHWSx5jfYr/0g+1WwlDe9VYXlyCZtnbrebyDEwJsMsrLBSc5/+23FrLNemJ3
erKm3FvjD4pBFeiUeZ8gzVywINgvjMbWyjStDuOJJM0o5P0ttyjB77Bys4M6jjpI
FMZ9dd2R3KuhWLhb3miD+iPVmSAl5sxdaI8gooamL7MfLi/cgs3HtP+ste57HGM+
TMsf6Q6tBgL6qPeReOnZQx4QCy/lRorfVSg2UlHdKownRsmix8QhRPe+JVuD69Jy
6x7aHduBHFtnbtwHnZwUwSFSLwRb9avA3ciNorI2iuN8Fibdx6yz4EEkTHyB2S5S
Y3ZHM2EJ1gqzOgrAxkkHocQGNGzV+qe/8VtHAVxhG9luvuojqst7PJIUSI6t8eia
54kjeq7R1w3BYgPBZ6NXNI4l4Z0kwuuZbzP1l8x/pNagGvELgeD4qfw7/p+/94jV
mgbdvB0rAw0vXhUhJxWS7Z4+pQzSZ1h7Jd/n7VI99yMdv8EYiOJ//aX3a1KNYMbG
tNITDT7KBsHd3QJAPnb/uFLoTxQilZiu/SHgb0O+OxNbtUY7igSh2OewliuNih9l
E6Q1rdyHWbihtqvfK4OE+UGYm4QG9HSNVYVoX51TZrUNlbD3ZPl5eolNwJEYCNt6
yKq9Ifdu8L66shRvlcJweUyZU2kcHZB+ENo2bD2YhhmupGeeDAVlvKpdZRKVUdt0
BeZGzxFQaxl32SxVukFaeLS6au8UDSYrKJwqrgDvEyT3/wXyRapgZ/nLdFq4IZnD
tPJqqCD5R1ktbBKI3p3Bwk6gU4UiqE09NG+YRQg5FWwJWXwgvX0otwx5z4LlvCzX
Cw1EyU7EMKT96j7bB4sMnH0GkcDY5WvkRXV8fIocriebCzD2BQaTkV6cYijejc5a
loJLcFUdLhdzRU4aFbFPLxQ6Nx82Ki3enbj0ir6tX0m5q0pyAqdZjyfU56Tu7J/Q
xkMNz0nxFxU0KV0ZkpySKUDnQssGlWErmCwxeb779QiaEnYJ/wJkJhQ+SsQksZt1
OiMIK6jla3t8zoWueOdnRtjrWzGJ61nCdysWS9IPtgcsoNCh8thr+cyaxFWrLPDb
gn0d6+dgEzUP194Y61UdJqxXBRsnl8gIWHuhQOv05ovAyh4n90JeGJXsHdQLeSk7
hWHgP6SifFkK4lbuMTt0PQBxQ6Scyk0AK1IWvxwK3Gt0vhDdhEX/zqHvS2+tzMua
lROhn63zcug8rXnV6/j2UaWAcOyu5yHUiUUzwG26CEmrma4P2V6csu577kulz4QY
4wOHovcoqW0bVlpeH0ur45Fp4TcLEgLeMzsGVXBbQsdMPUT+IGEdDTBn8pFXuwou
/Ef582J6aRHxtSR6HQR2i67Vrwev05h/ymic80gUnTA8AH9sNfrim+zw97EQb08J
pT86gpNklXsdZKvIOXPCuw3ig4vskGOu2usuU1t3/xoTULQRJ23TWhR1mc4iphkr
hY/vUBYjGKZff4eggPTfM33D4bkZWHHHFSFKCT3o+36lvvdzll7dTq6y2YlIpzzh
u9+3SVATYvCZkwRUiOxSmDv30P6GfAUCFscrilXvyeP7dE6bjUn+P6tKyrjhWPw2
zSN9caA8+dfqZdQctocs8naSAsHSyfmILn4uUP6MhNrMtoR+gVSOSxuBo1WKFcfj
+zNOpbrQ8PA8KY0OnmfjPcJh9Vi5h364FPdzr873A8RumrckKZsTfx/JVaukPdm5
oT8Mf7QroKhm3UQ7aCraB7UT8BX7uSaqVHsKH24i7yL1RuAF7P2dP00hIuCWLix5
z3CbOoRWd901Xz4BUaz5knB6BpwYc3Mmw/dWHoZCy0QcRNfmZQISyBBGT8GnHcw0
gNSnXDVwoM8Z9vvEN7IQLXCd6hYFfPnJo/3B69bwHJilY+y+hpld98W3z2oCoWMG
DwcolZka7aNW56RDKpdodkXAEh/PRSaLJALKav5wE6ReJA8zZlHDTVaEVYH8Fc41
E3ehzsbG6nvJTAstQfz7/l2vOf0DHFqiylx/eP5LeIdLp/FadfQ59z1L/3gVjUm2
U+r0ZiSa2LzW9z2gCjlDiwg0mTWnpYL504g7cuFTVN53WWfQREFrNn2ryPtWFQn7
VRdOtZ8T7UIDfLH4tdroq/kcKt9VqDsZGefNTQQmNvVVUdvPS1x6bcHRGbjDyPxM
twx/8fHLHEJR5sD2HU+HetH2UWoZX8Pp6cK4PUA+wVlg5k8E0FRyBtdiuQFWLrqG
uIp9PZTDDT+MBuN1rmmIv7jF3xkMXz9tnvJIIznKjHcekwG5iNgya9TG/Ir3A9ve
enSi6KA6qk/PfSSA5+jhCWRt4H1kvULy5pLlEWy2WT3JUuMueT1/gSCKK1ArpF7R
fmXJA/303mZvlW6pE6HR4THnViTp7d8PxleHX7VkgVGQ9xDQMPGTfenqlpwe+eRU
2OmHOSK6picwIAjmJiKrGD9SsY3DeG3y2KXWzp3TDzQBfBr/Of0pE7PwEfZztEwD
kibYR9wJEsKXrAs9QRalD0mXIiVCMYoKsUrBUCc15rzDNvWqRpJBHib8qkCKpdKE
njhtM0l5ryOSPW7m8gw2V8CqXMcI2gN3U8cCrcNY4bOxZQQ0D68oU8RVxVtd8vu+
R1EdGtbxkUtVwdrbzkVcxOclfLjVwelzPcWKESioIjjGichIik3MHeGlRbEsD6PS
wP95NWdgWVetE/ILd/VP//ss49b7MyNuQoPLzxG++YLTsDhGTW4QX43T+0wqjyAX
dkWlPGoNRdUVkpEmdxcnEzrG29Oow4garbEi2xFsMVW2peoL01H3zvhjGWzgmJPy
lkk4XfwRfRkGKX/UpOsN1hlcwyzeBoXYL4eAYToJ0tdZWOYo+8/d/QnQVE44RsVU
Uos11zI6CpAysz30o0wUCH52iHNooRCkSKUnj+beshUPdRYyHeEcrNVPVJKjNaiy
LSaasSTpKO4mjyOPJM7xkH239+Eh0W8S8ASltiX+1QTZeyZI7jAxl1sBNGiA9ne7
l9Q/WUFNkcDoBVBUCncuf/6t29WjBhEh8lVvjf1JNizLYveImh4c0Z4yykc3UxfJ
8gOzdZgYxUlk73wZ6vW72Y5My0fn66VS+yPWjt/9rEw6Ewlb8+CsDMMeFaQVrfch
ABb4DgHfyPW1duzE2rA0mXs8PlXPIwu7st4r/Wr2q01/mCzwR2mY2JQI9u20lOfS
tm78PM1aHVcpttBXrEed+SoCOavMJtQdj8W4sW4WBecr/reFtciYmwSz/zV3eRmy
yEX+nkDzC6/Md9DmwXEaNujfsDZukX710AYDwjOjqctY3A3j74EYQOFgMuSRYW7+
4OMqxx4+/P+VfJMfqtG/5sLz093sL1zRwzAcilh9CWVXlAfbijkDijqfmW+ggWqK
f/qzqvfgBS9sFfhSNMgEG08uwGyNyQ4NzhQMRfUfDo2rdVtYCNP2QIsPxDQ07J48
oGuo2agWc5zFL9VB22X5P62d3yPIVHeD4FpAQ9AXEmmMU40mWxGbt2OQh/da1tVL
HTHA0Z5rw2t5Jh4a6rNpcb6JGftN4LmIeyzuyfP6KgrsJwv3URnVJNqtRlPKaJwP
NpMH0HEaQvtmj5f3RNyWsbSr0mKINzOK9Ar5VgaVHT7mQrNAAL5EwI66/UByOyj5
XkMJLFNVEb+SYfmRsVgHauXatA3TQe33ZIuFbvOHQsaqrPDWdVmcvbsgLLF8y72U
xc9ZDzx8QdYX8ECqrHpynptXlMuage++dhgIRMdLWgB7ifpt+czVKwi3+Tz0zpg3
AuXhTae9ZSvk54sOTjBQoLQ6U6krePrLMPgmDipMp1GdzfPrnq7xDuCuixUc+9NZ
r2kLYeLEKLMArsitlBV0XAlDuKcQ6vcFbCzGt5JoJIYrO4MmZNRzQW0hfhLNgTH5
0oBf1tKbKTxltLOD65PyO9LWz3lKF4zqI81Urn5d2+OsqXKqc/SeiAfY6hdm9Nik
SIO0mu41ierZldBvsp+ZEd7/y7+CuH3h4r8Scx2rOJND2c9GRShna0j5Kz5moUPI
If7SaqdMy6DHNBCOSJFiLFJBS88JSDixWZcl4fHHCnypja1bOI7tGNEdZkhii5F1
NK9NCd2NMoVTDs9gNHi9joO0N7zgTn4VCxfxpolJj/V+IZVLZarPkooNonAOs2Lb
n+LSDAAAqpJglSJHsfsOMBOpTieOyfnh9EB2U69zvNQRv4N85HvFiRS4BR1km3wO
JkVIjEMllun9vgLhD5Ha7xM/NwR81tY2dvUaILlbNSbPJ4+3jbt57QBf1Uds90c4
fz67k65vLJMowWdGhs/ltaWrVeRdX6hUxRweA63pMo2TqZFfscXNO4al/fzoPkmJ
RXQekMCamjh0tyY/DMfVeygKJkMeViCaE3oxgYB1HrOGNiqgHqvtfTYYzfqDgvpJ
fSQn5dPEiE+PQvW2tkEfLpydxetfJ2QAqrDzZqZdqYrUmtgcAMVF06lotTUacHZS
VrzP2Vh8oW+PxDxP3Cj1QWxn6SR2N5jN/OFiixmAAeepLIa5Wbj4sePlaAzhuZuQ
FK9wroL93vTQddGE0CniLK0Dhkkb5tiVjqvA5VI+6lugyD1OK914x+YthZk/99tb
6J+MUXMd2DwdMKccmbRGmy03p9Ym2zbr42srIEScVHqCpHTqB8Wqv/qhQXIY5z2i
BU64kTr4Gl6v9Aklv9EYzdkdjRsB+hfwFeKe8ScUqliV+87cUdDXRI0ChxTG4SDl
Xw2a1Cvc9TXDjesJaFp73DstKfyKm3/LjQnHuHdNdh1cSsivf+NKVTjy12BXZZGZ
RdUAxGpao5oPdD8mcl9s+dqF/b2qXVQtQaB56LiDhrXk6BRnGl9z2T4LQgm93xB4
hmF8h89CRe6G8QfKwpr+LX0JK3bI9PDvlsmAYOkMZpqExJX6mz4zc0pENTNpY0jD
s0BYIxw0plucFxnn9qs98MHTg9wH73+/X7CS/Wn345eRI3SXG24AjT710AzPmcnM
ub7bAgr5zNR3z/7tvOiq6HOVS8JMxvlAVJlNqoiFhR9A3OqTwgIw6P3VK+Em/e3N
xPw7ayt6Jdb+yGja9byeJolNxxnS1fCC3Zf5svuCLLLmbs28eGlTTBTvE4cNVOz8
1bpb15f1j3b9Zpipt3sHriRHNvfTPpl/axkV110jQ8MxCVVOxsZ8k1VyY444Ewhl
gjcDkFKKV8QTWN+Fahlxkg6kMhyxNOZfpG8EH1EazzSCEp+O1D5JdO/t8fyG+ejs
t/x66CW1OaG45nJx4J2vLk0+10hS4LkS9itGgr6ctEISTFEB/F+9ldKrk88GAnWn
0FFv2ARHxk5h2hXSVT3/oeKo0+JUUdjDcs8QUhI5n+70JXaLM72WsYkRQVLGPVpV
iczi0P5IjLJFAwt26HGNIEX0RSPjiRWO8A43b1gmbMK+ZlHRFTqA/HRZVvyll7+A
BIUYRkI7ArqjMNME/TOsfw48qJJTBt8tbfFV2oh76LjAsjIeTh6zIvX0Co/IFdU+
bl3bp0Zi4rzDbmxj//HEaj94cmB1vnSvsfuomnz+40+OMJTmpMIkiPnVKgCLQjNf
BWicCKY2d6qpmntRXG0S5TljqdFjvSTjYZ0Nr+2UnXSeKB1XtMTKV9XWJQooQSeI
XY1+wwAi2CdCfcAuAmIEpMqnSA0MLDuw/97csvAEiUAwq0SIFAnHt9BsaxOK1aoN
eoslkBV1KHgBCwmie5TECAC1jsDKjBDnDlMlGKQwbT6qKgRj01l/qxJO7DQ0ubcs
kJiTFWR9EIf+OT2x+mOQQwe6kajRtIRLIf+RvM7m4Fuld78ehpPjWbl9r5RAWjRS
SnUN6tmrHOU+LpvD2ND7ZDHHkUWUS5mZy2fDWXLvo90gFNw6DLhlUcZLssasTggV
bMqgD6mNO8SZR1rx94OHv433AFsXz+nD60QcnLzTvu6+81RPEM6uT6+Jyd3zZWfM
57+O7NUCQXVO6lHvwbmcyqsoGcz/rzf7jhDtTq9doHXXfMTekFhEltlGQHSxJQ0/
TWFZ2Bxqde4YYAco/aqdMc4GiSsQ9HByha5/UUxXrpLToFP9tsanY0T92XWFfVil
Q+S7hFZkX+u35Pa4/z9ELYzJDurs7OY16GsD8/F/5adFdEU0a6/1i+Sb3cMKwh8m
WFhr6zj9WOth0eK79qiobuvlFZCm1x2XIEg7FuebgPWGj9KVkaRmsDRDZ794hajh
kETnI1qWkIsWhhQeGVhh8sGUZKGak/i0iT0PkEmYjYGMVj7SkKMkJSiTd4OiN0t5
+Mf2lzz8En5VFontYHIAzfCrMmTF9EM+F4J8/ekb7C2dCNGZR73uf/IdZMwE9Bnq
WYCBtVcWSrkCM+ZpJYpsx/USLE7ce7zMsN8t09AeftzgPrEBiY7CvI4wm7qxBwfy
6JLBlVKYpzJ/2ByEVW6Am77VxILqbZP8znLhtqkr6fMWR2oTD3DDjnVgbIOGK/zR
3l3h/HyrI4ipA6B6tTim1eX++D/skXg+MSdeoytljz4Ip7eB5WjWRP0v9nf1oiC3
TZKYtl1KbjOczd1V0r1L6JCtVwk34tyVS8XWDNq12zymBdhhdxo5OrwKC2lGWtHP
J/QoPVNM/aLnC+MFVvh/QYleqK1842vl71MLMpsQ92v5lBNxZTdz9LMe/r5qWYvz
nU9I9ooefroEAYRU51TMUvQ4XZn1/jOwLmNDQM86xnSCKyj9sjWWQJr/YcK4LHfO
0Y3OBz3iOWybpTDXkOBT7qgbmqO4g9rfNLt56mcP00rtTUKuRqK5H82y1sUul1Gs
oC+KBK4psUJFQRjKdHSX/fNUqrseoj1S3jeLuj2WunRq2BZplPxte+uRSz1HL+9R
PSfNDrKZWtUCHg9g/437u2QT42KQktBU2dgZzbbneHtMCggYemi4UXsUI7FHfdTg
pZXR8/SsAQ7Z/IkZo0CMr/5u6P12ln7Hu4knQRX6LP4EAHsOvDH/PrrCHRVmCuvp
X9WYeLCHmqO5yuRtYiBhP1sNlrnUfwFr+IcthBZAIPnW8zlK7I8+nUPtSvUbYlck
TYOUKlIOdIM8ejhb+582TBLRpziee8+1LYSFv1wFUBp6e1kIzGVMek3zqOlNG5Mw
DkFrymnd/zxsmkv3/BvPIfYHc2kfVUeFe1ayUFp83T8oZC7te6U42m9y01Fwdbea
Sdn0hXZ1xcVMlb+F9NDca5Ph9OrNqg5zHadZguGSy8bRabXQ85yVZ6aWFryOBBLW
BEIiBJsxTUxBfmR7jSZITIG83tAX9rr0C8ZKkp9oRQH+ZBucLVb54AuRJ+LQf3h4
KZbMLq041mbZih7P9ckVeomDKVVJWaBhYcvZllzz7YhG2xslI24MJrlTvYBwmOEw
IS25BAggmbxssjOKGrMAdBA64+SrbWohEDK11jY7weqtkb69/711x/wTNuwzRFaA
0aJtQdifhdAYunJGdtClciFRv8VwMfT6DhEShxo1NsQ7DwCed+Vd1TjwWXaRQCkC
BKDk204mpzWg0xGapR1eQEJyQTCiBNshHf/LKoHeS0njS0d82YlnsRgePN4ltxHK
PvFJd/gL44ulTSNMk+5QbuACe3cfSL9XkjxWC/ny9pf4WZNVcaNntZZEzhmC2JxU
YabrM8nq6Fajvavtk0kFQhHYfAFhnU/S+hhnJIAaiuXIq0LXZ71aDzRPhYqI7kkC
+O7+t4coYtoYuUt1YHPdV4PSL9biXdEOKWlvwlNd32ISi5tnlTtW9b11hNWIdAHQ
BFKMdbndvxp2lo5coXMYGvGxArcvoEcFh447g58+gUx+cEtafdpy8jCJ+XGOAcMW
eOlbBbu6XbpuRlcrL5Wl3o2XtYCsr1BUBKx2GEqlt1stzH6oYvS1z8AURJEZ5rNY
V7BfoKMhim//lKrASHvC1wrG7jDrG+2uyx22vICgws+CbPcXuYYTjH0WbzsBo9lH
z3Xl4jjaG0VZ0SZayDaKmFS5BcST6ghAId7/qgV7oB59vpOGVR+5mwvvXYlzYaOK
UdMlWgO7oKknODUEqOMXQ0pZdSRqZMmKMY+lnShMJqC/APx4Ptek3ooxtkEPcSE2
LOhla4lr4nP/a5+QHz1ECstWSDMwOTgVvp0yjT0Cjen5/ecN5y8EB90kx/fEW5y0
Z+mOjvzYGLlNbR7KSJFrqUxzyfk7Adsv2mwQHTEe/auOU1H0odL7a/hN5+WzCpQi
pSTxIAAWb0vMovXYanvatctbgaCHNccLo8Io4PU64uZrUQFNYwFI02xFM15psgfy
JD45ReMLQqT2NicTjtPxM1cr/+sYjdMS1i35Ga0ns2hIEbjH6YuoqCl+wJqIaysy
XfSgChyGcFRKlqFDUF7PV3PkjX/EyK1B8cj2V/reqvLNGazS6aHMFQ+rWt9xwbv6
mAtAbvuRKM8fyOjUWhX0or30Zn5hUYp5BgZeQclxN9RKz/n6LHkYcctnZD4ibimW
A50gR64VyRjtqpvvP+oKvAA1Bwjwn9jjigbw549Av9Ga0FuxC2276kIe69qVbezy
1YiAiWUFt2HhtwuDNp7stlgSBqrZrb80gi+zIIhxDE7geLI+vIgmf8Ogqa8PEiUF
CFK8Qa5vV89OuEf9gV4niY/Ak7U0Teez01RUqkLCIn0d94m4HoTf/T8HrgA5sTKd
fIlALVMDRwn8Nexe4gzk8GfChR4b22v5pLdniNsRCjmdKVoQm6x5sHTdpPzg8SnV
4cC8UB0cPCiH/eM0oQK+jsHsC0Is7jJ7NNGr6DgIa58lj1Q9zLltwjty5gBh5U8E
zZFcubsMyveOE3lp/Odo7NrjWUW0HPKKyxwXgogYZnNrkabMwMSDUrmbC3tFONLD
vZnAZYPhLo7IIxcl2YykY2ngDHxaVzSYqN6uQ9LaDaNIFgEWWELSO1waiPElS7U9
ZAs8wx1s5zIggd4ZOCeknDo4ZwOTVRkZvYJmxj422DDKI84Rc2z5R0igX4whZAfQ
kC4vk2c5cDeFkLqfhe73Tbft+jERBKtZYsMuckTpgXbbFkSeB7LfLYQKwoolgKgF
a3C072YZ5EJnNsexOk+w4HflCNPCocQbx5K+8tIijNkJuFPun1H8qR6Xq+OnEJaI
9YUi8lIyEu/d/diKQ/i+fxcTRwR+WSltvtfmP39bDT0bgodUhuDUlK0EaqAnUtv6
yjQMY/Wyro9C1csHPTg4LAXOBbfYpyFn+vxQUwU8BqyNuB+Y7ulc2NK+tBgl3KoX
CPFZXFmtY9lCGWumg1OkL7HwLwrsMV+n48/5MLN2rWB4JdHzHhQxIo+qRvqfAb/e
22MW5R3hjXdDlEBraOI+8hQfP2ppbNhLI86+20P+Z/BfZBhvlA98ptMmC6pNw/j9
8rM47o9XD7asV0PydXy8POs1FOyhM3YcOMWqEegEInFwiLZsaeM0He5rEGc5hSIe
jLcoyPNXu0NaW/7PJg8fGEeYs+VltLDNMocfhgGED+I54vXX4D9h66mJ0p6QV/Ro
MToBjDGMpkUAIsM8+yDE60zWAm/WI/QKvMSz2YJ0ByH772BMugJvWyrIP+A0O3mF
rG4+PxWT3Ir8OFfPQxjQRaOmHDAvjFCvAC+oPCAWhCdop66WobsjNGRwsT+EaMAR
QVVNYwt3X/9cgZU6sY3EF9jxTy4ke91krqAtLYSPPO6LS5lafuwoY8r109PGF+eK
kVovpsRaktTvyFTkvkR1frWHLHx1n6yziN2GNF3alX2pZk2Gg3IG3kgfdSCCBo2m
YxHjCEiMm7TKasfYXPSK5AxgqZ8RTR0yIuHG4uldPg1E1UK1wzvfbvzWTXsgSXPF
OOZI6O4mssJkchlnBKfABaRUIeLNvypUp74VldpEUCN6Zt1mGsOZ8+mtazymY+ns
qq7Ml1CVI0bF+wpcXVzixsyvAbNVHURvGUPiDXbfjkqekAC/4h9tcVNS9WeQrbLb
/OQz48mA9FR721wEYBJXjc4+DVSQfALV3RD4lqSjl5B9v3YEu9+3RHj2M6/0c5JE
ywk4tWyCKxDcLsGHZjGkGpDtd0I30u8RX/4ObdGv/Q7jlmLzbPrST5Czivvk1+28
pXUDGx6aY2Ht3YZjxRCznQEZefZCf8WyY6YUEKNECMuMxKY5lJNvyBFoMrU6ef8t
z3V/eQdmtYixxqOu3EbyvOYbS3DMD3hsZXqpbkyMXKhL919KVoWhBBq/ZzRenQdz
YUhg2aZHmMfzDwhN4fcDrO3+XHORsYIjlQB5pZL/+4qiM7P/I5wVp5czPI5FUtnZ
FES8iabCpgYZZDktup7BSoCxIOEkWUhUnMzGnxmpNVpTXNMRKyMn9qMptpTTUthz
dW5h9trPRuwE8XJzyTt/FHoUow3ekSFd6jdw0RYebu1V5VMicwpzA6RMscLYTnYb
Uj3CmosC5C//JLP9T555Srr/kcZosyWEJ4Vcdw2BijANnj6oYNabYk7IT5+VbuqS
yVEZv9GZj8xpME+Q0A54iX+GD9WVh3/ZJQSOXdfhgG8/dXiRqJAqDoxc2/SUkH9Z
KPalW+gVwVf+vrRyyiJyTYMKy0Y8m2HP4rjVnuQvegxMg9mtYHSSwfdQiljvnfHA
OrJ1XYvwIZdWubB4bvTb8qh2e9ZE0L+f9glsshCLEIxevpF4SHjYC7isjBA149s1
7ZV2H5a1xTaafPwFP52H9Pikg4czRvQE2c5VpBdJDsm042pxaQtrjyjDqBF78/t6
Etskk8/8XbNn55GCObM20CqD8OglCZKNPEpfxWph0uvwh60Qr54r+HR4XolBO7p8
Uef1TDRuXTWNkSlt3Zb51kFq/ERy84Fs+LAyl+lQ1g5yU2TkSBUCKXRRz5njl+lr
1bIXaiy25fQllHTb8usFH1DcjQCchjKg1TOqFYXiHmiy8c0FLRGiW559mu1GrNa3
lsoLpCLPb5bPPAPeOafr0JVwC/iVh88iZ+JMOkwrGH5cZ7HrzEJHR+MuyxbMebZi
RfbQJ66HAKl+YwmNZgYxO8mY8NMLmDR9kYbPyJDWCMsMA6ciPMSW+UYiSWVynV5u
NQfJPiWAPWSu/Ia3fIZv5wxPT+tld57vjw99Y2ZhOGDbHo/IuDbXxRvqo9o/GlZw
iTii9LGTRoQhFrQ8N2iEywYcouBECvjU/1PyF6O7PBNAXK+U6nB6y0ffvXkrWw9X
yBeRJJmBw5mXPMoUnYf5NB5yEHd4BcIJUClXldpdZdn2UR1v2Ze+bdVjKCpyz7hP
nUCVbwX/qOKZh6cb2cZwrmwbcB62bOBy0aOD3zB+OGralnlbv1MCk9ITcAQLkXrX
aEU7BV78PzVoapcqWIVg+sog18X+wGAVYDQFtUFac5J1MYPENJ/yHSeLrn39dTEG
9SulzvbvUqi3/Dn8oGvq/Bf769L2tL+eYuUN4lsyZ7HMvKq5PiR8lHEjYEKnFUZR
dHzSvSILHnN9NXMzKX3MCUWDuZUyXW6jwKd33/g5i1Nym+S+tfzPVz21A09PpeXk
F0iumU6QdVuGcJ8Psuw/CNGlgJG6hueq7u4oBKourrutok26/9CSEFxZ5Mmde2eC
znfCvJmsWfMbkEIoo00DxQ5YIgB1HKaJxGfWgYG34d7aUzIaZ0Ec7ECrv160fjSa
sxUR8c4vnY7ctA8ElhIxHHqv+gM7FJHmt8fcxfl/aeh8WN1igt1vCRsyucrG9KAi
VNAOlStuIBDzp6S1c6VH0yq+Au7OExVBaTT9PGVVpJ3NO4DLLegxo3jhPFyEt3Af
m3OsMaWHzFHlYKQNHXOtJG2rTG9HdNmVaiaH+nPGasNXKEdYIgXQm24DF9lY7kVd
Ir87r6po73LsKkFo1vrGDsjtgYhYakMkPPkvpjorh1qynXJg3Da5hE/tWB4ZXkSv
wRPTDYyx0i2zuzc4KzsRYg/ObVS30rHbwShcQf/NaQtg33i9dFLVLrmmicdrpQcm
0rM+cpOKXK7/a9meBhLrxkYrF68iLxAGlBzZ6QaPlKeJOgfGcYCpw3+8m9WXZIFR
r1tgNkAhrXlIjbV25XKOILQCgVj48gkqKttFYyYSetNQ0i5q36llFjv93AkyRFFG
LYbs1OauBUZSSA2C+DMaSdB1uRAN5RTu7tvdwiLMYX81cvcAfHfJW2T/yYbi9/SU
AotVCJVgtqSzZJCq+nBuTP3uNFa1MPG5zJioBKxfzNnhKXviRQzvGNHQg4htl/71
1GUCVkbeOe+4/Y1pQ2+ev2NykWvI2y69yJlzwdhHFifrDa85bNH0IO1mGt0bTBeF
ymAEdwdxPmGotN3RoLMt1H7IeAmo4WfsXtwXnNl5QXdzXQRwe82lfgkEq6dBfld0
EBiVbL+7Ak3lNmoetZjubfab3B/2vGEpVJjS5acErVkemFlKyewnufQR0F7nHhG+
GStOQMztq7Bb9FW+UhxAwTmmO1Lz81buTSWhsQnbX/U/EijNcZLE6JL729MwQaSG
18PCOk7zgbI+OIwSF0o9BBAJTQ0AsmrHLQzosv3bHbYWhLGCdrMLw4vr0KBtdrUa
dVpkqmOUP8fOVoCpbWYndAOEnTfw8YBe3MQpCt/08Dp2wLG32BDr1N/U5tyfiOKT
hq7n5POGvEOdgbKbS9RWoZlGZU5Eoco4vB7CtCI2doGL+hZIR7W09mWg0IULK9rj
b6lpdDemHK7Xd13VSXSDDJG76p3sFAUTz4RNtzm/3dFTRjZ8A4THpRiyRU24jRzg
aH1OUi7i5g+DIH4pYxglb2qwzGf1KDKXGHM1CTITQ+0ivnsw/CdGF1cDk4/Ls9/c
z+bjTpuXZy2mDvt/Vbx21KzA6LQTRAtV0HHoWlT/YxCFMHrCJA2l1qZ6nR4jz1Zl
O/qOki7Jiabt5WFetD/xNhWMdUbxuqi61pionzGIke6xZvhA50UBSLdv0dY3jbLc
7J5hrICRSO5yt5A7lqooYfTC3CTdHLEY+otfX+5znvbbMG1x00IZ03j7AjLb4qtP
ldmJ2ijt3PGL7DSvPhsKNV1X/2IxMXZNkAFJE/ABkHLoIugJTBGiy06HEepLmgl7
GqpHy77ExzLFuyQQtezUq9AGHXFpMk7NZ8OhyjhFLF/pZ6L4ay8eaxuTolkpmTRg
hC0J0SEP3M6dC+29U77trJaBkDjDTRuJzID1Iw4DGj5EaK1b17BjfoED2OvLKf1A
HlOibDYJ1WKK9xUnDFUySewvQZPlc28mGmbvTjxWlH6ufmQUkwyssd/DlM69Ze9E
hfDp+rQNP6iqNvwVpYh2oBm+wBWu39iBWUi38nJmlQtXv31GiDpRKxR9hAZd9JIu
6vgDDCbdd1idRbYzt4gO2Er7IgizvknSyBUQImfUpO0TPGPRer6yMQDvh+kaIWqD
sAEeu9BTY6IRj63YWe6VodhO0b+ox94WtrhTavT5IjQKP+YaJLuousjXArF5Vi/i
XlKMVukTOK4PEhWNYM3sggRw5w28kQ16Zd2CUS2HRw2N43J7PYShbxvHAiOFqF8p
VUBwOKX12InhbvH70lwLKziYBfMJBrk7ivKyx4h19zGO/Hw5bMbZcCDGcCXwh8Jh
SuMQgvpT75C41J44kjUG6tjxLjOj/JxehbPCgCTvJcz8S4eYS3h0ceyJ8qdHzyhe
36EFxYSXT24KRlb1sDbh9ATC+uY7w+Ynir4fDhIpwhrR0u+CXxD3cHAFm2MTafdA
DKCiSFZAb0QUMsajBfZmebVVAMhQsXFCgc/DHibU8g5lJiWIQbM3XOD3av9Napu2
JI5pP27PdUJSNwTkX8EAMcJXGuJjeW34RA8JMhGHXVhe+IreQc65E7EZRPoi2x3y
+A+eN9y466YueJu2d4wUJBTWyXpwzSoX28y9kPtnQSpF23wa1M5kIsQfQWl6Zi0X
FLFLfX6kvwbpxuCbYy90yWrJRQgsZ2LITGT4ZpCbbX8MCgI78YpxJrQBM3nxh/Ad
M5kI0ZTp6HaZ+oJ5bGSJcEpf/ghNnFIZyl5U5fnbCf1e/RxJIzBTbvNyoCyLqK2g
GMBoaHhWcQQ/8MJiBOPF/4g4dm6Lhtj55ksKAZsqMO26gzrZzPKPg4aDnrOb6XKk
haPy1/wg2NLLNiY20YnVpmuOezrDiwLI+yAZHbBJ++5aN3cPIordrdVYU68W6Jtr
skg+TeWOuoW5AO/k1HRl2pE4j+8uzuwTyJrwZcItZpGPYX9jVt9lDtaQAGfXZma8
IWPNOHJt2k1pxr2DdNm0QfE6+8rroP7/7wTjx/WgbhNcQeT8cQGj+FCTBIZpBKCw
+j22676kvCaijiN2ut4VCqKtrfOaqF9fy+QZby/eiFDn4+cUcFS/TqqnuhyH22E2
azJFUkfpQ9WvsLPOD3X+npbsYjE3y5ZRlZsqfxGOyF4JiGUMmkRPGsEalO+gF/UO
E1NqKhGKWg/Alnlz0opsSPUdR9LsnmU6UF2zjhEfdP0Ilo06o3Q1akG/g3m3Sbmb
Ycym5bk6HAkpOcgkooiPb3C0NUJdUDS0USv+egKwBQn1Li3WBm7MoCuJLhOVZMgc
eQxpr+ej3fJLIYmFH5OaK9zaOhAhOT6jkhw0kV8xivsuiFJGeRM0/zamhzZCxJ1p
AUG0+0ys+blSBsFrqLnMAvdcDyh1RC8s47/4DTbJ4uKdVN8Be66vOTcSliMMhVoo
A+pimtSDAViErm+2y0oa+b3J7rJiJez+vErvGvkMn0WZW7DHuR9BpJRUayWHGxXQ
56o4F13ad2FPikTzrexxUsWRB/Jlb8YRHFCU83DVLZMQA81KFANRC17VJ3Ntsxnt
UprGxBR0BX73HA/5yf2ZDB83ifOXT2mDM2GDQVt3FVEHua1bXrs+JgoVH5OG8i29
foA1U0WT3Gaz4DKzpUoc3YqdOyLxqUZ4mtXQhKZj6gCixKK2skqmCWXIHX+zpZnF
Je2bgn4aZYUvmfsw5u666B9GzHAZ5gKjxdKAdTsKIuDmJTQk57iV8NJDyBgwI7CP
lcZILiByGM+/tRRlcPyS/EcPO3i3OeFl5Vvl0Flw0ADrSgllrUzf9/2u7hxVO4hu
KgqDcgulfGk1PGp4qdySwutt+wHxTMCuRAyOOhXQyYxRQNZObj+FtPap8XYVSx85
CDdgUq2TCS1U802L0y91MOsZ+cdYL9palzP33ltQ4f7FNRU8xZ7mvTauZkx0buvR
29b9okVx05yDiwa5okQrhBdJuDKvFv/hBuU4hYUINgATMYzsBmAv+I006uKYClyI
sOASUIYQRl/nQS/9D273O/a4E8QRpWTqwj/YVuBRAQ7V3fprSPVM1I3uVjqn0zN9
XGSWiLsKECkKfNaETeaayz6FUBT4DdH1JnKaqwE+LGxqtzRne8Lug1W85pnHdM2X
DedAvFkBVc8a1hxw/OunO0Wt+S0oqBY6VlR6OmAojmFqZq58OLJ6gIRa3tq4rgwz
Gv7ZFnUix9VZ2+AE+wqdMEzpURt4ntC14GVkQFkwHgzOna5RIHlhsKGGOMVW3biW
y84TWSa4GjLbmqOQjnOnzFxkoCWL20pddKYpkzqvOuNi2DlOgRXef+3xLcSmIwO3
I8b7BpAepBF+6OIdjXoo3LC88y7vjPu2CnltGz/tnYXjZkn7YKyISuw3QmA3+5tb
NGWJO4vqkYTwI1Zmzbyb6ARdZJctDju6U+Md43Xy91McxHM//apELaiGaBO2V/2c
0rR5e6urpknNzemj7ie3YvyBwHwJeryiQ70ZhzypUJLVg50o/vjRUSyyaf7yzuHa
JJ3Kn7ja3UN4xzjrKymVlidU30NyiMqm9Tf/N+bWLOobCBApP9sQB1LJuR1iDNt4
OO4pIXBRx1xzNcDJy/Vl0cP/Fiq3boAQ8ChISVtyCvE0FxGbm+bTyf1BRAJ1J++a
ET7CnuyJ/Ubp3sGKrlqvEUQksBO5z3VPd//GiJ9U/4G2HbK+a++66dfN4IPNxqDu
w0Ef9AwnMDA2tOMiwELGzYmDq+iQ8EuH+SVrFg1WI1aCmz35wstOgvXkK/mvXY4I
MbPkwTFxEq3yf1sw7wn1Oows4c7MiCI/g9bIFncCaqDBmWLdpCht8BkDbbEWtb/i
1vOxTgV5RYU0XCqdr7/yiOAUCHkaKINlgd++p6sDBGOHjqIo+eYo1Hn/eu9qQeM8
HCu/dqE4D9GoNuFd8L3ot2L0x70zmA/Xkmj92DMK8glbKQOgdYfoUG4LHxXMA6eP
o1s+kdVSMUJvt+F37EIyOO1Ya+wciekzDGUDYB/AKf7LjoVTxE+1p/0uF0kKKxyI
kUA3FY7RljEb9fKyoYBLvGOGxeL4iBfP1Bfsfizp8/BOzmHeBGJOJLz7+q4t1A8d
SHRmFImrX/r1USL1iHj2IRmehliaS17Aae2C5/0qyEwMyv67jjUtbu0ImO/GtUfG
dvw/mIeH5jZNJKTUQWXtO71iQmQir0a3lrvlTyedf1Mt5BwRhLaBP1ECSIn7xkbM
tl+LqFwoIiSN6utI4AeIlx0w2Wnbscw8ajxX2omY7ouDXlUefIOZBUwgYyHt57vf
88DX9BS6kqBSw/4O6kHLm15vy9Q3ZlV0PTJnbrhPuncm9RIHJwgX2vmW40qPdc28
uyEq8wLNwFsawdmFgzebpkENz/WZXd0HeT6lXN4UGIlOyV/P9ufthYrYIfQbgxrN
vswN71pHyDa4Exdx7VzKzuWc5C2rz28FIES6FvkUoi7BS5n7n5qRYOft6i6Pbxaq
uzjI9xGlolXjDw1uxMlmdTrpFVRl1OnErzteSYfNXcMJUn973DJimCR3TCEMZ73D
o3dPyrc8dosVZj9M0/JjdXToVC2Rwvi5T3g3W8z2y/Fcf8KvFZMUhPL2GGKWHAeN
sE69EjdOkaHArfVs61mgFjr1BcxuGguCWuNoBIuEs61qbqW8/qmmOn/GIEVqHx00
akMGrts4RtC04UpnvazeFhr9nweJCBPHa0ZiAdzqklGqBJHoIkVR8O0OVni1QKmo
PovQjEnsjMmjzmQsztvXmLpUY8CtphlP+N1RYbjHy2fTmruGO1WgDE0pFMm7GikC
Zg1ugbFUL6JbxdJ6+s8Q87TwG6x+JJBHyBsJT3e24RKj4oU9DL5DwUuYgZGD42x0
UJ2YD5Cxyy/I5X6n8uMYh0X6wcma2qyLH6piQjJsMjxgP/hzXcyQ3kD9CvN6CQ7B
DvSI/279CRxAK8q2XOf2QJl2BdIHF+Y57SuXumPFDfxeeXUmujPMvuQntLxj/6N1
+/utgvz6SF57ZmgWINXxQyhyaJp/LG0X/ProJxunuXNYth2Y0jL4SOsOBHH9NMBe
lTH1GKbdSd/u6KXupbiA8JlMaEPZxAitrT9vv0IP4bdNYy2Kior1sWdH1ek7h/2p
/zkeuAgNCVBMhqe3dedW/Um3ZVGx/lLoisAukQLQkd0oLghWsKulCZVzZnvBPEDx
XKc1Tr+KHzUn0FlwUB89/GNZTSI/ALyYgxDlbrQ1+fy5Y7c6LmF5CqxVuXhcNzIb
n60NglUGwLKSS1QSw48IAAIDSAF+71uTfuwU5YE/dfKzEeLP/TPbiuK/VdMTd+fD
+82FYbpu7gF1Nxl9CfE1xhlLd1TPKwZGeMGPVM3Ap2d/fcOlbIs7t3WLnDc/lxjo
bxpE9BY6f3Y+5xQZd84JMM6wWZOegiDnalxRL/w7nd49R4rcqLR6G61AuyrpxIpc
GTledSowo+XaSBNpEXY/fWHFw/bYw+83171PYPT+dv9DcHC3iaeki2696+750JQO
1lgNX78VOcVSmcEEiaq2OX9/nkrdxAmgwCD/B/BtOicnIvAVpgLEF5pA83NM19vd
vgnQnYB6th6WNbMzuA0Puo06Mk9iICIFBp5t4S+fl+7G7WdrVA9bBMhtMgjP2JaX
LyD1c8sfSzi/69/B7S2Zf2BVbroCYDzYHIvL/XzODPn9NH9y0yCsa9ai7MiMh4ln
8SFr7ZK5gFKbNLwU7BlfId7+T0SSBR/IOAYHLKdB6tPPS+Fv7fs7t44LV8xVIgmr
1eh467xkzsfWLQTGynmF+c/BTpvRIrpE+3ZoSyByrTDr20BDogONKrGl4N2pJpfX
NbeRoSiIqnIvsPGa2qUzjzKTcsAQgsJgErE5TOzMr5PU1++l8nXDQs6UF31C4CEN
zaMPmdORwHgasyxa4HD19jHP2rhDXw5d1plCt+X4Qdhsl/G8rA/mjWTkZs8G9LLe
H8DRZc4HmB0YbrIKSlje7UzVwsf7yuW4vgq6JM+dNaguoxhxZwnUhYKBfj7Esrwv
qdto0ZYUqXWuEGK1nGCEC2Qa7qiMrmIkiJHcghpaiqSdxpirjSWyf6g4WjYAo5ho
BcCBIMUx3VDMQm888JXPXDLP/lgcKlFMOyIOwCqDD72TrTeqpZDUcSa5h2ObN7V+
FF31BBLyadguGxd0XAnoLSbShjvj/vhr9yAI0hQq5lnnd5rVs5BcNFEx73+65lYm
Lp/Da6Z3meWa01JpAWaZ5BL45muJLTYPI1GHf64FuAFAaxwgFEIfx6TMCeWBpMnx
vBuFadWcYvpk7MSVJh+iKhaOWdPBEqi92SyeQztuPqziH8V7492rdXNeLo/HEeYN
98es/AY4qw/rYhoxXvXLHaLiOWalscjOiEqASkhFADIok8B7bt4sFzKXN6Ma9HnD
OzKkKVm300GsoFjIZHDL/csnLps9oNebNsbBlgS8nLuROatlYsepOAznntsAGz/E
0gKVYqIa0M6gtPcqdT0b7BscHKsuDeWdU5r2rEjY4PAbWhqyf0QiU+uLoqgYSDnk
AAckiU4aQ+o4w8Z/zTEe4RrCcmnYIOmXzoKT92PULZaLSNAyCjA/yOEvQUTY/iOO
4lMqUlSo/DCXXxPfHnakCvklDqO/Ye2fecKy+t39Q1yrJpKi3I7uktMsRSCXz4SF
X3FJZ3o2ntYpmqVPxmGg7Bgh4YeYvbMvS/vvO8DB/KQeVwL30WVxR+opVUjzCRVb
t7wiRH5pdXe9BDx1sw7A3qkeBJ69pZ5mTesdakz14zg4rknJz4IwCsFCP88B1r9s
gMZOYE4QKXuuX2rL80XUqVgvdb6hVH4kukuokSW6YXn4jAfori1fdgkVB9n1pp5i
sBRuZe0J3GY5vrYmWY+xTkVtgSTK6R3fHlt6goNt5pqJKK/IDs822tH01MJY49Co
2n2VtpzpCxULj8Lf++dFX+GLawrYLbD3DMxK7Qy/W+EJDWwY4qb/m+CAbWPotXNG
AzzddG0NzjvxcMDXjhJMXhnCEwNUC+77I5CRv+PvKvcq7ofcIMwPn25ySrS+h3rk
SbFqeitxQsGPBGWOMyQaUIcqf3Q5DfG4bN/LVQihqWEOW9p7tP55LA6p8dglu03W
YaolRrg7M/5zBBBAHHfgwIs+Li9mlR57HHN8MkbP+WYfC9cOdG0TPAyiBlXeNptK
5/UJ0Os3rsZGG4xtTgyLAhc/SHuVoZm6t5zBihFcsZ/k6UZvTtVj6oLP3UD7/C3V
G9fAV1SAcd9CyPk1KJ7G4nUK9fDZHh2V4o3OFqhysZB3XZhETurFH+ivaxK3bpMH
zQLZ/59IyLY2YGVKdap2rrlVfOYtGfk7H/jNLzH8gkRt15xDduPqZ4ljifdibGnG
zMVMWBaxwQcqeC9rWlfVQGaRcUxV4h+Q/dc3FxrDq+iIPhw6gfJmkCPsVCO4pnZ/
bKBibg2gOT5B2YRlwBYpviPDImLu/07+lUfP8KbEoAzvnyIHoDUCQEmNb2xYYilZ
+i9SXSAHkfDxIpqcuml/+B55MtFVBP73XD2Y+D5e9BSIIfD9OOzMZ/0n6aRZ1tYf
1738TgLhBgdGe06WX+zIkiL7rcknhFvhyCfdvQpAZbkBXS5s30m8tEQXJQWKbeI+
MoCapkfZ5N0uVwnev1TcgnmUihicE0xk4rOzQI7s6zImrlPvLyjyMmdyIqCUo5L5
36AfxfgcTot1pzlbUvPbvA1cd+HPLkSaxRaQuFBGkRn4wbc584jryPe8SkKJklSs
bjT6a84cFGfBphuJ0r5vIl3nRbzed6rEz1JweaDDrht//n627IusDLGJGrppO6IQ
cXeJXSciZYv1DkBG3fQxpfVTbbp+rZvpGNlA65HF7b3XYugkpjqJdmJVSOaLqeHj
XcTZato743ugoLSpnt4OY1mpg7sfp3qUZFZY+d5+vU0cTZcsNiGISXKsgnnNyF/v
KC/BCPVJL9nhUv25W2hHMlsRvzhcNsEdHnwGhqq70SbnGRlT5pIQrovnOIhMxOsA
dg0Vus+ETJmkDA/ZtJNwOKpX9U8thoCxoPnQaq15aPv+PbZD3b7H28q7D9sQpz1w
PlINs+xyoivTpbA9Vxr+kb1w5bVwZFIpoIzdhc+rfLejjv0MkWFqvkmR8WJ/QCDC
AX9MgbYylOOQBwBcV3R9FPQ0ybEA9nuPFFFpEl4N9M5HrX9V31jgvc/I2PkOBIco
ykLNeOAXp1FK9KzqDA8dhUHjlRoJnekQnmbmow7bF2ivhAr8q2R645NInnk6nmcl
K+AKLQU55NAW/RU6cux4t2apghMAwZ7K6jzPI5ovAl9G7UYpgTGuG8KNDC4ZrJ2v
zatQzKHZbsXoobuJSoj/wTEM7osauqNixTPKvcwsPcCo/NdMbmigIh3M+OYejkK1
t0Q1nh/2sbkU6/KzNjTuPpyIe8Jjff1H9ZYyXjf0lZwo9P3la/h2L3F046wCPiBS
MFJ3UuVobdPWdcjaNtkeDywjeHvMlGI2NEoQf4JlsZiUPaH4PL/QxniBDZ87CW+C
JveZcNMG/5jJVnyFIWpO3tHaXv9kCn1phrxEMOMSuG5ljMlvGOdU0c3NUa/Nhxar
0mcm3+PfamFXwEGsvkPQVCd+hRvEca1Ibgy5DcqXHvmtxhwubVFwe86iohpO8Ele
RAvtDIzyTa4jHBVHmGxciLmAUIyhSgs064obIVGw9wQ+fPKq8UX24F26ydlPDN6C
qkz7xpWjdlZfeN8nr55lXj4gzmXg7SyemQtYhX3FyMrRixVxaQ/u90tTFPk9AocW
cdeVlcUEKkFZkfzh3NvYs7UF+YTGU8guEvHecqbhP92mmYiAdowQ2qy8Tc/yIulJ
h25urLsTNcsC09SgT1GDlTpXfnRaWSg4Uy55LclDvpXhIauVr4Kbb3COXZatt3K2
r3lRpbBdtxdfNH/8nRwKverXYrIoYrAIj83QqDTv54GeH24w/Gzm3RGJCO5vydWI
olJa5p94tMQ49N4Y3Z5CheBLfXz96TG46QcuEkoxTbO08x2go/YsXWu47ywtTtcB
KOXrweQ5UrQ9nDRZISn5+W72j+y5xxJ2xYK6bXb97HfP/dUZq5MLxB8MdTTmtshI
9BhTwUM/Q9HLGw3Rwuh8qh0s7CCD4iJUQ7jl2/HVBwNbwPtveQq1PzG7d3WZhZhm
uUGIto1tCcQFWM6NZn7D5p6njthkDxKb28maPa1vcmGAtSwuejCQ/WGjOpO2p/mG
JR4KLFpHK9V9Y/i+/x/KN8Zj9cIMKDaXtDN4GHGO+tcmMOq+h0GYk556oiW6D8tb
5ks905c8Qk0KaADHyUSjz146y9I5T9jeteyljGy7fCYC+BEeblYkVORmXaIP0S4I
qjcmZotjVfGAd7GDseUyYypUoYTVQNn3Dhq8JOoOKpsGnYCBat76BO4mKgiJYsDI
k/JfvtTXKQ2w74D95pp1DmRRUl3wKD7aS/sFBARpB6z2thKJByMAPeJMMiArOSMB
PfQBZ4sP0F3b4yAo33YcFA0nyigUxCl1pDazhR0R3YCwYxSEa0kuxT1lmMn1fCUl
KJhXt02vHdYq9lN+oYKWNZA+nYcUUCZcy53yhjkrQztTXucwW7ojqjMuoTdlfQWh
62TUs5oEavw6eU6xKCPTO9nEaRc5pPlDG8q+1e1CrEoQebEUUAy7icdSiKUQfzks
D0j28Oozzx8/wesYWBBJ2zHkrEIfMV2p7fH7sxW6WFbp7DlhiV7F5dD42FqhIAPg
cNMNHtQKQHxHIlNbHmOQQqi1zWeMpoJW253RNa9Sv0XrT62uyDvXkiO+hfZ292YM
SnpVyfdolxyHpBdU2LeEdKowC/gHFkkioyXoVDZeeAI0uibLSP4Z17UJXH4g1Y32
+b164ScnpQ7/WLX8L5QkeNBLnxR6UIZrJlKAfKxOkCRS48RJjqAj/4zlUeWo8PVK
1Xb3ppWQ5b8+ZE0oCM1LBsF2GtnNk5vFhxLBcN52Ell0w4iSMUZfQyOziP5RvJ03
LOk4/iH2c7P3ide9KBYv9cHUOvC0uh33sWQsXum00hrekGKiRhlN0UgWD+ZX90CL
BbzzeAe+0jpTG0B6XsWN6pwL2bSwj3TbQA5QJmxIVIa+kcnroOB5g/LO5FgU+5FR
r9+eFXS/MXLb5LGF/NOqN7vJxKZQW9rrs0GU8B688vQqjVQVUUhHBrTAbR7KCVFJ
Ms0b6FWMcFjJBAkwew1E0pVIBpL0sQKHjKGUbt+lkmu+JQv+lWNgq7W4KHAnV9gq
iSdYGwUomn7h3qWKu9cLg3bcpFRY3+6UNzr9sbgiNjJ5B+yzwqzWaUaLm7y2v86X
yHQ9hu71vDuMOHYaCWLMIO0S0yD9NugIqb4BjvwP70LgRYdyMAoh2JPnrjMunjQ9
vy3vNIYdN+MQIiC7yI+ox4Bk+natjyNYoGECNdoK/4FuTJs887LMr+6VdCi0E1aQ
hfwJEeNbAT2jaZvrIQ9VxIKEk27pdIIBd52TXgHR+vxE+8SsTcx5vEtdO3R/o8/I
miAAQlyoMapwR7spQrSOD3FAWlE8KOriV2PtY9DBquEwrIl91rQtJtgFNrTdsjMs
UVbyeO394+korzU3x0hg2Ph1ea3JH9yfPhUfQsCuj4fXHKzWuemCH4TprGh9fEmh
ZxvC+Q04HdFdBQaaMSekyOZT8521rPDZaOcSzYOY6aDiHlsrvIy40HIn+7Ub59c8
SMDHrVtluuN+ZGJBS55wvxHQbl56I3vqAAOhFHQrYx7JMVbPQWG+GpgTzO1N8WOa
GBybL1ZdOsF979IJbyHtqiuWBGk/Gu9An0unBnJ3kzCudHWVyEQy8WCuoK2aNgSW
MwP5DgdYH5hfZn449i02/gQsnvb8UlgQQLQvLHDJRkTQ9QFJhYOR5XBSOqSANSHm
BuMCAF8qF4VtoYCVPC/eK5CrAq6DsRUc6z9hbMLZwjtDITCmI+LIKhWem5paOfHE
j0bMQfFhjtDB6N3GdhxvFS1pWJcha3kS1xlKm2s0UI3vLXl8Fm9OU7xEvaFt5v3C
XrvG35zZDU7l7EXIqDdBr9Mq2X77NB7/HfpUtVeMjn808fIrEe1JboVasD5Zf3dZ
ZmT3eXqKhX3cTIey0y8+IprqtM2J7Ab3SFZES1XO71uU09I8sHU+AenhnEkoTL1k
77KkWDxH+ELngjXsr6zwMdG8IklBKdhJaAFuFN9qJheuZwzkFjdPgg6ml4EWjWbJ
CGs4kIHlceA1RJjm/jzc/B8TChXkLCyAAco2qtxhphn1r4M5dQk2HPGfCeOeUJbZ
TKcP+TEdAihhXfE1JiKQDv7SE6iGLNXlBxJ3f3gYwXRP3kSimmWW3YXVmzI0iXgL
TiUb3VOm7vrdqhei+4U96u5O8OgWwIJCObgYMYzWLfIlsVEGovbL6HTHlKjkd1We
huRihYWTZ4jWu8146Zbs4Nw93i84YPMzYzXnWcKVzm7srUwYKCKbm7kBmV4175py
zb1kEtrIYmHC6H/BxLbt0wUlK+Hdfn63a83rGWYwKQxSxcxKXl4114/6keNgrOZt
QJcKBMYsmdGtS/7jWfapaCr8Nf0nYF0+98NRwbbFmTqXpZMCZ/XZGf1AO6duGJa9
OT4ZMN9Bn9lMNt9Y83JvntddCxV3uNL5/jJeafqPXE+FNKgogRIbuk7hJLIFRM1l
tyuoXDf+6OPSpeo3mCwlMqR8+5Be/L3/c8g+++XofuAoM0lsVAclamLP/4W/wok3
T+JB3uPZvYIhI+Nk/9mpp5qFxVpFFQNROqZZL/uRwGDegXQV/xbjT178cvHZlqGK
+1OW3VJiyrscqbWqQB8EP6W+LvgN5RlTmDtS2BlttXo7RaB7lnL7+WL6RqDBcpuj
UqSSkP8ETsGmaAHo5SmHB3ZWJkL1eHgByJ693YzkLtzfrEUVAWzY+5fun1BWaRKl
NzPqOdyc6DsMdmRuUkihTmKebT3gbfcfwwn3zCs6BWIDL/CJUn2k5BzLqTbQ32yN
y+En8CEbMxEzlc0jFVFiYp2VnDTKGB3GTTFlrVBZ7WaLWZtqIGgW0m/vzq05MQz6
qTtxUKBBnMlQkgTUeU54HW/N4fgdPtILNgEen15Lji95erpwe5pjJFSFPTRBXrCe
/jxoSxknBd+Iz0QTgybl9Lp3Hlld2Kgw+ixavPF/WnKGSc3YIUmk72+tcImE4E+y
PAv1ihxWIuvUqTVUZnMSdL+6kbixRI0mFCeuc3gNeLfGwTWNqhJR7Ss2z3qxX4VR
XHeoZxKmx1/G2FxIc4gU3B4G+bV4rIzGwzgWCrh3OrsrUjeOai7ziiQi76Hi7pS/
g7vU0QaNEd42XuN4pUOYB1sEX9dkqfS/mWoh8jr6vTeXlMzb1AROFJZPuFJxGfkV
rZClCQV2FfHabOgdMKXA2O7KkXVnkmTFkN5V1CcKDAlUxcHU38wOCHmgEraanxfe
HI5QH200h6rWnnfbeALtrcIWBTkwA2Dovrn8/0q6uyJ5a18mTi2enekDyOB2JOPa
vdbKGfJOoIQCrt8r8jfoMqdkLWa6IESB53RHplRGNljjtirhLsv0cszUTkTd09dW
us/56Vn6KJHC7rc6Q2UCR4grgkdJNW+TC1G4QzLI3N9gVVWZ1gg7GSAGfhvAZQjC
96njZ0oDva/IvID++XKcFo8gEK9Ktdu7691GPzJGrkJ3jCNaHm1DFk542yz2yD3y
/XDNjOREAPUicDL3yUd/XPtzEoKwXln6Dw1DoynvoJFroPWAVK5iLiwzpl+CTeJ6
r0lFdukkIW1tb75oNL8Z1HSGyQievgBrLZ5seTI+bJOiW16IO0C2olUCUeq4Syzr
1dbz9JDQlscFJo/L5PHVEuF/M8zF4U/syjtYM7GmVkSaoDQETOeJovI/lwNb4lzq
hTv67ER9bMjakyeuOnG+MM66GEnBkg7UXWXIxVp5DBB8G5Y2McreT2WtkyUAEnch
JNK8cDhG0Y0jue1n1S+jPn7iVKwz5MPluAA/EGXdKHiOomw3q8OLLER4KN4/OH6G
kWWh2MZMf/aXT8zPVxwen2cB7zU55ETyDanY2hBELPhl7qOiWsQNRLaeXHSp8f+7
iRL8XNi+tJX9jXpqBtck/yxrZHw9QVuBkSDYVTgso8ikiwIOLJtxqn4jK6eGqqOd
0x/oczAyNULdPusPHEBRFELnIw5QcyLFFUp49M2DqpfhrJXwk0yceyJ2PrKG0GN/
WyyVjqlzkurREdBbj63IxHehxwYTCiP+PPWddMIz0UvnmqIKuv+Q7e4neJaK8ux4
4+S69qGkjz7s15N1Or8cTtLVeAgZtyIisfQQf8A61n+07hpgCK7Zbgy+nfeTP9jB
pzCR58u1kjSKaitY9h94Uo5KQiZYrYz2nH6eKz8GdMVZQ+468B7pEpW+L8bmWVLL
zW1TqnDRmpaBsd15PZqCJqmshh3bKcOGpnt3V96AZdZUSD4bhtpUnuZE8VpqtWI2
keW5Ft/XqWTHyGlEWUvNV8f9fWwyTcleRezwurr96HsOlwV74D3fLPMf8fPD4Rfv
rkwUuwjQXYoPIEr/p/uLBu0zTj8pWiffy4so3FwvW2Ay1Jt2DQa18zuqm1DiPpDC
d43s/Rd++eFJBks00lK0Bab9uzRxm5QJWX3K12FyzaL7dQFTqhZikhj2oQNHqKWk
37n3nJJl6X5pLxFb7+03MQLm9D9M8+gSmvveoH8zBMEZ14zHKONs1zeS2NJnbeuK
6q16m73yEXlEqIblx4/oM3ZXu+H3xzV76OsVMBxpczp9/1p8tr4DWQtqRo9+ERdM
5cGztnQKut+QmIctCGMXYeCtBs7GRebZWJZYkXTcH7KnXmK3Llgf7D0vuj4Lt6kx
PxLQsCgxvrpEk7SGmaA0GNg0Mf8Y6HtIKDbrikjuJn7TeWBtoUPc09apJVZL6vKk
iQBvSYO3Ndt+sVcxv1VSHlWnF6YE37qIn/Z2J/MlrCgxWqIlhvyptja9LL6+jLwH
PZbEzucMOfgVOs16QMn4TkZRb85rgsaoUFWmjxAKwO/V8oPsjreuTzmqhA7T6Kvk
mn7f3w5owxr3pZmaXs3qjTZ9kEnGlRydAa4Y93FDR8/T8OvMoVEf7j2g7E1hwt/C
e6iRooWdKeNiWysknhEpAWSlMR1BTw4J5B3WnzqbE1Xi1gaffXQaBU7BPt6FPDR4
uv/D1bWpIc/ePzbb75OSIJTLDNNhk81fg4DPINVIvu0zlON/e78DB8xRuJ7m3BjI
mHYrpmg8G4o+F5oV1aQRmoPb2RLpptb7/zMXfhvtDECwBMZQBb9586GV2xFzpZAh
cdhHLcNdDCPjJPavZYbv4v7J9rDlfK/GU6OrGey3CObZHy7sXwTiEKu8y00Czhn4
2H8ch7FFqXa4nAPg0SBTzKRpwEISY/tZgFGnlvnSD2FA7pKyeyBtvoZw5F6PweDC
8s0Wh9KhDExL7Zqxr/z637okR8yLcP2443LW1EhdjwV52qSXlaa5IKvkC/xn83fQ
uXKpmbNXSlWvHsfktDp38udq9E3648Ng6C+6JuaUXVnldCENmhNDyV1Ck1X9cFlU
/oQAbB43TNxdwwh59BJ2zny37LDM5+/P1CxXukFEifhxQdfW32vmKrYV615rUrLw
p7Ac8U5ytY+O3X3ACEShmfThQAvniBFJLDbOJoHmSI+0xdsPR+XJiLfGwam6mc20
id3e80W3GP1Rmzpk9s2DgG3rTRj3sPis8+rAMDsWvOQCpq6iYQR00AVawLQjBbJE
iu5c7bq4BRIYaA9IDKlptfrmyzjFmp7HPkRmpVaikjJechiWl/NjatFLKY0vGvkd
x08eu6T6gAuGww9m04aBqwbYJZsLlJnDdwY8/zP3foPTuKyPNKfM5LJZRv9qkDYy
3CeqLwLrIAeeNSgoTjjRnXbVUddafNhcW2Qn6xuwMHH3yxVEEexEfaQ77ktPbGBN
4y9G4NVeiFfo67tej6UNqPfhHKHZDIr8qNe5lpELxbCGxrktcr9KJPb1ueyXZEBj
h0iI+7ifLAIBKn8r0e6EFYVOBT1NxM9fPyRzSfpofY2VpCeaZO0qR2QopRgdjoEK
J4Y5yhnEcIvjOSx7oe5aqjZtl4EDovefbZK+a8qvfL+o6MwRi6ihpQwZybOwF2QL
YCYzFzrfCMPT9MwALuaZI6DQonMFRT9F+x9wGzt2OxEzEKVreB+xxrr4omFeS9cl
U0lRvEKEDzdAqaFMJb3Wivp2qUB8jF/PAG7D25TNpwKdLmtC+HGyZ1GHgwNg6TLQ
QgxDQelh6gz1eveosRZ1PqwESBqUqcx84mdyoQv+NOdcN2wg7ZwRXybU+pNtOJUx
Fcp6wcjDCvETYNRV6gWwxnGiK2D54KgmpjU7RMq4mQpXnpF6TTp4iJ5BKbJpqDVl
TUvuHhunhlY8AMf2FyGWeKzjldanEDFVbdChhLIPcsSlmxEYIHSz2gQF7Cs0ZWOv
EDwSiwWHQaacXhMCv0aRmUUSjXKeRv4wtju2APYhLDsizcUodiin94QiZK0dkTsh
taX/DWOXCT3BymP/DFRVMlUkWbNrcxqTfCVCGiyX0wVewdZNZ7DwxMrbUnutPXbQ
6EkxFBxuibGgddWTI/1mihjRfPz+r6RiHVeF7jDFJDsVimt8rrv2qmT/7/WfzDGF
Vjq24zCKznjHP8xEFtRj+btFZeIfCJJGnwj8UWJP2x82x5LMv0/cAjW2AbhjOP1V
JkK25cWuBONseqwKus8w1V6KwOzcZw/xrAzlzq68s/JjWjAYlpz0pYGvsK+b2LFn
RQCctFEu5zo9SHPw3BYLGjQi2ufgMJujKBbGDMf1QzaQCDwSGQfz8hWleY+CSNYX
ZPFhdbSPX5F5fvI4CNiaMLkMJgCpF5wb6cjS5DcVDcFtxLapYgZjjtawNvOLw79v
QX9kOfLgxqHhTBMDsBIHwTUw9D+fXbbV9NUwF2I2KYAPZ7ObGGFWnhYYDYqquPXP
WH9+ycECHt8gYRGTFKFs5cR1a3g/lX6f37DQGEVpDY7IUTyLa9nWqMD+Iq/oQy+t
Z6Je9TMZFIMZiDZTfiryacT5oeqHmPV9r/KXZzFLPI4PYpqWmmW2rZnr6u5VbTR5
tiz3DsVrfujfHwAFjKQuRzvJh82c8LWIAPmsoeD3sB9dyNYaeOKmsw2BSjPFIJ4a
svr5pa7mJ/9BIrKOn1PVy1Cx8YkXsspWFJvLQR8cfZYXUV265qGwTACAiAN1zD/v
3+kNO4q5RYolDPmB1HQJ9OP1jBfLKWChq05g91tJQ7Or57i/K7cuwS5G8qMeLn5Q
rbcJvMS8WL3uPLArjpj6x1B6yOicmJEhOOdEtlESJd4/uF+NHaQGmZm353n4Zr8o
XqEyfXfLp+IVKypy4eOkOuMmhP1LW9ix9FrH13FBH85EKrW9UJsyVX85Z6zDAbHh
mglLKdOsrPthPTz7n8+BdXVgM+2K3PJWl8906oQNrFQDuB/26P9pcz1e2AlXVaUX
1f12CeM7nL+kgwxDOrEGu2CZ5cGUAYij5a5nA+X5JYgrtfJIdxk4Uw3GGNpICSAm
ocy7AcB2gRNzhWPmazdOM0IEx1SJgQCaky3LTOofSjm9pMpHqN1FT5evbBQxRoFA
w8ysAT1ViT1/zZOqTmmCTjmn0eH1OJTFXs9AIrv2x9vLJ4W3O6WTEa++rKvnjdOw
iKEK7ZPEgnXmZI7WoW0wjZ5JNaQU193cmQc64mk0Hdiy4eBmHPzKWoqgpCIUD15P
2+3YoVxX/yWW/XrQpcg88fqFnfQhU8/0pEyTkqwrtunM6aSI8hja3kd7BPLLqwS4
uTDDpbDY6HyfKBYRrrQ7pXI/7BJB1WiQYHef+W6iBUg3CU4JpfufIPeql2iHNNzg
PdShhgai/ktWyyDit9NFhhOJYk+3SJ8Pw9UIdn2RlhROeVFbV0RFB1BX/6Igd4pU
eJE94C0bIrqaWICgQ/VYsQgtVPAXOUzZHMUXgScyCdxlasqFYY4BssknUIleCKeh
q85DeoEDSIJcoMTKMK/92dIuDU6Ew5HVy0wj3X3ea4TNATYthVU1pyjOCuu+pVDz
qTi02NeJ+FDF7knLTXEOKnv7zG67B8Fa6yhmrrZYKAB+KHRqnH6o+x1j475GO31G
ZuQ0UaG0dpRzq5XhmP7uywldSDr1Xk/XlRxNa26U8lw5jdctP0R60bsV2YiooNld
j5aDGJGCUsHY6PhMvyilfFgTRr3XupE5IDTGDXp23iZJmPA/AQR4j5JFf3PtgvOp
Vz90YRmkAx50nk3QUL1DRrrd3yBKZQ/t8rpDKxS4rPOGP/ggLeO0a/uHYpSlPaXq
fca70kdXQEpZVBlY9Q+jT6CPWRVPG8QfJOvCqT+ITVGwkCaoyccQtDnxRK8Nm44k
g7qERRIRehj1MMpcq3SAXaUjTkTOXYxP8Ala/SZfdAqg8U1QLD0/anpvYicXGD9M
kcgkDGC6lQ5VKVxtAy3tY3WjmVtlj9PkfiS/ZWjiPkq1A9rmoMTPv9plot9qsiZE
F8uPk4KRtKqKyF+XWpusDvbvit3xoxwNI/qBAjY788H0gguOlX4f/zYo5WoF+/2/
7uKRSE4Me+87CBPn4RvckSSb7anHuXDPoSWu6yS/0WHHiwC8BUv4OjHy5likOETV
JZClCuOL0f0lzPjsLxrpEAjrx735x8DNzXmUDW/wUnD2MRcHYEM9FS6fRbCmELhW
/Gw3g7W0246kU0rLdWJSBo1bXEqdhTSnOLppVcvPk4hzSILC3TzyGuKO4k0DxL38
zglZR2jAK0GGTxy5EzFIPq7ufhNDgo4Y5jYfA8KjpCb/2bvaX/z5Xyf0Pa5+PiIH
+PUvUCcCpNQq9PEAjYsGKbbY+UGAzNp3ZjXBnsMBd9BhhblT0tlGbdM3WwIGte6K
MVBGwRL1hosP3tdRN4HCDw7IA8j6iqpqfvcC+1dqiYqNlY0AChQFV4ccLpWSfgva
FcqiJLTRsvBFOxozRB4xpSA2htua/PhbKb7VZoLYANp/D4AfJhJBjblL+7r+5vDT
bISGBwWXv54El64qv4vklDmupHMbjNhnXiI8/0XY2/FRHgf6RH0toK6d4AnHC0wi
M6zzSKO2lmqRGldfM0zcfbF8oreowOcs2+mrqGQf67GpMO40XNBn9OS2Bf//B4F4
dGorCecL2d7Yo1435z+AbI3yOugtph/KIiFw6JOgr4lK+h1A9b2p9kqciWKkZg0J
81rtSfKNa/J7tuHjXYLmE98EQ/wJpPtDplirBUvQygw1/BCU6b7Fgd3yON2T18PB
KsYgHT1z+r7CqLjUlmxx3evOrvERMxwR+UXjPczys4mQEIgdxqh7jdg22foe60l8
MHLuJqu6OzX2IzegoIPST/opzpD5Iui2pLRQzwogKFLCMARj+iSBKNXPO+Q5RVAC
S5X6wXOOb3AzDuIyIZqqzWsIoA+XUwl7EUXq3L2Gd6TzKYCmcEJRhO6lLtE9wyaj
xgL9HxLwdQjGXIN+QvmBvfekV03mc2qkNcJg4L2WBdOmgFxCN9EEDihlFveWVZP2
TWeXDU0OfaAO/ieWDIIPWuLG3OArZnFL6lIkqhoK1CyhiRy9MiL17Jbg4yRAEGsM
vgtuuL9MHewp+CK3asmeSzNN86SXuAUarKDbHl5x99EvxPnfGbT565g5RqQSmGn0
JAWo1fKt9EiYtJYxogJzuluyRVXMfAWPMn7P4gGVZ0yO7siayea4VzXnOxZSFkZ4
+3sDpB1DcCiSr7q7YlQLMfIAqUCjXcRHY2Ggk+6nLQvSHgy1L91XRml3Jx8LNPFK
JsCmUQ2Lf/v0tokAsyUPb/FxNBYr61CVAY8gwc4Hx0nSg/J3ujpxW48dRa53Xi68
pEbC5pKypGqoAJIFGNNRAGaoZ0rBQdIF4uu4ihMHLo13oL/HWkGUJtgCyFrGFijO
y+//CLhykbLYqpCK8EFJQlpfKESgNbvusZg+HViPOIZMyF/dR7ZCSjjxTdLCgues
oGTk9z8HOO5Q/XDBfxULd+YBEMLEGFuc/Vm3fbmbrXnt4gFnD/CFgTLArWPQHAAf
C26mMvvojH5KuANaXOGa46OhdkgoxlTS/FkkagGWSD8NuhF+O29KJf4BvAlmXeyi
t/8CLl/zRJVT/r89rq/qmvw3av/KkVvFeDIs1NwpAqU1P4tUc94+jSYGo2U1u6SQ
GexcIU5vjP3BqCoffpW6SOSTbEhjiHYI929UTopgQeNNgU3bg/EK72klfOrPPDVA
fI0pqdNMLgRBGLCqHm+S7Y4IAMQ3X/jUq/VjQ1D+g1VDwJZug8D1TKOWZBILTNJq
uXjMkAsoS4g3WQUsipANEBsb/+ph6YiUZd+agFefBdZPiFHrYL/cYH+3HC7EU8/D
nsnLZiGRGm2asrN7uJZqsZ5QfWLf/9sNLVYJC7vWpW9Yjd7EZ4UlN+rzf266FY/q
xg72gwB406uXLvoYV9HI6B2FlaktyB/uteEyj3l56wG/jP8EvWrWaEpMOvf9yI1M
XyqwyNm7hGQURB5in/Ljz6ITbiSCOl9Uhg/QtSjJXIyw76Iw9iGodNyEY6ptGEXu
pA4cGnEYkzy4F+ivOStXuleXIwTH9xsVSACZIOjbpPAwMhB1TrvWUodNhYFzmS52
cc4x3bUMyAxrz6w7B5au6o1tMM2d+FS4V5iq8Z67ZAsz8pxtHBMv4r+ZHe/WGunB
wFNL1jbmjyIGKXubgiOkaQUAJA0p3+Hey7tfjnko8zbvQZy5I4Ys0r3yOEgT0pQ1
CRGeYrEPcD5JomPPsimU1KGK+Gek9OZQ28qJcJGuTjJUeSRiokfyGviGDxLXNPOy
J0phzOWTfnIksShgPYjJuy1+J/NOmKOHLLvjxClLtCC6+AxowXl9QouzqGQQgXfa
5v07HRVyyzutFkbF6XtqS7QQPefSPNwJ0YWPV/Ynch5kY7bXu2s84aPpRSdToAyI
vZKvL2oUMLXijLZG/t4Zbnlfq4GoVZM5F8JrK3hwnU92luuj0I+RTlgA+QdncDSg
kfCVnAhHY+cImAg5IxV2DmhR1pcZr1rzD1weAqyQUKZjO0KiMzGm/l41H8RKb00d
xyCzrf9smr7bBeRgebXVDyu/8u4pvjuF70RHRmF+7Yva19bopww0MeOIM5Nf6eVs
keMm+2QhO6l/6lBd4FLOfIFMLKXvqGt5Oet4as+UbFlSfDDFDA/te4TV0xMQncwR
pJj3sB3W8/mH6P+3jTUGHF1m3zpSZ6h8GB2QhguHkuj72ED1nVaS00NEbr+pikJ4
9NCabph2Yg1KnG/9cCYPgBEkkUkdshW6rYGAbQay3q6Q3S8xPn7YDj3V0c4vymIA
8xVqvWCoIY6TzRZfvQsb9TJY/DOODN0uPoR21w1XGhgkzO6GSoYXZV3M/n4SvyXc
ZAQI2MZJtmS75kNcSDTnIUaNnadf9vqCN2sBcd3scUX0hn93JYz8GshoQ2cp4/R3
9/maXnRHnznAsKcZst23N89cSVgAlwQr39b+BdgCA1lu+/UOltX++K6EacqHNGJC
EJmMhJI4X0qz2u2gEL5Yodr6aj+vwuE6bkaDJLkiIY2ZIflH3WS4sQwSw0tklJfP
7ZX15YpzQ4w1KH3wurYLw4laobrJ16AzHolih/dpNFEE/Mu8AHU/BifT0l0TnDbG
2GH7NxmxlJfag/tFib09PYdyvmIyhpzOkF3SqGxSqQF7mjDz1UBiraLJhqcdpLKn
ZWPfpkRfjUrwGKcttjSwwqAG/iJhxSd+o7ft0sDHKAso0l1YmUO/t8c0dcMe9zoy
8cAQADxG7caXWykiwTv/+7NzNqVvIBykDxJu94d/wRNFsiSdwlED/eoZK3OMjFwj
SwieFX/v0rml7BRL9nAzVOJfL1lFEJGigUWd7WB+ksXidSpMkWsQpZWxEKKQzqgm
dzUTSZLhrIT65MGm8zZXB/lNEQXKLcZbF6Nq6dLGmpSJUFgvk4Yl3RnQuxqo0XGn
IWYdMZyIYlN8nWAfFWZ9DXuoVHJ00c5XMvTK5SywbuhCAja40jWFWa4QXM5c/TQ1
9MheF9ScJ/Xrxv6tM4Hk6b0CibzLjMcv2FhEN1rwttBd8mrhz7sEb/mirMJ7xQJu
vjmoE+PdpWWjpZaPggqorQ4GnVzhnqCzWpfwAvwpKk1pKOOYpqwuNe47Z9ZQYoTT
fDRbrGtP5D08n6qDxnrH8wvFozuw+cTAtdf/WK3zrBIaycUdFtpZxTV8qMHiXOGI
ZTFB5hSjgcQKDS4XpWA0ni3Bcs4tOHTxEvIB4GuM0Qw0NPXZq+g4l/yXK+NOtGjK
+nsNnnNFPUzZwU3iCJh/m/suyngdqDwPO5grjqXIs21B20tDFy1zasGJij2uXPkc
WVARZNZkaFVkT99QHbhP0tE0lYZdJXJHz06ivoMMC3CujSR6XKI2iQ9mrMdtLpmW
PDhLZ5LP3eBdAlorejW+b8pcooAq7No0zjA1lsjYhO8wc8l4d2Au91yBqANR9Wds
ODT398WKfCYyw7mWbHZlGDpdNPhhIQUvir6CEemwkza9AFe0L9NkFaVHbMcT26Zs
7mWFRuBjAJEAagJolWc0fNF8BIUjF+Aoi6ydhwXkI2OceBFmfzAOH1i+55UzH15T
8p/oy7yOtmhHUPWCilgwHa3eksya277sZF8NdfSjVakIMsTyWwPn/3G40lw2epU9
S7PmLSwy7BnLok65cXamNB8gD5qIKYNJ2s7scNrqT+iFeAnhAjoH3bBPwC36aGSF
AkLtxDp0G1nsLP+usyhLHKQL1+qBluB0pI2rzHHJjXinmorTTF4eDoWaqUz+QqAU
LvgW+ExygyentRiMhqGUMBFFBS9JPzCK9GI3gbmanffaoYJCdw67bCECzb0Z8lZo
mQBrAFY8bvnqQ0lIu31r1PhPuV0Z/TglaEnwAwRVS/QyOHT3m6cHhR1QH9sm0dNq
pDOuo3FBOZXz/yo3P0jT1oZsv0iZDwk20SKtuPJ0WB4mtLmdIAR4m5nFJT2R69f6
3Ch60yDpEMr08A6PMunPBshjc5/eM/1JuE9q+S1UOq+wqx4Mu4JYw6MU+9hzusyi
aJ0bfYfFtbGs2ep7r9Ri/yvzd8l5nFxhsjdDQ8BIaQkDI05Ln1zzYWgF7zQj5bk+
28o2ytucb1anbrz3TYofHWNWDhi2hyrowRQD7gXPa64FlhVTZ8B49ARr8fHJCpgk
Ip2MCcJh0fMFAtUxmJYIrMe3DJbxe9ecLD/vlr817DP77bfD7Q1ZYQcXmJhJ7R8K
ZMwB9IVEXG/3Ijr7ba34s0Xb5RwbMN9RttCbPV1lh/JMcGdfvIdWHNKY+prwpSDS
cgWW9eIdxp1tGDUUw/yZTKD8yRcJWl18VL5i3+q73/Htv0YGsLuKWBzcYIHMkw7U
MyTNmGClY4YQcX33h2zDPZ0/Y02haH0s626Xo5ZADiuQgzOlvWLg23DSgF9enmqV
3jeXJXkjntbH5vfZXYqiK99L+LOhjnngmAqaJqjTwZiy6o2UyM0+dQJFB+84QlF1
IDJsMnI9dmgMHAX07xv5pNDciCMJ3iPJj4f0u49xvcQQ0tw5yTsKcIm5NKgO5iX0
lDRdlaso5qE1Rcs5FgXS5VISaWR7Yr022oWnXsKVMQNsQT400AHYSYL0bcf00XzB
/R4Dep5jdKyDCpH8ueLeeWfWWZaGzTE/vsnde8NzzJKASHv9qfFrJ+Z6OjXL9feJ
f4l0yDzC9w4Yi21INZzPBAfboOysEksVHNRRBq2aHNDcSqP/AnsTitl6QB9SJ1H8
6u+JsPeycAII4JPkEEYGzfnWjXtRahiKHArIu8P6pD8vh/fypR2XV4wkhqq+zmhR
iHefbXb/K0OhN5uq52Ag7acVA/NOLlzFJ4N3wyVcH7KJZgA/ZBXT0hTifTmF/N+J
1SBg3byGb8bgIv7t+slIfbYloURovQ+ZzASkwdYBvvcxO+GX/44XobwCOgci0+et
QjSqK0m8DOwDIVL6GVEbtL7045qGxZIrtnbq7N/mRy6xKZz0Vnyaz7FKFrTz1rtf
KWxn24pxmsVOqbvC6q0gAQCHvJ6a0jAo8z/fUyqtAcYXf17JjTEk8+Sp3TaSIrZq
CpvQ+lmxWR1DEO1h7TywT45Xn7fprjpsjnINyQs2O8xXiI3anO594XUfE5Y+8YE1
QhsECO2JDXqL++/thQP/Rx68IbKY77SAgyrVCrIEdLZC3Ky6QoPtVgOv/Bc17i79
lCn0nfRPRdETsc+Py7CRka0+TM5L16SO63TzfnDxeuTCmb9YBx8y6Xn/WKgQCvvx
+ioT8uS5WtM0wHQ0GVEP1pS143IymnGpOAcF7VmT5UYWKta90O5aLBqsh1CAvjiO
/O2hSGs8/RF/AAEyv/priGdm3GzDR6I8HteEqhcqKpAt6PUyf7qUt0J2UduxurPl
J2lbdFXFdfLeXKUbqb7woWXbuWUCC1zvReK0lk0y9uOCdPz41cWOWtFjt4ozFFZ3
rjZUQ9AYYHTazo7g02BqwjgeP4FJMtfSJYabFy8ew79Nv+pyT4Lsswn9RLnwv3/N
fOb5JylcTD1Y8QAIowDGpPcGBErC3gwQ23FYxOGhEQuGhOgOJxZHucb9ePnJczFP
sgcNIIlqh02l7ihXABtB+W2jn68WtX6i41JnnJmcFQtJIXiC5a2nFVvRbPSDBnzs
Wu4rNdt9VjyDwF6yIIpRMJsX7iELY85D+jkAazzPqZmI2OU3vK3z0qCPP0WpqaLj
yxwCnnwIIVTuQnxUR0Lphf3uHKB0J6OdYze8FI3e+p2oHqlN0MKPJ6dP5NdXiioH
FUJnS3fJ+lH5X3jXcWzBe9tEast7mryKiDKSUyIiQiuH1HCgCjhENcH3Ueg2HWsm
iVr6t5UouqEcNHXwlbgXe31iSMpSnT3Zg66lg0xFuf6QA6ENdwYrL0/DmOewicz4
oyBNWSXzCMxHCDtM7M08ptjGmnRiJfV81YnNLj7KWpgbn0uMTPE7/7IezcnVgBOV
8r5vLXm6njfVRzPIGsvoJ9cmtc616NCU0DfBUVUHvry9iSLHXFdoyZsBs44kof2s
1MCcFCfONbgyVnZU7GAB4qChqdPdttS4j3aG9SXPwO/bgEo3xN+6754tdt0JjCzx
s+lt9kIF/mjqTa3S2IMO/WtlHitsP17V0YklM3hx9y++JOQmfRElGFutJvakQsei
HIfyBfOrndBpRHLPAnDWPBGyaUCqNUvy7ligMxOM9XXSMnlRmBbnamH9Ev4ZqANM
RrDuczaxIMB42hzw9dNJGU/BJpd970nlwa37bTwm0NNowz6GAisRXxpHs6CYXViS
H8P+p/ufzVocffn6Sz6l1iM2cVKv2P0BQXW++lse7B0UCLl1bd1FujDw7eyB6FIU
k7k39eeGUrM5CcAoIcKYIQFjZNf3JRXrKumAGyxVvIsryRobpBOOgrzGA4ppZ+Co
VwRKKDQaCpLHYyPHZ50bVkxX+xqcTB+a+s/o3BS2GC7l025j43+mQU5KnaEA5+e3
5156h0ahOitC24vtOx3OOPSJ+ESpiDoMpmcsQ6XL3FEKncUpGgnYnqFcsoH9U720
xK+XjFpfLmCiDDwo1aAfGWp5IHp+DqP8h0DQ7M5jZFE/IE6SHEQjo11lBOSq/uW2
tilav603GB5xWwPifThcKNe20PGlXWPY+cHJJZl/oT+lJroracLHsDT7i1jWW2Po
2hPhNg23nQB2Ncy0IOuqhbY+Dh5Ca4eyZQH31RwdNuwIUVS0joD0VeWQVWTBN7kU
bHPlLtHKWkt1rtP8ihHv06F+f4kk+oUqvjPhnobSRYVNRz1f1X7L7LNYG1H5qEx7
VUTLQuvRGZs9omDNLeO6LZPhwEAyamPqntFWF2RHUvF8jJ0bnVdafPdLg1UxKuiX
RPYrEpExmXeQ59Rh40V5DTjvGMlLPorkevvzUresT35NUkcL3ZottXGAHyyX6vVM
8+AQOnPbjct8OK6irXoa8lh2Wd2S+ztKYPKEdhRm99lPX/ttsEZtG4I+DYkZ6Rfm
MQbwS2jrm6MefeqOpkpTI36HoO7w5Bgad5rLpzU9OTpvqKLN2Kf+Ks0kJFrpmAaW
eFleYzJFBeUvcEKnLfHJE5+U3Atk10fedaOmyA2Sh8E94O5Ywb29ouCPZbWcWTkz
wZ5sW+4j2xKjzJqVMf1JaNPB3pde1i2CQ63W0uOzpVvNltrxZwFwnGDgS4LNxm5I
cZ+949N/TshmhAHxgGk2k+gOjnBcOZiH3TdZPwHuFn1v5oqopskND/LTKKSe6ZcE
FztM10l8GKHM75WV0vkvdS9A9L3E0dHwfYMPVaSfPRtNu+WSyOLyKtpD967JuPbd
otp1wd6wk2O3dvzTcqhkkVNev66xnmhnleGjosQYCQMBbQiirG10Tggt4r2OlEJJ
EQJVSVtVQatlH2zMJTPSHAPdzFztkrYUkpIOW0H0I45sXH2Eb1lW39gDggDdl5dV
ao72lMANbrmrsACQXckfJAO3kygi6lrIT90R4ILQvslpz0iO6ZCS1/sm4IjXo/sy
OVRiE5QVtwqGNBJq18OGOLAKnOnMjS1hFAAI60jNXrn/Tt8sh4/P+R43A3ZXI9QD
oGwoQSSJ7z0mhuIrBYFwkDtdbnQsnug5Zf1/V4dgMzIOc3mqtt6hzB29g2plr+/E
5XzNvsB9+54iw63LZYUcWqBDXwLWhI/pK2uA+nEf/fShUy/1/42ySxsWqfXD0CdB
qllISB0CCl0NK1aEpEHQ4l+Ap2e0QEqt6Lj+H6z8czXbfZ5Ww675Y7nAl64UgVtq
2svG10655AZT1T8+OT66aCkJ9LNZPdsEH8dzPRPqwdeW1MCCu7JgWQievNxPPKzE
Bm9FC/Uutj9TdZe4/LzB/yvXLXoOZy6F+8/TXn5QLeiZ6Ibg4gdqDYguXzQ+Ub08
B9sjrMfliMwUqNWZu2Gz87DM7J77JnBaOB3llH92WOhCeQNk7FXKpFKhkvavkEAG
vzy1MYuvBYMA4WGK/jItaYxEBDVgVRfj4F7tsaCHSjMuoi030Z1Xja1Me/haReEZ
vQjH+GlsiawhuHYW7e0yGaVxy82SFsW0y3YBK0TDC2GQAI8cEr5YrSPHY/FLuMxa
a97FkempCyf33nUYIPpWn0nqeKUoW1ou2r+FyDat7KVTZ+5dOCmoPKDk8SGhIsoD
srJ4s039laEBohM/GKyqutPhOzfXSLe5o8d6crO/Cp2U9s6B2DUaGc167M37/2fl
wGcRqAbhJROyIYGy7MIvhctcbHXw1ywNa7rx+IFNvEcxr7utGW/t5es3aRF/U73u
O8rS7z8oY8U2q8n0XxjNFRBMEXKaCuFOfHNkIyoWi5rSaoSp7q69sbEjllTEyJbW
4inmiVm3Z1fqa1467z5l+bMWVhBC7kpU00lCb+j/RMlsLkEUMmfpED23844GP4eY
MLi17MCeIC6P3rNrsm9beZboGEDb5D3+tPjyLD5DD7XhB0Iqkv1Mic0PT4BUY90C
JmygwnXN1HOQ0wqT8Rq76l5bOXDe04u3cVdzdjf1oywqfWA6D5nVdO0c8HP7vp99
KHS5BzGvAux7Hw8iJ6q1mvuInwDH1L9RTYhnmeQmiggIxuEfOxJMWiikWXy9oBB1
EufvgzrqYuhkEBQuKJ0c6tWMFzKc+0JToKaPZdguAXNL1jE5/qmYkckiIYNqEMg5
PRHigZPMgV2M6VBNAPgm/Zn5/O/GA4HJR2B7VHYhtvJ0UnS5Fiup3043A10vOhIv
1WAJXyEcHlbne1lyOgcmJ40J9YFNmQwWGhHmpETozFwsvs75e6c36JvQDjjE3J2K
p57oeFfYfulA4Lf5ZX6Z4qPgkiznrby42KNAmMkeubnZ02lSwnrzDMRYokaXVahq
4bklqq4aml/ADLcTAHz85bJtcfjcA19aZwsDjUq/8C3nV/1u2UmVF5GD+E1SaMvm
k1iLr+C2EZW4docrAXnX8RUVYnn4hlLn34g11qSv1W5CG6tphOJgTSot43i2DsAg
7EKTfWYI3QEDcksDi6U9ajwJeUoh95S0eRTc7zfvvmdAgBvUWBF4BnjbDcEBi8dc
EvZhiGMAWPSHrVzPw2+F205kuwUVQr9IMJcbC4GwdhGnaxiZnlZIvJlFqeuqF6ym
5Ipgr7ysv/sB63pZ9tUBQ5OMntQ9h9Xwkagkl0mOvEb0w8ObziZh3goQTw+/h1nG
ZvHR3xT8OCNBj5t8QO4ABf1MTQZgoA9NjMWTeNirA0APCW+tDl771VreonK+QufS
W/+B5p8ZYE546KuSLyhy7gQASBFhcSwgw4N0dGZNYd2xaS7rvLN8m9ViRbbNAsrv
fk0MvymGOvLqrFM7trbqAjNH1R5iTVMAQhIe3Z3u0eovsKYrrwP/r/PtErJvPFYu
ifAG39d4NL0uoHDdxzPAGF20OKyOgYpMsOEFK3mYNFZjEaefn9DnIIHl9ivRhyDc
8aIhvXo66yCVExFM7FnQ60SS59SYHo4cBJUDv2q3qhWSPOfEj7KZQofOtgvw6JW2
X1GliusD0wlay1+t/48umL+yJgPwVv3EIqMhuWPDmL2K9NdVlt7PTNcU1hHFYc91
XIOH+9Ix/OkZvmighi72XwPktLOM/399DG7OGeZiCuQT1UsO4bRbF/vyfpqavIbL
LVfLypsVr+Y0wEdPdHFfbSuOuf1Dqo3/zSuJyFlJEMM/lCge/8IJHNLtcmGRZu73
yqudjpkY23vOOfAyHWRbMLxZ9e6marY5wzS+1H5x3lLAr3pExPVL6drkZppqFxIk
FRzD7D0wC1xH1RMKkzkUqGDH1XacdMYP7PawsxYX/7m5XHDdgQvhdTXImdur2Evu
erKC4Qstmf8uBCAhvQfgwpm9oxVX3becmjt3I33ftBt7hEYRBhCPXfNC6GOSiWIJ
c3auSWRtuGzsw4Q+NM5EjsaD4hekj39MkCUmuDLQTAPrMfiy48aZDXlTeJsjSl7r
iYaJnDlDCw4BBUnF4RXp7VUlr8Msn+uqGjS4JCrpd7GLQWeYq35As/mGeR/2U3B3
S3w2kIlwHRv9IC6AqIhUthTn78F9ixjMvx1Zz19ZujcI2Drlvqp2C2E83NbjpcdL
fyqP80jiEW9O9vLdEl/Wv0SswTPuhiJPZSd7EpRfR7ondbddHApS/tl/MJ4L2h0i
zBbBvyX8iCJbq4l0c3pn4mzMvZoKkDxiWaBA4ekNvSinclrkAbm7N6WIzSLIcjMC
iynsBXU0ZFfspBSLRiVCVt6kpvjpvD3ur4epQ6VImj9CQmBNU7CUREjjlOJaq7gQ
ZfP5Nudlqh9W3ur7YB4RmeWBNuQChlaviZgRi/Y2x/q+KgprEZijOL+RNFjHepr0
Hbtn8M1G9YtsBT9A+KZgzWMfcOTAHAErfRIv5n3lNrFqC3uBO98IJy64VerRazIG
6jeRmCwpuecXKcbtcl3so44gyJe7GARjiA5R8lMQvkG5f2w4mW92IMPifT+E8hJ5
U+KY2N9YxCp29TLTmp/BmZuiz9QG9VissB6HSXn7IfX6B4ZVvZVxxOlTUF9dr9g6
TH2MkCS0K/TwcW183UAeIEC8JLGuGitd/hv6M/tPKOuNMjTqCLFVWCbStA2hMOzs
NOKvnJMyAZSJgtfKPa1DHODHl8SD7qJk/3tTcV+sQUe3XA4jWznz8/JGONa2pNCn
Uw92Pj5ikL9Nf6LXuWZhTHWagkFsvx7S2iQE8ExRVoTGABzE1DJnBuAsfaOgCkQ6
YI78pqdYeBeQhncerKOCIvy3XnIy2Ob2z7NvEBdIAiK5y1XkA0vrXPjjUIZ4BL2J
mAKGFWGF4O5QGlowVzwpGsDhxCLduroZGvA68ohuNhd8Kk88+M1/Dn0uwo6io7T7
6nBAj/Q5PglIBNP8dH0aRa1m/EuYESgTd63TPj03YMZpqBXbT5lYR6DN4cZTdO+e
okmRSOQ11+LZi28MRKIX/kQuaJSBlZZN6cpjejDyxiplWdAMhRd2QGChSI1lfA/v
v/BjN6ZtS8nSTtM0F8b1XLtc1GKHztuL0/B0ZUwXAu6KTQuFNRKJJM/O2+QgZhve
ixOlxIe/v983FppcpTZXmlQPbxPJllR4l9y2jIgA/5z99LQQQzkp86DTjV7F/7jE
h5WrqD4EQuKyZZIEn75WhQUZDmV9rP8lRO9s8XGYw2O+6sPDnTLWq2koSVzK7FGg
kSFbiTSXe3VlWhRD6f+9ysZilbgPhbT9ELOZs0G9jfaBNqfBJ+VnNuIOIG5u4GGl
WgCZd+i8tWLNctz0wGnsXiPl8q8p32wRI1K4DwKg4FWRHFmRLe5gIc96yTVoVdD/
nnFCTnxieGji6b/kzOFlQzeRr34WykcsO8Ry94B/kRO5R8olha4c4zARvxXSdJTm
0LDCdJXb4XI9msXRAT4SGODFfGQHW72JhDJSKwIE2wIeSDCGkcDPgQo104rrVHSk
7yqu1KYBqgtFYrcBZIcPXPyXSPKdTuGq+WLLxoFCwL/alQxdnBvg3/bNdOYULsZv
/l5oOCoLm36h37j/etcSFh2FGTLz4Vn51S46sFYIIWmElGgNsPlJd5BkngVMl7pF
TvN5KzrqUofBu0LROiWFc986cnuQCvOzd2iT11YA/zRVLxBz5iWaEaX1Huo3lpXK
6MyzDIKDhVFDo88B4NuSYeXek6xtjZ453EC4CxMP8Z5X2UJ917NDTlU1dmZlDe+o
SP/DeGq6THJX+k6NhIJZOBnCkoaafFaS89ZFB+h0pZLyF8fBadWFGqjivguxp35g
gMPVrq/mST2Yjz6/ZdAQ0OnPeN2s0kaOqLilXoiCbePejhhOpLwGAabPaYF2+bB2
rWVvX0ZWW85pr2yGHjVACjMj8j6qsygx8sump+7wBR6KAc9snY3nwL4923GtN5RS
/1bWLb0Nn+1nwyfUSak65tIbvj2zGfKIyRdbmq7s37GQJEjLtRboWEMJDkccBNKL
+ThgdU3z4WoOtU7pl2WlsmrXB5ST3IhBvLphK/pnxSSB+nw57FWOwHEtnQyt0nZ3
0HArR27AQHQMeHCHxQPqRR7zrxsvHOoBKPlmBKh92IT3WnS8JMbgoOmaeDCSeScH
ZHUz4XYK/JTu21yLhmvDg9M11ZEMoFeLhwwvWRR+A30p6IwRsIBWWFCKgPJglWjQ
zPen/IxIhQz7oorUPJqPYGLQoO8nFh2rFgd4p0rzCtoE6rgpHbylRZ6SrAvjHHt7
pErZAl9XTZCLC5269R8iUIO4M2trDv8RDTcxDoStFx2sUUdeRQ2oUn8p0wHa0mRS
XAcR3g/qfsVcg3w+mEufgK3CTwXAnQKED9BCIjh4QyuUz9SdfuYBB26tDNoQJXsd
MXrKETy755avcjcpHfDRDWUGB8W8UvNUiiv9/VdJysDqfy/zPnKdE7PuQVHqN2La
d1FYXfCVXMlNVehrB3H42eZIG8eX8tU6nUbu2BRePRPVU1+K9unniGbF0hcMGoUq
mnadwpU1WicQ8qKrsnz8RYWHsrXng0ySA7SsHZufqkPLaQMIVl6JRkgS2WdfaOP7
WB/ZaJU7TOC6UM4PPby9M1JqUwA4iPtBXBZL3dHMP44TB5Mudl0W2EjYgAfr7NNo
lKYxi7osw+4UaGTbGaRqZ+FX3Gh34i8t6Jrc1DkiaA8AheVwDH8QQ8R+LfY5yzfK
VP0V/A3YkC2HbuPsd0ommHahUDjmb44cT9xXQV25NwKaVMbwUqw3VBdA2OWJXIe0
2MXzxqeJp53qDmN9tw2HQt5lJq1RdZf69rKcA6DAamy2bXAm+lodA6R0ySajJJS3
M8w8zuDwmL0DZFQ1QCEmWboT14Mn0MHLh7sTKg3s6KsIhSw/2vpx+KqjTTGKAr4N
2qAsbP0CK3LwkBrv//hwO9Qtiu0EWgm8Hafj1IEoWEXBYZCClbEgiFu3Hy82twPD
Bm5tPGS7Dnrc5ZGoFt5mj/2+a7pA5jsv8zDjk2BsC9INBfIACIgkFnP+c2AV/aOL
m5cY9d99dO20m10cN2LsqnctTNDZNsp9ruW1Hz++ga+rDqzssS4OV9QX6j6xg9F/
3b06Prc+ETNIvw7NlqeJ5GM17xAIP+8GIuaXWMOsefKWm2yR9fD762W21rSsRMiJ
YdpZPCSUuUeYgZzGTja6Lp5bc/UyKCkgDzW9Jtz5OSZKLCFOwNFqOtqfqIR4J6UK
bWVzGej6hvEYV5OOSbF57JFoSjlYWEnruYnCuMeaZzFbeeEa8VGz2PEeu/4Ssp1H
Pl/OGOPf+1sVabeG0HjHe52fKJQNlLGg5TCyPfNV8v4fh+meUqI2P+v9PdyKWSEy
LIbJS2U9+K/W8h15yR+61KLeL1FLJjF7oux1pudttoWX7BpdyWwhXkfvVxnMfkSN
NceTakTeDFKQcojppTKy+TtDJOmHh5LioimLL2RlmLUgjbdzv1nm1SSlYpAc4yWC
19ndW9lMZCEndZMVniSiTSp1cllA+dk8zQiiRh8tmFxgiAmkPp/kr0VDbUXwZwza
YvbpZbYBMkge7zzA7L6Wl08jYRsT6uaJsgemrvpjoo9O0DwpHiEZOy9EYqWSsvTl
ZbUBIc0BxFuIDvt6tmJwcekAs6WU5oDMgM8fNL6Jhufy8Y7uqwkkuFh7Wtm4eglH
y09ijvY9nXvRXedHhvqmvo5PdIOaLNI8vlRfk99EY2kOTgVFs5Je/GNWWnwRHSP+
HuyatCU2NzsPkmRiJBbSYF5vSZSE086eVvpnA/UhX865wtwOEwQyCr/QYPokchRa
EddfqeMl/IV6hMA15JoY0CDw3luF7aNaJFmQtBQH8KkmZiezODSOX0VU1pqODy5D
kXRp/jAnJOtxmaf7xecWyNB7NcCwpePte9TXPWhkSGr/i5q6RZAGr4vrJXMOjkXS
T71sDSOOIhfe6v6ahMg6O5Zw8dfOmHO5R44pu2OHgbvE9j3bD/eK9lfjTDTsNAPH
IWURb09p4Cl472jDqfihah5aYfKDQ4w+kq6x4LabEHUFF0yRuorY3ngGBeMfgBB0
zIhd9VBsSkA8ZSW9v4ADBggS1/2D+MBGZJhSjkoeCZASMZYkkdjLe4rGa/udbu1h
4my0OZdn4T5IcGusSE6zlqZdUeE2AHzqQKsihvmzG62Uvz4Nhsgv1TJctk+t3D6v
ubt9H6qH4s55qzwBm1FbOIEOWAVWSiXGR17wC/LO+RBfz2EChb2Fhe7YgOIwFs2v
pavKL/cXpPyYncb0twGB9wwLiOrYcB28xSRmEmS/QhgvRA8pdyaV8Wxf9X7OVZ2y
J5dosnCYYVQ4hC/MwcHCfYqQOA022ZZeZuHS2dWkER+zuF3ivcesHISHnXZ80wL7
cMPn+oGgd+8H4tLtr43Pp06MsO118N3heYsuRdtTaZyniaXx/pAmqILwJlufDxCw
1olKHknE2Nk/o0nV3hyFMNpJtpBQ4D7MmnoKSJe1ijkFum1MWVncheCdk+E7/N0s
oX7BlzORLpHHQRAXfKj3JY3OUmPy9f2NtgYp5HdsYtBvTEZuQaF6XG/25GtI1uBZ
eS9gOSRW5Fegs4E+7cMLAEwhf2Zma8wTLHFaWyLoQlSg7gz/22Q8YvJwg2/FF3s+
0FOUGRSZ69tgY0o/OC7zoDd4M0ifOt14zM2OkdQ863AVbKwV079INBRRjX4DXnKo
I+b2IrlsA6Gr1iX6RZWjQrmtCIk7Ysbpb3YbqeTNvZlL4TQfylU86rMeHpAoPw/X
RZggeYfuDmLrezV1ZfSNVTraukVwbKY7rp0kfs40ukrAo0xPw4/Yv8bWl6NRkKqA
PQ2K/jPvOlcC9JKnwQGelOm9R1l68BTdbAjWHCG4Sj64JMV9uTfGo2/grrLjt6Ci
6cgB5xq05srWOnTTT/6egTD6I+h2wczJcsWMIiFWXxLHLaL+wkPYmwO77CyPyypX
5YYLY0cSzzyfq6Yq58gph+MqaLWRghizgGomuMXiT0VxTKQS7+9kf00Bt7GBChKW
sGpE/f2tLsP77dLqG+i7Hz1bjqJjf16+wR7N+X1+gPMA2WJuQjFt0f2Oo7YRSiTq
Js/vQbirV2RCYsjKq6D9BovKo347kIAwU4u+vmkX17hy17wl3KY/dWDkiBAr23Ak
DYnLM72u9lOEkLJjJmCPDFzx9uHfPY7rhthUw6u4hgJ17dZwueOASb4TqRIbvkD4
/1pp7ydJSd7QYNglZv+2W/rFZW9xteIMhj6QjBruDkTwh0ikq9lGOlxBsAmzsLuH
zV0OoEdKAQwmlbjKC7+EbS5sCkYPlmIhJMjLf4MoNJCgrLeY1Y6VLXlIUmaMqM7E
24USBPEofVMf5488hDYHlQAdNsgUw83pGSgV1S6WuNDG+2dXDoAxwGG8twNMetbo
H9IfpI58VIvk1FFPcm+Ev0WO7MWyBMZL4pYBODzbSjHngz5+aQwfOwztTyg868v1
ruMUv5zjXxlFYDznpvhgnGjNbXkFJth9IPaPzM05msnFXeO+GteppM9gXMJrKwnN
Hu+9bz17ub+troOqkicdtrCWuLIp7HBWnqEI2/qNTHxeZQg+aWHRag2283Eddqks
g+DjW0jVy9KFXaR+Cjd63v/WwxeeulzHQDJ4YBBVS528LO6JDaIPr7e1hpt2Bn5P
BkpaXFjbvzr5xx+p3jDtEfzYxpzDrHbbgoZWmJUDB6iIfRvaAZQtPvzEwmlSKJpj
ZYqD6A7yNwKlC94eKTd2IDvIWmKgZmlCDT2gJcihnKFKjWpYYFBFvU2bsp2UuPkm
oI4s5U/5M5bCdnqOlkCKfsiB4X8pHqq7jilH1ZMJcJPoMRD2CXoC0Bz/wglUVT0Y
fU/1uZSvhpOaGmNpauGmhfve9hu5+7c70CmmVFfkW7HapulwOtKeXmGrLMpbZK7x
eV2ApFmbdyhLrW8HlZ01sckxjuVDQYCXqh6dur/yG1uvI7TSGSqqfncm1M+5/fwR
VsHHCoiKxLv/LzEOMxi6/Fy8yj8GF18RPReEXk1ByPI1175uyAp9eIJ4btWcs4+3
a2HwEWv0Md+8PJV3+34BJewyr0RzNThCK6oey7zV2oF9yU8Zj36VwxSi3to3QheT
wlK+QJmm6IMsuBpTTRWmxgjFiPPUYa8T3Vgdvp+4uuM//5IHnfE/kLjM7JOtnt//
rwJ0gPZESW9ddlF3DP5VL5R1/a2a1CVVXdvkx204jMyRejgI6d0GOsql2OJOoge4
1eYYEo8ycKzAnDCXkoYZCtt6dwX1IQ/cq4MB7Bsbx4fgLv/+fNIjUsrsb9P79hKx
qBwj5CU1xB8LACvIP3h0Gerp4pRF0hjignHA5ybpiLx9SduzN8w7ixPwFrMW5NSU
1zZp4EKSq2iEUPwU2k6WrfLzKUubKz59KvkGzwQ6W97E8Dpuxbzrl9aTQ1qFJXKv
nNTLILJJVsf+Cso6ATYKTs2DQ5iFujXWATPO93WeErgzMmaw7jxXIzfBBJDqhdm5
hqEj2HhouiVbWt5QSEXqyhX8FVMaeokAaOUZXfM55ZKuMWH/lodJ05gS+S0vjSDq
r1VMX3ySDJaajO8tVLbXulE/vVPpsOBzcPS7fT92tvEpMdNKZYO+OLANRSodt/96
SEmIERd8q9goGl2fp18LUR9gb7UB1ta/lZt7VkYKwXcK5LZ8707gXn3CDl6sDOxE
Shk06myCUFcK+lMie7nwltT0wtQHDDZmfGx9uDkXq3jnAuMXdFhByb/jPk2VU/zw
9I7Jjgot5DswubAMGoqZXBhe8eiJzozXGlnCVF6WgiqJH4RQgtt+bJkvW1BIO82h
vg0R3kfxyAhpuc6BUgrK7iPTZ+9Xs0TfTB6SriYoPVvkOT2CvaCtHH+46hKmGHEO
lAScIu1S4rJWlfo1CMf5V3t/vqazln2Bh/2I8/R/DENyOPMH9RH7LsEAf2LbDTf7
y2MBCrdrQ4s2hqHeYD3BQAga7EhZNGAHYGnlZG88xSYebpfJcIoHVND7Ac8TQonc
kE84ohDY9196kTBWMnfMkweZxMMEiLE29Xrj0X0mgAh6UvU3MWeoKDUsW5zycGJW
H5HelFMpu0qBNjs+xKAjz6tJZyeFDASnljjuPxLk/Agd+v2+C9xS75Jd4/1PAbl6
20pGpUJnqD8ejUR8Q4udAm+uhCaRZdbyXhJ7vYUKprLin7SaCN/vcRsFDTX3EajE
RHSpXgnFqydF7cwnW+jwlaq/n8Kp2q4sT+8bRnQd9suFKlRpKailrx9hcoleD5OD
dqTM3SbSrch1IQ4uoNa6QZik6l/lGmbgYkK/4BrwVy6CHWgdFRigJFsJDNo2wCOo
wGvumG4YDfwxRhzRzQOjv9yysNRxZHy+rY+7RGeHqR53dnU/TZBpzGUTnUTBN7WJ
hKmP4d8guC4+FMUqun71frzaV7r3brz5fuBLAraFCXQCeZrn2gV4hr8EdrvJxtRZ
GwlhEycLqWZRuMTPK/KHGbBAthejCSCTkFdN1S20EON/gSNWIP9q8U2s6FnQ1yfF
hqVcG7JJr871LNFFacvZXFinMgLwgRUR4W74mz89P4MyH81l86cAY0wleXCLR71T
uKlkeG/JtzbzjQGd2tZRnfnkQJ3J+h4LlGk864tMohu1Hu2+8P1gJ5Ylk8+V+Tlk
UtRf3wSVdUTnIregYxX3vPiaMmdSq06yYh2Nc3SgzUDe7np/vn5xsJrwPzAtOXHe
0O81Tx4nVhxNex0kWbN0SzRGW/H31MxuAJUNj1zP0YKE0wZtRJ2Dx6HGlGprUsxZ
Yg298+rqt4Hz3yiG62GyvqikL29f3+geFvveduoTKuDWw7nu9T2LkrE/KPTI6eCB
h7ZeSH8bK7/W2NmMzDdiwzPIJ6LOGwf/PE2JN2RXymRLSmoKcM+LYQaNyEBqHaw+
KGRLv/AHVsHbVaYeKmzfH9/KhgFfnq16ENp1P5mPCIxtrfjIJK2/r6ZOrGD7PQ+7
Ps3d2H+NTJCzWIbV2MHtGm4tCT+s69lNhV7yueyVmycVP7P5iRKPxFYXw3/nD4gG
4b13xUQmLPvMNGnvs99gIYMUfHH6qiKY92XV+BQ7OIrXcBtnztXxIo+Geozjiah7
zm+LQl5IaUvbOjAqaoalW7rYPxF+MTliHe7Q253+2uRRZtQXzLVoSFpth/mA1I1U
kyDPdQD11VQoKFi1GVCDiwMc1aFrp0ekM1YIdc0QEOQzNrBnA7HKMUeRiOK5x9SG
kSN/P3FO3WEGT3u9BUa+Kvazs6JAC4iTtkewHypS0gbROkycNszKcEkFIeUDY/Ga
9DTapAc9Y2puRQWpFnpnczEyBQBqMEDtJF8eof15mqwDQHQn5XvlBxlihtw8P5Sf
y4WVj1TnqafewcowI1FCRb0WXNxqFkozbYl36ogB/m8eeIEwl5PN7VfdzNbGC24O
V4hu5G8vbWXAyvks6ns9cMmu8IVsV8xHk7cDgkQP1Zc8DE1KA0BDdL8UQ24prvr2
ZEh99k6LEZ9iKW/1Syg50wKvmUxqbbLRGT6olbh30X+DWJgaIvKRTy/2uYkOWa9/
RWvrOF82beAEDuQgOZCb6ZTijhpJCmUub3UYZ44vd+1x8EE4We7LNAzIXON4v7J4
VAd1KgkTnnDtOWd37EHn2uow4XF+AK2CMVTMvERKtsHTjs7Ikv13d/FuZg4RgWqs
6Wg/B1Ve7WL806eQ3ZaZTHnqfpLXS5iJFdH04+VlZ6YXf5tgN6AQ3rFrK21o2Xe/
ULy0inLrNkSCbthcMsljZDvWPL3X9QdFWkwey7jsa7oSOv/qqSvUcCymEAmp+6NX
cttjEyfuUNrxwzV6UosGKdNA/gEU4TxXif5YmDicJ5oqN+2l5QtcpczXWt7mCo15
3UmffVpHvG7freWBsKh5NVE8DF4+RwSrRWLkPdwJ1fRcFXlqGNkaf9WPCvK0+FZp
gyhEEqxAf6FhBzdyjwgL5QdeMKUBPlcY0BeFofoUaVrGMJ4Mjs3SJnle6UKLfdIr
2tlk4GLtgoljduVBjDUHPZ7vy/CR6u7L+fSTFiXyoeUXyLy+dfDZeZg3fOa65PaE
o7+Gp2p5aaTcVAGoWL8dq1+EVHdKL037YlSMvAkQ868fNFB0p08NjI69ZqdXUyM7
Flo8fHPmgGzzk0NfJ1YHSV4uixq6HXxaUwyscmNDfV/gn7lZ3rGSzTBaR07DdASS
0zG3A4giG2Qejomd72cWkCAECqRPOTzUDV5/ALxABmamOmhYJg4DRamJiYp1MlfY
EmcnIyA5j6Ro+BNDIki6seaWwGW0Vf6k22+Y7AmESYbu+CzyYTROblfragUNDOKN
MZ2c4DfeczLh1FhHImYtBKbWufTcn+fLqnTJqMorZSdJz+iNCgLjbchvvd1ld5PZ
dBsV1zpG0OL+5EeBuhlF/DnLctEco9I7HuCW0+WhxnqUX4aPspY8G+4qRiwcC7S+
aE0BSLn5LQW6xSXfP53t8LzeFXfb7xGTUnrmCX/0p5kn0rVqdNFKbKNLQ7CTuInk
v3F8jCzCyEPm33i57lRilpOpAUxMe4WQocK6hfUqnWQSV5XkYMAO46XOaX1IcKaC
6xpdNUqs93d8fzUxs62j75+rizAVUYmzRH0WK7XyhAHjkAJP3uxE3nG1YqKxG+Aa
W+A3rBa+T3ngVPKfYLlubvvgT0u07QSsPnsdzIsRoPbssJSHHgOG8soY6YltdQpH
uL+82b9ZFs+hgQneD0ha7SMD4VubwcUgkNQ+hanE3n3htG6vfSc+/tPNKB69vfUz
MyPB85KvX9GE7QDodZQ28c/91MHmAtiwTa+Xk+8hHaQhMfpCsh2rb0FSeH/RSEUz
Q/Xn+zdgVTb16rAbVQsKCaOVib58OV6n3kAnhRIZ96EkU7dRmKH7db2Su/y7raGc
b6O/sF3Ej1CE6rmQxY7gLHnOYGMxCUEYbYpgFoaec5otud0m5Dc3wwi/o4YSbJbs
Wy7g8TD1NPqI0PiiG1yzgsTT2atMxsXmL8b5EoALKEvgHrX1+O4mPOs0RaKMhMrN
YCmv1hQh7/8aM7lL8qhfYDS422qKhRb23OmkJx93nSjZDiij6oS0HP7qAh0ny3Cs
EpJ77bm1yidjVvvZ78v3CoIYUZN3b9U0FBiS/O+2jtqe5wIC+W4jUF0vuLt7menr
Fp5MRsAK2xsVr4MABMx2ucB7ukJi79yYuzu5v7Hev+VeRGNsG2+a5IYt1abFpICj
ACDvoB1HZUb2wyn8R+D4HB7ATMqCEgMm3iiGnZELnH97lFBtKu7Uq/D1gQouFUdd
aBMLIr3zi7zo1OHG9BHEXDDT0huAtFhGbeTtCIWKR/MJsUJUrSl/pJqKQy4EoWco
RFq9pNpEK/VkX4WWaHXLk++RDbSbeI0I/A079S6Rzg4+m5dpZzvrvjtkIWVlBZ/g
acCMZxLSvnrxHpK1obC5z5obprf0CjeGmi26Xr9YYKXYyc6WzPOuqHjvONs12lmB
fBBSui5OltIAqWJGNmzXZ19c8EF8zRPwSHdvnWj24nqrb7aqIi2HyAY4tN/ObrGq
/sBoiyij0D53OI2hUf6uB8yIBnUhMyWUSIvjluRm+g0qTYpuVSPoDUGWSOHJGfPw
X8DbtBQ/6TFxQyAtkzXH5juF2F6ugf/rfL1UUeDi1CPU0TR1Yut4Kwt2kA+hPzUC
+ukTJICAIzFxXdKs44Z5I/WpE0h86iz1X2SUqZXMBIUFOdIVPFJKwOzbfmSb4Xnh
W/tS/o5fTo8Det+tijSY8djOeO3mMG1fhg97kF0ttwD0NHa+9qIexZIINi71IR24
6sReJ7ZsH3XaFdqjGXwPJgC5bBVrZeIYheE7qecfJrOp21RJm+cYhiZ6IIkd5gQQ
cFKxfNINZ5aG+7SSev9DOLamGLTZ7wKug4FpfGxEffQT/WrWpD8YP9uaszKuKX2z
RCrzrwcbPl2S0dEO0S384dDzYtaXI5z5UFJ1urcgA8jz5MwR9LHA66hcZFFekObS
vrVnGv5RH/vrdyskR/ibCgedcBKMpX98EgAhk/jd7I6KspvyZHzXv866oTLz49/T
4YlJZe3y5DGANi2Fzzmq97LQWGvemPEBdDWvxT4UUG+2q2Xxlub38VS+TUZFPnnZ
DfK+3Yfxzu6QuwpGmmQxFcITtJ1qo6QDKTewM7pFrRFMwNqhPnqZMAlbGLsPFFZF
RPP/pNsYUBcI6z84MLXNAilLXAMKCOI6CjrFnls0EdijxW/s0v2C5jQ7SBC3xQX4
iozI3jO5NXPIHYFiB2G+NvUJzHAtBukr1Dze8U2d3uEUlK+x21l/6A/9v6EMU1O1
h/ATBw6+i6e3jOLbCRd6dpGdIZ/AH0pX20tWIeyWoEp7ITUJXBxcrxcUq1ms9b1X
crcs8vyLjlxGoiYZZnEqGEOQ74t1TVU9LJwZrk+S3KNdSin+LcsbLW1GzfkyCebw
mVZal4oXQNeEmFix/ZSXOToMHAB4oiQMZdtLbdTHTG5IScrvdMRvjz8IYztFp8MF
183MkYAnmV+feEvWLJShkAvZT4JG8E4Rbcg1acuRNmFeCY90g+bMqlNs7K+PlEF+
wHKfviUXwARTGS+eK5Zq3/b1YoeTOZGHN7jRzmUPTu4E6/3LdTd/PQER9fIt1e18
SmgXkeEfhdwFYK8aQkVACJQUrJGibNMvSr+3iLN9q0mEdPxZqxFKOPzPNILdsND6
nG5F7Nnz++WxKK4PuAqO0W0fWdFVLalzpoPIPGGHSBZKmk2cw5Zf/4saao1eGqws
SyxQp84BEMaUkkDaJLwGpFgZoxkVa2kRT02ww1vIJv8MQsadmFzFNCbTKnO/5u8J
+Vmzt2hx1iyI2KHs8jM8wg==
`protect end_protected