`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
ddtXksX2+yylW5zu6QL2Lhnb2d1sD00763mmSITNX595NcHTEkwn0zB1Dry37fOW
FufOhVzEJp80NC5qZ/+F0Vk7Ik02dIR0elf3clrjeJRK85K4e3Hoo4xn7YbFUIms
l/8VZSb14+JVGURjfswrIyCUotIzlzVYZ6gzoZwDXIi5gQIBf/gI+KxNXPaKV+PQ
Ufys/12rjO6aI/pPlqSm0hCvftmBcnezN2hk1UeXgOIuKZnogjOsf0iJVX2aOOWE
6pD/psybjbnsNB6kH5uFTA5frkzIzkzl5d9+YDm9OyC+k84E83I/7/j+rk4L2dah
QJOvksSIzN867/4Qt8qYTQ==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="MvBXkzurAa5VTw+1JJ70nePUfoQXBvZOku/SMmg4TwQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
oRtzZL4VJ4iwysPsC8SXYCzXS8Fw2gtZTOskLcDV+1B9Nzn1zTyNtlo6lNICRmmK
ZRVu2BmCc2G+fmzynYlNTnSa7C0Cuel6FYpxCBlOuk3OF2tzAmLAuDyOH3Z1Yjzk
a0aHuoCdIRKv7BrZCdALt03JeUmXKPdOmIlkVGFl8yw=
`protect rights_digest_method = "sha256"
`protect end_toolblock="Jn9CQpRhJt4rnzZPRk+dOpzAubz7omckX1MrFd4p81o="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 9024 )
`protect data_block
gD6l00tciPUa6pDNTk/+t0OO0nC/UTtBwLB41d4inuAUA3i/ALrNyoJVcBnAmEQW
ptbcNp5fxEUJjnOxnedyZEuEBxWRieZFQnkRdF269oM9AG+WxdR/X2+jApj3WvX9
Nm/hq4iE4oZB3bVnM7fmqCP72b1X1Ckwm/nzFV7GxrIBA2mVFAR9WhjqT2w3Qilt
9XCtPXJxJapvsrviFU6zNRHCzeZFfrQU16pumKBS4Hr5ELQsAWyRGj0sW+sq4Nfg
MaN2dG2sXRVp9pA/EIdozRPO+B8o+3Kx7yH74YNL1AwcK5vXI0imZ5DqWFOPM68O
dkwSJGQ0qWQxEwqNJTDcg4nq2tCOTLVMSvMsMKDsHFPIi7UbFXUtEmMwbk+PwNtg
OQM+f87ywMkNoad2L5gMH2vXVFqCKLGAcBjvIYFMJF1ZLJNzbYglh8sJPuuJYaAN
yOWdP07wknoA4t/IR4obF0mkL7y0HiRQy7tbubYeHfO0jJAu1kUwv1GTKIZR/QwF
s3gYXdThNUCmA846Lv/DVz0USoriNi3bAfYhzkRDjKF4RLTAIOLurc9Quo+lJ+wp
kVXvZH/UxsQFROuA/1v/ggH0TqYxRBBcs5dPCu2K+iQmtwbrplXZ2KMlze0OV0Nq
xOjC32kI/9I1IoZcOFeHwrxzWcudnkpjQCQkrCE33RbRUXBgVqo4bvLFaUj3UCjz
bdh3Bg77bvoQONeh4nLaYDXdrzq4N0hmu9qfMigijm/HxinUZ5ErySB0YffhhJhq
n9dhQL9ELsBnPYXF4pBOlqHLmw1bqRvu0ugKZGRWIRRlf+BHZxyV0tWhduIQFcNW
LjcFx1iyQbwvXin5Opi8iJirUulKVXqkuETullVDNs/AN5s0kZc3LBNoriGox0tw
bwnSZ43rJq83zWtyElZV2Gjlb3UoOQBMK7+06S1bVKtREnw7LwWzgWsB36NUDL+h
gQgwLsAV2kotC8xtEJ41qJOqtLSeijRx9/7pHE0itt3nmhVO0OtYvcz0Xx7D7bkL
+Mq4eRvCA0xOe0DHRf1XTr4juCJxH4TfdNPDRIu3tHYO/ltxkOuP1kGvmQHn5z7q
bafRJXQiJoUf1bq9K5dFOZCyRI71N4raQhXvsrQ9k2WmYrKon0He5YHxmgUIUmtY
SYvm70IFstXzZB0XUwG4e5SVlugP3LAT0GaPL3Xf8ITJqGwtphF8DdjloOPenAly
bMUVqXyKot4Y/DC2XUWnylq9p2ZdmqKisfOi/S/YOFeUaV98Y9tAr5Z3ktU5tIEN
PAKTNdTgjHLziCtg9FdfbFy0vifLlekIAMYNNo4zKKJU0KVSKef/139uuEYOZ0Fw
rK8S30qdocXg6DwLUoHdxy5J/sEYv9ywy2w6lQtkxG3LpTKGMZhv41hXTWw/RaWf
hI9bpL6KFORiQIOYXQV0hkHR0fONYGp2ZNb5nP2Z3GcHAaLYUHPuoOpE7zI137uS
YdGrXsYvIYtN2BZVAgiA6j/sWFzVESPvvXU7vRH+2w8UUhY/ihoNsDv4y5c7uvuO
h/KeBBDaxkQAfNufH3s93LlQFphlC41coYqI90R5Zn0QoK9N5SgfF9zwCcS036TU
5Y7/b7LDeFMAAKdUWH3uvc+1kCCZ34pnjLu42YWynPu9p4kH5kXRzVPSaPXL+0Vo
xk3iSM0A8AhpVCATuXWYKYUXMm6PwpH2XObVrMbIXfX7a8YDZyi3jbi5iGONuBJC
gpH1wW66tC8Lv2IkwFjNyGt6d3iq4ByY8hHyNb9FKk2M9CQOoWyOGginx5jygGC1
2aIAF1ggpH8SzvNX0ZloCvlkAgJonS1uwPgcFYOfoEe4spceIESiChXyRw1JmF8q
Zkdz5vtZVo3B/8qoarCEblN6dyMpHuU2QqIz2Pku57zZqMFupDNIPbSseHxOxltA
iLtzfI4Xs8fRdjxmUYkneguWCz4M8r3p4RGol5dDpUwXAZvvp/k5o96bzYrDQlhR
M0D0MNtLLm0a3hH+tBnObK2KpWB6fg3JqlXsOlSHD5Ec1ayPIIJ5ApNtEI3BM4ES
j5KF66Z6AxiMcPlBxFjn2AqV1bYBzwQ6sorOUgHh9sC1VmD6vT5Jr6k0GNMfZ0l6
uVMCiiPnIqu0J3q2vBzeehinGLr719aDtB3GRYe87eggKnKvxF6t8CMECtrnJ53b
0svbzyu9AQgJMIAGjgtfknRo1min8x6fu8XnM3Z+Xja4gwS2wCirI8edtLyBe92M
KEyDfauaoeahe0HSttPfS41b/QVd3bQkCHs/ldsCh0IE+nIurwj5TmJOcoLmwPMf
WsC2aZsIGUXNEv5xCRUIZYQ0Hr3Wfo1zDxRT5XWjdw5R8wZlH2i0In/6EUkwi59g
truNch4c+hCdx1mqz+5GtVbnk4BJ41bS5pq5AFDWcibCmznDGaxZmX/4CCcECTUh
A08VIhwdhA/CwLQu5ALSWGI2oXiWefDtF/kZhQYWxMfxNuWe1V3QXfzmazvVGhhy
IKelG9D3GHXrovOpMTYLklAVQDxasBq7oA90LLF02nEMh3obNQcnNrq6eebgfoOl
quqtfDJ3DzAg5NgEyvihWTuk2dD4sg4GnOmKHU65OouJGKMNa1neZualqaJv4qZS
ReffPXVY6fQoLTOBxYiNWYwsQmUcHqWJ/opa0pSGWR8P2k9BdpTXhW7fCi26htfX
X1COyHbrMAzjN84Ddce/GCpx5QxcyQSn4BXUo2+3jJ6x1RfWE4YJsz+NGntL99r3
EcTF6r7IdDRBcwG0BOMqyhpDjmes5GBnQgYSltduV3eISuw6TL30BdVfODoEsKBJ
7MSPiZZDrsZx5mwR6KU+g7VZcx4zdJFJY/RdR/GCAXdkBLkbvTq2Tje2vtOlbsAC
oZ1sY7PjpRzQjoaTMfp6+o8S0rZK99YlT9rGlluHXXpQvMEoEaQEzRlFW5Qc070L
oniQ1EntAIcGbMcNJ9b6JVXPlIrT8De2sD3SOrQo1TfD8jjkA2/CIKOc/SuuneEy
coliS5Fzw+LjhMQAyXwi9PbcyaAu7ErPlAyrSSxA/tM2GzBwwUItNIKf5Mi4i1ik
Zzuv/BnNHA3CAczqydC+QCK5yhN5utjAZNYDYI2HulbwkgWncMNwIlrNfVmvUpGf
k54nIByfOqw55u/si6OMkvg9mHu515iW7zbLbnYro9l4MeG7ZeURqtVzcU5UhU8U
yIWHXD+q7qvgIOYxCWrKyarxVMjcmkDunhPRf77Zg4YOE72x3UYYY9MP6RBuwEYA
DM+6TmHitn5qD7YwqpVXbpVQGDOR0FY8BiuEHpnOpFcTbK2cgJgD1529PB3Z4QcG
UkplzIJ2i39E4WwlfEgLE/Orn2EcF9YUPeGDDytMZG5XuGCujLimDeFW01E7mULX
9+4F5jpsGRhfg140U3wL/2WU63Ly4BPUFTXdC2RuscQuTi0crX8v5GQ65fnYTg3l
JiiC1Lkc/WY3Cw52+jwt1IufXLPw/2+anHWZ4KEtV3yT96HguwF88tey9wyDfkab
ckqElWBPaxdBH7tlh560V801Rm9nKXeHixAyLz1aTtRD0C77km2HZxoVR2qSyhO2
feW/4IN2i75rrW0FGBU/CNEMLVn82SXeJxzqE3vep5/ICWWJtSJtmPgEXyTOi3+L
nthMzaSkalIQ8hOhY4qPEXRiovy6xmdPHZtfMOEJVBjZz+3jKWGu+QxHUdzYBInR
WiOZUEYaasEPhIaIH5xuuPKCC3Ij6W9sRF8GBSdVSkNnw1noZF6/ZAnfu3mVD5qO
veV2pQwyfu1nGcWruYVZmB5xzAUQMw5mGFn4YhcAt6JHTbL7xdplngW3EF9Eifkg
haTxShGJ8aeVkAeQrGCTHRz4EB1x/WKEnO860KOpMn6LJk6/8irqKSf9sMdxJi9K
CToS1KgTqp//dy1s0xCfHUXhvYnGVzc0WLi63QBGfZ5Th0u3Q3oHZtl1EJe+mdex
TBexFiRAdpB0tQTZUVDkPDHhzgYklN1aoc+bQpcrc8FkXrhy/o45jRF9GShv6+DV
CY/Dg9tONmU9e2DeXf659mInDOakEytDATLfg+dlQTeCISi0QYpDFqwKZRWd+3YF
ZSU2fJ2qMkOeYMvSd0i3letV9oCAYxNQmxT4YqyATSpj8ubEuyYWNDVFiIndYKDq
XFfo0f7ivYSDiUxRcvmdJxQsIQhMw+mVcTAgi+IAMHB55K5GbBKJbykH0cTpYtpE
naGOqS1sY4gttkCawlKAqtJ8waUjdBrqai8c0Az88h6JotWDgyrprnAk0sJ7TQXk
FKeZ3oIwl5hszczqNcumh4ZzsnSEMuKKGuRuOgBSusMdkeu1jZIw1v/pzgNNpGKX
OJ9t29MhFcWawOWWUOvK1zXq70psc4kLeYG2dwrApAtoHRWptplJp0B/n1h8OxrH
+eYC6YxnupK6gnT/OZk5DzydHu7Doh1alr5X4EycJsZdNbrSSe9EbdvzU+DXAT69
uW+2uwhbADeqVpjmKMlqfi0e73c/P/jCyJekQgbIwf3X65jrhg6J3lP5+iVxmgaY
YK92jsii3x1cLA30A5KNFPXehEMYLogzv0T67HLFEhKBqZxZAJOq/C6vJD4x4qJn
XdDJnfV1GfN5Mm1RQGpbt3ASJrXSgbcGnjDyEGRGlRLS1hO5W4AFoSjTTBl67gol
2rqNjfxLxBGZ6+pct15Zmkilkm8UQIlSVHni/FzHXWBp2fhzojB4SPURAqyJbVjB
m5K0RcvIV6f26CuykFMZp82QB/eZMGQogYY0JADy9Nz07+SJyKf7WQXfcFM4F7YB
7Pc8rQKzBNrgJM3VqC/slFE8eNEOghYgFv9XMgBzdO2H4uVcWsbeJa75tNnzXyyb
OcD0g7ezWGHWDGVAQm4tTFjaUWh2447hRS2OFeaiOLSTaq4i1NoHlDs4iGY3LJps
Y39Tedpq0hyUtF3QsCSojX2RE1Q26+CCXZtTzu4J/Xe6vHckLEJMQm67+zg6+Sem
Al9J1RwBwoWvrHtVl3F4QDLDrq41v/NHJtK4qtmuSBetkFAybH+HvMvs0Rgf2fai
GPc2fw4KPwnSd02Vyh3mYZdj4IEX8/ylSKUa+7qEqUqwRaw69pGAZmUOad790aA9
42r+0rM64VKdVGbK0aD5jdFnFJa4Ktd4llb5fxG1zMIyuKzzQ1d2t/O8Mf+h7wsh
m24Br/fvo8+a6pPKQxvtNkPqBIxe2etkIbl3EuRv99Waf/Vzcwlj/lyggRZ7a5gK
y+kFDh2967HwwiVAKkOUpBtW67dx17tFT2zhsl2eXzKpnjieC3icwKoq1YYM+aXD
J9/neJi1vGPxg27gcRrVeTjFVAxsbtnH8gaceKY6/KQV0HFsSW8b7jh3YLg76SG/
w/q4+pCpOfmDk9pYqugnPBqgcF0dou0CH2ykN5RCFcQRMWwwLoOKJmXpSkgR86oW
w/VxHp2uMYhoFhYnKzji5fmDM6yQj0uzHICg03hlmYrS0o8k05xsrcnTlmrCbaqr
jOCsZ4yeLn4+Zgf7FRxQg5Wt/c+tG9X1egejP0F0EGbeDk1I5CpCj5Kx0AdJL1Ib
EAfcCJ+Zv85b8kGVDEDX9eqJW65EXD5cFM3mB1JMykpk+3rY2aVZRGOUp0iu8+Ww
i/5vlXAMc/leOuY5/vlO6C/LzH+qjuhK8QgTc1SDseE2zWROUTgh6nhJ4N3qM2ud
vvGOIaBM6L3eQcKVEaQTZbwa2T0l5PYnYoc2aniyNodUPIorQNs/gj3OHGLz0YWG
FMIk341TfCWDsWBjAnpHwhAowDvTbIWXvKnCJ8TXF2TZs3MovxsFhG0E8jPG/Ts1
Q2Gq+QnMcs8o4c33S6kbJr4+lKMM2cPxgssqmXzVKeppABGsVB/JPtTl44huoo7o
LtGZDO5pwPXVsWlat6KGPXg4FupZUobIYHv2xcMtkzkRpR1UqqS+waK9xLkoSpPM
0p4TJWWvH92t83y1AdzXHfnpWx4pWA1nqY5RXw2VPsq5xJVV4qvf2TmDyeUx2fn0
/DuaZd9Q55e4Og1ZdTb4DRm5lRWe0aYKaC3rUl4zvkMVaROgukZKKDAxoEWHTutv
AMWq0XPdztiE820Y5Jvx2fjP8k5F37cDFZNssKDAZXxYpIJu+z7e6AF9CmfKgcn9
haYmtOij/I5PvR9x1pVQ99/I//5IwKhnMoEXYdc0zm8lIlKNNoCe0jSlavG0Zz7R
j1zxbsRafg7M6bk86wQeM8vcuskQbEuxbdGbOMy6vzv1/atLr3FWtnIw+t7pX4db
MJQLyZnp8kEyvzcuLhcCNUO4iZA4ofp313tjhqdxqcixmi9Z4Kiz8apjHI3uIcVh
i1kplv5H/cMYrU5SS+dOSiziMR8nh51lHWe7D0ixvUIi3o7xrj8ZaNAYOfQM+EOJ
S2k+ZxhRNpEj97Hbq/bV6NAvTQuS0kfr4kwKZhhk7a5m2GAzFNKNPl9iSBun7TsP
GG+CLAD05oYtLjinp7WP9M4hYPkoYiB7vtqtNTo8Rk+R51VtHQr+GW4aXTHIf8Pu
E/bRP+zVZWCd5OBEIZsXnENwqu8EXktK3nhFu6R6QhExcrImnjiihf05rIu8CUra
O3eMtWWP55HHQzqTde54Yseb30qjEU5wSmG8XKsp2jtQv89k1emkDGA65CKmVok9
je1ImvfXSD/f1Q6DtCtpxl0hwjG5OXyhq4fMYyWZdcbv8cww5xgRE6bIX8jpSWfl
8acF6rN2WRhuOxwvHfHLNIbVqZFWQt6/2cPHaXIgWjyHKfjQZ8wW2LlrNIEg5WuS
cDzFyy0CMJ2kQ2rlfL4nETbW2ciWmaO4KwkgW0NCYZJerE49RfW9ak7KbTzP3T93
N0/6zEohfE3ZKzbH+Lr/ASc1LndcbMHiI7nuW9IkFDk+pLjggjbIHHKjfwAB+Zq9
hdDvkcUx2jg9kLlatuR9gbcIceap9gZy8z1QhSm888cteukrK3jAMPUF/g3POSI9
19M5ply4vkqWWSHUiZSBLxGWuPSmGmjk/gGIJK8g/wcGu3fBHyEwAgh4jPUzHrwn
iO60EcYWIE1TP9PNbeK9OFNCrLST9rmxBFzbQlPqD9sDFdbQx25Lj9/B5aY20Vhg
iNqH8TvjBWqiRE3DtinyKh490nsEKcX4iQnmt/ppOdEiE3Jw/zWXRXI5SDAJzQD3
5iV9xrNi311UagJogWn7W3lMaMJP8wAgF3ptlCkETd+UFcWsN/rTjYjvz0pgB1kJ
fmzXnpadxk+V6y7Grhd9GWXg7OJsk+MM49X6gVoRueOBkHcNQkorXmk0YubHc4G2
4fl0ukRLHOkpbN+OVVEnq2ntidhZBZ+t/Gx2Vn36hd9fVbcHsOKD3ALNY7cpB/5Q
CJKfu0nxszA2J8foBC49sjnkV+Durqw3yJupb2MZqvTkGiO/Jnt9hhf/DOdwfJAW
Ii+QgNT45Vwm+wwgBI8Hdz6gv22SUaxrc6784dbaZTVMpA+ZS2opsXztVXf9wd1R
iCFzOY8pu8YbeA850Z+pVbs6JjpPGbZ3mCJoerwe4lo8i0WBorlLPXh4QRvotSRE
BKDZesL3ame3vXiOrcPMYWOzNh+5uwjd0Xo5G52qjcWKo+rKBmLMw3XJxYqnkSxW
2Pry2ukTfrcCoyo7BuKdXL1BbJVLGOT/6K8FPuuVYqqjgyM8KqxnVNYdiLQLwMQp
PBbXycUUIWZjsi6aZVq4em/3YH7Q6zBukllz2SRhgmMOh3LGIwIRS4L8AfMYYnUr
jBlQQKh44udqGw515DJzU9Q7LDJLE0dQzySmVKZyCDAzq2s3FRkqZ3jRJelK/xYW
ZShkr70SM+Q7f7GsK09gkbqLAP+0U5YQkgsC8q96Vl+Plyoii6jrmrLJrbUcl/2G
l4IgsAhCxndOmQtIen17V43K8Pb+oLnVLeqBALPt41CZ34RXnYFkEc1HwqpXjkXS
XEzHuZPwYvE6ruAZIhi15G6RjZBoUk3MK7ODv6UElxi6xtkwj9sMZRp7JdUAnqmR
0NV5lakbHwbSwBKK6gn9u7Yq1/thjBbjR2jvO1tYUBlSJkkC6ui85P8oN0qU/+tE
BnZGQan8pmRzRsltNElKrgLB6SYWdXgCvOHr/NF5K86EYRCCVgdjiY+gX0iszSYx
CTUehgjpUd7oi9kRdqb5lSE2rESgrYCh0UaU/5P9aSG3EfHEexZj8RDkDxt1+6xs
BBkL4Gn6BwGRhtpAMupxtQL+td9cmyhpqGhyUdUtVQ7HuVFO9Tx1Y1Q+dezfJdTW
pCU5Ynh9DzvSbOmBaqZuWgeCZH5qAZJcLJu87HPlFFr7qeY9ThbMLNHxuXRAYw3k
3QWwzbfxCR3E88hd2hrRxklO50MlnfxjvT37ikadanyoAnvpRJ2XA4fMShpXryeS
hAA3Xv7b9p5MgsAZ9UNTFnR0GnjOvCYmqKmSaG4R6NyJaW8qRcISzSJnyY54zkcY
fYRBFezq9RS2HRYBKwjFNKQb30LJdp3UKy7rs9NH8LVvfb7/lou1l2Uh8IYStwTc
OClJFxEc+57XIJsY9mSloBwHrbZIlrbXmzuhBy5UnOFHA/wpRsjsBkodKNB1dU7B
CnZxxUMjcjxVlM0Kn1cwYSlKsxlBym03mIDMOYpLtLfELZJmCG18W2vqYJDmtb2A
EdV87Z5o7y89CzG8SOUlenHkoMnFimsaYJP52SGw3qXMfTZl6f+y+DNIUmG+IGss
8eyQd4zKv1dftyJ1DKdx22OPUi4K6WzrW7Fq3UrxIzFD+oMbMjtLuSKPhPi4rfew
uAH66RknFjuSpykFR8Hhjm/EWRFwZXVJ1G7Cx6sBdiH4rdnDGO8VARgJ35mUrPez
3UCmuetA+CoKrKgsfb8iS5fylnzjlIIvLsjxxbqakGYcO79KrH42lOkryt3yJirs
SwavpXTCMejYN+gsTrBowEfIFYh3pgtXbEYvHACPSNokMZGTSES/2b64be22ioHt
ZtOXvACLzZ5Q++jFuzCkb8FWOwhYVHDaOoIxYHJUwkjPPWntwXJP0Bqtwd7RQiUc
bSinC/48sGniymuu9/GZ7sXTEGJD2Fii8hJ+EJIEqxBc7PEeCV9PO7h+AOQfZdjo
E3drQTAld5ZEnvoS4tc/WoAq7NDnmFlzt928jeErF35ierpsqV8Oi0bLlvQZM1PR
uLtWVK5lyjcV6gIcuuS86YpRQ6OTpg2aESbBrE4APjjoItR0AJB3BFc8gtceExZj
hxuklwqfqy1m/bnHUdcmB6WU4vtI2C2kmolBjAQu9bnfAq3hRIsjdTPBZ+RnEkOI
ig/BRtLOVQIAkJ238V109KXjkwHh5s/HOVTcUgUaDgO3ZbSrjaw63plo6w56bQGB
n9iMonqrZgTWPHDGEBAal8gpLuGWzG+E67kfDOucwGFjjKeODZQ7PAUwjyp6cnO4
8oH02vZByXdQb/fbOkr6178sJ5qiH7g54BOl6ZDew49j6poe+IGGc908Jc/BlSV4
3ZB22dmz+LJg/3UDgtzbSU51LIByMHOyePbz331/EQfV9nxa8X/ODJ3cGAbxNmtD
Aiw/oRWn5PAN21Jg5WsOhjhSuC1ug+cvu6bGMuGmU/2BfGoJ7bIhS90eGzRXx4Vk
90IY8aZSHMmRYTqTd90ROl/9T3csows8dawUN03lNMY/0OGJLLpN15L/CJVGAXDk
yF4omyapfDzudFk9TBhzJCwwD+cxE9/6/ZFRVzNX1Pl4HUv299AGMm4yLgEol4mS
XXizGn4YQNVnfz03ez3kt6yPxqQFysCR12EKLAaaMb6jke3qToZcCTzXcqQjQeGj
oJuYfySjbKkNzVGlU8UoWhIaEXlA0IL0szVTqJMdcmBXQLtWph3j7YhX/iO2XxDp
IneIfLXesLiEHRkx+gEV56/+CAS/A5/31KC6TZZv7D3W1kxvZs6AZuDWEreIwidC
q8TLFGVuyKMHuXpiBu0zUooAALQb8IxhLkD/iQJSAgbxWkTxtI0toIPwru7dGWap
F8C1AgZcVC5G2cwiw0Ay8Cte1ifUVZGVYdQlDcAPXolUMpaNnoo/5RhdRLr/HDkF
oX4rvU5U9b9TBBEgVHqQ+uaAY2V5wqzZB9oEO6f/2eyOyezXbJu4SmMdCDVWU8PP
SooLzRk8YPG0OIfAAEgnc6Cvt3CYiIgRy9aOF1goQp5hmCjN4ope5cSeyx36cvBq
ZrKq9IBWNQ2fVz7trsuB+1fyJj9WgumI26tAI4znI5iGXBS0vmo2wSunxsRYGVHk
0Qq1mfHiT4LT76tkuvKoLyyMi6DfkH0BektgSxuJNDuTB4qfIKskPeiese2zwH95
6G8LKdMRXMCIpEeTmFMTPANlxrJLj5xQDAqZ64JDPjhephgaufgGp024Zvtqto95
tkMfNyUKudmvQRzAFzMPG/bJtRXGDjQZifDV8DVHmGFXHoy+afERsr4eK/toHBiR
HC8MkKD0r6Id6vMjjzBcMsvAKtrbWeT6QNYv7HOF1RV5XRhFmv4bEH/rq759jRav
zbmdiDFPiR797bCudl4Ikxx+YtSTO5Z+WGDkizQK0Gd24vdWfD0901igKIj5BYGN
zZ0PHZVNopFKD2GsLcaeo2fhd8qwSrCHR2Jn8oviQvK7HjlBBytzNjr7DmMYBlRp
NUq1xmcAjuURz/NNEuV2ady7Qw86du9RFhC9uSSDD0cu2p7Lz3AW8c4CN7PLcg2B
ICKGqvTmVXAOYQUMAWt//Xwocd9brOKRlkXEf/pDfNIOF6dLdQp8l0R7rusgTRQL
yPGmGxkUfsOnv1kNHrjEn7sW5jdFHo1G8vmFD4x0TPPn7AOkXHOPfX80uTQ8Rrsd
k2LmH7aykAoCOD+AHAAf+Ce1AG9/xjylU0ezBkYHM80P2ChvJ/icFGsHLrv8JvT+
r1kfPUycsQe1EnR+7mvZ0jFM06Ip6ePFRIn7q25hxK+zeIZ8iEG3kp6qh/NZD79T
f532BX2nrLyUBivPFZQKK+9GAgHUfrvyU8OA0rNWRNPGO0lEvFcuIa4jaXsn9Tw0
BwygLbQuGwyTNFLwXNJ2mwUz/+RXVhBXopL6OOr2hRkgdz24I86pnDUk5aRvW+Aw
z3D0v5KTFJlqz9cZd3LT7wGgGfsdK71a+mAHeA8OvatGfh/vbFSbjBYE6BtJJXzd
gSpRSEATJxy8FDJo8K2PWg7QDCxakJS4kedpuqyLpSkTL/B1FaO7aiwnVgUy5Whw
DbFs4MgzsXGGiMJzfmfQ800JA+DL/MTgrA56P25soEUqgvaHQ7moKetassgDohnz
E9NUKGOc3EjO9j1vzNU6oSAA/Q6Gf11UmB5UJ+7GH3kxzsdRCfTfH8VEFBKei7S+
yFpFprdRo2cpbTXBW7JxFb7kQ7LIuevkiVFT2TT7d4naZa0lfTl8U+k9da5AqKTR
Uy1itW+/6fr2u8DhQjKgpXXfG1/yjaEEEBAahGwnB4tucYYVZ3bPliScanSZ97QO
EaQFHTSCWaGiyTz7swuFuPSi+2i+4vO4vQaGCUhXy0Uww2FNCsRetgDD6+N6NTuT
jTrlvoTEWlv+X5T8iO6rtd/R+yipFpLZ2nfYQJSn44+d/AdPBbjmkmQsvwIeJQ46
lSCSAK5ijWldvjOGK+YpTNWjbbjixNYNfpJ9g1lLJSGt9btjLqoLocKzMAiMKckY
wjMY6WP0t4wgA+m3BcwA1uvGFy1DF4Q8Fm98UJJpWWndXSIBRMoS1nlKpK33rzPV
go3rP+iZ7jG+QjqVm5yGAH72/pavJCeJE97ZKcPRkDx4yiNhLwutuJrkMEUopkh1
ixWj5zCQl+7vPWcWz8yonkHpJq1OgsKydMVKzjb+Ed+vDDgFEMgpdpQ3btMN3T+t
Cchq+KWyBR8NRPovlmG8uUpbiJNWq+ZvkM0V+2tAXikEgkOffL7HfTr9CevmC79R
IHv7rh1L/iEhdyTAYsiG7ZGDQ38ziuz8h2picIO8z5JP4j8VaPEH/lTuOmutjtQi
DuvuSKslVXrqVBh9S+W/huqTfMJyHLQJaOqjQFVXhL38Uf21a9wnHinYR/yflveY
`protect end_protected