`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
ddtXksX2+yylW5zu6QL2Lhnb2d1sD00763mmSITNX595NcHTEkwn0zB1Dry37fOW
FufOhVzEJp80NC5qZ/+F0Vk7Ik02dIR0elf3clrjeJRK85K4e3Hoo4xn7YbFUIms
l/8VZSb14+JVGURjfswrIyCUotIzlzVYZ6gzoZwDXIi5gQIBf/gI+KxNXPaKV+PQ
Ufys/12rjO6aI/pPlqSm0hCvftmBcnezN2hk1UeXgOIuKZnogjOsf0iJVX2aOOWE
6pD/psybjbnsNB6kH5uFTA5frkzIzkzl5d9+YDm9OyC+k84E83I/7/j+rk4L2dah
QJOvksSIzN867/4Qt8qYTQ==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="MvBXkzurAa5VTw+1JJ70nePUfoQXBvZOku/SMmg4TwQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
oRtzZL4VJ4iwysPsC8SXYCzXS8Fw2gtZTOskLcDV+1B9Nzn1zTyNtlo6lNICRmmK
ZRVu2BmCc2G+fmzynYlNTnSa7C0Cuel6FYpxCBlOuk3OF2tzAmLAuDyOH3Z1Yjzk
a0aHuoCdIRKv7BrZCdALt03JeUmXKPdOmIlkVGFl8yw=
`protect rights_digest_method = "sha256"
`protect end_toolblock="Jn9CQpRhJt4rnzZPRk+dOpzAubz7omckX1MrFd4p81o="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 16464 )
`protect data_block
gD6l00tciPUa6pDNTk/+t0OO0nC/UTtBwLB41d4inuAUA3i/ALrNyoJVcBnAmEQW
ptbcNp5fxEUJjnOxnedyZEuEBxWRieZFQnkRdF269oOCNMEPTIWFoKq6EnqJqNJg
q4JWiobxVRxQqdzMJNnly2rICsuLSd2+p6NGrGFrOlnp6L7PU+N4WOXGwbrPrW+D
p3q/VPOolvjuLtvFw8YASphsJ5K0dkPj7ooLzjdlbZWlCRH/QunngIwneIHCSjVg
/HTaNE512bs7Xq4E6rjWTJn+hRe7B1CUOzndmRXpRxDwZk1u+Dzf+7UM/BLvEpFu
VjJSx3UIvDpzz2CF1BWvmxRdTxKWbN7GEgQLWjvSqeXXZDKUNVnn/ExNO3KqQL8v
RuvUfxbjaKSgXSEYZK8GE7jduNhqoKC6+vTysFT6ce/9caqMuk6hy6yqwNBPmuVn
yjds2q/AtB7TVnJ1IvcEGo1cvVRMf+8G6XVzLksJz0fNwfjOtHVSjiME5SwE6goP
aXUkIFc4k9wJUU8ucjEEoIw3D3nLwS7f44lYXuHV/wkupGk1qN5bKl6vj+gS9+HY
aczqdAnYzBTBmMNi5KGyN4IounMlzsuJFqPnJ1/sgD4s4kKhV5pywhU65dV3FuZS
qpRJeQmcynMOw4cpymzxhOFmjy+6XShMvSWEcNEyhTxijm+be7sF2RutFee+XUlk
VE0kT9O8vwLIoAsluw+kVGU9bRnvtEGP/q34rmGKqzE0XIXZqdqvpUpueHUNdFG2
Z4RFEhxNUJYVZSAUyNbva/nhZG2o34tQpD/PpNY/FmnDbke3djfCICXyeS7DlgM6
l+3OGbjPjae/qjT+MByi/j9vLfOAVZvcgIEPb7iLTV0vi7ySQntbRZVRWVQEvWMg
QR5w1FY+ESP849HGdrdem1nmOyYd8QjF2Yiwp5zT2OimFPpF1ecAneZBY4iTIgL1
FqXPxQA9U7v9bvfE6ecGFjfdxf6zYN4CXfEJeg5wMNS7KgxL+P3W3sh8uYZquEYa
RS3LbSW11nZnphvoC6l3mUNiRPdCcd90G5/pqtx521hriV7w1kvo1xelDcxo+lOG
hFWRShGnsGrwoxgtlFq+ymfjC2T7Sc2M2c8DkIG9RAiW4DoiK7cDhiJoXIrxHLqy
6q88hNvRbnaK+0gaudvIBVGvi0L4zaSqnQJ4xwwf9VCBAADiGE4JCQeRv97Ef7X5
Ckz5ka7qsgY46DkdBwtuzYM/PmtVw2IIEKhJ1SUVf4nYnURYGFTA1fBtVPYNCwx6
jLjKjd+DBteakdu75dE1SQVfWshlpwFNzCDH9TiHg1vVF1hDeMpHcXUqJYU+bNXg
1uMhyhamUXo8FkO7JWr7avhMBtRgvw8cZ1CIKdWQTcCZonPXANFiEAQP9RJEgUeW
JZWn1lLe5VRHjYXs7oL/T7Q/hQv455uerPVx0Axlan3vsSmH5zOmKihLsXIG7bRe
nzFN3qaLDiBG3Lph/XvcxjNimiuEeluNjJ9BYCNc4z7JPqUPupXLZxTa076SDA7l
qxWJYKI0N20xmcMe3/ebWaNmlaH3IHusc8uj49c6GGzgCkB1hLZsRo69efgEcYKq
fCAisr03yK91oUGPAxU7eWebaPZr1B86sP+GOOJ+eqrVATGYlvN3BC3PjAs9cOXi
LYlA6wWvJdsPDMqXwRubX5LBlz4bJpCu6eEPa4knQ4DseoDl6blZAUjs8Q73W+/b
7QGI7LLW91zU+putmiBtU2MSjzKUJm6dqjBLaIhxNxRHcp58XpT+JWIZYyK8YNNU
6IUg2hU2xF6PMcGxRr2eY4AlE2ZgZlNDky0AGqPmR1RaC6nTOmEZELicSaniHbck
Jc5JED8CXu8ZyyP51zZNozqPmx29sc/euaoF99UfWP57F6vZ3bqFqMTwLoE7XrS/
CoWwcBTUX11KnuLNXgzsJEzLwqpunivgT8BKYemPVYUtFfEtK+Omd8F1aUNazW80
PVqfzOfCecjNlMxxTLyQQlQI3yMDTOBMkIYTt/mPKT6Yq9TYL3eNhTxkEwBO6/LW
q2RQx1XAn5sa1JTyP+bAwontnh2i4hD+gL8lC84RKfbiuBZDhWlaUe1ZdxPGNsnf
0m9k/igbxmOk6DHZ8sYNY4sXtqN04PN/Yv3G4nx6/gdmuCtT33koa07ToQu/gD7Y
UFuAB/UufqLC7V0mtKp0Kn5rvydwS06zwZVgNlS0vKsrVDv98RMNY8S60+X7krfT
ISMRLkhKKVO/KzoTcHpz3+YawsFt1qKfinn9m9wSdLQ0l2E3y60aftyoybEJI/5O
Gr3en5pUCoGaSo4FTZW+5+c6A/VUke4W/UquKX2Ct7vm9e5f/U6lOXpJRz+gfTKV
ZBSwKqlPC5hUC60WeiuHOiAeVtZCKoMhBLYtgpmhKyYSzM/P6++iVoRwtLAjVSj7
qJuv4q1vyVnWIwC0py2YGA7qzi22AaScuKT0XyIVMhmQFzMIQg91vJ9RL7Iro75j
nPF4Wa+a96Eysa3nk5t4gqUo/ZmNjcNXMfF0e9lc1qNdmIXkDAcyOhvuxRK36VHq
FB+T7DPIfOazIYfTUphdNvnbKQOUXFuPRfQozwQ8Cieiyz6FraQi3rfL+zhTgAMW
Z1yHgR8HO/TuvBRGCITIL17MtA9mBaL0EXtRTNt7ydgPqfQuw2vYwXxZCF1ZmCaR
hqJtvjbb6MFAB7p075i+wT8Z2+3Ozn2MoVbLdhSGAMu7eVvMd/Wy7LAcLkHxp/CZ
fxTSuXRAUjiBipG8jdUfIgeTgPGuX6XWHgYfYsc36kSAc5ml3zO3nFIwpJxZ1vFC
ejEQJLhSeUIy98xuI0TV5N5RZpHLDXtXjgXWosEWqqjicOTpCHCtGcu5Li3BrrBi
mebO4YCJzUK30OXEJo9oXLKcCVPHm3KZtWP0ZK/b67SBiIATx4OKZShguWCRTeFl
DZ++YpN3usOg9hFbtS96gu2ZAfaZq1gIMqiZxAgVFtm+acwZs9EQ4XCllMRR3vao
1RTC6r2PoKUnPIBceL0rkWCNNzC4H7cTXxrljFt9Rk8EOB8OMEdt/c8cF5VlN93t
incpJXYjWV1uNhML3DHCWLLRzzLGKxN9lj9sRutw9x5iBHuQBgg1ZB0Xf1qxvrym
hM3KneOvEeYz6/wJ+6svi5pigBTy+rMb4P6ZgIn0T/xQ9xixSFijEbUuF0DBbYGi
BsxNVpLRRn39eYi/8PXsibkjwp13oG841hOOazQoVFsH0NhvYBSl5uKOXe4ODe7H
vqFRFVcEKVbIk/+BxT5eOEqGsguVTqPpQsmyCl0G1bFqMiBl3sXdiMUL7L3qQZHM
i62pFokPUILKeDSjdT/tT5Rnn8GjeAh7oJN4a0xwrMLKiT0508aRVBLWRNeszQDt
tDpoi+4V3mZsRxSg2hrbTuC9Elg6ttVFXyjny06I0TzFtTsRAdn2R7fVqv40yo6N
i4pD8HJbxLp3gHMy595f+AmfmKvtQbs42XMCExpS6QF8/Cu00pbyHMcuDblDm0g2
pkyfX3jP1eSKqPPbSXFaJJq2c1RG3zsE0vS4z7V7V1mP+gxwgPb90jgMiL4PWERY
r64X3GsNYN7B0fMEq/zXsFeTXwpI7c9vGwe0Pr2rNOOhJ6yg4NpZOSpiSitglvqN
GK/RaI+fodhT1nqFxblj3Q+Jhxfq9B/PgUx6UctX+CV7oT6tZMY4y/Jd7LysJZzu
UEJWEpvq305oHvOzRUqKL0IExLOlhCmYM3h8noyjWy5VntiocCsL8pN5yECFq3sU
rd6zoDGOfEfMZJXHTCAFS/JmH+Z3W6DkTTR8zJfMglbLsqFfnjIfuLQyHP2RAKNS
N+vdZ3CKviXSg6wb9kLtRWMERJrmQskqJewOY+8sj0CK5U+epp8ewzMEfOtsPqQp
Dx2jxL7In9zsUIAbMQGzqG41zrWuxVoE386SoWEcwExJ5u4cvTpo4p8kbwt14Eio
eZ/8CA+u24+DUs8Hif74l3GpyTIXqjDm3EGo58pHuQWrlN4expm/2e02JJESQN8X
43+/isgHdIzhF+dBkfSbp/uElBLzgzUxdF28cYrBt9qFQJm/trl9ggJFekO8wm/1
Mckkh3Qbu5jc8DYCID7i6iBJI8lPq6TMVcpXQvFFTWfcffqbFHrnRE6AEtTgUoyF
BITbmb7ihJrOh7jXPxAHpDSAqUTK/xhpdETeZKoJyKkwzGLKCP/RC1/ocfXztAsC
KV4sF0FgdFvezm72XeCxhMe1kuw+EDA8pUCefI5iT5uIoezVyAVImc9E2vjyDoGc
ixpRl64WZICeBJOMJIkGjSTOFbEPExD4dkqiw+KtJKDc7CoY2Y8dVrxa9Hwwgp3e
DpZWyc/coS2prHJGkmHsHHrvqCJIljx53j88pfrTbbsTPtANzz4w3f9iS77e+3Ji
mC7aYMte2v8YVG80vzjBBCslqoyiZ5LBNN5wQEC6r6EYnrQ/WFJaNc2ZT5yNOIrB
YZdovkWxq9KTSDur0xBJ2qdes0Y4hc3upuJJ+gyXVXPMmSLrsjtk6h296dWtGLUj
ZcWgNsDpwL/Ere0LpqALLapbs//ZDkM9QPRQAcsk7gi9XTT9/x/11jt0S6z2DYF8
I6FYlLbHn+xvwyblATOwlFYDyNy6V/rbj9JEMd+T2WOgAwg0jL6r2MyUDd0QmZwU
YXLzFIR0QN4OHsy/D6k1c//kE9+s2o6HXBU81DTj8o0aOQquIXwSwzFMQxm5nmCM
9AYmAUaBb3QuUI6g8R5llE17kKUE6dZ/4soqvO0K2B7DbeU6KyigrQUcAqNIledh
z0f0lM3Nq+Oij/B0I1bopdt2SSncI5wwOt+5CklkHMMM9WHHoP/KYrGZP6U9OMFB
7Lo5ZLWl3kE5u+WcrDSkoFTkp2u758rWwvtwF7mdWirvTlFC1IV0hn7CmRxYttPu
ezUViSFUiKxgt1SN/Jfj55PvNJ5B4oE2eID0oxpN93J6J7/U3m68858NaDeW/Pm9
bUFtWSiC47ni1BjIj2CpIfqsSoSZSRhXCjVEsgfATjgDaobS1n0/AfbVQH2yt4fE
lovNqYNxk3HoGGlh+J3pUuLbWqcPSTmOQAoJxnVZ29YW5Dl7AtTLwNo0c/3KSEFj
sEf6MtgsYPxwngPU3qL18oh7ccOJp7fva+Z+c7JjUcHqskZqG9hGLCFndLVmaKUa
UDNw9k98cUFILBKIdgVB4BxhX5789fHkTJ/hjJm4ggpLVA3koQgzbux79yE3C6qu
bQxXqM7zzv9RKiqVCJyG5SIk6yW8OUVuQqmY1HtwSk1l8aVYUKqpFeAiLeMBpoWs
dNAB1jkrFD0DV0n/kGk3TAR7f7QhCexMIvYc2HlQVYr1EIdt6L4LSF1L+uxfgRPU
RBp7MokypKVFuq+z2EiIROfGJxgBbVxbNY3+LY/+JNC/qP91Gxy6ejaQgVMEyaMI
o2OiXo96joiVLEgi4nJPPot0Ihyk1J+MI8WheHwll2ojFz7/CmQ2I5R82IV265zU
uBLkfcjvvcgmoBMDNFdFt+riDJTXNbDuZU7+Wt+lzmlOiVryZJuF0FGiEeqQLftw
aSFBBEpy5m5U78MOfCj1ApxgDp5qkxwfhkpNKv9wcshqLRXWHCSB520hWa1Yn+3I
Gs4TQiBtt7In4p3vnESXCZuZDOqKkS2VznfV0j4bSvnOZy4Ge5hBPc5XtTEoxz+5
iyc3qNhGQPMfRXr0YdP+hGpB1/FY2taGaVJ/HaWy7zku6FUkzF5ZYz4esCWSTzyj
R9QXnmujv0kmZiI2Qu9EjAYbHJQiG+P5HQorFVudsxp2U5vdzWnxP7jkf6j4pwZi
alwoY3Mwe6YoL8M06icIGT3eZlgjqmNatY8IEZQnatwxp1X3a+ZC3Hofc/FyVvRl
xa55/azlqw5fXKJIfeOVkhBw1PqvlFVLUASd72f6/O5tXa2GBdaU6DqscbP2bQnx
Mawz6QM+q39IANVm9BsP3LC/1aqtg24osUqCRxNDY+9+PpK10cYy0i3AXBDCeypA
vIg+kwKvvULxfV8r1rGQAXxRPWzQfxB9x4LlheQh3r6MVkZS8Vmke1jQe25ECkvu
JKtQ4548IotyV9OyeDwQZQ8sCF+xyntZ99457GUVw5+Z8OIKszZ3/SeUo+vDzCPF
YHZlHyORJ14Mwh5Q7YuvMETmjAx6vof1aau1UFgyS/4q3aXJDzK0YK0+sHtIhcrW
+6eIdjsabG9Jkf9INJMlWP/49rxASgPHcTeuLE3JQNu2VjIcMqQd44XQ0xbWmgaY
V0elWCPNArei0k/r1NwWSnK0iTkbGhroBLvkKZoekroPEThccxfqQ6lS76+G2EVl
LfXVGl9QsSfEd9v5sGe94+r19cYsFrXb9rYuNbLBnbXlAgHYqNKKGeADMrFj8WEq
8XxULXnguXanTI/L4TNx6+Annx4kdIvklpWCEO6blIT3muw3TFBrgq20ptaAcO2C
rYKEfeqJ1tO7oiI5F9utKTVguRzrf3HTYpWBskHv9hlymT9HtxpAx6NOlogEHRL/
DWpP6/8qdMiUUd0ImsmYjXdands0eG45RmJPSj9gXjqYHWW0WIS+5joxrhZJDNSP
CsWAzYUoYqfEPCJ54VCXjZafzO/mH/X4gCClOLPSMcE4vyQzI0/tbTDcnNfQKNCg
K7ynOprG1wgjo1vw9Itz/rc1xFpuvTW/+gTShExGXQelQUzH8djNTfiHQ9dyswZj
BYIAxad62bkHf4MkEweavVdbj1FjFqEPGyKjoO6mk/IP0mmTFoHyokYb3X1Csu3w
W1bq+eDtRtlgE3JdiDw5BuemVMeo3JRrqE/3W7xPSm+JSO//rvOmr2uBy2xCZ3Zg
VOOdxrdCpLnBEMiupXYVyHWpOXnAevMBwUWDH/gA6WwGKad9J6QtN3arzBHrQz1l
KIMnBHVlAj+JbGC8ZLar/5/7flKO5R1WpVxCdv1nfNu67XYIpwUyjWZZBReaPKdF
ExZn23EZyGJSwVrtle69sMHIKu2NK4CdQB2Cd5e/5PRrTvVypR/es5iVzZN5dbmi
dDJJnz4O+avnnH5I5AtuD4TmOTKkTPXp/naKmf9a0BS3Rs/93YyYS2L4LGhuj9hk
E288hG1fMX4C7uJ1a3V4JK8j3JEUtickryThy+GZQWgguL7GHq2LG4pf/k70Fl2P
ZKUSvJ9sM1ghsZAJbdBZsuazb5t9H2Mwd0Q9Wt70ei+GfiRLEN6gIOWyjajanqkV
ayYcX3QWb42G+o9ePdsyFqVgosrQFi22WSlbAzfrhTKLoNcLKWDt0RJE1mA8vMd+
zy+bi7XsdYIbMosXax0sk2sbcYQ+pRknMfxDUQkMO76o8FFY+tHH2pJXpR4BaFn7
TqBXye95Tvso2FoAwwz9E9wQkjeGvKMPBqoLP6xq6kQTcVUx4bO1KXyOR33qVhKh
pHYqcYU1wDC+91pN77xTZ2gKMtGb2UOjoywgVgO9NVW0BiGvIZZRledE0+P3nWzf
fiLop8p8PZ234lgEboH/Sn5+1oY0hm3xylOo0SmadMWG81/fbKFfiaMBZETlxkgi
jrtVPkwo/1y7iFik7+kIOv7EF5tyLlrlaLDvWrbZP4PBzelhIFhEdoL5DTwyWrZd
9V6Ox/bNPHq+JAzt5zhoygXjp+a1oHzcavS0Y5e2L4rzowW/dm1fl8fIYp8W7niu
ZU2kIxgwTnBLAHhHP0mlP/j1WcOwqq54qO+Q1TuO9slfK+ilJv72HKVFo/dipoIq
ZyTw/AyPnhsJ/WDPpIH5UbGp09qWv75MUu1fKHypvvDVHRxflDdzB6BmBUTcfz1f
xNIu2tLqW3RnVXKEEc1j8F9cF+kI8tym3ORRLJXvupkU4n0EuvwesuCyP24BiTge
4NHFuDlPP1Aujfwxan4fXgcswt2EwEKtNLNorMKmKMdrhX86wKUChQRIEq/Ft+i2
3ktBF9P2R5iO6u3Z2e3i/8Qp8r1KhSdaxnRE0uAr9Zk9C/cvSRJbOGEwB3QWsdra
5TWs0uoimJESiTnIYsR37momtCJT0Kkxn5e5/x8x4dessj8DIVc6gERpsBCFH167
5+qNi2X2L2J33GY81M+3VVLGiWuLLrtbMac+aZg8v4dv5LSpPKZ3ZnnQYK4Mg2IE
2rhikBxbcfLBqXM4Q7hYFPQ+g1hFdhSrZighyCC56VJNYPHolS1h5NGnaJJULbfi
puao66QR2Vc4BlDB7GNK2NU4bqAHeij34B7aCb+jqaswK3OR8mdSNjUun5NfPxvf
yHj5qXKK+opTEu3Dh6PfMEUT8tdOdPFi60QjFC9j0mME0BmROxSRw5aqDHGmclrI
tJE/dKuWvf92M82TQ5f+w2eu38g07NY/G33KmwFQq16+qDkf68VblJLB+TZk4ITb
d6vjHieW9YClJGCENRIEpwBfCAT50fzyhrpJH+vGrkubXedmh2dWTo5H20KnBOjG
Ws0HoLbvl+EKXZv2IHJgsPH9njQ9OYFvTZ5L1rBdzkuULUvDGDrbDe8XhJlQBmHp
A3JyfXuS1i0+G/9/SSO8YlKu3J7kcu5FVRBVqjBOS5vKnnUdpFLf33Ty1MBOGgD/
5htPilDdlRH5nLzqDg3FodO8gtYgyfvkv/a1k4kTq3UYhTEuSNfFA7eKocew9W43
YF9OyaJ6OISXiPpAf5O4OqM1YUl3rQbLrP0VO87nL4AcbgtYu9zIldRr3lhTrBMN
640Ued+vEJjMZSrswJQRf1Dr3KfHLLIK/nsihxgmuY86wTpxmMfGW/55JWbKCokE
K3loWpMqKw7v2pH69/TwPVAtp75/je7uN3YLrlISrgbBts4RbeBBFOyc5aB0VXOh
0T48c9wEz9haA25rGykpbacp9UNn/E5gFXW01HT+DSJkpIz3sptY/Xtir7Kb8yxr
HrdqJ48BSLpQAFlWXBH74GKlyWO12OoYs34rD/65l6zeCtsOqk6K0Abbl3kLzCXF
Udwlpm2afSY+IclDHBposBvlK4G+i26XDtqL8p8GxraSSzIoiTGh9w3pnG8H0UhJ
miDQ4MtI6eEyrcfNyiWumRHaLUhsNCsb6dD16QT3NVc8KJQQrJvSTLFyHaeX2UBh
D2I2v4KZqtGCWlwErHnpVuYWJcAzjKfPNulCIYos5gqDQsDMGhN26GRPvgMgKmwq
FtboRmyxqbxTxHJK/J2yaolAKu41LAUcmkC06+Dtu3pGRGsOcS3gGy3Nc7+J0EFz
a1bHNXSBsEXhJz7dN7A4A9lqCs50rTvJJO+n5r8mfv9FrRfagznsVsaD5zP97Gwg
D4IptKknin8rfWioWxhsbZZ2H0mJMNqi6pNIsT1H598EYlLEo10zS1wrepJNO83E
jZWFKoqDQSwvHAB/rB8tMfLOG5ceRjsoiubzSyGADVDrPzCERcMC7JVwlVs3ZIUS
SDjFILl0vU0iBJ7be80hKmwzORkF/ChhIU/snlozBVQ3AnqrccO5ucqVhlV35TPs
Dp8b33UGSLtEUcKCpbQXA5nXpL5HsSy7sxcxHcfdU+tsJ3IX9XEss55MboMf7s7H
cE89aFnFzzTzfTmcmPfo8/s34M9bnWPCLPKT9fNy8OhXtO5n7ZhDQs6Nt+UQyDpi
PNVP7yohd1CkMV/Mu83GTPuDkP/sydD2EOY6961NsqZuvuYCofDh/bWtrc1ZK2jI
oMVRhmWiRf8c81rEgGQmD1VejndxRlC8PVjzm9g7XrdUUgTtOMGiLzWohybqN3vD
h8cyCyJ+CLbPElQUyttoAkGpa9bVDCMnNisjhDCAmuhlBHKi2d+V9dAX1In/WgAq
XHq4ztiag8uCumTzv0kdzb7GOO7Rj988ufVqdcSinVP9z0H5aYxOUHgxHhhSlq0v
EE74vaWau3dCWBht+WPjMUDXt/PR+kfAgiNMUq3FLJgAHhPlxHa6r+BnhS6B3/AD
P0RWSWFlVbRzdTHjlhLAjB54i1toqikbToMzkBNReJ/2z4KPsxxvbzj+DpnoMZe7
YmCmdbwwAwaxY1DLCgPEunqcrEwovAHodDZ6zqotwnTEr8F/FlBdHQIGdpAM4zSp
9K76sarYPPJYXaEFzui20byKSRzQ9btiWJG7M3sMX7XvYQQ+JR1aQ/Ap8g3Znj55
1k2u6E1v/MNzF3kh5BqskXiZ06yEYWKsS2buj8yp5D9F6287DDIn66TCzlxhmW4g
5+smY+Y/IUQAApDU5GM4tm8QTk513af41AM/ma6dD8XXH3O/uKjuvZPdJPa8as0m
paiagRFUT8PvJY5LUyXtPrAviWlsYawdmTfYobaqfmwbkmBFMDXRIpGPFhaDE/I3
a33H26UMWW2sLHFYFRaLqrYbVphFYBMRleKHo2xvk0bjOxUy9yq4wKM2zzZLHMgP
R+qBANTCjmXCzLMTN0gOkeUCcSlgCyBYkYHxz4rT+5XBiCq7pJpUxsm93kO1V+E1
ofKzvOIQecD81MNqKxhjTYpX1mDogsWdMarnpwmUrRCRu8gquedFZP+4SL3pLpvi
PtKno8MaXrP/qVUpK3BuaKfdTweQcH9hL4kklfaSC1VZGzZ/i+oCmwDWOncucKRO
vwoQMSrTGsg9IqExvfi0+Kfl+XCOAovp7m7tALOtcNm68a/JMBkCi9ydBQEtU0Ei
LwUZxG1XsCwVZRRdx5vT4vh9n0rpG4sCnjy68yK5k1ySfuUfacFp2j0EiYYQxyDB
AvPi3VZgcwHVbXliCu4mxU+uLjzjkeb5ItEbfIvzRTqXlsNZ1QoKHFp1HIsxixLW
cOmiDKU2C9APCztrkH+/ub2Ui8Y0X6p6CcJ//DT1fiWo+JvCaEPsCwJ5mgc71xh2
FntU7jBsO9BS4DYBCbNcqxSEzhQLsKrW3yVF2UCm4RA+rEEcm0VFHkuNYlxjctsY
/Js0vkX065a6cPQEj8Ab2rsxv70rL25tDjzXVY8Ixj44fLv37i2Cq0V0mjKheOGN
ZRkSjiHxZqjMbJI8XLNGTAW+DG/lwJmf5xxSg8zIUhjiLPZ7BciBJDRnVd2uK6Uo
Au+gvO0dNH3uJpu+Yjvm6fq8WAAitgn+VYm2G888gwLc2xRYOz1IC2tL09uDc6HA
hThPB4kwcaq2S4K/EWir9/2Fo46QR3ImV6AnixhRYHtqMz86Q75KWrNf9ZPU8VM5
RptTqzOvnPPBYOd3zdc9eMHzP0ohAdA5MIjr3mbF2biKf+mIYn+SovcGGV0f0eqM
/VwemeUr7krnTRj5x5mb/TanH+hobqssuyKJJv6uXRXGqHnaPs4/YIYHleWUZpoS
cTxAlXZGyrAjSj9G1CgRFBNa8nCgP388bVJLMiSzVqbJ9lFAeSsU9htZTzkXPFM6
9fubW84QiDGqDkX5pPF6uwRMcHNkUHmmx+h1iFJK1H/7HDfdq8skFmpY9ry98yrw
58KxaXbyQAQx94eM34U07xBKH+DUrmQ6ihbF5E1VzVKvktn/6G7SifTs5HtYrS4z
vXxbiqqwJVyvRJxCUvFyEqR9X8yHXiC1WilJ2lJIpLAHo2G7/ns+8G3NhMjx0Dow
SWUDXrwYXSI9IHaZLjFodD3gSKpIMs0zywnoAsTq8N3fJuFrN+M6X9HhjwS0cWTb
kN/07A2WrbYFSOdBdxlHR2I8/2VlwXGmC0OxdAPbOxZLbjSPDjlLyPwCMQhnlC64
Gax1rrF8jUfCK6uC3j8TcrijeRZWxE5jfWf9Aaf8TLM7/CZpUbvNPcEjxi7H3UQ1
47oLUjIx2FuRx8rOkKNMX1m39syd95YWfczACJt3SBaqB/+2RY0RECvycb2ke6Gb
+NrEC/yULyL3hVfGnOqFSH/Xskag9NCRWBFKQszwUUKeKrliuX3Byv0yFA7YQzIJ
tjFrspkxkpd7L0qoj4sf9VFt4bc3gV2JdoowZmXXJDyJp+zWyETWBtcuU8rcMI2O
PuSBFo0Vis2Vy+H48pWKfFZI1gOmOR6XxsN9yzIi/XNWMb/lcIMCYRTgmpa1tZzb
ujxiMHLuihBcO2EYki12ZIwZaMXDW0+eK6nabzcXV7w5T/wWjBiyWnCMnW7LGMea
DlK+tTA7E2OJVCs7TdlsWVKFls8eaJFC5Ka38auQoUBE3oY3cCx3mrFq5dJMS5Dx
TMfkQChIdA4ZUnHnqNHfEgvn+syIzaAT3sSBiOOaAhzY694WcpRupKjuYJgo/Fjg
DOmRebi9SnrhIyf1uvPhg7bZ3zEeRSuygddttdmmMrJJh+JubV/fbfuqt+BQf+9U
1UWjWX6xPh1x/4dshiwD0+L+ShG8/kNwjp4gkTo25jBZ3/XddN8vD/+RyQtkcLYR
Xn5FXZ0iB5kbpBoWgC/2TFwxhGHpjvxji5BgC+vUh46nZWylQuOLWxAWaZkNtm4G
me5zBmfYK7ik1hq/zs66OUwkzp0+D+FYaY2Oco0dsXKPqLf3TeciyJGtfgzCKiHZ
COOmOnRudA2mMc55l8lPN47rhuUf1bfIz5AoCuheQtxirMzIvKMPg6rRKqvcBtON
Go1pfB27H/tiDv8TSh5QiisNJcijf+fYK7TekRjeiC0guvqjXeGAa67P8pzptS0T
nie9xvmT+/Tq4wPaeXLFyBA9sa7FrQpgoZruThH6oqb9gS36rJY1GfReDIPX17qq
ZM7ApME28/7+D/UYzjXtGwLAS2N0NtuzDd7VWCDkEUN2Lkwr57i8KQj5zqQQ0w24
9L2rJbaUXYwk3vK6+50MCrEsm03I4Defb7tyTdpbZWaAZ/BN7OydjnYAUaANb2s1
dbIvCGFCgBk0OrAD2wDh4NazfcxMAL9C9o8wJlG1pGMMeBrVLOqBKhUIAMg6Zufe
320JDYSMidMy4VtU8b2LdYXKa2CKAN+/2HUyX149kolmAASS5VM8Px5mVTkcw88c
mAuHOCHw+ry+RnerJdSuU11qESnDnbBp7AbNiaziQKUTIltooNddWwvOs8NRbQHO
Crs6r/PJ8gqkdg9TW9ShfkCc6caBC6Oijxtc8A0A8eWlWWNwd4jsKnF7Qb9y6fdC
tqrYl8kkJvjVvbkm0+95TaYyH0ZGZcY61ADv7XJ7QRyd5JPy7NEZ82aFou2njTtT
cxkNcIJqNq0tyWe1jhqPACkRzO5Ol78pNUi7RvwFerULWUpKdeOEbiZIaBifx9MC
Wf8FN/MlQVn4Pjh1WoeYodkIiW0LaoL1N4PW6jYiL/KilMbgkzPyj+gNWY4pdBbJ
HmFIY0mbnudoO9LrOeaUjSWdH4cFklcXmdXgmqKe0psnL08g+rv6LXEjK9QE2Vdm
YMSXFqROCTbttdlllBY+F9yjmkoaYiqXdQIyKAijVvym2UKMargHA+Dszxa7nP9z
8uLd3yyoHkaw60AqBoo4ElzsrtJIVPHfmaQLUtm2pAT+OShtBgwXUY52FgabJdS1
qbxh6528ta1XhPTTo1j/kTvf98p1YSJwlpjccXxXULg4niI6oQ/fvvvhnDe6HiQv
jVVz+/VB4JmegD+CAq5q1MNQBmynIS8DnC3LHkBXyAGnQo0vvVf2KtvXjIrIhmbc
xsJXO+io8phKIqOesv0LpWiZMzS9bO+nTgOTtbtvcJJFb9Hc3KPszqKIL5W1/SNi
kjKTgase9YS9wPVVrTTr22R1vK0RGwMFsnaBz2VhHo/5SHwa5hHEd8J4dwFSLW5s
MsR9f/WGuJajaW/9e3KVqejhkWd+R69dsTQqqNpxDLMJbRJpcHyf/g86GNrwau60
sr+Px5N6ntnvjTom6/9yKlGXjMdph9oDrqDJOCp/fQrvH43NzITd8ievQD214kQh
9WChOGnJNK/uxEitxQfqm09LpJ2Y9cQlxskNPuRSeY2JFnYqfY0R4ymd1KcloI3h
7wkFXrE7l1tC0p8tNeM8Hp+CORy0EgLefCC06/W0RZOTeXI3HA8bQQ5+ta//thFp
1p4dBJoz+pWTAC3XppUiApyN35qCDWEgFoytfJrk4JRJMGWr0lQCMrgRWCeFFwsM
QCMO2zksLTElSHKKagY8Pno5yuIxJjzSeHAUbJZ31NBXa+Kt3J6oLK2pS3hpJ728
U1UWLQ9C4T7dJiWM2ZBqxv6Hp0KG8Uwv6LIhF9/zSL6DGTkOEppB3nw+qSvo+cHQ
hHWZboKwViwzhGWJIc4XhucqPaRN8PqKRSZzBR4ncC/kC97qF0E6BHSla56sKxf5
hh8GgWYXAJExLMa01tmsTmvl79jKM0YXfTv4+XWemqftxYaxq2/75Im4sGcsgg29
KiSYnbdmmyHytABZr1qPdezYRvIq+optV3nofDLv2s9igN+Piiz2cvQBlJbHHUpj
xJhGUhPtdNzB57jX5HPlynXBwwVqLyCbPeTi66mduzs0EP8OcejXI3nAEWlgBoQC
yGZGo3aq144+/LV2rLpUyT5hdjhE8Fjc56DmmcwAZKNB52ZrBpFyz3nzRCaIbPwp
aX6LMF9VxG18V4sf50fl1rpltttAki4o3JdGdxe670202W7qfQLXIz4/Pvbtdx/Y
ZHuvKfokjVGRAjDK1GFIDCi0HDmnq+I+1Z5fydKbbgqbSVBHRo62o9vfrZv6t2xH
HUmo+gCPfXC5Eyy4rsO2ZCNvDrHtzggUdQ+IZ67ZnlVtNvIaNSMDV8CS9s+WoOXZ
UjuRroP+Mjm8nqqjDznhpU6NSJzZ4f2Y0nk2CebVkGupzxFObZQhCpVaNKiIq0/k
7xkDpFuiPH/IcDhxkJLiP0yA8wVmF8nRK86631tRVxlrygYfbnB7n6TuyFL+P/xt
Uc32l1jr/T/2yDlL0NSo/BRSLMJTmOoq9egIi7IMHmjiX76tP8xLmWmvoThqv4Dv
popfhAai9gwD+ozD7XowLw/S/rUvVwUXeQrOhkiFZxc/opNbAuAtyGKGjq9pxOBo
CB0yioeFmwEG2A8Hxz3f44RHPRSiFXIl1wxlOyubx3PpgX9nrb+fdJirs5Lyv8kS
fOdFLJ5N7d+X8WCEGwxGPM0y1MKo7lueiWIwZCUp6KM4Z2OXNYkyf3qVxqV3amWr
ysPlrLT9qHmr51aovQfxHodK0hpwqVc88HwnMRJnO1pDVDmSlpno2g3TeaWUGmzQ
iCp2y+U+IobORCRvpodO2FokfgKAUuYV/iLQJWK3l0Etmt8iSZVUs0nI1CSAReuv
f+UeNGXYZlIAtCC3msxaFzvcK432FWIs54ZSoiX3rUSwdBXElsxXUGyJLQRW7IzS
EUAvoOxYCLw00us7OqfFq0l1uoXzEB0NvESLl9ZZYRPrFFP7m4A4HzVfH867szwP
HID364RQ6ryt/rPsLFsECPTIjQsTvUqh6yx63qH3TE0Ep09Pj1ECc75l9Q6+O4eM
VfvG+zeULZtppKgiA2DYv4fqngc4Gb57QRCySuahrudqZqxIBeBA1oArz9IE3Zi5
wai5rMdasvFd3NYQEe2ufqnQz94wFBV9ILtf79iAm2yVOpraevMm4d1UkQ8YJNSW
nO7ct3ZXARvafjcnW1LFFc0Rqpqi3KKV9RpVPlrMQ8E4jpGQNY3HEsWUP4fTWvSG
URRYa/NjUEAqaCzL6vu534+F7dnacOnF+VxQcO3nZNV0r7LWLzbj7eRvzGcVM0bR
tYdH4TTyjw1MDey5WZaSy82NOE97epzdR+hbaijTqEahxuvXqSbtoQXPEthuZJBW
P0T+zIZ+WG9IV1IHlhhqDrks7oTeYiZh3YQRgBoOh7iH076f9W2FSgKmqs5ON6Sm
p8cVp/LlWd9AH2jR+zPlraTz7YNuBKONLdFH1KpMkl5tyrjOAF5WfctehgSTTllt
0+nMed0yz9/zTpnVsUP58WxouE0sFJ0218rCbeCnylJFfn6cpE4sy8joUBM51WLE
lxiwxt31J528iA4V/4DT6WkYTekryLyb4VXwBJ7JmTlyRmB3hVoJWlhZghVt+DHN
K7d24s6WfcO8krO9ZipteOUuMl0KvTIdxsbkhV2t0gSAFqdcDTcNNWoPEfhEuQ9z
L/57wjGrbtWECUEUD2DzZFSoD/aulqMgAiClfRwdwPBa7AhCT5AKIQP8BN2IVvhh
osCivfNFbXUzPPntXiB6smIXjqa3uQy4waDX0WnR7coI1U2QmBfvlBx0lCDeFfPV
87plUjZkzFwLD76ls40/zbL2l+r6oBjz1ywY3KFdj5S9pExKKZQS8v+7wBLY/bQi
JT/ElV5nw44U2E5r1vVVho4xptTwUZ/7g6f1WWoUHGXwbcH5MFr1etz2oa9hSmr6
EEumZFV9xeutt6r/hUCmGuZzN4hmmEoLCbWx/JQpiWbHldhhnpKWlD1OWyAMQaZL
TXx1YA7pOwTJOBzW5b43iEXnzkd7rOnRtvyqvgTSVH93o4nVotqbSxAs9HWmoMB6
GJs1bFtF96ssLktm8nUFDGCC/noDl+qYSNZPAwftmi/lodPoAyUHKIs9+65KBgc2
d3xTGoj1M4aYAfKgU1E89PjHJyJ5CfXEsxUM9hsHJmGxXBkPyOBK+Ik5aa7Jo6/z
hLLekK97BLcJ1TBRr9VQ5fxpmmjpFCqYQXSFemYBbjYs40lU9p7QzT9fdM4diGBo
s/bO1vmA/eWI50ZbUruca3gaL/hnXHuSEGiu/LXgkVIbXGwsJ4TkDNbxbf/5a+6K
f3NAaUCeLrHkvsvDtVKxjcZ3a51IP40Ma/7+Yw7G7bvJs4phN4v7qeaiDY+pXt/L
whF1IGB+FeTF7f+CA9vXsFijBCOsXIxYvIA9dyO58+nikPZEffxSrQuE1RIkSF72
XwFLBNsb5fEQ58Rs/0EQ3t7azP47qA4/a+Rhhs6mRDeBPGu+vmN7ph4AjhA+JLcf
PjR9C7Dt2GrmT+fl4xwm4k2AsCfyL+smcCsIQuFyc4IXjEiado4qk/SCugIsNi+R
HA4bP9JVYrjrPV9iTZRzrYBZ+21zh81Q09cYEP2pVK0ZtIu1c/aRQmVFzHnyuceP
P9hEhRpULMXnZo8PjAK7iEPwCloKAwIwDy+gVl7UJmFjTR42FJo9A7T3BXZlMnA2
+ZAqbTapDXXLnUaPd7udK+h9xKumBvRr6ubiEE7WgnOecd5moB8z/+xAOEQlL05l
8Y75znObFeWsiZD6DB8ZeGKIoTaLEJLvKagqOP70qioEK8lztAGNTA9sOnkiuh79
gk48tQnGnmxyfuZuMhWjysHVzIRxSjAdY+/N6p8c7TDMNXjNNDaUy6+/8ONsP8Ls
oU7RoKsdNRKynOtIaITeXo9J6d0tFa5tSykCREVoxxfuYbuOljNTKrhAnnH4yS/S
IPd1x/9rvjfaKa2wcAKQzMEEtwpormrV626B1WlVM/cBRtty5MtLG4bZc5rhUYaM
G83tpVM/+OJLS5TATScNkX3bHw4iV0Mx75rq8a5iFKMXnktYlpBUX54dgQG6/Bwu
8/JoP75OefNAfg+HFtNwMCNXwpjgae36gay+nVKowiQ/LypT7vtETv6zvODjNW69
DbSp1ssAFallnXflL4+EnyYmWrRep3ZDDAh3oVQ1w9FId5yx+To2zZciO/u2O6CV
WAzw9Al+hg6q0OGdS2YambJxER4hYRCOpCicaFR8r5qUY7tZ4E9HWM9CG+pcPlMA
FO5f2KbMupYJ9C9PyNx9ZUAxHLfTrOvB2PzRrWB5NTibGuKlXpAcx4y4GKH5TWar
CmDsMhL7gKMkqQKIj1sH0o9+ri52oiMvLbiNrffSLaH+jx5fAsleALZWvBr6y4RP
5n6YSYD8yYwPmVgRd0uLHH5SYMW8OEAzX94W2HpRbBv/RMLgslkjduwL1Zo588u1
AqRjK0SuH6tpABb37b8M8YAkdFkkcO/bne9jPz4Nr/JMnsKHfZqXlwrDCNQ/XzSL
mpfmMGT9H/moS0IhMGaRk5Lyq8zj1uqWs3O+WgkhFK1Atrp0MiPaS3JYWY2gC2BY
+/aLp0LVC+hpbq5G4JGiktCD0V7410GuSWDopTCAd/vp/XpLfy69J4vpbcquG5xR
lKc3FVeOBIj1vqIvFpHXiOUrUl2Q59HqO2rNgFG/FZO5ULxJIFusWuwINaN1hD1N
BLAHpvyLvtcmIpO8ayGm3USkOLNTUNmJuv7JrhSHOUsuBFns8W7Eh9WL1apWKCug
HL5equ1fxMWovlRgiN59XKa1JaFxwokpzdm6rJtXHtT83uveQPIT8RxPP/Ot2aA/
jEQEiBlRf+lw0HxKKhAPf5jLh8drhOCPah4hAXB43NQzK2O15xaNscFFGnYE/CMt
latT8+Ft/LG5Dn5Tt8iJtsmwVe39VPNpvTu1/kFP7ShGls95aaBqhK1w5tYoSyV0
0MSNByWjUl9+G4Ay25REfgtVIHaj1Hk8CQx23cNAEhvA1hpL5a4XYwd+OZFp3FST
x34AwBAtad8BpBXku8IsJQ675Rirfhata47GBageLj7+iBMMfrCoJAgdygJrIYO/
caBS8yXNHXaY5KMPoceOP/OtWCwi609fMFsb4+wKHZ1LIKG8KFlp+Of8dPB1Ykgv
M4je42fCLssJjt7hZoNW82GdT0Usx4xOKMu2w2iE6dmeWhghILadD1WHfNU7RwvM
aNYyHKFyU2nm+R8MQgvcEkA5NfOZJoFlW2Cz3cFR0Xn2TwW38adN6cXyoa0cuBIS
Pp9WvsafhnvjR7KVfa6u+E/JoCtsgXw1m5NYePS6xOQtx725pQlwgdCBV+xcNY7n
PYjH7ej6L//IxiSusG1i2shPlfWRgD0qePKJ9RCf8HIAZMU6T4R6YOYDCzhr671d
x1xONwb0P2iK1aOijQwrzYyASJikmo2I6mjpljoGfWpjKIUMxtGmDxs2KvcTdN79
R+CoR9MUs9Q2Y6uP8upTVjkdc+J3Muy8Iv5hZyJK+QaRLbNnxgsy9KmtxbAjG13R
pOOxOLFn5RzdWv1/DV3c8+EGYRuns5anPLS5N1RPo9v4xlvEapg5pEGhyEum6ELj
EkZGnB86ph667R0iOVt/4KjSe7RNzjpr/B5JjuKaLvc1whsyWJpi1QrGYKR2h93Z
UDKoVukXgK9OL0sz7YywQE6i3ZNlyeGOunPwTAiHlEl9TzvEs4gVCy4yI8U++m0M
epoHKj7u4dcJiE025evXgcrB+WYgKOMb3J0rm/6GMJbPeysMv2NSsZsv0i8vMi/x
mY/xR1n7WqsMogeKtQuD5Y1cv71zpyYU3z1680XVGh6HY4Xea/SMN/AQCHVffTvD
MfuDRKqDp0a52+DVfSDbqBKR4w4whoKKhUQKQT0tyXVMQIgGk4p25PiqByfwVxt1
4FuploobjuzA7zJdS6BV0bq79GvwUNiCY97qL6Ql0DTNL9STwfIWDx2ZbFniAcOe
/Emb81uZR5utgP0cdE3Y2aqWUV2Immgx6e6lX4+VAoaeJAwOC4cP8A3lrBK2XybJ
lwIA4EXKYzdIZW+pTM1PxkFLN6hNq25qqdzBtXMoQlkQtTe8xX9UZ7tvLI5pRuwJ
EdUJExLZfNBOMfDN8YWaCvrdD0+KXv/kwQEZRWdnf6UG69s4GpWbMIlDI+WILsjr
Six/IrD08SNBAc4/nTeFYY1gzVkspT0R5CqU6HlRcC0tSUkCCozpswWF+D9pUqUo
PQrEYN11s7Y0xY84HYbwiO1u6cIysYfySMcQ8GkrTBYGiIDvu0jxi0Z4GQ70eajv
wDQVc9U3+yu+irK7scit5b3hlqO60FOQQijexFxXup90/0LcfvNPjuqmTdiGysBH
XDilEMfsn2t0Sbea+qg0EA808QX3Ep59pCLzZkX2em1pXQZdtWnt7RL3G8UbwK+g
c6qRCq2Jzf5tuDFctwqChnK1VeGucMjWHZerVZ/Ygrk4ae+RGm7dBhh50rWrZ0iD
qoj9fpq0Obug80urB3jO+lf9139az4EyrL2IweOnLCGEHIJsyrECZOmLHRmrVVMC
CJkyRkzoaUj48HPjDeIeOedmuMNFX0g4T4hrN1hT/8GWZ+VK4zO9vNe/v18fq5Wj
go9U7DwNoWbQ7ynBSM4o9SefZugXO5SnljOaOT2S89n3At7DXsZTkWQRfF+wceqn
4ZKFbXAZZhznswuNAiL6XxETuMcVgc3yvDJQvEEMivi6uwcGp5pDPmMfFv0UlmW8
U93Pr2idZC+3519hUT7GXDWTcv03PqVUd6LPFgDFHKjzkSIvu/0PUI/IXGNW5cTo
KSbQJqchaGK1xv0oGZzTPpL8qvme7kOzY2cMLgGq75Z6KnM9JrqdzwHoeTYkeDCp
VDWM8AY3AopuueE1EsyHuvOt7Rr/R6eAI0J11uv9VuD0rL0WbhWTC2uKgJ0cf7F3
lAUGWVDch2KLrs3TPA8V9lEha6q59tfBB4GvhE3lF7RI4505Z/9l8wpz8Tw1HTUO
gJGz9HpIln5VhFKQfvr3rj6tZVLRmMyBBCFiC7SyQbOIm2U86zXmbv/wOWYlmCkd
HarlzPoPLI98rg2xkwIlBBDNm2M763D6hrGbGAaZbdr18tbqYalFGz+nj71p1nbX
/RkCocTWnw3xF7AC3yvQqXZewXG0XPQDZjOFpT/ihlSlSfsj20/R2zHJP/3fZOdT
jxpSVqLVWu0TWI3cAtAJ0YM5GfuTlrPkTG8AB71WzOYkf1y2h6XFj1zfx5imCgg5
YXdkNsumuPq31WGOF1/2tHJ4Si5M1ex0P4FIhnpaTN/YZv/Am4Kjpg6ngh3hfkR9
aqGzS2/eCFy0bLyItJv6V+p000EuGak48U2IBARZv3ovClx4seggacKtBMS9RmJq
7cL7Nse0IyVq1009uyYQlI9OTDid+RjymkpCVpMFtRLRCIMr4Ij1tv65t3yVHhSW
ijUwnvW3smjjPqZ1xlE/PzoRwFzdrRgLml55SUrX1tvpALBuoef4E1m9TVbTdcjj
Q5n8IfHGDcFXCpmatI/5VYLWMi08OQDAOVpX7s+jEnpktVwpdlUuyQojWumXktpO
k8GA2UO2cGYinUecihdT8hmG9e7VV1dAqa0PqqifuTaHanTkYyDWu/wE32uIPF98
AxPmaDo3sUvDO8KeJ6Q9IF0/w7jP3pYhXYWM6zttsy8stFnAsywRrf5nPu7jEemY
xEgmpKL+JgB/GF8MAWdQTWjrrbs95GrC3eR/ycWLd7BcNyxDgSmXq9YlN6amRrZQ
/rtnIuT4KoFmizOZ+j5u6sJPuRkPUsJR7pnx38MojfIDFMGpz3DQOfNLFdue8f+N
8FyUM7MgnBnffl8TrJ2gVpoaYx5jnoPN4cfg/SdZ7LoofhrLvmP0HbrveDcZL8BT
Ph3IUX+au9N9c7yPt0uCFBsFgG8WEFtoq7GHw2ynDeZ2rljqOHjxDTS5NG/GuYVX
a2jFS0Dkfl3zo9Z5Q+TYaGgmLf9/79gN6RPmO9iWF+MzkDAFaRajre3DQO7yCzFY
0Jd6vMGGNoodfMGFWU7dSdlInvbu7F0APMkeKObkC2ngp9TXUfbR/UOGACJ+HyQf
5X7c8kr6wJpTfqIaXKcbpqlIN7xs2PD5otZsmv5awc19kF9YLfhHHfa6NHrA1QfS
BGBrFQeR2kbtuTIxH5rVGF0bpzJPQuEyG1Ialcn581kOm+gUuUXBzdD6nzxfIMux
ClbXy0cI/RnSFktb65tx+xLhlqKqqjKDafbLfFI7+I+z15z1QRCd+woHlUJfS2F6
zPz6gPuy5goa046dNghgEifTy4U/+UvJZm38HBfvUtFeKhXJFuf47hxrEo1FHSBb
cUe7Cwtpx5gszm87h7FRWctU6bi1cANBwYnFPrKrrYDwaIzS34oix0MMzMOuORET
j0y6dlRuGEoTPsLhok08umHbNCQlnJ/lo7gQX0n2raZhfrLGEKNBnd4bVOaJMP90
Kqaenhuvu03/25g42nqBAfy6swsV6Ctu3aozEQNiOO9hFCNYS1UE4IxhUOsb97D7
vYKnCfwbeZ+6+YpvAbhs/ddckxFMIzsOs+lEy2pLQgzIIGuEwJgW8E5AKmOIB+5G
4NpjcUIj2ns4FX1HPp91Ef36pTVdQTAO2V94hjg29halwLE4Zuy7UW+/Epyfhi08
`protect end_protected