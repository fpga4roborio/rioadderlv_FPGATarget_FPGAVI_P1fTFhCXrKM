`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
ddtXksX2+yylW5zu6QL2Lhnb2d1sD00763mmSITNX595NcHTEkwn0zB1Dry37fOW
FufOhVzEJp80NC5qZ/+F0Vk7Ik02dIR0elf3clrjeJRK85K4e3Hoo4xn7YbFUIms
l/8VZSb14+JVGURjfswrIyCUotIzlzVYZ6gzoZwDXIi5gQIBf/gI+KxNXPaKV+PQ
Ufys/12rjO6aI/pPlqSm0hCvftmBcnezN2hk1UeXgOIuKZnogjOsf0iJVX2aOOWE
6pD/psybjbnsNB6kH5uFTA5frkzIzkzl5d9+YDm9OyC+k84E83I/7/j+rk4L2dah
QJOvksSIzN867/4Qt8qYTQ==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="MvBXkzurAa5VTw+1JJ70nePUfoQXBvZOku/SMmg4TwQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
oRtzZL4VJ4iwysPsC8SXYCzXS8Fw2gtZTOskLcDV+1B9Nzn1zTyNtlo6lNICRmmK
ZRVu2BmCc2G+fmzynYlNTnSa7C0Cuel6FYpxCBlOuk3OF2tzAmLAuDyOH3Z1Yjzk
a0aHuoCdIRKv7BrZCdALt03JeUmXKPdOmIlkVGFl8yw=
`protect rights_digest_method = "sha256"
`protect end_toolblock="Jn9CQpRhJt4rnzZPRk+dOpzAubz7omckX1MrFd4p81o="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 10912 )
`protect data_block
gD6l00tciPUa6pDNTk/+t0OO0nC/UTtBwLB41d4inuAUA3i/ALrNyoJVcBnAmEQW
ptbcNp5fxEUJjnOxnedyZEuEBxWRieZFQnkRdF269oO/csqYH7by8wcZuptbJ7SW
k/HFn9///u7NtRnno8uEFQBrJ6cA2kYcktw79RZv+syq5MFBIhgO7bpf7mKBCnYs
gOq1BVi2050LYT/9moH6EvrnxT4rMw5Yuhi42/n2kLEKo+mMYx0eeWCZfr4x/msJ
WFqdoyQeH8FPBssIx9+W2eP13wG62uja0ZwdgxeuhTw3T1PgwHSPcBqANEWVj8jb
alGVhYk/qHYdqKKwkBW9BenBgmTau/GTMj72Nr9RtiZ7VlNcIa55j3sMIYeRheCo
ypAfo7z4vmTW4jFzl7B+lWtgPZJ1gOsTbHrDXnDr2PgNYVVBWQr8dt6l9kXXAhKA
N03WDS5JKJ+Dki9nkKMlKIMLc5ip4BQivKKta+JlecDG2A7d0Jn+O6ldacVgDdRv
AUjBZcuY3RUf0iSALcYHnrWsn7QogiNPZGVywraWmSa4pEFh7QRyGKeHu6Bx52z1
p9KVhVMPsn4CaWHhXuD6z7p0qNUd9aR0BYfl7WGBwm4wE6/PKDWANtJD490MRN9a
ARF0wVvbp7b1EOgnabhbj0tImOxFo4HhSR9KfCjQf9HVsR4IQTJmAwc14IK7dzzk
wSsMSGZ2Ibdw4DvnZ3nXPSOsWD4SMwNB7E9UohQQ1fN/V9Yx0xoBFHtXveKSsrWA
uBKmYLbjX0lRjVjLeRDMrOLU5LcmFhJtMmicgpDhTMcqRZwEb0afBT6ZsCZgU2sL
esM4YMhFzUM0IICYRl7baFAxYXvpnvUaqx7W08vStUHZteLwew+uBDr3XzMir//k
xd5mgamrmqyk5FnohjoEUe7MKX0EvJLgwgJ/iJ0GlVUnGnyvGK8bBlYTbs8/giOH
V1J5Ye4mDW4cPmSJbkcLb1/20g/SGMUOmHJWK+9+rHaTytKga1X8cU0cSqVxyf9Y
GUQ8ZlTItPO6VAvpNM+DSgXLtHPNs1/xD334qLQ8o/083d1BFWfGHCrJqz79jeaK
iOjjw1VWgAMKjXEZXAOuf9rRR0txRg22oMjXlpoClXrWOeF2L0ZxJOhUGx0h7sh+
HZlrI4+7ruoyVDzmp3vhkWKCjnQQkADvQwv7JX7+hf6LroS3Q8Ev3PizGjE/2LxX
P/AKvfasK2G7PMKiG/O+/S6dh2YG+5gj2t1hgAAexhKLIrxHW78tf8cPOIVewwbb
gRVdOURujgP8SdNVZptFw/EW31d6F1lOIS0S1VRJyHd1iOw8jl4UqsbGCtI5KOhT
KQBbwBshDscdZG8uYGWKywFLqMZwqUAYHOn+GDygh7KovZGbJzQwEpG1rYGH9HL8
937pjfnpiMsbZlomf8AE0Uwxl+BKMgYyAKY/DN97uk+QI/LSVY1MuCHCQ+b8n4Da
FFMTxT3dBqXOCAyfR6H+FcwivP/Ejyb9kEEeWddhoPd6dSgSucgNuIo5p+iUfhQu
b/qeO0vwaIK2B0n/EhKDb9NgItrY8Kzff5R6mKhBiNQOXphsRj/63ZsdWs4Mc4Ju
gblkhuSqcy8hd246qdxox+LTWE31HZPMzJx7n5nrgtlfZCsl1y8h9OnMAI2LjsPW
vjNU4NQ7snmCc+1j9kWz4g59osl2fyPFYxeic6sSyoT8MiNprYYj0AAYtqpKuzKb
3MmNlW0FxeZY5zBz7Qs7uL2vrmZyIOuMw3PmeAUpignAEPBC+z2Op2J4O7rR/pkb
qLQhfs+hzPvi1uRwnyAdtFI1HDoMqYTu4v3uD/tWyyoSZ/RUj94o/2od2EWK3tU1
lYJ6w8i64WZz4pTdP3T3sBHvpjbWnJymaydXYguijFVDwXNWmya21W+eU2yzkSTz
tUtxCUAXKv5/Zn/b087qvBXCU4hoxUEokeRdBsIZ0vlwAJHkwkLTzu4/Va7hB2uA
/RUTBjpjce7ClB1S6aIPZGU1L4jUsH+4g3MrG7+tkDhsBE17SLJl0iHM/cbD/m0Q
ALCem+MiGFb8vX5sjf7K8RCOWgDc96K1GPqZh4y1JxhkwPtVsXTqLBLINakRjq34
GQPhKQoYlPs5bYHMJO1WXJ+1a14TXf1HNw7nEdENWDBSH8rHPmAjpeozXhFGi8XX
LUI27oikU5fL90mv4wczjIVRzc2rEQoVovXogyulsFL2UIqA6xTVoa+FIKZJwTfa
FRXTjJ/+NVArn7b9eR8g5LPsuVGTpXqaWFKHxm885Om7S8VCuIJ3AVrtaP7NB3ll
Ud3Hr2nrAreyCtM8HOWyafBclAF87FKdokyQs5I18qlLsTZtN9en55mJ4DcOLzeD
tb/TTkwL5gA63XDj3xapC6GWOeIIc6T+k70cvKRrgEhbi3ptf7npmX5lBo3aWKSN
SP4FWl4GFR6tkdzGIeYjY6aKuYJH3XlhO7iKM4WHIcVK4HbR/8NVWlSsBT553E7g
8CnTP2YMcI5qK4G8BIWpoOyDo9vEg0nKJ9sidwUxtgxpSsosHU7yCBDShvu5XUxO
QP64ZWaAV8nxy2a21VfImrIMQnMXAQGLfTRQVDKIMnSXSe6bEk1KbM+8sBkQ8u6Q
qU4fPODhSOQGODa+vA8SlReeaoSgER5TmLg18AvG9ZnvGHpztG41csILWN0XifhS
F4EPIrlY7IY3PpcfJ32HtWL7xvKbO6Uem/uA2VZICIBcyUYvMUZzpphVJdukfcc6
jKB9w8PJIDbJVDaCpWepymRGwjR1zITVr5NTicRDPIZGttlCWlT7k6l2p+EEJj1W
2BbdXNpimnsmCRZm+zOZJJpCWXyALrYFjtCYmWotV1YrbOsxeyFA9AQKRS+FX0Kg
W8HAH66wY1OaSIT9GjioAczFL+yXWBDmoCI2ZqkdMe+2lkhwG6HiMjBXubluw3iY
iA2QkLFOuE9jkt7eqQNlikEeZGjaUz8YbTiXLUtYALrCMgCNcbf8Db0QpPcZN90F
tdcY75BD8vjeiTNRHZ2Xv0p0SPmR91moa0LaEBgK+N+5kNhlvEi4XYeZSZxxOWza
tN0S9ni3MlqbcVnneqWzJUqeNR8RQwROlnOlAlb3svEUiZVwc0+mwZGxCc5x8hLa
rfhRFpGIX0IP7e3f4RCnfK7AbdVgXlB233xLbEbCOPDBO0yWL+Tb0UzwwzmO3v6k
/UVV3IzBCyCsCIU3+QfaUFFtEtnpNHmGXaGegqhVzSwXAa+1Pf4nTKjjrkEllGSI
laAMNQc3uXRvSLXgb+Xg8MzBl2j3BHiFW11sCOQA+QW9Ep9x6dF2CPzaRjvTGU9h
ea00Y2LhgRYI2jL5hVhUJi9s+ffKh8SoI3GsHhtzhibZtmR8IeDXi2tbjq2pEgbE
oylCgjcVq7iv/wDSU00fBufg2ynMJ5MoeTa1C6/83ZM3zLEbcaJYyDhThT5Ni5CZ
ZC0muiiBBbIVVszYohhgmQpJhoEicA5yng5DooAcdF5r9gSXiq9yvx9w/ij3HK62
5H1WK746TOklWVWC6C4mahZwWuoyqLciZ/Uu/khHxqrZYMGii04RnQJNimLhZLs4
lOf+YT3U5LJA79SL0hIlE18VhyaEt95C1lv9ufo5PJJbHb5tXdbEaIlrh4XBdS9P
B6y8O6YvsSQoqdPsXHMRBxnpJoPXcZCPlLGonsLimganHfP1CrId4etpK/YcOVC3
rEWPttKYm+NUt+I/cFPJw2W6IseK/dO1Zg0OL+0l7HBjZrolA0cBiyabTRU7DrWc
sBqt+5SQ3djsn2ITbnLkXPxrrbVvRhmH9nJBveVtyZXk3y2aAIZv3mreS8qaaeXV
FSjSBjFVjzvwBAYALdZrXS0Up+JYMkPwtgRaYgH7ZQJx4CohqbeS4FfRACgSCMS8
MmYXzrNqpCjEuespoHejK2QLWKVFS6yD4JnMSB5ZhojybO0m3m+1/VDfe0eFmpnE
lclSjBME4TYXvr0CsasRwFIG2epVGa3P1JVtNfEw9vUwz/nYrscFrrVeEwsrEUR/
Hykg/VzKIT5x2KxpLeIHLXnCXL6tTvWIV99GBNPpnYDHRVHbuVUqxYOc/vqAZ/eH
14NqGtogIIEKqdgt0B66Bl3yNCdRZgdGUrOwGT50ivwybOCBTyleqzoF94uJb4Un
DuTnyesZ4dDxC81KWkmwQ1q+KK5g7QrbmiilY9VK0clFVC0MLcmGFYG0OpGoCDSZ
ZN+43DQpG7GVsEucBUWE05hqBXO3AhLgYywQ7RA0gq7qayqKz7jYroeJLqEZaBZT
iyNW3Tzz1+wkO2Rg4yGu2h9T4cNaSQO+aHrRxSqZAq9mNCGbd4+nQONZ0BlpmWkq
0RfiaEWmL+rDcc2BzIi+37t/aA6VTEXiwUOzfANTgAV++2+/vTjdurQ+eGQHFY6q
dYWL7o1bWRsoI8KRFPS3RLEUzeiK1d0DUP5FT3qZ0ZsNgKnoV2NvXn1BQKUrG0gm
CWOUH7qB3uQuujsHl1caPjKPeZJvMm9/+jTbQ0p9NO5k+vav37H+mXXam2/NpuZ7
7ThKIcnrCtZZ+CPaM/4E2RG59dWxS5cT84fbDGtdet857Y/yAFh423LPE3ajyHV2
pJiofPMK+23JlSA+4F+5mVuXxy/6TB6BwYIVajYYnz+dmEp59vPhFxR0VJlGAaUO
8ga7WnOttGRiEaAB0CD726y1/h0bsGiw2CJ1G0AX447fguO/bYDOruUEYsNC6E6c
T69RfrtZ5lmepFgDELdtcNRYVmJiGz2+pr5xkoW+6bhr/Gv/nkQfvRwVPAKYMB+D
XEUuhZ//91V1x4LBQbtuER+jg7axrMDBsDgE4RZAwsR0jigTbqFmjBNk/fjtpHte
0RrdJvRCnEkTtDkmIHjrtjKdN6uUZJ9+oE8lZKtRZOqhlTDFS9HdyDS4goYhsAsB
Mxlwwngda9ELqDCOkxEvcEnIuOMqQffCAfJVebE0+R5RsLDBjqUok3XGsm5hgkmV
qiizBQMc1ryWxOZ1YHBimNWayar+DM1/NwG6fZ1JW5eesCkQyaucxN7af9vXLK82
L0eA9gdI5UcddbkBI1lTtDkJQxwZQcVBUY8egS0c01F/IR6s8/7jRzzmeuD0B/es
wetkg+4FqZiAL6gxYwwh+Cw2COUFcTWRYq2ZIECGRzsAwZ4NUFPelEsIK5fqMQFP
30Ip9sd4LengqnQovCEgU03vpCCC0xXMZ7UhFxFXlIh4N0Plam0D4eqMr5EH2SFn
IcdR50YX8998c4FE/DDNXju0C+sffmvP3C/ow6YMso0msocGyQOdh0svd+Jmqx3k
Z1fimUm0I3JWeeL6oQKsHHqf7nOGxUiMbsiJSDAIO9WJ2XzV24ls5pB/nnkuLors
c6sjNWEZnudcS8XyrnSvF0qRuwgm/5T+6VvQnJZq23lVUuLsMM4FofqM4m7T9sx8
WJaqTTkm6et+DIYkzcSnMgzPvfZAHh1MmS8rZekPGnK0nsQ4VuyZwoHyZ/dSlFXz
0X13KrMXYtQz3XPq7qFTcYcKJEHe6tbk2kbEhEfE0wBswHZZ+EKc5oFSZBaFKLOp
YD2znjqol0AEGat27aAsEX0AkBxCuU4uqPWRIWrAOk7BT05KJZcQCL5KSEjdMkxI
pkByYKzyhJsNnF70sszkLjPsHV411lPqyjMx2eIqz0PnHspYGoAWTkCPFfN45MOm
gMvRn+ASE7AlHGfAtj1ihoKVEV8xhnlggeI/nmae8GdbAMiyPP2opDqjFq8xzcQe
VjGQp137Cy8g6aOshsm5hZEN683Zf5S8M+KsVufSDnw0A92rMCoxlivq6ixJmbJh
SOPHUOFMKFnUCTJEHvb28ORsfnbZt8850XHM6ug3g/dLvrntrxl/yQL2VQzxCwyx
g2aWw5n+n9vrsoH7+03E90bTKFUO9sxVMe/GJQYrpAcehCjJ+VAjrw2aCK+7IxkT
XlDfNLw23STxpwGetCEEudEuNPuhy0nl98xR4Tj994B7GRL70rolqclSOCh2HbHo
mX2y8qYNAyXIwEIBxO6WVGe8SZFC0V8m8PTzuPS2p6/bRekqCL0nZeBNORRnzBiQ
f3FapQgkxXzfKDSccangCvDGw8seGwAXXwfeVvdaQ0nogw+7OupaRE3S3ad8nbF7
tH6K7Auv1O9/nZhHU9Nu8VE+URU9b+GxaJjSRBU4mrfffQ5z4eHYhKCeAB/a8XYF
GEPwyWOq48RQdDNt4okdpIVkIuL0pAYrXbnRCKgN6MsXzoqQs/E0o30wcg3lh65S
TcHBxfml81c2iBZAEaVV3/GgUDBblrOZPEdfIQDexZCgMfBOKJNraYIEXrKYzi8y
pf25kK2+F9U11d0a12auDFcjkSPcz9VFhVGitcWaGKFvRn8UkL98d1GSiUJ/ENLJ
cRDyVhTF/XYSPWfIPVcllldBP0d6z4DFWDHPBpHDoMuKxrE428GmgGfKOkfBUyJI
OSlgbUmE5F5kuQu1b05uZxvSfVPcM2dEFuLu8tDiR3UiHD6lXGGyUgzkxrDfZKkd
Z4KhzM6JebnX/F+waCkni7M50YbGXdGvLchS+hk4kDG3m4La+M8k/f7TXqCbyjWi
H9s/uIGsWtCLHcgfQKz0NjJBdLAtdAf0VrWm+43xG5uRj7ZU8KSNKsApyfNV7pDf
qu1wwfaSd6iNPIhp92vqeC4AyfBuX3rDt38X/MAvHb56Z6elmHUR1AANiy+DxK+L
CpLacKNXG/urZOvcVipU+rg5yh3FvhAKcizZOhA+SxmkXZFELkdl6gLPlxXCRqGA
AyBiRIFXGNsHJ9skagxUfLKhD7ZEoPZFV+7j5MKbQOstbkI4gix5ovzsm1yGnrYx
MKxyzBPg06rJp8JqLQWcDOLZQHxuhSce6v0RYcmB52pZjXV7f1OtfNPR3uknkA43
96Kgu7OhBQVvcKif+mQZXDIlOqGg580Lv8cwTm4ZlWUGrFNWeImHsn0adaOP1KIL
O7RHq0nj+6VydGp+N1jIjh4tztQ+U47Alm+fiTxfN3FbCaeqObFKSz5mL2C37QKM
jpIZJSFlVbnh/0zUUgAH4Gh/lfkNv8k+vQMLNOyvbKnAMm0IFYgcVmRXUvLpkqvn
i9cae2jnquhPciZWqFknOHZrnoTFyQUPDkIk2K6P5qYdCcT+LSxRHC3MlV8jhdiq
F2jnAo24KZJGwZ53E9/LSkn2Evh87rIPPsrlBrRIUahjIa7TNaWmx1zB/GGIjnCc
qdc+B0qIMf8LILlWvcrIn99a5X/454UcdcJzhkN4/bTP1iiDV2JGyal0NLPmy2gI
ixeEKBe72V2rec6ITMI48yy024OEzE9Az/0bTsTYXQTX0cD1KEzZ6uNKCc1bKQ/U
Pl9cQoiIMoXveLnhx62cU0qOrzcHDYYWq8jOxjVT1ScDTpD97Xh596qc3RW/pzuo
f+vYQ+HWSaIhtDK/78HcfiSY314K5w2+gQjemxnR/2Cg3SjhtIYnps/jZ45Z195p
m2LESCl61FNHJrBCEr2zoR5xzPV8HD10cezUMoPp42LnHMNHKQC7ZqNTavzot3DC
AXMZAMQjVRarDGiwRiASE8a9tN6unYEFLqjqagjMp8yCDJhKmBoSmX+x5m4GlDfr
mrPB7iNb9VB3wWIx4Ud+IJGn4J+1kuea0pGeHJ8/ZJrxQMuP+sL2YooqrfDUefLs
1xIBKmxlDviWFcH28vzYGkBUJatSifdyrgZmfUnUlm79cvuj0VNLR4T/OfQspIF5
Pd4BNSjslYdpHbX9xJahGWWz1O/nQbz6/02DecoMCJ/1DgR3KMnWDEVES7qgJ2dr
1Ha+xySAgepivkPwmM2wzcM34/4I9kXD9gjqO50rAl0M6zZEiFOzGiDkqp4F+TQd
gaA1ObmaDdkr8+XB78vdtpc7ozXlcy+eybAOF4AOlYe8QI/MirXEJ2+k7STUirJm
Gcr7sO2jFTYvTHoVBexH7DSxTmgnKh+flvyi1KjKZW2CZLD3xaCbBqH4WzN6nJBU
dcCB+Vlmd8K5XMEQzouG4+RjFE/i+sekL8hfmz33zZniWU6xXiNgF+RxY5jbTmQb
Z6GaNuxd59+9O4PnXzHq3K+7kJvkwDpxE8X+uZ46zzRx9Uq6rPYZ/SW2t13qmEra
uT7BuUIiDAKQXMbrzdXpM4xfTRtYTfsI3BvO3W86+lsZx1b6UMrHwgFquF5zeKkD
0yrgcW5nByddcdsFWutvJUUqYFjeZLorFjmJ3Q1A9Dl/mk+5ezkmbwtLuEHC5Ojf
83CmNCGL57xR46ZYuZIRO6olNTtCNolmqogO9peP0q6SUIES0UuQQUbjYdOOUDTn
3yBmr8oihKgTKBFjykrV1oJLE1HMl8XpiMmr2hBIIewN2sx5tnqasVzbmIHH1jt5
XVB3jfP2EniZROxL3shhUj1bYMrUX2hfcKYzrYcILyjyyeLBgRzfsaWzpLjS98ZU
LWDScpDMed+otRlTSmHusHUhsAgr7Q4/ewBCzbEAScwuSs0QsbFmhw/0UOWbE6vh
TTcdlL4bIy0gFyIR32skz4e2O9ocXE/FUVtBX4lMCqA7LsHVaFvo97fin4U6q5/E
ccJ2J68yjV0HYouy0pCFUSsGvmaCuAKPlvwFF7/GML8IA8BQiivJHObZypjeh0lO
+2q1eMf1sDdwfzHPVaD20RcqNHIxC3IOGRGuJWZ69QR4DavxZPznIxgt2+cu5hBG
sr8A5BoV+97XcZg7gK9P5lwJnyXkXPZl8vtTy7t4pO4WOkATV9PXUK1eGyzmOfJD
MgzSsS8iv9WzeSRO7PsWAjq7AkQ17gt6HwByrpz3V40/MXzKClwqsJHcwZLj8ysd
R9IHpwx/HATrscVm9GOz+N69JSMX22zwYFwq/5jT8XUjKBSHWNyrXGvNn9iSdu/V
r0RBOQhGQz/AdsQLooe8kqQdZEFEBw1a0qx9eFS5sc5ZNFW+jbdFaCyqhVA+LkMD
XydMk5pKLY17FoS6JGYcYzhrgs5H+jMTdzzh80OOgS6H4z5GU3mbJgn4U/6txKUy
K9/C2v8p1I8x9CV87D1chwwtBfVysHBtMZZWVgh9TrXlCenGcK0qCMl9xyDp6u2f
SEIq7eRq1WmLn4Q7qHfm/MGfAdx47BZfX3L+SuJYCbSkzv7LmrkPGl1BhyT1nzIZ
zFjHea44m6UM0BzdduHuP6rG698Bz1kc6LDhgqJ2TL4GxU/eBviH+mF4tLLW6+uw
1zfgbs/TSBTV0TQSfHpTn6Rie+wSjmabzabVxBC2M9afZILIyjbFCvJ+3eGFQuN2
hsOA9r4Hhc/2r0aPAoFFooTdGiCFrBeLWNZKvUaTruU69Y2uWrDLBW3T2K9GHH/D
Mz23SXVyK68uU6kFOjJUPwWYZ/IjH4YUykm/UA6VCnS5uL/ohYLlXcgRfK+9N1+m
XZ+rm6RvJZ6PtPJMYmtTljpNdgIjywwgytz5+Lss2blkOc9uPMeexJI8OX/aH3NO
R+ax/9MWv5f7JX5BtSlKgaOZR6k+H7lxmd6gRxepWn/BowTerdtMmx7s5Y8r8Q3h
k77d1VK+wsxbSjGaOJvHmCH6LSwLPOrKGcs4WIXPIzKtkuXhfVtlOd3wrzxhrk0L
+wcBiWV4hVy2n9b4Obwn+ebqTHqLkQQv2txZIhQL823pfkvBdNjpzYkd9YvGGL7u
LV0s1NV8eKfWU3jwCDORJ+oGCJs3imum0YAPmkY9bxZWNZCD+COdw9zcxVgqtCRZ
qgkG6Jfaxk8e+a7UyXAAFQSYqTPJG7TyT7M3uzVKrtHONHr+h0r3fPJq8VU88rR1
3tiWlAiK/GB74iEQp64HZDUs5fB7zVU9d0cE8xt2UvOYtyKYuoC3bgWj3iZNqMLP
E3hVXdAAjy+5oJPgQ+6Fe/M0wUiJ1WrG7I225lJMAs03M+WzFxR5PokOMv2vex/l
sSkJqzrwcbmWPo1n8GnDD9o6uk8GPPvBTPjRj6rTNMYz+QLSBFcvRRfkEn7i1bUQ
54x9w6ry1Zl2ZKOASwrCD7MvozICK3gdFuleFY/mVH+TkCxlhEuozY/OIW0I/z5t
i2g41FH442fPwB3YkyHZy4cP0r5uLzePJ2Rnz7k7HE45wal3GRl08ZYOisgOJd6J
pkoYtJ/Y4yaZZeN9XceGZjRDhuqB8cMFvf3UIUz7Q2OQ4TVxU7SLxcpO/HHSTM+K
Wmjg9GJ83/jaIBRY6DR5kcBdZrj2RS4bE8oZhEAyv3o7+iGQ0CXAvlTfl8s2G8x4
eqDoE0OwckGHS+qbsUvU1lzUC6lV1wSik0zPLwX+j3WBZjXJAyd9MLr8xjBs7kZM
bfB7goi0dQs+Cf47W85/g8etWWCYP9aJ+Ukm86o2OCxCukdsKNIwkjGHTeqEaff+
e+LTsPWs/kznfX9H2qvVRomp+ZhbKXEvFsctWHV0kDCMAr/79gobEcvkI2aAJRgt
d8W3iGoKQOuXqadGg05VLY5lD0QvgWsMGQ6rv6xa+4t+COODRjBwAyrFoBtzdIvb
t0m6HF3KsxkuU8wClXkP09gPX9DOv51Tn7dZoQA4LVo0EsNY7zQZ07fwxMzmORqe
M2c0LpoLiBtSkMSmR5+wFhHoB+fje/hwOVHMhqbG0HqLMpMWGy6ETo16eOA0+JFb
n75iqvM4DJpWUyOLU/ERQpgvTJykQqtrNiwjYpEzYJH964YKyT7kI90wcKHRJBRJ
dBR/80mYUxqWyf9rfT+N4F2AxeUN4GfaoWJS/bMoPKeRFl7lM2j3Bgwq5lHKW4kQ
7e2jdhp1DpLld8HbkExsxhIie1OiAR/afwdD5ezVQ9Dns08GH1vzM8ss99qCJO2N
e6auncWM95e9ZpVxRdytAG8epQnTQ2cKcW5MQTK40CqtbqyfXBy95R5olkN4vCP4
pyK4znqFvZP65dpkEaU3aHR/3+5uoMsHgf0A5v91hpZ9sof9sa0Ba880+4HgNyRu
dRq7lHzKJ6b6KEDxTPSKt6dnKFIJtnD7w8np19MtRpK3yHvxkNbgT8U8PD4HaaLI
aHsF8Nfbprcg1IEBv2lot7803j5NhI5nTPQ8FU79m9eMlnSlyNHzKbI+h5pfT/BP
bd7QhCaVQveEwG5YXpjsIYYkiyr+Y12PUkAEpNgAuLtJuC8/FdukbNOUBRzKEFN+
MAOgjni+gyFU45bdOTDE/2xsF+VYfhNUICUmoCZOKQJWIpyDObUDoQVFWsTizSwu
Y2teEE94Ht+YoEUz7GUiBtPpZYbiWl+pTbqhsloOC0IREpcDgYe63e+hKKEdYdhe
/qwyGMu6DJ4Zf5O3xlzoisFjMN0uU+fw5/bVBXo945JtGBnhLyCFXq+3FndmqbZ9
nOD1UvvvEiR6MoVTxKtxv4c5TTKt95Q3jBbIEw52s1Qnt67G7xWa48UKKiu4FxZb
2bBD++Y976F4BpLMaxyHLtH2hB5L7G1P2y3d8/ImcGiyUukWNmLEnRX23MSEfIVx
6kwd4M5CnbrCKe2Wk0vWtDTGuRBRTsxgIBMka75R9W0CbnMZN14+fURiiND0zuew
0iXvTDNjmrdc3FmMxLepqhb4t8z8JXrR1ROjLfVzsbuuBl1lMBL3qx+X3BfFO9zw
J/Tioiq1zgUg63MYvTAiT7sQihS1IAIjXHumlaQbPsceaBCNFai/kfad8LnzJLwK
WEwjnWS5ppZO5woSkKYKzR46eufv2i/Ng2cH7TO1X8Xr49wcNM+Bfq7ShXaHaLL1
TpE56jnD8vjIyj7YRVFW+DJY3xAiM2uVIPK8l/1UTcanZavY0qjeW3j4LSD26GtO
rRHScsl6/JTccuODm9rx8sFD1k8V0QPGoiXY+b1hnPk+n3OzN3iXVDkdhhc/TBy4
Z+iBQ9fHq4MIvRgENd2E6pqNmNgHaaB6IItrITeew/28BYXE29OJPmrn08tpEOhc
Lp8ZjbBKF42/FyigahCy2Cl8Tst/HfJi8QrN+BvSxB6ao9Uxd/EgOZEfy0/49Zm4
+3BLO928fjIboNOn4gCSUbODAivOvzVakS8xVhmZl7aModDrKKukJuFVGJ4LzqVG
CpenhZnbTXUHLLVcwIQWeC876zQUuI1CnYGb38VVazCPOFZFzpdLH0Bf/4c7ETfe
FwmPfUvokaqpWg0lBe/mHL20YHhhlF2VUuxaRWvB5zGfbE88xRAJfK46Ydm6OWKb
Kkl5Y57I+kXSfytAHyN9SsfeY3uYmflqWK4JOvBdCMweMsd3YbxrJQ2jpNlUlpCx
qbaajPOzE0ftHuOq0vubmVXNiVtvVMw65SrOCzRMU5mgyVa57PtycAzBl4GXEssd
OBHkfj7fC/83dGqWbhI8/xmDzj41LoQNl4KId7vKaW8w9h4XwNVDkGJjbmA4dbpf
0cRzsnvt1uWvql1tpWprjHhTIoRIBjv6XmIDPOrLwUapCrbaWnPLiHC/kvSrUwH1
aweQ95lrABcGgNTL/zduIjutSQ1QHsBKRhPQRmImxP8DuHdEsPdfA/76JXykjaqU
wKyEVvaVXyN3kVNUN5SGsy5k92FRmlvxin4wo0HCQmMZV8yG8aEVtjOpoxuRtRR/
tmqMYcmcInb45YuX1HK2aR/Kew1HCjPTy+qdtol3MKniQYTHfGgKAma3rUwhJ8tO
NxDN6UPhlwWHz0EOq0n7fGXiyXsa49Y5pirB9c0DaJs98YvF1jtoUIYzTx88jhUm
wK0k/wWUtU9SRQ9zZsE8OltcrgN5pchvipSPnoHYa6ieX3CDpUlp+M3wi4J6sc8f
s20JR1K7Qft4Tj5/fu90lj8Tqxq4Yspqjjmyyz1ItSnCtCuP+lF9q7utt14IE2ZH
M2TgoWYxiT1yOeDZbA1OBSZq7CNpA+mLo52xDikR7gDdv1EKF7gPc34+n8Zxj+Oc
2/xAgBJe2hDVb1zaAEJysch7TD9H8FN17FU44T+rS/Ny16z/bflWa37v5EIfDMZo
SrCoQOCtowt3mXOmv/wrcEw51woEcH+e/kfKzC5K3rIuaWRXU7zhR8/z/XWh1XV+
/+4H9maTVo+w4eJYhGfjRQaSmTNKo34BEtwRbBHp9oPyrSvKr3UKP17xPuTbAy/i
ScOZeUcCoEVGTroTwCcUmDALtDc6tx5lQYDDt70XfphKLZu3eLpYifap3GlEB42T
/Q74ys49nW8xQulgDDtEBglg1muau+sLZc4b1DJmULu181uMpaIJs+X4aojwIqni
GzBhY3x6PcWap7oAmDr5/0RLlEl1IZ7F2OVYJbpEkUknl7PqAHFdkKcAdbCiJ8K3
iPuF04m5kzsqC0woPLyklq2RLHAANQpPtpUStGiTZNtsc+pS2ryZz1wUVYCU7K/a
MKOvPvL7vjWp551+rUd7qmv3ofrurqWWZfrqa97LVBr92fKXUzOKq5HYhrbJGXtK
XKwILnktaZZS2b+t3bKsqKJ3htlwZyFTIgiiwzu9aeTS5+NC6bLt1T0NJjslonRl
MNp1sR+eP5oKrQ8WnO8jA1BbEh3PshGOq+FliVBJADzC+4DGHhviXetGWkNl7cwP
Be84B72Yf8RsBUDtjlk70qiQnX6ROGi/FcJYH+WVyevboPSQWd8yvfa3Uo9a8PUj
ssifSZFwii/Mg0GQcvHFSitFmSE6IRLYSiIPpF4j75tlEMAwj/iZ0Ust+S+xRsgp
jONgaIvjph7SOxBXEV9JgQvGdpqLz3KuiF2gqfHFvhpMafQ1k5dJz07AQrhpMhG0
l41N2b54rziIpWO71/b3WVTAgPwi7wGNkMQz2w7gy29yJ4TxYBaFC7XLv66QAswC
3q/iohq/FVzwZkW60cr1jCFNVJCyH/SHAsSJNtzDjmdBDPedDj/P3sSSbxyM1bwf
YBN3TAIm1hC0xH3dcucETMhmYX1ecRoZFnIBkiE+hWY5CFrInpUgQe/ilJeyEFlS
/PBEf2g8MZ4NcESeOh52OdXQDtFtk2XFofyQfFuSI9zRK+WZh+DIsZsJOd0tz8Ts
jf5exxgwYXkjbJAzOh2l2jDo9KBr3yjl9mGrbLEiDysj9IbNXc8x3xTqzj6Ns15y
pwYyYuUuVQck3aCTkdPYPB6BDbuUEKt4fZQEm+KGvuZ8jX/s9aBgkIAW/2jeqQ8/
wPHwbk+paYND87dSSn8KIxLmNV3pkqWflVqW3UR1tbBePbxtdCj5pYxcajXS2bJQ
8FhOH4KdbD/8U0jkJLVBw5lkGpnp4+PMk4Us+jFROVxLCODS9THyIE9YanimCYfQ
17y0bXan6eFaiEtOv/IGe7/6dnmpBIqHYQOVMpr+JPse1w506iG4wgUOKSrCJFIn
T+4enWKQGJDv3J1rDTgYx/ujqaKgSI2q37nxhOOpc8PrJWN2GELwo7K5cjPdVMHk
x5yVOnIhJ6/Gm+XcEn6OCkgfhslt1CjSkxr7rAUXYHds2cWxVXnvWnDNgeOEq+lm
jw6GUlmXEpOqysyPsnHd8iOx7r2sN3FDQE3UYI8QDb+L9fG9V5bLcYXT6yL9fPjr
MUY9u9/MPHKZ/uMcnDSdqXNzHYkWyyav1XRL1s2j3RBwCLR7t9ksVhF62ihyoiYq
NUeoo0hgeIxUTfkH6lnieQ==
`protect end_protected