`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
ddtXksX2+yylW5zu6QL2Lhnb2d1sD00763mmSITNX595NcHTEkwn0zB1Dry37fOW
FufOhVzEJp80NC5qZ/+F0Vk7Ik02dIR0elf3clrjeJRK85K4e3Hoo4xn7YbFUIms
l/8VZSb14+JVGURjfswrIyCUotIzlzVYZ6gzoZwDXIi5gQIBf/gI+KxNXPaKV+PQ
Ufys/12rjO6aI/pPlqSm0hCvftmBcnezN2hk1UeXgOIuKZnogjOsf0iJVX2aOOWE
6pD/psybjbnsNB6kH5uFTA5frkzIzkzl5d9+YDm9OyC+k84E83I/7/j+rk4L2dah
QJOvksSIzN867/4Qt8qYTQ==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="MvBXkzurAa5VTw+1JJ70nePUfoQXBvZOku/SMmg4TwQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
oRtzZL4VJ4iwysPsC8SXYCzXS8Fw2gtZTOskLcDV+1B9Nzn1zTyNtlo6lNICRmmK
ZRVu2BmCc2G+fmzynYlNTnSa7C0Cuel6FYpxCBlOuk3OF2tzAmLAuDyOH3Z1Yjzk
a0aHuoCdIRKv7BrZCdALt03JeUmXKPdOmIlkVGFl8yw=
`protect rights_digest_method = "sha256"
`protect end_toolblock="Jn9CQpRhJt4rnzZPRk+dOpzAubz7omckX1MrFd4p81o="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 4912 )
`protect data_block
gD6l00tciPUa6pDNTk/+t0OO0nC/UTtBwLB41d4inuAUA3i/ALrNyoJVcBnAmEQW
ptbcNp5fxEUJjnOxnedyZEuEBxWRieZFQnkRdF269oNKlyfoVnJteCMVSE7Phj8j
ZKkIlQedSHXQMoFEZLWJ3KuQ/MXU8yLpeoT3A4OBdNSRRm9gNseXcfQ03B7hQcZW
kjhH4RxkxUnoC/T8aFmnkOzsFUF30594UmcgM9tf4LArPQ4ipZ090yUlECZhpNnf
HjhOPsjEf9fqU/tWi3bXnrAI/7L8TRRhGb33DLwF6bBuvPK2tLsC1C1CdqtKIw3O
ptVboPE5OxQUs1uK0SFMwPb286c1urIZPywpUtwCje0C4Y5W5cx3rO7mmrlkxjxs
ki3nH77bkRZiFNU6ZsqCVpI4r68AjwFc5mDYpTxNPBZxLgRL4qOg8RKtIBNqQG12
gPGj+YoArhyegit94+ew0y7/Duyf8iHBmI0hQw5zNP4q92XCoh6tCuwPLTZZ5zVK
ST3E8AqDRsY0kj6p4fu13oewTIYYnjn3WLKgRR24mvmSznuH9SQMlVm4uTdr43QZ
oZkUDeFtqz26nhrDaV8OGEeg9Nom/RKDgkbRgyH1W6AT8NT3RUzeuNv22wF7ZHsW
g/EsI+X7dDQibg2xossWDG9I9FZH2ED6kRuMCt6gA67L8dsi3ugxLqNWY5UxchHB
9aTP6S6vru922c6AJSjugGQJHeMZRC/JjHHSj0hh3LzFZcdC+H+HSIA/k4vdd5uT
gE4kNR+/mJvXfangQN8eGfY+0UgXWQKRU3+NJ41a59/BoS3V3EAr6/OXuVZuYRYO
Fdg4mPrQUTy3eERpITzTf0X5WuYKQOaWZve/1raaOLQiZdf0/ZG4qx2VOU9tonQB
IgGLOsP7ZQc14VgdTKO/VbOWpXY5jXidLk2ombN2FkwkMJ+vt2J4G5uGVSzTwbXu
fktvLAtBuiYIRbStSdvs3+S5TYiX0GDxZg3SWnz/qJ2PFThuz1r7ahxfHMDSZJPu
XTOMXn8JRXYP6wpN+NSlQckJcSBuoV5BOterWPo7HioFFmX/s10gxwwEARvzu5pX
XgoNoAxS0PpvKVfU/rtb42CdDMogyPXwG45a8Xk7DMx36sIGjhP36NrgiIax/9t1
AjKhFBDaLmD0qkpFbVI3xHIxkoP+kcDFozlglShmgJCNPhwzn1fq4FMKuA1HhP1Y
6dXow+dly6SQ1LQV3HYaiTVAEeczLrLfORHXky8L+462wWrb96xG6bTAx8xMg004
wsxCxNcgq48RTAtJXdG49B4Vi5TRYpYXE8nJRaAnBx0zY1qV/RNhiL+ZubCJqMxP
9Na8Kw0ISerD08ikajugRI5ehSPe2r43wdWrR2N2NaoAxEWpj5TIJXlkWX+dSDqu
eDLMPpGuiUFG3hRPdUVOwKNCB6/hn0NVbXmfiOdoDMuoG9X1qLiddWpgj71CgcIB
NYAeWwatXHqD0bAoKOg7OCk4D8n3OWC66BwTEqdDZrW8zCxnOM1S0TfzJIYYLpdU
Z7ykRD5ZtnLTXxYlHWTIPSYRyDGlmNS31S6lEp7PtsHdF0HA8OLotwT3RhcR8z2y
4/pA5/1RWNXJF1H6Kf0fWfiw5WtTL1SaOa62yQXvlzVsKHw9qPJ8fEAaASJfgrqx
hDVVgrwzw84E7mQwoRzRwuKTkoYidv/oUuGNcGnOK2O5OT2IN+0kMrGS0H2ySva8
qRjlLcSlgJ6inKB3RGCC/Qv9YhlK+KK8/tk2dzcz9rSejSBu/Mzhuuw8G53Zli1N
9kiaH2HUpc61iHZgN0bfhh60LWM1BifUUp95LZWQcFPOVbDmkAaCu+SkSgWK9n5I
7j6m7xtwy9k/ccVY+G5dz5fNSCwwBYGnPQ7Geure3T0ZmjJeQhWUeLDewbp7i4d7
TgcmZFDZDTLFR9IFeL8XjEYs6+MFQXlTjhFrxharsAqes4PwacF6OErYVfRww0bC
BJh8zELOtJgPYir2MZ2BzW9KiF2mTpKNk+XWAEoPGhCubLRiBJuTABttF22aJW77
xWGPkLAvSAIcOmuIB/tvYCWB3PBHiw/iRLGyyyBDKD14zXitNtjrS7GcyyPGNgNh
JFsmAoJ21vOV7rTg8r81YFDIf4iGOUDyLJVtVWF0P4q9D/LmHInjrLlGXuHRT6Sc
z4i8ev9n4RSKad6PRExtyxYblsm61F5j3ZqTSUKbz4kTu4CC1mFcSbU+SlMZzsbI
s/hTArykj5UBdWTZ1VNbVHH0PhIbJU/xMot3wfOStCU857uePqw4/CjjPM0PMyMm
hvsHxT4o2pzBeITwIg6A+S3dNVm0zLxIgpolYT0SH5pZ2AjeA0Xv2zltyLut3FJw
SAfE7aQc+UvI94fpQArijqE64knG0AHtMykEbVGcYWkQUAI7OLg2qTQN8qapnOl+
SpsRJhkDfAC870bejTVlsUv08jNQ7MJ01ykFt8YCcvtNArTzsrW5hlDBuGVQpGZp
viQv2x6RA7qoI+nV18r0vDOKuJu7PD/DRRX+/1SA6IzLWhreect1pQzxXGpAtKCE
KAqGsfqCPsKyu/RVhrdoYrSBBRAUHniViNM2HRuXKzAQ4iG2rpCjzJAWVJ/p01tV
DMxN9cwRVTtvEsp5jJeeMJDJMK0i7dZyuwxDcgsMtJJ1q/my+MPfNcUwN1ka9KFK
vzutkEzb6vH3SFc3MVz8CDT2peof1r6w3X9YOss84srhTpVtCSNjzbwQ8XBBH0h2
h9Ar/AnR4b4qB1Qf6BZ5uY49LBJh1twQAmfgnc/1CwDjGllPNbLgOdXEZOvA5mIn
bOEhAaEotRqdmg6w6isAhFFCkVh2HgVjq9Ijy55dH2IOVDcKRlBZ0cD/9FJVdVjJ
beFIyd8Jwohe2UeE0hMbsy5k+1PmciuYkW0Ern425bxQuf0dhpzfLg4Y4N16T354
+fxsZTC/wk8IXxcXV2CV46vudrfr+m72Wsr4wenxdPvRYPzYFNBK1JpedHkQfhP0
QudhIc/2zuxfBPo1DSUCDjDyVt0CV6/J6Vv/djZuZcp78jWHxUCf0PNKVp5NUtQb
Kad8m1UdwaEycMDjlw17R2e2V0VsLKamZWstvWIzGo7/oIYcWdTFzEMFAakZycDF
EXKjj1gHViM7ojCJl5564ldNa2AD60Nrozvz4ypKkCLYqURNsk8x173VW7bTxpgD
EHny1tlRb4vYgWKfT2wOaKXzEm7u683l2PD4ZvMYtQJM5PkbOxhkYhAgsGDx4gVy
6VtfWA9YypPW38k1vjLXEs+246s2ZOXGxR4MmtB+A5qqp9xIiuG4CYGJc3rDkMOx
dO/+0PINs/fiIjrMrk663lnk2g+U2Y6fTo5rGbOLIEOMi1FWcK+gUhYy2ZJldGQb
9w7XHD5+/1DIFXsjBKmuQ9uRpMvMM6FNGGaZW0dcdQ0+BcxPUX5GWAB9aPGDvRXf
gj1FmhzhdoklNpdAUkPfmCFZrUQy+BJKclV8PhAJEtjDT079iQG1bdJAI1EmQ5Fi
LRYfY1m8MTxmbVIpu3TlocH4n5iBcHMY2I7RvXbKkWzbKSFpwB2f1dGAnllawSJR
QNTuOZUq8PGVB3Us+O9Xir4AZy8BLf40+XiFpWnqUYFf/DytURLyGWaf6++QC3vP
H3dJvnozVS1j24yEI6Dfr61l9lySafeE838274SINhOe448B1H/L1rHH4q1WDma6
BMEAPa9DD8ISmIdRXL/pMxa/lJO9y0u93t16DvZSd/STa1alltxK1+vEkctEYVWw
9gK+C+J49daT5egfEsh9eL0oQYcHZKUICbeSTVuib7l2lK8suflTP6/o87reaOcA
7JH22yrAwfyfzvfLYStNyxJs5hvFyB9rMg4jUKNtKPoFnTCfMQxbKDL13KhzC3G0
VeRQvVmmrw4MV/QnFwdnk1PS2yjivLHzD5z8lHNUCnjhKGaNdbQoPEa04ekf8bSU
HG4SRjtrk07ftFSB/pruDablFmJ5mCSUm4+jLTSlzKq75DY5VfHdiI2ywuiteV3J
3qfRx8uS4aNnXjRRM3hQOrqSJad3wB8sO6gWslqAT/rr2lvcLPGK0FVKtCipBEz0
WVA89Xv6JEpKtqPn9A9IcLzTwIPw9aYJf5j4UKW6wh2U6eL3Vhv5PLaMHnr7anyQ
T/jYrJsQa4V9unnBEw/ah4zgrZvmXjU1lLVg5klL+nyXKH49EB+RN9r0uZQB0IeP
fB1b5bhC67eXL1qUhM5W7BjU9tIl/sZGRZyQW76X8B8bAcWSUPQtbBWLC4EpbI7F
IFk0RjeslQ+KjlX8B1maeuDPwOMe9Kb/Ewa0gXbU1EWbIO8IKITvGHxjHjwntZNz
qMdQb6Wqhh7UWQxWUFMn5bd3V//qlanKzrhvc6J7dF07VcU+5Np3dmQzXcS4n8pJ
GUZxYBFePSqpaOlP2PZnbXo0yLhvsMBcgrEovjmqloTuf6Snz6R2yRsVEHZzDRx6
qrxd5XTFjLUvhwDQdhOf3Sfb7BCpUBiubyghB4OdEwndZX4dnyU8pdSmmeiSjs/A
1QBTw35DQ2rO1qiG1P1VidK+8ufpiUQh+ZI0/HseLvuVE8ub2c36LKciwATnlCV5
q2HkmzN1s3kC+O0HCfnAQxRkxwJallmTJa7cy11fWgZaZmim5BBltv3y1ZfuKDwO
ScIiaRg7LoiNrzIe52lNgE1glcegQIZfFxR8T/DZI+EcS4pt3ZeSfCWwpzOGvwxg
smSTQypDQZnWuzMJPERODVIR/MAurJTOcgwYHcxEX/7pwkwUYA+x6lbiSImyBgAP
zzJE+dswlz/ntIqrM8qDLXaX5HQTyzpJzryw/IVLa/PFH0hSeIW6U4e+BBfcZy3q
AI8R85uAzuB0EKYs3nPpSKybULOd/DLodCGWzVFCLjYy0qWW47GF+w/cG3hAIUbh
lOmUFn7UbRuMWif5TjvP+BQqT+g5R1bgXo2NQvSm13BaUDRDBC62jS7RJB0MtYF2
I7MZGB8j1DVkt4AH2vOx/HFgPaEqRDmzLIERUq7ySgwE5nEqHNnndeUoYZVjOFU3
4sW7bwfVhsWA0DiWmq2oRKmfCdG67pk3xFn5vrQOP90zASOWQj1aWIKIePPDFJor
SpRSoyt2SJ8NxOHGX2pm1roRARyvwznR+pAJ3+TWVMP3MPFQCyATF0twkRXH33d6
4a3VlhQlthudOjC3xZkydss4nJ1mei9iJGoo4ljOPA01SH+l1GhATU2B6aifrBiq
29DH7AOyTfBqlaudjXudGe/DbLpRmJ0ftEHLqcLKKxqz61XMBURRDSmw40mOyEW+
8ZgojZp8u54eDMQ559B3/bed+V8cGLhUVc6rA1j05WP4YAFPDOjRj6s2UKsqJ1+m
LM2DMgK3HeDo8c5Oo3eb+CYzt5CeQHD+Q/xFRx08JTo9O/lK+rxVmZHO2URIveJ3
o0L5nWSMhCCQIbD3sXXRjdlMDnCpwyCkHGZg0RaRA0UXnQVENT84qwtdWO+8nyMH
NdhmWbtwSGYUtrgCPNFX18WNsD01BcLkBvUn7dElpaDylE/N5dUX52GAaDSnnAd6
U2BLHPCm0DVXb6GESq131kuVjU50lqqN9zV7pTBDPKFFlWvKGggF2bksunFnDA+n
Djh1c1GmsH3YXUpeTjzm9zMj3PGlyOw/Qr4RiT/CV5PIKKmPCTSolgjdmJdT7LFZ
hRFUHzfmhb9yOYXIPp+qGHoXLm1ZeL9Crv4NAKTQ/xxzzC0EGUqHiGHEoT0t/tuS
yoZZFXk5Fz0EPTspmq8lYmi4K9wbaW3c+ggTUoK/mJ6uzCwiGDD/DB+zi9t8iDGb
wQ/eJmGqmFzi1ymoFS1TJuM1W2hUovs72/GhHWn94FrWKHBRGUvli9GK6jAfcwlX
oKozpUSyHgqjM//gWqv7Z0Sd0o/6+/3agB0KX38kxQAcRQOUkkFFqcR6jTDavciS
O5JdthBmqEFrBM22WyI8XC5I97mjhw9VVoYTvY0/R1WDNdBi0wZmP69eSBAg3GhA
7chTD9S6RyC5kX+PAquXBXcJjT9fjj+9G3+20VLBOydto+o50UdQ7SnZeh2QNBSa
jVhjRBXcJmQRV+lGXkEc35T85N3z9XLbJ7Z1THnOZF7ya/YJ6FsRM5yWLDe1/xyN
Iw/IpAWeKNJX4/j047JEf4TkHr77/ltvUfWtbmt+b2o5q3JxX7EaZgcRhDQKvHTs
58UheUWV3a17Q3VRcnC26HTWj0iohkyHiIyAfibRd91S1lnjxY3JXtj0BBrar1ia
OJLrgTOPwjOIxcN++TyJ+2S3hj4iBaqoH+Bp7dapo0y7E3N2y9Z8T0f6DS/SF5Qs
kuwYEx89CsH7qSJI/sFqYzj1MKR0iZ6A3jF6ww/ed5Wm5V6exodaBrSOUikXfL5l
CE/ku6BeMFDqQAjYC+AnXtjdXKuEJ7A2/0AIoZ4FwFF+4KAFE1KujN5PjQ/BgCo0
BTdkUFT9WGdFtwMi98iGFQxChrjLG67AgJHIZoPH9LzM2DTbICgJTKmBc5loASR9
CqplDcIpO60snwtWkBo0rw==
`protect end_protected