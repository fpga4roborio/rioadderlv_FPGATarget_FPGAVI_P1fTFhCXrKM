`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
ddtXksX2+yylW5zu6QL2Lhnb2d1sD00763mmSITNX595NcHTEkwn0zB1Dry37fOW
FufOhVzEJp80NC5qZ/+F0Vk7Ik02dIR0elf3clrjeJRK85K4e3Hoo4xn7YbFUIms
l/8VZSb14+JVGURjfswrIyCUotIzlzVYZ6gzoZwDXIi5gQIBf/gI+KxNXPaKV+PQ
Ufys/12rjO6aI/pPlqSm0hCvftmBcnezN2hk1UeXgOIuKZnogjOsf0iJVX2aOOWE
6pD/psybjbnsNB6kH5uFTA5frkzIzkzl5d9+YDm9OyC+k84E83I/7/j+rk4L2dah
QJOvksSIzN867/4Qt8qYTQ==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="MvBXkzurAa5VTw+1JJ70nePUfoQXBvZOku/SMmg4TwQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
oRtzZL4VJ4iwysPsC8SXYCzXS8Fw2gtZTOskLcDV+1B9Nzn1zTyNtlo6lNICRmmK
ZRVu2BmCc2G+fmzynYlNTnSa7C0Cuel6FYpxCBlOuk3OF2tzAmLAuDyOH3Z1Yjzk
a0aHuoCdIRKv7BrZCdALt03JeUmXKPdOmIlkVGFl8yw=
`protect rights_digest_method = "sha256"
`protect end_toolblock="Jn9CQpRhJt4rnzZPRk+dOpzAubz7omckX1MrFd4p81o="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 4992 )
`protect data_block
gD6l00tciPUa6pDNTk/+t0OO0nC/UTtBwLB41d4inuAUA3i/ALrNyoJVcBnAmEQW
ptbcNp5fxEUJjnOxnedyZEuEBxWRieZFQnkRdF269oMbJYcnsRrAgKSZL3b2PEV2
r5t1HmmOpZ9xEWcLAFqq9ZVedZRyAt5M0EFckEjpqO53lWs7Trep2QP3fhBmEOd8
Jqed93tJ7d77nnd55sMhJMBv3w33o+WB3Zdf09cxXT9yWNe1X4R2mGhsQ9ff8X5Y
T+E/doPc+kl++GGzqStiFrH64EaX05Hha84tjt6CzTnE8vwRzlVwhV490fd2zNiZ
mj1KiLhPEnRjvkc0gtdD9hmqh2srHSpz45TWOUof7kpra0TGe4qn95pbx1ZKPi/V
xUT75mY6sPwNawpEHkWhyrMdybaLjEwZQCQyWO3kCNv4FfoNlZk3AEME1UdJcziv
sK3XPXDIaDboFcauG/sEjhYHZvfTFgjBPxD39UzRDQc33TFV7dUvxsiobUb0CLXw
gHlD2dZMkq0gWvCATEAG/MtMxJydpMkurNcBeI2sQGq5ATXZWj7pVrKpAQC1Q9eP
Qpv6IOxP97TvgfcK4POr+US2oKcb98UGNn/I8ggf/qy8DaIXYQe8vDgZSu0WNr8g
Qg5KCD4KG9E06AmI8jVJUkUyeJUqxfmNp057kouuFghGp48U+c6pO+zFXgk1RrNW
4o2GEB6pkzruMXj7IB/dZqkz1uZ3oLOMZWIzxtlmqoL+8zOtffIBQ5YGAQk0C1gr
PxQny4tEJTw/o3hqWSlNzmmb1s0aRxCwnUD2oRIi5bnYH7quBaEm5iq0jH5MZhmY
4dnsMBMqSxoIC2xrLDDPUIXtygjnvVKES6FsnECZIMk63+hG3dfyWhIsGnsomSEW
nr1MXy9rjWqj5G0rRYNSt7nq5zURJaoXiS1nRxV4NWcgfVdOlT7Zcv0IGkZUMYJE
3l/JTXkRqVFXRcAqBnKqG5oa3brVxxffcxFEWOy4v4jF6aqCv7rvjtBMnKqY03O1
Oe8CHVLiPqfNenr+iFVBVGH85xbYDH/uE49tJCLFzY9OS8QHLgSB2hYLW0ijsiug
J+MALhxwAA+yOyRNBvrxEXMWLV0viLwLRZvxOfFX19UzpmQY9ae01g5zfboGucuy
TrZF6Dm/ae22dCVGf2eyuAn1Wp3s5fVUIkIomeYj9vqWOzQK9+tKFcm0i4hjwFHc
bJBLBdLMV2PpF9DVi/9jyVGhuw62BOemmgP6tSW8eKEXCJovPaSqeYoRULDJMbMX
1LikoHoj1m06dlimqq7I5rv+A5xJknas5j4JIjIKUnkHCMFpXaQ3VLXlJDttSbO4
gpCEiXeA/wXmgm0sKE8QQootp/bTrp/sjzMfxD284gQXuCw2E8ki2xiTIFO8D3YX
JX05rhOTROOV+3UEEZmne9Ut/IzL7Us++yo/0s0tC8mdMi7tvUqX2im3KEMUgGOK
+ON/aPOxNECN87EMweUiM7czMV6J3galVwoX0rkOGzIz29bL2tx+piyiEDVlTCCt
EcFrPMGort4+338ekdQJWsa/WsIZyXGHH6EDinIJ8K1EirM1d8IVbK4OUsxjFwsO
ocJdCiPEcmrmwKf6mpdZK2SoB07alX4eA1ykTsF6zMnWhnbDZg43VBZZ0xbPeiqm
htqvTBsFxzqLWqLDvohQt9F5kWi4NNXg4VGMyBCDm0qCYm/QPUNgtMhrATDwfnKT
b09kzO4zAf1JDCytH9sxDRN4jdpiR9J3jLhBZb6IQCOL0ruwjGtTiqExhDyls8kV
+xTCyzBy6RqSHu+DswpVLmH8VfUc3K2x3+CAfYRHf/R3ajV0p4SNOnIi3DSBJ5vj
n1a7cDOR3pG1otZMhd/N4/lRTOi+ekyosvJ1Q03w+IZdBZOTR0VngkdKBQ4QMclz
anuUx8VFrmYYxT1MBvTLb2qlBk5Pr1ysZb6a2TYfTFjT+dfIxHmy3hQ54JXz8rZU
pYQAhI77joWieU5BZwdB7sRYdAXcSHlCUgqC/gO0TEIabAt3ff/JBI3CweF3a+iX
YSmcyTYYv8xnqQgYz0IbYnlCaqtMYqAKfXjH3yTQFLTgZrmvVPv4c+ZYuAgDNdYs
Lkpcxn3bu7UXErW16jlHy1MIFhrOmTeBGggU3B3DOhpc3vFItFmcjxM9/lgt+oTg
TcvHTIdtsxTMtgh89yLw1LOHhAYCExPFFHZX+bGPtzE9GSaqIqBVoIAnJyM5asay
stvBvSQjRwjPOwggvS+ibjz2ciCpTI2ZU6Hr46sf9dkhdQiLT5yIsR8e0Uuh7D0f
YcDHIS4ZqqetT3+YN8LDEUT4b0gZuVLPRzm9ah0GF3U25x8mOiFnEzWMA2onkZwc
WMEtkX2ypXVDB1gbhosuwzpe2OR64O3q1fOWrq5Rd9T99Rh2BVK5j9L2FRKiEOvH
R2eUOLqQZKG9o0Vn4dcojBp0ZMX1saQCazZERU/bG8rd16GPzOgHqKKDldlwKZj3
HSlhiSuFRjKWBEmwU4k0ffA3tNUD3TGbNK+z8vkJg0jXQ5e86a51JwnHYC0RFYAO
aVKDqz/SGztm9wN+0jM45HjV3xnwB3Se71HCQiENCHRFYijKks+/OJHKaYp1E1PL
0pWwj3amYtUW0kR/x0uIZHdmiN7wmIoLmOW1KSioTEf2CHY+drpP+AcvELns6vu/
89BCfPPeF9lfbODwcn8ae+e2wIJz6hbx9rsh0B0BRDoKqiURstVIf9lqX4PMYPLJ
StHh4gyTvY2PTfKzzdP3z7rd+Q7AkozeoRFV61fYIhqPuh0GOkxeQXS9IGQAboS9
ol+XL23Fep9bMT0F5w4VAr3GIvjTNshLBYF7VeUDNzpE1qG65MrS0dDSa7Bp8a6Z
uiT4XdV9aHVU19ZSF7Wingl86AJg+yjM5XIDEoH1ZgLfEewsTDjtQyzOTOGuZYQt
nZ7sm/ZW5/sMsY4SL10TpQ5meh3d6jpqQ65KUIsQQ5zctJaohoAUAB/W2V79TXBu
qNBB2sIeqVh7DP0hhLz/X0SDGtvRB4dWshE3YPHHzXhe87wlRkDxfIlrKp3rMkHb
UhPwCuy/3U8k+x17ixeb3oFAY9Ra/fFPqK3BPs9usB6l6z2F3LnboCjn+kl3p4bV
+66nkfWk/CqEXHl3izZnYHvWzfECIyXdChew66S1AxDfL4LVnWi1Z7EQykR+6X/p
j7qDM/ejHdVnDlRQv7m9mP0u7G3/CZOoXkhgPx2Kknf80po+6VBzV6GZwthD54qc
w4qAxqsTSXVsioHYZuZB3wRBodgZWLopqYE53uIer8pX+kH0uZ8LovfUWdbwzc85
SVIpDipWxKx7eW5ideJzPNEWxTeSP9+w20DrAxSOFhL4Oe321035AbvRLJ+WCvMl
RUBU4tPY2+SgZVEFPMRm2+mquwXKGy1rF1l4bw+372XrVjHAHPc/ndHz0r5Qx/0F
Bx1ii+wAHO/6MEFCwHUc2q8BPkA7WtBWUquimxHzdHw1+JYnebxZ5cJdBEkxuqhc
EfyUOpe8vw4YfRbih+i+hhibYqudd4dUTd3XO1RbAbLVADVBbxcofL7K0NKmaEaP
Pd9nQVG/743tPkC2gZlVpOkUb+SCvFApoa/EyfKmPy/mTYx2Lk8Mpf+W5/9jU5xa
oDeZ6yO3vJp2k4RTnYNfen3BlKom8Mq+xEoeBOjD7A+E/GYoIHle5I2qGzfx52LZ
i5LCZtoqZD0YIp4/V3APrC2mNbSILiyox9PgUumyc1MzSnjaplmTodxJpnF5x8Z3
Fc/5fUY2Hj6PGfRtNxbJfUe52Yj42oLcq/zg2Za7U5Avw7Aku4KllnP3NZKFUaFR
yVnhH8cegBS7my3Jk8ETKiOY4LChSvDYQM/kUxLazV0L3W3NaXvwEzrDSeX28G0h
vlSNzqaZedA5aPiWzqh3Ubr4VBk4Dw9zB6A4z5O2Nzl5NxYmi25OT522zTXRSMyo
VarKM7HqOtLSIxXYI3PdU2xDhbf5gcNfmo9OtuSlRAkbnXR/QJ5x/jch0eNQwLZJ
cDKH5hKxKL0yIo+D4ujgKH4FUAjy9cFVcziELgp5VdWsl5lYolcRGs+iJdwpEkPR
uw4/79LJ39dVqJrJUzQevsjcydRiOzX7jhxpN40Bx8J6X1+pWkzPpIlJqvl5NdVJ
/joZJiV9TG2DZ/v9IvFBe/vjT5FOfpJYWnjUpFiLYx85ONL2Q9P3g5U5pXVrRuqz
MOlorAhe42n5j5zLjcV9SDuV2uTH2Oa2CMx/jMz2JipAIGUN3qPgySdBFAHieSQm
n2bRXXdR2A/34RflC1NvcQxE4ANdvvWNGINweaoMr4K7e1DAoQfLdSO6Ts5eoLr0
uQDZjdtChvuWZo6/Zqz7v1ABeC7xsAijGasjk017DS8jkcRnbTZRkBYzv0izYuvg
q5U/UnbBHufAkVqmwJmKHqeOEKYa4c6kdLxn8CA3grXb+aZunP0iHTfPWBRV0EO5
8zljIKpupMDZQ5Mwrajl6ti4ytIGQYfC/kOgXNtCKBhOFJmQX4F9IjVczpElW+io
FzyhXpOsDvOrzdSaNY2PM9+21luk0C/2IYUJQnuZzenTplRxsoGzqUpycK21snIZ
kzuJsepfu7nyXKcwoA0lNlnyZzmIIX8e/rTi39mxXzQ9awndp5n1vszy01rB5zBd
fvP9+YNDj+GY1LZadeHJPMO458sKufGOKgu0bBVbo/mJ+WAgzJi1N0pOqsGdFGD5
+KPAVLPLqhCbco7SLeUqFFNapDKvQxPQk5G60I/YfwuccgPRZrxPrSGQ7RWXaYsq
8aVgS8scj3MioX7vPAlN7wbOmSo1NOcidzPRW/vJo3dtiYbu4X5K8HMvXCplnBpy
svgXpSMfm6/JD7eNXrhGmBfUwYi53GWzZgifJ8QbDOt3yincRjHyt0AjVqSdtjMF
lvRNuWASTUkj2/Pr4Tdzo9Hazc21IBlC+TnSQCXeqdwIAMg9XWOjz2L+uUtl6ClN
cjkwlhOTERSws5CZWlPShRJNXifHmd5ojCFlbrE73a7O3TCkGTv0DD8i43uf226u
jFdR0Rha5qN8i558OrOq5wHrKgED0oQxnwA547VjtAZW7ABB1IqNx+v6cNLGLSzK
mIUIJ7uEt4fYWajLdm6ulyRCjNJzH859a4L7cx6EWpC9yKyDPouRNLU4IJcpl6Hs
1VjbG8qRafrtYXTwwk2jRRcxrbMdR+HyTUjTrY4e68+fWsoy0mt8290u8EWTpHiT
e7P8Xz4o56PsiiF/T2awT0AK5ulK0yiKc5f+xJfUDTi9Go52aQ1pKvLiROO1kPnI
XRtAZMZ04BuFUm3FsVCRIS0A15Q7fvZAe/cYrIyXViJHFGcB1TI8tTajPGno9/ic
6pk9KjacIJn5np8XGpXYHOV2krHOMeQDSPYZhB5GRkWEFsEGqaXXacxZ+UI3YFTK
gc6jFbPKeJSv1RJcskI27pFHJaeQhqKnf8en8VfLzVmIahRcdWG4JNk+5ZP2ISI9
u+Dudy2KENexSYKcA4ZSYdZ18RF2CNXFKDMC+deOhRvS8cxMLxGm5LaLyZoYcCHJ
vjyzZTT3cHmIQg25F7GocXcIQ5vOE2dbcK4p29ev4WBQeTw80VVGH0sLzmwZBruy
rckC/y2ZwvBCdIPpFdQme7vpvN7hwMz9T9yA9MvVShhS5Oa6XUV0oj0uLb59YkGS
GTURVWu9rgVMfHBr4iNSqBP3Zvgz7kkmAVeinrYJLEeRwHDIy3BEPrwIMk1owQHC
45qN+Fl1mEglKi/GqhCE7hCrVB7ueft+/yOpGDR8ZSthS+ZOZWSDjPLfAE/aOcvm
UfoSrYpyBbvEp8Rk+0ii93My7d7fN5LwaPTxycCDbqKFP5jH1qhafFddg03EVyBF
UtXiguSseBMqJQBprlqNZiAdMO/pHM5xlAalVUCQQoQbCDRZe1s9zajtZeUAZ3ht
pZP92Tdwfj7WZwaVwvRAAPxojN4sNbQyOYfgVd3NMC6ybX7W1o2bbycG0bDrMUl7
CMUlG4Gq4eC3TWsuPGLUe0GHt0mP25cVhWFbW7pDQgmMEu30IS4/VBUC5B3UI3R+
iuTKtohHpWZ0tIXu1/jtJXlVt+TNrJZes4JupKQvCpO1vFou8p+7rI9tHXGgZ90s
m8+C4Q6ztmdA1J27o2K08j5Imt5AW/GNWfikJZY37GFBC2Lv4A3o9edWElch4d8G
lUuyWliEcLUy06rhLxdZp45fi7oCdqd2+g5cc5hBQWoG+NqFQ54rsS5VIelIecM+
K+u1PujzfdOTGZ7gWu55eDRhRuDdbRyXdKFK5SaJwE+oS5855OdE5i3HOmO8zU6z
Te2pPwOZnWgJ9y/aJKmbpbwfR1aG37gM1e7l9Lm6Y+f09uqw26ZCRvmJZee+u12R
HHdH0l8Ebwa6glYwPx9BdcfqcJo46fMzn3jhfwyzD/w0QbyGMRd4vjEHq9lmRNFq
2LQuDdrt4/I+vIqApZN3DKxZbVOMCYSxap74ktcuV8CpvBBf5vzWur6hRc2yohm6
CtpSGzy0+0absiSuxjrANfTsSxVbtq78CsR9p1NpO7xgiU0Gbde+M+YCX553R7WS
7zqzQZKrEnL2krXcJU/xN7pqNKoTSkvsO2b5I8C2DRPlBSfLZI5EhhXXb/5NWcoE
`protect end_protected