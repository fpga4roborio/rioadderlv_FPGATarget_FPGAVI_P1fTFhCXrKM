`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
ddtXksX2+yylW5zu6QL2Lhnb2d1sD00763mmSITNX595NcHTEkwn0zB1Dry37fOW
FufOhVzEJp80NC5qZ/+F0Vk7Ik02dIR0elf3clrjeJRK85K4e3Hoo4xn7YbFUIms
l/8VZSb14+JVGURjfswrIyCUotIzlzVYZ6gzoZwDXIi5gQIBf/gI+KxNXPaKV+PQ
Ufys/12rjO6aI/pPlqSm0hCvftmBcnezN2hk1UeXgOIuKZnogjOsf0iJVX2aOOWE
6pD/psybjbnsNB6kH5uFTA5frkzIzkzl5d9+YDm9OyC+k84E83I/7/j+rk4L2dah
QJOvksSIzN867/4Qt8qYTQ==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="MvBXkzurAa5VTw+1JJ70nePUfoQXBvZOku/SMmg4TwQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
oRtzZL4VJ4iwysPsC8SXYCzXS8Fw2gtZTOskLcDV+1B9Nzn1zTyNtlo6lNICRmmK
ZRVu2BmCc2G+fmzynYlNTnSa7C0Cuel6FYpxCBlOuk3OF2tzAmLAuDyOH3Z1Yjzk
a0aHuoCdIRKv7BrZCdALt03JeUmXKPdOmIlkVGFl8yw=
`protect rights_digest_method = "sha256"
`protect end_toolblock="Jn9CQpRhJt4rnzZPRk+dOpzAubz7omckX1MrFd4p81o="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 11728 )
`protect data_block
gD6l00tciPUa6pDNTk/+tzLxvdHE2s3DQL3/JqqujQBC/Ei+vcAB8wM3doqg5vTg
mdfn9XB1bLOis2CVSfu295W2DNwHfMSTc/8BhCDRnTlLIX0UCJs9Za0+LoM0rMrV
T7EjVWppbP+Em6PkVKCwlmIQ7JKaifJ+Y+kjw9HCGboYo5074hY+K/CBbfsBQY86
DFekqOo2vgag6ud273wY66IsUfUmcIL60SAgKD4jrb73rrvIm/ZCe0qId6U0AH+v
SXaV0n44UeB+tjwJgX1JeaFfn1dA1CqQ5TSXbj0CizRqk4wqbTnh161OlKURAnHx
qxHxRQ0FezcyHYr1HyCXHIuFMh20Eutk0V/WS9efllJm+iofxwAsDp21uYrgrKwk
dGwjEbc3fCJhXpiyAzbNuZra3O2l5nF2G8QCH6iOoTMEIluy5TlT4EezLjt+nKvh
Uz656uIwexmutHIBGTsYx2Z6sI6MoCrXX7ZqUw/ec3kgAJ/oofxCOM/CkKI8L2iU
cce2HPEqb6MZOdnUDQeTs309TqxzSm5ApW0z4NVgn6eR/6JmhXbr1raZUs+FhkX0
s6moK6AKdWX7J2GNc39vDs+bba6V+Q1n4Sp8Z/tVs5SOPeJ8t3p7uY6UglFpge1S
UmVYROu3a5y/afaFzEx4Tr8pIf735fIm6IPfIaOosy7Xz4XtXCR0FJkYgNd/Y1jv
CU6nHU9zaddOgG2pn/V+BunoUuJlneuUMkpUHloJCaxsdTjKSQFrEu9+8kxxDfwp
b/bB7cHRgCQKbOIjKYB8eKD8EHwi4sO8KRghuR3vxtWCu73QFkEnMrAEgR8oklz1
UWLeDdun4k3Qa2Fvb1oAmH7vnQ6pNBVRugSUv68q3s9GQys9/mytBHUN6pxuM1YT
QPsf4lvSSwmBhzDi5YKGoOH/12PHVCiVv1jNShwJMtQ+SD3RiXFIJNCa+nL0/rHZ
eXlEAGu9dvCQHcxCQDyhNJqK08E2Tey5v38Rtg31FfPilwGBTeJw+qQeNee99m1d
skDdImJ61aNm4sel4xH5gIOx90Hhe9FdKDhqkHoLV3YnPyK3RPvSqzfSDtkkY/Rx
tJGDgiq3cgSzExPEugWQhS1JkpKu7hc6oawiMe3ok5rfFlpKKr2Linh9rQ2YBHJI
XfWuDj12u+GuUWxov4GaEeHxc/F2+G9jR+2msBuj4AwaokR9YZaBQqU3IC6zjZ+j
ALG0XIqOVbwy2wOyrsRTtXrJbe0kdwcvjbUx8daTcnzxV8m6wnm5K8K0wGqVOyuA
bEJj/VXs7Hd9t9hJXWPCFgzYG+F44fLoFy9yS9W3kCjFfRPBa3B10HLRuJI/dT3C
zR/8vaG1V7XHl6qY/fSr1ezqp14tuxvWAZ5Ug/m485NBWGtwomG+6GYySvYPd6sq
UtEROIIm73Z9ngDzaDwiJB/441nvRhHX8Tkuq1/3ytbX1nylREaANmsElO44etnC
sxULhzZs2b5R8rJ92axYuvBxYI+z0aB1ETj3TQELeTz6i7Po/9FZB0hUWinheNm2
nlOFE9sSeGqmTed764TpmEBa8/IuKSE4yb5l0XN7cBwktyWN/6QXrXQNzp8Kbfnx
UuLUXlvG7498FrTEe81lJFscQ8Slnf35JA7L0t2Q7QRpLSzIWJX4DGhVMAfoOmUJ
NQ3VJdt25CqxX3wP/5LWRmdo5IyINB37VQZ/B9BoBE9NQFt7gCfaoEUjd2aIGHaN
MrVeU+IAHOQ6yEusnsSgAZYyK/rki+bjWLQiPLGeNm9COfTCB6b3PsyWLRQHrRAv
PQpTMZhKILNYJ6ychosB/4e1AIopy+3b77mbiW8ZMuAcLNKR+hIeUqYpqYv7ia6u
sv0U1xh3KkNonhmnaUVpQDuCDFtRXGOLxXaj/K17iHdURuFb35+yyl8ke9AtPmQK
YOvnmLM0d7GtNYRaY8aNfzTmRZ+sgI+EvZezkcNewF8M0zV3UcClKfDrsvtcx7Vm
WWWfXU5a16u6CKV28jjfSsQmlG390twyPiIXOdykOed00Sfw7F9LrQzODUfYZsze
3sSP2QlQYTOCK8EFLCHv2PG7WvrnbwyWftnNtpuQ0iTsVKmzBxquOLRbugnHRTXl
z2SeJXMZiWMIyQX54dKyvOnTb22grQM3NFSO5sRfDyMeUBBU+Ar3IbfJWUdGGFI9
6CANwDJ3TE67G3lNf5QB2TgTI8lioPoaBxQ/qV3r93yLq3gawlWF8I7jRWZHfQ6p
QwiSpHLxFwymrgsqk6aSbRAkfiVcRrsdAMaCmx7sNN5J72jhYJh+GVZA2OxBVhcY
X78dzBJ9lPrY+oJECXpczR/CRzifNwt3VmeJEbBbxw9gV5XnUQe5mJEoTrJfA6zc
ScxaeJXtTZk1tOlBsRPYVYPd48qjE67WQYwO1Eno9UfSTcJFe/zZBj64T18t52Z/
zosRmNt//ygPrSVnsNR3furpC+U9yhyk+8beTaQKUdrnntBUftdm6W3bjur0mN36
mqt/JmJEb/U15l5aelTv2xvyNhVnj/mIG4NxIwN/FarvDQzFbArJCGSu6I5cbW/y
MggZ7w0U+5DfzjGVkKgYS1bIrD5Rmhm+1PMWGvRqmdrr922Q5ZXhBlUcWnZA37cY
eI1jK2XItfZW/4deJ0rMsP2fBXDmQJy53aguwy6DzlvJQ8Fg7oJcekfhzFmYvDo9
xE1jBHiD9lX4Pxlu/jgocmQB32G4X2cym+YI/QZjdCEbBcH8/GS1u77S5V9CApNn
CIg4kLsnWSge6WWLaipt60bKAR66MskFMKIuHi0X8PpiHm0gxn8oV4lkhm5YuPPw
WOPu+l10XDBR+aUlaxcQo8SZkVgxc59OIKdq4PwaQTk0TLsES3iYiJGYilCOuQhl
cLmYESNHj+Oou1dtocx5j2nl8tRBS9iTOEZ5KMKZrVo4DUhmpBku9iv9ugOrX/zx
YZcVfTV/U+ApTmJLu2rlpCCFTeh0zbmenpmZz/uu9QqlKf3lXfkHsZwAsLYtftJS
milH7fQtYHbgesl4IPj+F7ykLDL6kMGfhUISgh/e1TmG4LLIGGC0sFMYhL9o+HDt
diPtbv6mpBdvUIiZ7LDXeDQVw2/ZTno98yI15kQW5Tjtljw3hxwDhyFEXMgSsXKZ
6dVF6UHBOfvtibMajKAQkKnLRNwMJkMuBCdcLL0LfzcytOODNQSM23BzFiatP1ua
aPlYh5p9v5b9f5ulD8FUGxrCTBaorOsSNKy5UAclcJNeJCLu6hNv2rmlIkwraGM9
we0k6oGyseC+D8UK5OxshtkG6Tmc8v5De24lbw0+QrhPHhMYxZ4hcMowH43gZgcc
SBbIAEl1C0j1r4Vvy17M2LO9+mOKN3hESwIYDYBC4h+Ve2qb5igp8BMI+0A0n5QG
NxIs2GETGeBwxA8j7DlrzN7Nqha3wzYABvQorRfu5D5jh0g4zt305uMo5NQzm7HP
HS/hPrNDROW/tHPTUtvFjGWlIXf9zrr0BaV/5J4TTHfWFahC2OtOxZHKgoXmc1wE
KCETjPL4Q9kotqPqbMBFdsRK6EAkZM9fzP2QWk71zA5jZkKGtcYAVMHDZUzmru6a
1OgvkFHkR4t63v3GaUjAT5SdHOuBZiSx8bp6e/KssV89e14db2HckWwm32Nvy6W2
4WNUDLgvmFU4YrUtk8rw0Ph9ZnK2Q52LlNE46iWebjPKkj2kHNz7rIXcj9NoiFZs
8V7N73zbLMC8nYoSBUNkFdTwb0NjqTFuAE4yVClflxwkVBEdc9hwgzING2mZO8u4
hvZVoooy/ZYf4dfpmxWZCshQtplYdZUtYW0MtlfEU3TX6ny/ybJVT73c4w1qNRgi
LsIUW1h/u+Sk6E3Fickjga09KKWzmFbF7698KudOpOMhGAELTRXAIhEgvSibEoSX
FBT4DZb+KaEx41XuZ2a8YtQ0mwY5CBAcoB8EDE4c9+5gkbQ3DKYQljOmhkHIUJlb
gWIOftaL3OvJxTeF7dsDOpWXPWi++HAttqcKP1mf6yx4rTYWX7qhuAzPBTrAs6ml
ROo0KTSuUS2WoW37DJ1y0VcZgfa0qAGODWzL+uMiEknqpiwP/ileszidNIlnrUIO
I99uOlxLaQjoxl3upOxlN1npTkjEYuKx7Q6s9COZWvQ/qDVZmG7L+ajw1SK2+XX3
MNAWuta0E5y0GG/NJ6V5Mrg8+MFrBadb2pLRUVXqKReZsk8ij1mCqups+QnmOViz
JfwD8oxhBEq/m6+OCUQzgmPFUm5U8EPrh3q5rYksPUyYMFq7P8mmtogx8I9wcEy6
Ndih/Ilp8ZvJMD7zcocu4L80IeePW2rAj6cP/SSFAIOmUceBb3p7MySQ0xBip/VQ
Bs+SU4/yi8b8pO1Ge/CPvbuy359RDpnnHuh6Er30aUY6EymhVZ2Aqc/2bLrbDMM4
xkV+VZ0QzJ+Smhhaj1xMkeG9cUAGZm/FOnbUiMq9ri16g0feUvOEakH4cTLx4NAY
uXvBYnaRra4sBqolHBdzO+pZ7CT2U4Apx5ykc8xf6S4uJv4g/ctvH9qKNThPVlln
bGPqHb5KuU/kjcnsKLvBLnXBcFFn297QKTk5UVj1DwI1chKzCFLRNX+Rfk9uPzW2
RDlilFXqO+UuHhI2WDQqCSsnvL4D8hseOuGMBaiQh3R/trMxHHYwBBw2VqrOlW8y
iZIsqmlB08r1CsXSdoQxTBh6vQKxhdcBTD5ZHYVd7ROlDT46AtJNfPK5TLLjKzK4
20bZLDKMKB01Lb6i6eAfLHK5fMjiopfAh7hm8Xb8EEwFc5y3HxZ2QWXWS5laI0Mg
sipmCQg2jIgFmHatJD3DGs7svKIuwpEHspGvYMOHxcGRkBJtCKVkFnTeeZ9WPqGi
O9z3DpNPPX6zT+GL/md9SX3cPpL2QacytIFyujMDwxP0oivMkB33ReLOrMQ+q4iO
JFAlZDqM+bIUqsje/p3kKJV6Uh2DbUrdwgO6uOqScXGxsrw911wrmZAoAiCf9lSN
cqLsFS47nqdvajJOjo5QzZ4Var9pISit/UuvK6Eq1hXwfAWGTTNJOZOvSVYj9ZTB
mIZ7G33V0/ONqL1CHd3d835VLO0vVrnkmqkOuY0UDNQXPsVjebpujM+gRQakXujF
1tORIBkqKHEFeTtQimvj4i5j+h804i4fZjrH0qAoouhldoLw3gd+I6SIDXAsuOn4
LgKyDMJIMDPer+J7oMq32K+ApUtQwbijkNSJLg7+Rl+GmIk1O5S5BtHiOTQ6/0Az
yEZRCnsnxE1i+oNybi77/RfNJKqyJAGX4F9DKeamdkkdJbNoaBWm1eR9dGCRcRa7
eHxCJ4lRU8tfQW2Vvqe80LSTD8ZARqSgMWNJXz1oJjkP8DgSKesdmhksS4TN7ku4
W97+g+45FzkyKhkDsEB2XVh0MKK6498t0S2AwLgbfCCp5iH1Etgw1USBvupaRfUw
S4QFDxnW00ftCwFrgK6BNUrikqx5FYmT5oUMWUX0Ct9BxN1oRpm21hAxECZj3HkJ
kd0gCRDE2C1rvJWvhL8jx7alNMFlERlwJwwXEDW6P9yFUQ+OZley/6iOvl1qHQt8
rB3GToZ8bzZ2bTiPC1dQxP0sM8KIUFC7maClgRbPfjQcHGQ/46uKt2bBknywt6YQ
1QE90GAQTLXB70ozN3GE/rK/HjpDPA4KF1GU8c3ioZO78//OKQlP61hmX24DEu85
Ugmm0MlAllpt2oe+040hPKliqPhctiFQehmfwgGDJMeUqF6lbx5ZzCKQdCRu7ucj
yY+j+THCLDemgKeVOgHfnlnstLoJRaFA4gZmQeGojYGpqYG3cEjIlW61D3/xXrpF
ghE1q83Lasa0oUBZ8wnUjRMxlJc0+YwESqqI3psYqFbYVSsp6cfDmWJOCmkGCw4U
C7MhAUi0jGjGcclUxDSM+tgZAYyrrR/L3W1ntvAO6rA6SXnyDx0760Qbfeq0jrtI
G0dWnfZyOtO8zEKP5ofjO//TAOjluLF4He8b3Vk95FZDdRTpLDykij/DqS8i3W9I
yNlitmGo5e+73f6wn1EpI7obOgRHHKJ8IcF4UzbK0q0nBjGslWXU104ehwlsJU6H
C5XhCNlRcuwCmud97OMI2CCIUylLK3JSR+pjgJxnS4Axkm7e6+7iJRinBjCsUkMr
oV3y3lvHnIY+4eAQUWmNcjY+oWKiZX6u3EvovAcI8rrDnlTxvzOW7eOh6rzUdsMv
d0YC4nCr8l2e4totH6za347gFPLNgptqWwMkf5M4zJTKBEAW2scAI0BupxCIJgUJ
avdWoVIbj6S2i7l2gzEl1H+JtujNL+IS0kFTSBzqgTOrtCeiTHnVFwqc8KmpZYA/
soEP84fD8/Aji9nMuv0omqqFlIM3SjiwP7asGV3MHhxDOP8SDsqRLGUOZ8D3AU7J
1EqKqfKWfdXexPbZNHCg1k2lPRFCpBe/djJencD287r6zFRu0g/rMW8zHVdIiV0V
CscOMvDCU1VGHOHRMJVeN09VjjJv3hYyr+vD5QXFkTRamxeLJT/R8kzMsEYQwLuc
CdMPAmKEOf6r7fhkekebsew+zkVWfnRVWztcXNlUqJDFoulfPzJnqvp/eK/8NNNz
FQu6+hNrOLzycP3v86ajA8xqQpeXdnpLrUiJ3iyTaeJiOns21y7z8BcPdK8wlKPN
slC9484sd1kq0J0eabc3nUnZ0BQRL3VtNaX438u+VT0zKJSUf87iKyza00FdRNIf
tT04kjMsl1KbhlRPOBfYruoenKPSkiLBbRrtvm5/KS5nVWlxT76OsUo+P+dUdrqw
JQZdAGAwZc+AbdWeGjHSI2JkYQqc7YvhZCxMXehhk1U7HBs/iv+0Ss35n5rDLvwl
kEF2+VbL7huNSUM6bBVGJfR4uXPU+/VNolsqIfTfOGaLrJz5ErLnaDIzjyhlpMyk
krmzntCSZvn87x/XCfVXNRRU2l1h2oeFGsu6+MbErk9BpsRALwVXWzi0Zsl5oet1
CtORdRcVIFgKkcbyJQVoVsCOYzHyXQ4UuDsQjapHD8ejTZdzcON8NRiaY12HpMWI
DrZrkzbVV1lMrdryOVZFcC/wpsrLlHHapAg8VN8VQhlB0rMeAXhXshxv2630zPxw
Jg9mmzmV2kvI8oXHnADCZnDcvBTd8CF8hJeG0IDL3skpoGt6QUYbSDGiuAeKPrWq
yvxZxFIGZNpSiKtY502lWToXJ3W6ry4y5jGq4uM9ieeA01OJRCHLyaXtb4RULgai
2jeg86rs+84DU6w0zBMCn8CLLEnxySe/2LdcA8QLyqSIwB5035XzB6PpFrnPddJZ
vpBrN/pBP2LF+CGzlnnlmjwxRgRl2IkaSwKu7H5jRQz+iuMRt5GQlcfu1Db+UaZm
R5CbsZMsNDVOA5Co/2wXXOauPEgBv03IPOtKM6tg2gPBealB7bulIB0a30ekqd9C
ePoM83HmTBTRrBjnszAU8kFSxxs7suyB8vMlquL0ZUGzYHKZyBuEVeVTOBg7dvlM
aOQE8IcirxUrVcn8VZ8eWwP/O1ohml/IeNZbpCWo1FwbbiPaUtjMtTFDAMSjaTWN
idBTtANKmGTikZus6IVvIEF5DszWSOBOmyi6c+aFVqQXBVd51zAphszJlyQjwrAn
vv6E0Pcj0lIef548hFaj9XVzgfLxFi6F4jK6buOaA9ICjFEPTeFtA1lGZtgbx54Z
GNX1XFqTP+T/mjiGeMzhX8vcZCoxEv2ov+6sZuH3xFeD6pWllR4qxV/adRG06US8
0LwH8IYed07xo7V3i/RE9xjwbRuFdCBm3booL9+T0+Jv5V52yC8FJTrgmFyR6AbJ
YSwQryg5Mc3xOPnMmjhKucq3jmmiYMvJmmIkEhsU0WANZcos6G1LKx8kXYw/ckmf
kliogtOi32Hfq49sG2/iVBDZWrQVsv5PwvZSBiGpj9xCv/tVo3EiQxAEGa1Chakn
McsnuIRUGGixzc+Xa4VyCrqSc6h8DifzaC7zB/fFka9LzYjqAYm1/ANRfp3iDEU2
ht7Puna+m21a2V2lgC6cublNH113cf69UsOoof6ceSdqpaBfLHKx17dnflZ+3jx0
UgiKFCKOTAlAayl0MUK4mgRu+TqrJ8hLVoXsJXDgLJuAlS2ZbXh6FJbO8XdbJVCr
TsG7Q9Ld1lb1vfsNARwOqjsqGIv7UXK2IWh91yIGywFR21UQwc8+CsgATXcpAPUp
Afd/TSYbT20I1adL8w/z4Q0WciMdpASeS4yx0puPJO1hepl0+KCKMzhLJkhMj+sa
RuNTj3NoBFgFwjXb/7yoWbYaG8K8E/IYs4/azHm9FFf1XLxqxnZBrtoY10Sahgyo
W/LbHizDvgCUikGbwE9kiFmjfEwOSHdKwNVBSyabbdbT1Qw9r4oXZDuqQA7KXpql
EszdfLjpGGmRZE4qjrn0t7lP10vvY+HKrivDjxEUTla9LJGxBrZohlN0sNqlUPgV
yaTR+Lx9ZmjybRtw8ex+BTyPqoYUjVXAdh6ssedVYgPnc2XX6RMmw0GxG6aXYjbD
qxPexIwUTUOVEdWjhQhkvF7/GvTtjl0TG90i1bPdbNv9cT0A5+Kfiwxa9sA2xCKg
fHtWam1iZSJaHvulRIfd97BWjgE/6tCyqRWg6C4LDoqP6TDJViuDvb4+WpEdRno9
7PanTugRdfGIsMhVT2pDMrDuD7wE6YumhGyARtFZZpNkDn75Spvtdp7dhGb1rTUi
zrBNnLseohZUtD6BlCW2RTAUPeoXxl451FKeujfOZ2lSR8swLA8cWjiz1V3cz50G
ncmFeqb98vzgkssTviJMI4MM0qeDHglK4DySrY82rZ6fCWIPq/5k76l4sTuUmQvS
5KicpVWYsnjh2ByxMJm60P4t/BZfOzxfO+QRWyi1FGr9Jbm7+plxwcF7NFim54qv
xbOEd2uchxpxeaqFySbRtGQB/REs9rRh4zfAw+c/sPL7CqYCAK6vu/7kXaPadcps
UzkrbVP32xIP8q/jWgsxFHS2Geo/NoMeV0+nHik5XJ2YfHjS7TD9Gt9pPt3T1JGj
hE26ttIGNKy24mvR5rrZevMF5J4r0P2VgVjigTAswSl+W3L9y7G8cGR0FsiS859X
mm7MFM62ItpvJ34kG6EKzDh+d+utxuidOq2ycxxirybIxWSnG7jzyjFYt1IHjv9U
8A6sOoXTLGAZKDNz8MG8ZT65PY0SAv+9OtgOa9h42+xKrMXhRNjhOuB2UY1WMxSO
HBDSgWKbNEc8w13UUUOlZD2Qy8HRypLp0UzKt02Y1jsTHo/XTn0Y0PfPo+3h7Cx4
CJHRiweYINlCmewepYX0Ca3SYFC06e8QcmXHTST2OPElFJManMdK2ssTXevcyxVy
AyDl+ve2owank6deOvE7kkesd+e6zbGO86MXkBfHBcx9UymKrm2TqlQsBEeRjEhV
J+/WYPWTGTM3RwKsLQnXooEtvJ4CsnN5tiZpYHoYfvKwyWgDjCUgDI7hb/kGI/dZ
lav7iqYOFpL4nbPVYme+tsfPTz0Fjjhdsax/G4dYOT/JJL/XSF/uN1lzRaC89M15
Ku3Z35YmlwZIJu7Pz4rzLif09mCudc4hNy2arlgpntX1gFWXIUohgWKjqjHLlWEp
gJwdjlSZEzRFpYdlwg4AYp8ckiWYQxG+7n2PLPaBgQh/lpEKYkBz9uhCPnTS9a39
KZGqlONj1K+TjhVK2llj5lQiP9MWJ8iJFEcT09gPYABWAtWnpAof84aQh4jVeFFI
LYZs2F5TKAV0imoNfTe3mveNAGZqRFwLHAFkSEHNclS2OxOCZjpYsML62uXlXHOO
wM1Al1wH8Pc5AseF6WZX85fXlfqOQTH654ko2TdJbdMW2seDwsk8wiSLPo8iOHZQ
25ETYkEKsSccdGFsMIsPIGdAkcwEwaP1ORBlmLdIwYvq5/W4jcdg0SQkqjvm8DdR
AnLi0HncuG37VS9CfGov3GmOpJfuT5jVzhfC7Z+q8UzwFrei5L1lr2VQe5Dh13YG
/Mn9G+nE/1CJMMplviaJQ5ndZzAO7rawNt0jBO3LQ3+x9MGZ4DNXInIPavHsSRDl
sUO1IPb012Xs/CaSe8Nala+wo7gILHGaUpGyI/qSI5RJwIHbXSuGXi0bg8Xacp64
ZZIVPfdnLKCkGrt2FZSnttTFLYbT9dnA69A49zH8c5b/5NLDtAuiFYO1DZ4knICJ
XK+QnFGd7svCKxDD1lcIFKMa8GuoXaW4mGFI409OHSZosKRGcW8MTZ7jF5WBwvyL
pE+RWYASj0Qmna5Mv6tZzT9z1EECMKePiofeNj+3qCDbYiq4BZETydwfrt0+CY6v
CSuswVwUxsOurIcM685SZ5OWR42cg0BuoQLd6HLkvr7BZ8Lxgk6hqxm0R1/ggLE+
7bWDDc9jPe1q57BjDkTAO2TKYScTz+VuRnzfIwsNQv8rJWi3P72ReHNFu9aSdU3f
9y9hSSXUlrUsAuNcSgSzUOdKYu6Uq9g4ubgiVtN+YbVeFcblAi1F4iCoJKEzN6y0
FBpktNOrrjwIw66BGe9qhmXv977R1mOvCZaK0vJUQ1rTT8Fmvl/gm9qe8viOzuyu
mi2vN2R/jo7itzw3F/g6Ohk0/7Op4IsdXJgqqVD1N0UbdI2ZUPbICrHsB0GTFKxg
Kghbqw76KQuhi2O5eZKbrvk8YkYhIAOkeJKA7vbns67ml+3IkKjOVz9bajXYhQ9j
XhhVs0SQmCga3ixsiUs3KcgglaTBwoHHH+y+PGWs+DmKClJBaocXTscbI3mU5k8x
b0CDCfJH9QB616Pml9yVGiSx6zBoPd9XOkygEeu4VteI1y86wpugPO0RPHESwUFw
DBd+WMe9Wx1hcVKqWz8OPlzmhA5Z2KIKYB8OpEO2y/O6olbyAQz1hSdlNEi/UjLr
zBaRJsJYjfox98BfE5YDxCxYYQTa7UqOkwqWCAJCwewtcwEjKGHFKGLroqrMKsKU
p7ln2q82f5IZOJ4Y74Mj+5DfX2dnRX2R4MqYwCIItODJiF0mzOH2KYhEBD6jldDL
OXtsUFj41Vw2ySGC6TPwmDvB3EESmS4jf31etn2mrw49FYd0cOexeBLnKN5QijxL
LSSoRTj3Pgc8pms5c5glBhrF2WsD5ZYzhgljr2B/Ty6mQY7+6eZGIg+HJVgj4H36
xElBoCCZfr0EZCYoRx73I3+g2uC3Vp5WhLePZfx6BM/t4o3MUuqyTrbnYr1WMqbi
7Yp210Zne5a2J1CPOrmc07E+Ucpri1vUVs3qguWvy1iWR0c8avv/p30BX1zB1k1H
zt3d5UA3gQjhj5f9yrZ4n0JSRslLeAYBB/66xLHcn8/6ZIc0D05dIa0J298H4XYt
U9BR0yrQOeglIhTeVCXK4nloV+tYz3ioPswcVasx8kq72EYWVZaXSzC0P5eqmmba
ZkH7LPec4tedrKyXfjVEkb0cY0qnDf8a34BT0qVexOyeXDLfVuf2KfvrrWSG+OBA
5YTALGSzGB2TknFcWLY3m9iLpZHHvRBxuF+JO1EArbNga2ZRxERhRJGOTIHO7JiJ
bkAEEvVfY2MC5KAvkCRFVjI4pOD5/UKJiVR9yZ54J9iNJG0cS0vnSTBl8sUqD1tg
tX//BxwADrfVua90oltoBVow5yYpVal5qDW+fNmnxc0ztoyarO4thRvhsJvCMCoY
Z9PhA1CsPU+X0mJbQ7VgvsZxV418Ynkcs96PQ0zEWCn8PzruxGHwiL0uSwAqjgqh
ZevNZnbZYiOKYEoIvx7nA5IcXjkIM2PBEThrob2zwP+aZDsTox0GpOiyV6uoXSWs
XvEZ4GFuN9wp6iR218HPQzD6sciKrEi1qvKrNiBZ6Gf/uGKf258XU3DyM1sCxMXY
JeS69WSV+eR/zZ7cU67ih+UT7kP8BPzGl2Azb/fpSrg8aBYR7HhDRGlLnLK2Ombp
f4MOlxnmVsOQ+2/9bbaZwO50tv9emY256wogA5coGxYZQ7vC2V4SBYCgZ7gyP9d+
dOohAN1bxj8sEybUB+7Jfl8VVgaJkcJ1VMHFyD/yzbvj/oD3aQ108ieakDr8vN6U
04H80ntT+mGy18KUcWLM+ugKYp7ATmYALsf7iYLiF2wAZT07oFgDIay8tioFTKft
BDiSAFcPwQJYoIhEdHGnbfyD4LirA2KYwDw1L8XTMluSE5/zpMX9430Hd7KT0u0B
oRKqtvsHxv1l4rsSImEKQ+vOcqONjP9kvlAjjNuNFu3VA9NbYx3x+G+jJT2dGDKk
xMyRaJqBzBar6cTi6HDub0FxNVhwUjd9Bddx/u7QLRIDWl9SkN/7WHVkgdj9OsLI
UI1OWAWOU6OBPV9Szp6B/5biLLefN3Zjv2fdnDKMT2EcgRYQYH4W0gdVNhnPZVNC
eOpjoo477dP4l6nF5ol5MDdVPRp7zP2Ou+WTV8hj8QQsIewuTgQUqj1rIZIkGsC/
rYpctACRHeBN1UVl/PfOfcCxGg7+4mmTcb2+a+4XkEjx4CNA+0jiK7JLQX2T9Ybz
ftxAJV4mRquCloWFi9sGldUqgijrGiuHJMhw7Z9wyXSBDLSA4kE5v8kFqLpo9ITK
74ivrB/9HEtJALbFc/sc2b8rkMBWPtcYBHPCTXV27uOiqwqh/6K/EptWLYkGGj2u
b9JyxPYcwoLxrPwZW2RaQZyBXvgqW3VJ7alEVonM3VoprJQvOrrc9rOO7LaIbCYE
/o5LOaNUzybwUh442CvsNaLVZTPvsYtR7KToU+uUvAridt0bznuNpkmsRNn5m7aK
Xzd97ivjvLIR5mQQ3ZzKplc7hs5v4pPzHsWsaH2dZ0vStIfueOYITXRzjsF3kHCD
xJ281lABhh+R7OGGkQ939qwdNe2oepjahAiIlX+Z3PnrW1pOcKAs1NZKICJdgMfl
6DDVwYMmzQ63pDfc3VtiEjTSIcRKIvAE1b0HhApnmJgEZSZqm6Hko1BFOZHPLSYL
fKNHCNdY6yvHuy55JFEOpCFf6gP/Ov4vj1BcB4pD5FMNZ0PRgRZLFr9wbxrrGEr1
ePWXsapg+dO7/IbJ5GfsiOaDy/lCiBoCqNItL36/To3IMNObGSt6s4gsUe/XiYXv
of8ECNS2oFeTEK6VeEFcZY375MbDRS5sCrXKNGHXHalVHwP1sLLogq+URt07SZgv
3dMJPXf3hhKNUQOwpqLwakEm6+LEC4/sM116e5dZHIyZC6YaMbCxjBZ4xX4Acrgt
2v/QFZzhQEcNZVPhaaSKF3OS8czC996hqdDwTNFzp1KICzHrPd6P6LJGN/tZTp3g
HdeevRUEQeWwHsA4vQMHJWXPkQVkNoJMtynZ+AmzMBonQ9r4PiB3w+1M88nQBZhX
tGkWOgGXqe56X+PyIzqB2ItvgETB0hTr3dGvet+ybIxwlL1Sg9biCPWDNsRKDRln
FDfbDxFUiVGz8+CESKnmuhJuSosjyU+My2SsYtrN2fU9+KA8FZvzNRUcFBrzWxzj
vj55cgR0pK1QMO8JC2QsjyK+KjXAtvGqg+ya5xGO7IoVQlUt/p2xRalYCLW2NjVS
w7zdU1MyMstKnJREfo3SGKQQVvqyGlaD3+Hh/09XNF1gl9zKxEQxr7BfaYWSI57m
1J/+iP5OiWkqo+863xJa2powatAijWJp4T//2N7pL70+I7YGhop6Q/6nUw6lU2Sf
aDTAHTYDerIB/l3K0yLTu7TprCJS5By/J35NtEvfILXQZvBD0HbTXYjAg1x/3b2N
dYLdslsnjh/mztoDZ0s+aYqG7E/wuUIuZNUwSuTxODq/drcBC3PMezVRMZ7NjSz/
qBAwOMn+mGkXDZJLPsP3eSWoi0j4MWNV7XKkBGtq5OfiHGE9wTJ/uvz43eNcl1zO
muAMQrFWbFHTZnMovb7xG7mMOG11PnHSzc3FzEfsFQYLIn7ZgeSEsyEKCZIQTSq1
ruHvHA0QL8GUzm8RrY2975ibxVfK1df00i0293wSrB/3LuArgjFmIA6IfiMDTlEt
YswOcMouTpcQcjvMDpp7uJScAejBR6FXCEwhRosJQZ2L45+nJUsyCbTtaLIta2/m
ViKmuOzejic5fJfVUFdP8qgb8/mZaWJeLyQSHpO9cQZtGWPy7cx+Vo10mBQIoKl4
7d4J83T7lsWSYRcAKAwaShG8KqRkFqp1+A8nF+Oxp4uLWPf5z522htsZ+we86Cab
lNCTe1OHEyGX0EvyCGjajCSQWEh6e1azkDtQNqnVdQePyUdS/Bb+AAv6VJ8JgSGy
5g/CwY4XvJ4yF22xtOsdfB0/wQkAJmf49vX4YPVkJaXOfLIbHHMAgRXYzECGWWRM
nO54lkiOQize3/a/3WBvoSpzaPtq+XqpBNR/3iqzuQDEMXsYqBi3zIHq0j8ZMYRh
TzbkaFqUHjOnyPCEzIEKtY/cwGfe86S06zVFA+ZEZoZBC4NgRTBl01x/yRxREJ6S
V2xr+g0TfPSju1C8tvGKRMfEDdxhNA9QgoKLv13bTFHOhdZI5rO0GTbQDQzCaSWi
0QTW90EbVAeneUPXIAVnNzKXeB1EYuJNFMCXU5Ng9Wi1wn7jvFFw6omxe0IPC44+
TsVGVCMDOduV3xhKdQjXDAUYlO3Zi9bSf0XxS7xYhsRnZZm9FMVW0WE554ewxuHg
BGUd1g8hy43lkZNdELyfqBb3a4KVUOrUgrYjlIEsM3iIKrF1bYyVBst0qkcMd3cP
WH2tWT/a84yu+ymAf4z+HhqUvvWfAqr8yuNqB6ud45mm3G1yxs2uxDpcwzkTvlF2
R84eQJDUmCP4sYSlm8ChuawE+DNnclR7OiWY748MfvUhhnWEVKSRhlTcrvWAwZy5
6+lSuQaKe9IcuCIzZM7nGQk/9Bu/MiJBy2QFc8YaqCyOQr/3ByeQH2D6LI9oLL75
aF6j4u8ofVXY5lcYsoNLweGYT0+CJXmMURHmh0rokfuLFOC7rwaDaPv+jsirNjsU
N630/DC7Tjm9MGTyVy6e4rqJIpTAnl6/yL7F6KRZKBwW0Vknor3gF8vQ7Mgo3iYo
Iir9sdvpvkgrueuu+elrHMis+yT8VbuG71wJMgL1hmxLUkWzoy0hDDWn/Ca8dqko
dmzK4fumplceRAKGo450F69KaSTqfNq8mwlltd2ch6WS7/Pf7jAi5THeGQYUG/eX
Xkr7TOjjqGe90orlz7UX/0OtUJyZdephMvUg8Yp671yVEtupYzRJbvoEzUXDH7Rq
hrGxyCSXIObrtrtzYRH+H0PDHtnBw372UloaOs9svKsGjqW9AznhbzmwcQHC3XmH
JVnuGC3SXaBMoOrbXdNXBQS4k60klMJrlvWX/WWIXjz7Ha1XpMite9Tuc4yMRA4q
Yy0wFpPvYaGAtypT/NT49ukBWsK6FAByQHmaaaJ07MCz9yjjYQYHbDAotedNIG+u
PGmifXFfq9lAlbgPW4CQM6kn6qBGhrPH3Sr3y8loKQ2XNK5ytSbWIOvMC6W4J/9u
BiSD6Qfdu/F68/R6pzc5UW9NNNw8YIEOftXhWMZx640Yc0cYKFEOYdUndBrS2r2J
30ELLiogFIaajN2Tcih59upR0VxBwRp6CzVGAPYBHb+thalKdgMycvjieSp7WKzx
XXUlYx1WIruViZgv6SYmEZnzszGOJPZ0KydXfExRTtIND6pe1tV0Rlrd+kuURMQw
eg5rirhNgpWfcm5cMkhOYw==
`protect end_protected