`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
ddtXksX2+yylW5zu6QL2Lhnb2d1sD00763mmSITNX595NcHTEkwn0zB1Dry37fOW
FufOhVzEJp80NC5qZ/+F0Vk7Ik02dIR0elf3clrjeJRK85K4e3Hoo4xn7YbFUIms
l/8VZSb14+JVGURjfswrIyCUotIzlzVYZ6gzoZwDXIi5gQIBf/gI+KxNXPaKV+PQ
Ufys/12rjO6aI/pPlqSm0hCvftmBcnezN2hk1UeXgOIuKZnogjOsf0iJVX2aOOWE
6pD/psybjbnsNB6kH5uFTA5frkzIzkzl5d9+YDm9OyC+k84E83I/7/j+rk4L2dah
QJOvksSIzN867/4Qt8qYTQ==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="MvBXkzurAa5VTw+1JJ70nePUfoQXBvZOku/SMmg4TwQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
oRtzZL4VJ4iwysPsC8SXYCzXS8Fw2gtZTOskLcDV+1B9Nzn1zTyNtlo6lNICRmmK
ZRVu2BmCc2G+fmzynYlNTnSa7C0Cuel6FYpxCBlOuk3OF2tzAmLAuDyOH3Z1Yjzk
a0aHuoCdIRKv7BrZCdALt03JeUmXKPdOmIlkVGFl8yw=
`protect rights_digest_method = "sha256"
`protect end_toolblock="Jn9CQpRhJt4rnzZPRk+dOpzAubz7omckX1MrFd4p81o="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 2384 )
`protect data_block
gD6l00tciPUa6pDNTk/+tzLxvdHE2s3DQL3/JqqujQBC/Ei+vcAB8wM3doqg5vTg
mdfn9XB1bLOis2CVSfu295W2DNwHfMSTc/8BhCDRnTlLIX0UCJs9Za0+LoM0rMrV
T7EjVWppbP+Em6PkVKCwlmIQ7JKaifJ+Y+kjw9HCGboYo5074hY+K/CBbfsBQY86
NbkSLCO87IQEY+0Q2aP6txsmfd8pwVyLY0eKa12DqN3xoCerl/S909wxQ+kEbtEu
5aQJCWEtC9Lhuu4IFlwZwt+p8ooRUmuvRtH5BV9zjAp/iLVsi9JJOBGBCHCQymYE
biS+NPK5AVf1bkeALjR9d29VNav//xGssAALVDwf02ygOHCpYz5/cwJQEbjlKJmG
+PoUJrHSl4mZnS+n7VvjFRnXmxR6jz3FNrmOaXn+rs8Bnr1oFi+X0LEawbFwITne
5OxWgz+eoAzVqiEwQ5Nvx6jxD7/wj8WrhvR/hoOIth3eA6GHrjO2NID0JpTq3OqE
C3jt6Zrgapr0LQ2FtTevcunhj1u1CWbAwk3ES/k7Y8stn0jM7O8AIXZdr63zJpA4
pNH8i5tDXv/9t9MQggo3IMaRD7NFh+jtuXUKtmPB0Y62gd9/VoZ40QFVPhfHXVtZ
VG7ZCir/mISP2D9wVOegY2yR4acKrbDnziYPzqfWPWNhRkgAOLNJID5yA+9DIKS+
1gSjlsc/uQmXl/gmWhSjOmlJWQrbpAepKBTBA3FDOsjC9kceIEwkwfoXnp81IXJN
8YqQEMuiMXc3PvETWedHdiDOwOqW2u4APUC71BE95XO7VuK+wToiQawjKRFp6sWR
fhU/USPkUkBsn3+o2bymKzlGe5129RgsIMMitZouka+7+r926VP/V0vrYegL2O/3
4zgjWzNkXTS1qvQD9umxhzBqcRzQCAGc67MWF1x6yImEJZxk5gtDk0mr+09qbUJv
KZzNyIbgLiBi98gRqOIsQG90lNDbrw4ZAGMRgTZR/lAOevktQPp9lpEJ7PDa/e+I
BJAfHLIP7vxXOsUvMMEXepjzAunnmS032+bvmDRMS+4zldHB3+6EsTJN9dDUgbkH
gAwMYFWptfTliSVfTpsxXKqqVaPqNx5Bzu5pnKNsh+xyp01MjRvXx0gcBeS/6w7X
sSzEv0IqGSd0oUkaPvxSBN2UnLebJUXVEsU4vsb/iQGVeBnO0/XnGY2bqszPYKtN
zZd6P8AwuwPdfD+ZVap5C32RZfb2DqVqkzx0CnXm4e6w/zDU14KuB5KvkniUwIPo
s6d0R3YSJ4RPfewNl6im/eTImbgvdzkJSe/WVuuOc0PFq+W4Tz9JkOrnOQlaSEAq
zikwk6cPs9zgWmjFPRvGqQIxjHS7Az0nIc6Cd7PzSXFcYOuSzmFm9f2hsq/ttfZs
NssADxPyv8uiad8fvMcZ6an3IFTi7Hsg2yBurXccINOKol2ByqP+obhqTpvWybWr
IcRzqLRSolwnpj1QpNHYObg/3+FEL6aDFQlEKKflVDPQtDYBSOsUS6ssqqNAEEqZ
CXMHMUUqfbOtGmn6xdnifINzALdTJPmfGQPm7MJhlXd1HCnPkagEoZ5cld3oJqWd
B62ZD0HI+5BZu1JGQsvSFl6BnOwUU3Ad9oYZNr5sVN7fsgZQcFIFEbgk2P2eB5R4
sfMlcm/jRnzHnvmi/q2gYtpuNiL92pShReL6GYRWOegZ3o6fbujJmlkLuzmFVJl2
8d/rcgG/0sh50yb7Oo8mDo8jPzdzLV+zb5hM8awVkcKmKeStJST52rmOKGnInt9a
hzAVQUYbJZRXyREsqQdP9TxEXJlcXnNxrl7PoF2HNmiigzESkI3+lx8VqIDjD6aC
k2o6qBkqW/SCBU2HIkWrLonIDcKzONGKQOpo03/nhP2sk2vN7KG7lpntZkMhFdEE
cB/aw7OTE7tnSabeWYhtXi/XphtcS/1Khb0kn76zhzSx5w5nbD5db9cgzrMweX/b
cf8rFdBJFqU+jJkUJttq31VHBMHYaeHg+zIsweQzI6ZHKYlFfHhX35ywHQq+Qa8t
S+lbKgSELo2fKW+3OoejGkK0FLpDnuhm6/y0pOEdP7AAbfs3z9pirOx9lySeIOg7
2IOfFrQMS6Rkwm/khCxc6NLEc9bVDf9tnKcM0xJ0RWa3s6wlc3zTxUGHWInzcRgZ
RTPJRq3v+Y2wbgUQUEahl7qRISme50/RnwPUMPv9oEMp/bWGZkcXHiWRI/YuvJY7
EQn/kq6wi20BaGBX6n6F0h/+uNib2p8l5SqbhD02v+PdXheg6cblGaFID01kRWfn
16aJqFjdkQ1hKhaY2vBS5Q68gsLmi5b9V5zv8ri+0CGR0+CVDWNw3TkgxA1scik2
uwd/YAFJJQ2gXXa1D3gouwejmZbQewOdHcRCpvaG5C4aK54aVyUxvTKjfsT8giQ2
uWxW4zq8WpXz9B99GMzGlAX2I8vaoXxwTljikxK/oj/xbX74v9axbZ/lpnm2OnOf
CXVzpAK2R+SGuLsB4eXRwlgDY219blAFRraT7f2X9ehMHL5lVTiZmgHxUg9PHl4a
kblli5rO0CpUoxl74FP0D4uWnzoBPyL6WeFA3VjGJtymdUxEg9yg0QrfRzTQM0LL
JFaHAojXa1qq2AvUBT+n5Ej7Rt4QjTl+d0cGF9e9dPBitS/nhxpzRTe8c8NVzKFH
qm6kiOso95e6lMbUKFKvB6cpwUk+lEgzrw6TTAqA5ijikSIjnZhzlRg1uAstxTjp
Bw5t12hw4IOczo75XUAfdyn6AgWEqlC/9ERlRUU+/MZ7ak4+LhlySH0rkBmnYs7m
Umjq6DY63yWFYQq2k6I/veVoxU31nF45UdgQp1XPcUvyd89BYrfZYkN8vc9J8FpW
EteGVniEkgv5Lcad+HhXxdMEYTIfXwqTDHeA0ckUl+IiCSGT6WL1RcQiUkFtT9he
n1sLkKjWGDUXPk17KNI5G6L/sVZVog0Ch8NeVNvajsQaY4S6FWMa0SpnigH7Da65
LUlDBG9t7imy16YMZ6btfuDxsF8a08uNSUPC5I8wOEhBeJ+0QMcG7d2rO2UIZcTQ
5kMThoygcvGXgHHOlGCVMiDOL3vQQiOwKh8tZqOgqXVWB10ikiDGwxUB6Ic29tMP
si3F+TT/a8nkiJhTif8jxIDTta//o6xJeGWsctzHcKU=
`protect end_protected