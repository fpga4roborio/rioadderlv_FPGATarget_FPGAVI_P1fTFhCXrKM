`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
ddtXksX2+yylW5zu6QL2Lhnb2d1sD00763mmSITNX595NcHTEkwn0zB1Dry37fOW
FufOhVzEJp80NC5qZ/+F0Vk7Ik02dIR0elf3clrjeJRK85K4e3Hoo4xn7YbFUIms
l/8VZSb14+JVGURjfswrIyCUotIzlzVYZ6gzoZwDXIi5gQIBf/gI+KxNXPaKV+PQ
Ufys/12rjO6aI/pPlqSm0hCvftmBcnezN2hk1UeXgOIuKZnogjOsf0iJVX2aOOWE
6pD/psybjbnsNB6kH5uFTA5frkzIzkzl5d9+YDm9OyC+k84E83I/7/j+rk4L2dah
QJOvksSIzN867/4Qt8qYTQ==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="MvBXkzurAa5VTw+1JJ70nePUfoQXBvZOku/SMmg4TwQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
oRtzZL4VJ4iwysPsC8SXYCzXS8Fw2gtZTOskLcDV+1B9Nzn1zTyNtlo6lNICRmmK
ZRVu2BmCc2G+fmzynYlNTnSa7C0Cuel6FYpxCBlOuk3OF2tzAmLAuDyOH3Z1Yjzk
a0aHuoCdIRKv7BrZCdALt03JeUmXKPdOmIlkVGFl8yw=
`protect rights_digest_method = "sha256"
`protect end_toolblock="Jn9CQpRhJt4rnzZPRk+dOpzAubz7omckX1MrFd4p81o="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 6368 )
`protect data_block
gD6l00tciPUa6pDNTk/+tzLxvdHE2s3DQL3/JqqujQBC/Ei+vcAB8wM3doqg5vTg
mdfn9XB1bLOis2CVSfu295W2DNwHfMSTc/8BhCDRnTlLIX0UCJs9Za0+LoM0rMrV
T7EjVWppbP+Em6PkVKCwlmIQ7JKaifJ+Y+kjw9HCGboYo5074hY+K/CBbfsBQY86
h7FrhVb0BFNFA4lVvsm6L3ECOjjyTeh9BGL3cwmrYlQz2NdS9LcgXLFQ71OcgR+E
V6lGQbXj8iuQ9cS1eZxbkLRZiWz/mgf68Q0trW+S2/vowRwMVHwrG4TmAEeQECrF
j2l56Tx7EchkQQ+dhX5KjAkWgwTIq0SuonGYrIB8zWJe97DcHmldofgudleMIBUD
HE7LCNlmSOGwJL95daq8FzrhyLcNN/xTkaykqdjYK+EgCkOm+VZTTzj2KUB/I3iC
iCdrfMEY1DXXk/joHeeF1sbBjL0Js5Z0JMWJw8kfvBUZ65t3wCbRULCXn/ppNnDA
FucpYvgkDyHRBbWGpX+qc+Af4+S0r0avOx8Zx5Wh53nUMwOzObfZFa5PZzCHNpH5
gJnFf6/lUNaiuFX5tQX2txhrl/jf3JCvwUprC87YCBzuAoPF01WhoyCBmhDEZjm1
JVXPUfR+HZNZOhhWjtjPN1znH99CIN6/iD4inp0a8lnZ31xOBEDVNy306UhxdeNa
04ivCqIugEJFcHnu/xBmvvzfTSJC8Hf/laa4VU7HMdBcMlaANYvTQ5LWo3iwZvua
8INdbXb1aqk/mu5I57WxDg+e8XVhY1bEBgqs/xAEaeBpEmCZTAoEXMuAr7/wpiTg
fgFVsb9FrjplqTSaKy7zP4dxxY/56U/c183KTvtgQDSfhrWk+65VylZ4Qefxak0N
b4AGTodTeEbOYzuVn+o8CyCGsxFdzXMQSWTvsgu8OYe8YE6FcD4vcf9U+ZFAOuTQ
dGxoKkzQ9FfhL7rBAcEldsiyh69EGHp42v/CsOafU+ezm9TJEV7gGykCnEMFqQJ9
OwbmbzYnHkCq+/pf6X7vm9B5pivLIlaeDpNa3VeC9RBmAFJyWlRn1aSlV93k8znf
FwiLPc931riyoOtn+w8lQfoPAwOaC6pTr3ELxS/Mt6YaKF31DxFbqPFu2GKNefWY
dqSO/kW1c+2LvinAsoo0Rm7Dt+e4yxT32xZSN7sQ4tEofwB56YLlNMvMzJlvl7+1
K4r3nPVIb9Cm8R0p0rLc0TMG4srmd1g8IO5rPtYb8dOnN97e5kOlg2hlhoGlpegA
87F+WoL0Tm9aI5123e03EOzJfebxKjxpcb+abwIgEt3xffvNHKA9HYr+Tfsn3J1R
bhAGPwAW0/8WiqTNlePGNhNsjXDnuwU38Jpl3z66mpEhFcpDtOhcsTlx78cPyfV3
KOTPwn7QJv8giEa0VeB+YYFClL5lTtsXooitD/zqfVXIywCBTsIrDrke6BTeDUi3
o2OR5CzuEu1NeVNYnOvsA2CJqW44cbNF7gmVkOcCQ7DQiI7EV8u9kAVIDtqoGZaW
WlqH09v3/+5Ef9kXlwB6uOnBIN9mO1Ekla9q0FzY2uKcWXAC4Hqvf/T/ztHMTjT3
D1mfXS2PA43z6O4BFuHNnKepF1WjKYq7kZt+nKoP7YtLoorZbTAINiM36SC/9lC5
Ea2DK3BtzdtnyEIrEsZhF43crIRvdH9sUye+QpKLRbL4DLRQzMT39BZpp28iKS3G
mW307OjleSZ0UWOLSN+fbJ3k+iEL/z/AQlvcW7TVVGixb/qXZVQnUQpIZyz56er1
m/1xLEl95b5OPTLPWr+W1jUIsExUOlmIp428quWIbxDWfcMR6/l6Upc+YLaNlqpE
UfiC5296lVs7MkgY7xAjEJ29+89d0rMtgpoAJ9SkFluNeMe4EcVj0tXj1R/BDr2L
K8TnDWGf6749tESxSu7aie5COrxMFg7jfAna0byEHwFrSilqEm/Un3Cq6Pf8VB6c
E1AyIml1yzSgkJ2JD45YC5NaPcmEZRZfqG4mI99T7oj545niEzVXbKsbLTGOPS3t
h66yKtIUL+185OlLYGNN3J9J+W6h0JjvqAZepsLYE5jAutUS7uDb5hg4FKExxbfb
pb4iAVcen+HedPhUK28+3UVZ7svUrwER8N/BeejokPg0oDoVby27mf8+y+0jzyDa
7628Wpkze59OnGnKoPDj9Zb3A1Kph8JPBDwIOGDjH0Wv8JAmdBjLM4OUBCgYAYOJ
DUICWL8zUuEALwVGSk+/Lq2biitpcjMW/9Bx33AQWzSH3/Fn86m9CX4X8EReGSj4
LlLUpx2JtYrgOe3Di9YDpA297d3Y7ooU//woWqMc/9VnbvwylB1q8UlDjKFtCCqA
q61X4tWarBZEMGuwQsjtkp8qbWWVgoynnTRxIXNVQXxNJUahJc2gitYjy/1Dzc5P
KiyM9HhQVOOhlIP5fgFlS+XvIb3iLUITW3xt4h7QhFXLLGyJubqUbR9GfmgPe5P2
AOxcsY45CLyD6i3w0HRT3/ZxC8a/e0jtMKqO9SWX7LEd7eQ0pfDKsCDMEY2uhrxi
Yd1sV3TFVbPTsb6+fFs6nZAGVBtMoD9nQCzHHPYgP+/wzNRGXtkgkMkibUfnA1ce
uUwlaqYwEYX/aOFwJJR8ZD4uSFzjOAfRh1sjNvL6rXOmHBxqw5TD09N1Nwu6d8OR
xZ9htB0Hqe4aB70HMIcvYg0IbJbO9giO4K+21JzIUFOHAgIESHbEAbAcSGK68bBT
pYnoJC6aDbUFE50WfvTSLj9bwc0KDTX++QRlF1tb+emRjM3ObAt13hr9asaBN2Yz
5Hqfn1zoLhPQWybC88VpXEzcmSl3+5AoZvo3HdO6PoLsD47h9Mi2pO0boJh31AB6
zZ6kEKhZxTpj6F1bGq0LRtCQLJu8SOGr3UkLXR8UeKDsY1wNskn0/dIMJq4kEdas
IgIpgYbFAr7PpVUdSO/YKSfpvUxiEsd691VPtFuL4l48aaIrlBegRg1MmsEuj344
5C8W2ulXVu147H36q/KEAWkAacz4Nh+w89nPViab4k8q3rQeKlD/z+XSDQxXmSoY
PRJU+o8Gg0s+kSGYV7tR+8mAh/aY6aPVwZOJqrWKdpo7z8d30xew0zvF3mANik4t
CjYJifJ7/XglLs7s60S7NTDBfjjHFotDMTReQidYzMFkVfhvUx/zy+AmpJiKPx4P
gtyYBoCvW+GejyGYWLaq+Mtk5PWWjC6IrR8/3vRbxKeoPLcpZGSC6NIy40yETGOh
/5uKqZGhz7BgbTZwIsl90Q49URLPqJ1VfqLOaJ8y9qsh1nakllE9u8ouFMLgVGRX
kP/ZwziFEmF5g4BWL0eY7zBW0RC+46mhwwwEIbpKLTJeL52QiGqY4THT1UxDgXC8
GIAHGhIjO88dvR7qJo6Yr9XVg2+syvjhSRKNFByE+ib3EOFADgfDV+tVJ7815FyQ
uypWQgmlRGdFf7O17d18HtFwB4Hh4iKnkj3+JCzvuro4P6drvrz4w1DYnv2ZW74w
HjNOrStZ3hJmvId4appYWtp2PudDklb+ELuWaIDWuL6Yptl/lyJyF3Lix1XiolvA
OU9biuNTuAnx9Aevpya7BEVwagu5Ubx+Cq36GyxRFzyK+YjiLoMJR+6Be1xz6CtZ
ymn02fOhJBdJmIGMIe34cP5o1NVXb4Tt7fcXr+rWkiRfegFJgDqKEzlFWxK7RNNo
++VUgcZlht4eRSTtqJctrtlTC/6/S6QmgqWWHaYP9vAjGFLvc8lc/i2PWVT/yJNZ
aXuYvPJk7k2IxReOVgPmZZdCkx/SOvZME++cchHqfWFb4YcCgeQKWrbqykFPVu/D
WI6389dSTMjy/k7k1ZuWF5K9A35cJ2aKqgf5CJUwdB0FXCM6fiVLylFE7dXUDC/B
VGGrW7hqFhrNc01OKX8mhxVIwOBEMeGVHru79Vj5p3IyxH2J7naD6AcH2pgK1kF9
jAOW7xfB2iU54iTvSaISSd23DKCpaHixFRHGJuu+9xju0cfPZ6gAggLa48DjnzM0
YDX/7p/v6PgV8WAt/xmhyJ3CYWOyyUDEANwYBrxgfUGz9IGtqAx4Db8SKJ4LLmmm
DQ+4wSIRzRf+VLR0FXR8xS5Mx9UpogWbDMnyNsUbfRsy9gDco3/CEvwdqq8GSeWZ
RwYLldIQCkc43tKE9CHn8ry+jwyh3M94BWMrLA41nVvI1cPRHOr3GJkZt5cmz7Hb
hQ8q0al/q2svsZCkNqCxcoGAhfc1VU0jbTy0Pbzbks2loADkbWm+WBrRyDXHrA6A
IHB3WuHdGac3+WMAy/rcoNbQb2Do3/o9zPCLvUrF7eNhEYv/ZKJ/0nqqBrPv3qWW
XmsU2vSUzWeJxGbEtqxmB1TodNjb/eoMj2jSMmgg+1Vz+8G9gxt7/69bhmTWcrwY
ZO+FeqjHowfPLBkuK+aXp+gfKqdgqUc0nk45BVd49ue0WsCZcGG3fZYTMY3Qzf4w
wXl16SurM3ZJDjaFWAW+CDWzUHq/I3BQVkf1XO++qG7RElrNgXLJJ6lSypskjYVb
mo2Kt+7m7GERpKof+VahYvmNm0O8aa6yDMIpaw6GN5zG0HyBshKt+nRlvoRqlbVT
pyWC9X0RXsBCPNLfFQQHOVMQ9JnFg/94soMGGIinpLh889Z4qEoHyAmUPiqzEGHa
9zos3M6uHP4HTeKCRlptHzIT8bZCy52xfwUvqRefgfctSKHzjcRRsi/rxYwLMQHw
7spPPqMH+vTg04bXjrSiKVGasvwlJiq9s8zWXWtG5pKAjyIj/FaijyWenwMh4mC5
qNYZhNjFpCkfFgrmz7ez9gmp6VWht4VPPGLVpaV0ZPVkHEPe7csGvC18qS6XIFMp
CntLHGCNDL1EGTxKwfBXVLmZ22iQYjdgJCoFFi5BePWXpOKGAk7kfRNdkJdT2DbB
wo+6WczgrW+8ehmenGgRXKYw/ML3+6M7k7ZUZxxgJTidzQeIfayjYjRlA9PDGR5L
/byWQptZV2gCUsZgfuLe4hA5S3M14JvahDE09LeBmY2+iSpu2wADZQS7LS7Xq+QK
ryaFP95v1c9U8DYoROJ8oNsg/wntDk+ooJ4/Kao0OYnmjBSvqHpW08kSLVOvlN7u
gZNSVYX+KG1yUwSFCcrzAtAeJWA35nrRS/BjgK1h+f/B0abQiTeZ9joV4Oag9GCO
SToBC8GFbifK3x8jqmFkua4LKU+yYuJHjLY2tolMAGIL7gf1lvsPFTwgSlZXFMg1
2f3oPhWGx4Mas8jaBMuE5H9yABYZXKjpYPiPLhPce4C4E1ffum59JH3cylaLGalp
YW4hwCdiPLNxUMCxTNiQo/dp3TRNmA8dYnvnSTBsQRlm/VDlgLeDljJpRPWeE8Jj
3tQZynIgedWjTL35Vu5pJ1niyj5ovQyopekPLnHt79PmlneVh5C/6bZ5jHn37sxp
UQFzfZ/LT3i8+Is1nw1Qa2E8pRngpxIuvMLJ1VAIMxeoRgP2STcEGi58qndK432N
d1pPo7yyB4lwMCCmlWmTJPzHQ1bevclKellr+B8LF/vnsdCfbGTFaxgjDtg/iKA4
S1WdadFBTAetsoOn/nfiyYhwYq5sqbbW4MFA9+8WLD6VguvToRM7jBhuBdnlmiPT
+WkyrQ6ui+ufzUSqpW93dxw0Jw62zSeVDjuULF4YW+H97lYVyam1xQpyznfNWEoY
wIyAvfeu3dCTxs1b5J8/N3OB9hZDw8IGqqun/b/bAWC2J/Q/zu9qg/e3JZam9+hV
iUH57sEBKDeoMYAoQrkAY57ladOyroxmv9sZ+H9VoLrEAAkr33Hr+TV6MkNiuxl7
aE3bPl39jML+frYE12lJVYg4A4uog6Y2IuGbL2svbVxfYjwNB6SBdhulKRIiKocS
vPw9bzTcLUfsyMSGBAyhN8bScnDSKQ4fOqGPpG1aUlYE2jUKU/kMFdlJE/sRV3J6
bhcBb9KPTM5R3wspdOIOq4dPHWdnhojAxImTIdYsVJOx2B7qjewiRE7PFJIyrsMY
OJHNH3xkGFA/xuer3VHI2ekj/uFsOx6ibkHlnJTVFlMkvPbbTO9YbiysqBPqWpJF
2dkYZNOZyt4NRWg/OUS8g71R+SwvxskmRUP7i+jhn3qs0dCU8KGP6HKvlGp+YDmM
vapRac2Bs9LANgmZPQ4xzc5qGhOAQEXVTmqEpre/Wn28ecDvo3IGxW1SfZQmcReQ
t4RwWiCr9jrLHO5mT2jFEKQNy3kZiO5li+cCxDyM2TEmUu6Ad3H0IF1iCMG4+c23
xZVLujwP16qggfOl72+7rbqN+xyWuI1QBzZniaWOoOSYZunpPJhXdKD36R6GRG62
uaI+s6flyLRatDLGOvNSKhAWjm141KX7xphuS0rpGkZEGzYHjYSwUI3NsNCy1lVT
vlmdMaDJ8I1zZjvvCQRDH/b4ugWlb2hcRIbsekWHzH2QP6JbBEP81WLPwBCHln3C
2r+lJQv8evRVMRXBSsiKU06NmrzJX3jk366iavWl65PysR2msVFON0LT+oR+Ml3o
QTNRlmbVxdl+mDdlTA7eRU7cdMlfa20cwPH2JSB+mnFXmPBSsUcgsOsoK1XZxMf4
EW3uyAYxVl0G1GR/7L4pcdsfSRvFhLXrlrqaaizLN4Wt8gEcN5+QqlrEYIzM3N9C
H1ZkOIhY7/idrANJRt6aAhzowyHkrYj30o/q/lkbuc5A4M+CJ5F7i47mWUavXxBf
q+8u80EuMZhkDaLnuOsNbc/jzEZoU48xTqU+kWf0Y+OkqvG1yGDR9L2YSj5VPJ1H
YhjSaw1vUqEmvlwJeDw9c+23uSR/4mpr7LZNkNO4ik3ITb0ec57HgNOKR+77cC3E
4pKA1l/YEova4Rp8+g12gv0E98rGmJhu2nmbqDs0QVuXb+QppWFapyIdi/6ZBBVC
G8O+ET+3U/vns6vM+lHOI98WP7rcre5hB5rZAGbhvztxQ4YX/dc1JHJywW47Ob36
D8ZM/3qvKJYttrYa2u2lO/6i3XPN+d9QCpSjyiOAD8GywygJksezaFzHUZyBQ5L2
2c5J45I149OQr9bBvS/rqUvLB96uG8HxlHJ5j/2jHLFp7G8xexzarRMvngzTsKCD
fLIEUgBCzIBvZoKDdJ7Ux+Zge1B7MIHkzsFnFnnvrr9e3oIpVwCn1xURwrPs6YFq
G0wTfc+8qlMO6lPtZ9UbzL2OlGv+XTRZw9uqDUDVDGL68i77yKdZ+aENz7P2oJLe
bunhGDhQ1BNkqCgIUApBRbTnCALf+KrLhmToP9GxLEv55LslYIM0ZRu1nvUJSobJ
a/WCJRFBSH6ZONict1sYZs8vBk3FFaJmphHNVcUso4CwPEl3KI28WV4rvjG6YOPr
iS1DTJNZLfks6QwcGlO0iDGt5c0wb1KwBwl+LrCoLr/7TPb1b+sidpd/JV3uz62j
zrHDVz/yg+Lv8OTCg5/zmrClI//NYTdr6icCGmOFXp0JwgTp99eIboE+Ug8JSLl9
IJ6jAWJhtW7l0HhswCSjQCbgXa9J99QnLPMONL2xtkxkU/F41Y8kRCn7hYp/3U/r
RaqXsYr5injOLtjYxpBWMRNsMX6Cp50dttnSnOCXBPDBJwK6gvjBTF06eehD5RWX
IStldih4vCQj/mIpjsTIIhvMQ9M9ESqbLaSjNyqssYmLyvxVwTEHaLyV0df2kiSp
JtTKbH3FHDAey3BjpkvZGH0ZhTqnjnvp7Ax+3meV7CR5zt9fwU+NTCaNYjp17FFR
nkTGKJbodIm5ICA7gVAJD1+8JF6/cjMCOy7pXTE5QqEhvuMbNXgJ7AWORKa/yPbN
w9/BUfM4kdWL8dpYbw/ZD+t2wcjwwSRJcbxs2+7gjZy3jvEzJy7xXa9bm6x9ccgC
5Pq7jBJOHdXzzKmZ9woCM1w7EjEAuChyUe2GPRsQ1NlotjV6mB2DtZv9DvQ4A6J5
6aDuriDsDks3PqYFYCZRCnBsDWHWak8TiMaE4Y2LwkFhUBY7074V58jtUvEWs43K
scKNqb76d2JXRYvPOGsk8MJSMIFML+D6apDZ3UoX5H4sMqvLt6NmFSY7nqoWzeU6
PFWhaTHuE1QkLyJxlbmPvKxxq1rbmKts466j2K48tJE2JXV6sCq8ho/aL0pvDcKt
W+0rWfSLh8p7D9XJjL3A4VWJ0xoNyRPgdT3XDTUWjM1ui/lsA9EbVrVSP5scMO4i
kxvVWxdUkgZwk8NHveey//hYlOP7q31b4+msh8w7L8t897ozFgfYtMcHx1H+1OQP
4KqkB+/zPSW1sqaVjgdvdp6JErIRu0VibF1KiDypF6Res4TQN5JiVD4HNoicsumy
gza6/9tujj+Ds+Ppep/R6Cig8J2gmlKdVw7bq2Fm8eOqx/Llglv4NzqKu20uwhr4
J1xWZBNJZNEdfHkwqyVuDDEbXIJEmoC89h2XUGGRGHfQDZCx+vqwUimI0mDk3pyQ
Mz/+nQuDZ+XSMVuBmc5v5p6Rd6W8yoUI1MKVIBw7lWs=
`protect end_protected