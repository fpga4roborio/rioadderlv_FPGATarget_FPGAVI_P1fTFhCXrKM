`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
ddtXksX2+yylW5zu6QL2Lhnb2d1sD00763mmSITNX595NcHTEkwn0zB1Dry37fOW
FufOhVzEJp80NC5qZ/+F0Vk7Ik02dIR0elf3clrjeJRK85K4e3Hoo4xn7YbFUIms
l/8VZSb14+JVGURjfswrIyCUotIzlzVYZ6gzoZwDXIi5gQIBf/gI+KxNXPaKV+PQ
Ufys/12rjO6aI/pPlqSm0hCvftmBcnezN2hk1UeXgOIuKZnogjOsf0iJVX2aOOWE
6pD/psybjbnsNB6kH5uFTA5frkzIzkzl5d9+YDm9OyC+k84E83I/7/j+rk4L2dah
QJOvksSIzN867/4Qt8qYTQ==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="MvBXkzurAa5VTw+1JJ70nePUfoQXBvZOku/SMmg4TwQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
oRtzZL4VJ4iwysPsC8SXYCzXS8Fw2gtZTOskLcDV+1B9Nzn1zTyNtlo6lNICRmmK
ZRVu2BmCc2G+fmzynYlNTnSa7C0Cuel6FYpxCBlOuk3OF2tzAmLAuDyOH3Z1Yjzk
a0aHuoCdIRKv7BrZCdALt03JeUmXKPdOmIlkVGFl8yw=
`protect rights_digest_method = "sha256"
`protect end_toolblock="Jn9CQpRhJt4rnzZPRk+dOpzAubz7omckX1MrFd4p81o="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 8368 )
`protect data_block
gD6l00tciPUa6pDNTk/+t0OO0nC/UTtBwLB41d4inuAUA3i/ALrNyoJVcBnAmEQW
ptbcNp5fxEUJjnOxnedyZEuEBxWRieZFQnkRdF269oPJDhyHfcKTUpvysLLAYMgz
0lvWKzpw3AugUNMZO27LnW8Q7hh/IikDxJEoXWyMzSnFbiMQeBvIGulFIzPzZMv+
cUT9dx5d1/riwiRFDHslnPw4aGXHyagEla8Qia6tzX2UWt84G5Yn8hc3osdGdZPa
yl8Syg2bYnpM/+Lr+wT6pC62l5Y7O3JYyq0DAuqJKIGRjr6kl5VbaJXMygIfNpO3
JDlEaDGVRt4mxKVdA99esQ+pmkryLhzD2inHxFcRHCcvQkyDyBve/tHzSeBdE/To
ZfAgyvtJYfWNFlOS0wgKDAW5XWlhcj7gdfIzUPXZnMJDrw75JXl1gHzXs1hsFIlb
/sH/eEnOBW7ICeuBjvcOBo6ufnvjxa9wZnK5653I9+6sBjW8o2Rfs4HW96ANkmC7
YzKXBRiYZNT9x81KOWH5aUc3fCbH34+3NEtcd0KfPM2iFUtKv3P/Za09X7tR9FaF
mutg6wrcPUuta3D//yrI/HQOvouKusA5wjhiqR64nt2vipK8HztrCtAozE/aRraE
4BD9FbSZPFPcm2+l+FUoUL81p2XMz2/OPrQbgwCGpVIJ0YO9DdPl1eUYdWXB5S8F
xbdFwhtV4mYfOCSzbz/aYTxuFUGjyUhW5L19JqLY6IJB0Qh5rSSUksyXERCQKymm
1sh8vtgMMToNIFn1nAM0duKBekhfErWb3xDpyolB+gHcYKCZAd5Pd7JpQbmZw1Re
lu9R93lzWj1wkHs48YMAJ8dZbcCsWfy0X3TtwXwJBz0HV7SLa0wkNM24c1yx3sqI
4S5CfPcTGBlGh07/ma71M5iGrfwbHbhZTBFYEkDPzABp/CVRS54EBoE2KsO4G8Ce
EcjYFNsrQa3G+4lPST91i2nUKc42ID2ojnGbi9gKffCpG1pp+7j4qqkyQom/Ems5
CIszvJCuwh0W4z4zk7q/s8U3oTYVAi+LhH0BevAGviIfH39fWXKk3XFxRugMyC4E
PEQ09aAYQo1HsFiL6YzIFW+xr4gB8GCQ3Vc/0SfQdWls/wV2zSqF6Rg2u5gRzFvg
3oZBO1TzHkKigwYHyyG2ICv32jXr2YJSsoSwobAiBC4ifa9Urcnatp7ar9NuwSAH
9pDMszdCqbFZYCRece5s4Fdf25g50vW5dgeG6XzYEFDnmbt09rGZgXEB/JRTGz6k
8rdEUCPCNYxk+JxTmQeVBo9qSqVcIUeDTDicfAIblmTMkPS9rmYgBra2Kg5g0CgH
f2H6qUEWZW6P2Pzxduod036WVhjxC8MFHquDZmoUwTJVNONCnNjfEG0xYkmSf/oQ
JVe7c1ZIJMxJlWPMFzCcJpx/D6YCG+S0Vq/SND1VTDuMKgis4OMRIdDvLn9yXSd8
QaTbocgKP2rR1XfYkjDe1jBU4qCsK3CCXNSQ4dH2JNt79Lt0ugk9ePonbYvefdiu
u2xpEA51Ld2ctr7vYIXuqAareDjNKHGJiDz/90gEy1xuYqYNyuNopK/n/0qk2UTu
zrc9EDJbK+jbzi1YYRIECpHo0W6uygN1hdaUBEKLyQOvQy5QsUcurqlo/LiexND5
sL7sIEq9YvPGKScv1YG1t/Q7Os9CbZcDnTfg61LgvZsYvDiMsGf9SI2daC3U94C0
WI3Kc1iwsW6grUTchsgC79+A3AWUgbYbb2v3GZebI0u5qhcl5LHRgXNaYFsRSWBa
ESG0JpiUr6XBeYUFRHQ4ywXON5AavPrvVnrr4DFIb3wixSUMkPAwdkVxhH53I9/y
rC/U19ABSxz+HRYSBNY0mvYSqzNcPuRCYjo4sQRIVodWCkgUjUm0Vj4Bw9G98A11
tBD654NVnH79l6S1+jNku6DeKHCxaouCTdtAaeUWhlSHCFEqX0zvFaDW1qB9G3kv
0JyxquwdHW673UTow5PX8qQjwCy1OD/pZHbAT9rKVWTq/pH0zMiV+xNQISt5pKNs
+JVCDl7LJUiUg5SMPIQexGlNc9JoL4sjJtmxjoU+v2MGcfdu9mjXBLntr5sO+uws
Zj+CmSIGQejDxI8+8u3I6AQ+t69IPL1J7zM9+oTJkzXoMQ7ZvM+C5NU+9JcxlM6c
c3CUIoGvIW6sdUa5nX2G3Rr5JUJf55ikCNiMqXHLj7n+yrXHpA87Y+t/XL8Pvkbd
+zteA/QqTJJWoStyAInirLErtbOkoCKFjHCqEx649GSj07AgCLj33igi9KShiiaw
0NFwPV61Yt22qXprqq3nJaWLqw5IGnOyLwIWlxpvlBv2dXSLu6mVimKv2nq9/nW1
pBt4e3CInMuMOKMBcVgn20qAbVaaS//YdH0Xm9aex/2DJ58Oa71HRLiLKJdwHBAE
T+OkL1o1ZeiYvBXyniCqe/VCS7xdbtRJI6EpoILOP/b54IAWWxziUEPLzsPzkU2/
0qJNYX6YxpeGvbvNtBZ0xloY6ItUPp/8DVxgZMrQlBwS8NLthruhqes5x1ZN1PCN
ccWTs4Gg9JaztxBu0r7yBXhIHD6bwTVhVt2IIkQ8qANvDtljgFGyJy8kpKQHPx5R
P/SeyURYSi4Uz93B5xsfUE/IAUGl0Igeea3oMf3Iv4u+DRr3vyuH8MX73njGxrhN
gGGH+xmwXn0gSjOjU1anBzRwA6STb6ze61TEY2harxhmhR+eeHaNeA964fd8HxfA
hQdVY520rkDyDWe+4UOwxuFINiOOKcZTnRZsfT+V5DVKuy9vCQbCRPj9UWWyOC6Q
BK139LbVg7t7HFtSEXQZ7/YruWcmLRMONcNq2WqTL5r3qOPcrHdct43mp/D9+W4w
sjuuqne9rcQoW6HRHZGAN5hmsJ3Rk6moJVFVmfydlaUZdcDNnV8lbLKRQo/xNYP3
PGPEYGhiADXVVQKomFPohCLKI8HKtDgGh5dSJdwQC2973rKBu42bpnUiD92Mfrya
8UPLBcOUW24aIQBZGx5eIocV3vFmjfz22HxtrDQCymODYg6OOkweGVG1It4PQm19
pt6OZppN5Jo+/27NaKaeYGY912ot3h0/PeRClPAnMCk9NWYVmswG9tMve3ix6pBP
b+UnM99cdk40BRPWXAJTn02agxhtRdScWKQuSEW8Htcj6gNbZuQwXMIE6FxFBjO+
vUaaEhLNiFNIb/ZZDSj049WNFGiOlQwuZCmKOcmzGIU40eTs6EP2K9cwn/e9aYkU
JlQHnQPt3bdZM99c9B+jcIs/q8KjdtWKlz0fXO2R+jn5BQf9arXEG5Mb574ogwmZ
Nx5/7YDEIvIecNwzb/cjaLY0GvkZg4ZR+zMjUcZOHzugAVKhuNt/kELXImFIEMPZ
kZG+riczQ8ELC2fT8lokLMqB22I8eR3WGZEPuT9b6wJi6+Sk+kqawtIbJKFnYq5H
vbwyAyYLsISI02XuvqkBbDdK+C9gueJdx1DRrpdQM/XZ4EA74QNVes5fHrgAFtT3
hJKjQqnZsTOhaddWvQInou2zyQJoALmYwG1FgASP22ZxcfB7hfJ7uUlVvbGwBgW6
BmYREPiRdgBA2aDssZmy38Bxom7eYlGU0q45tQy05JfV3FULsJopqPyoLfzwkCIm
gmc1QHDtSe8HbY9lu86bD/S4KMTcHp/hgmkBPTBHH0+89sw+PSxO7zpMnLk8KHbW
jHZ9e7ZL1YBFQ0WDjZfWc9UazXgSJEO6Em6eK8MuJWZdvRL2hcwwplyL5QCk/1dS
0ZOVDG+E/ZonASqw54gtBdZ9tGTzgGm1Yio+87hqXKygKMAOW7zK8ootxhXdhQsE
BSoThAHOj6UYrhbrY33cCAr3RZn/ZpQjvgE4QIG8jqt7qCs6jnRLlY8/t2+xflRt
kabNkqwpDQgSrhzupCQXW5//Kafh/u63cnp/DH+t05SIAgLSQEtSp8W4L/nLAhyd
p8L1SJ9FT/WtS7beQXovC9f0Y0CQnTONZmt9wqTcPbhGf0aVzhEA/+xs6mLPISdr
9KlUfnDoSHOBCdBu7vqisJ/b2HYHfswLBulUzyrPCYkvD64TQfVk41Fy1omxSwy1
U9WsAxdND0Y6Kcwv8CMuR/BZ0+/U27KE9FKC1UCdVUOAbq7+m21wx5jsgF5FIkqg
BFnSppREoD+nFPqm/Gh4pwKFyBavi0HJjEhcyxjKJv/JReoOuz80Z+gAXwUYECzJ
xDhZ72CDDiaO+IFPyUGvTbajivKjF0uEOXLaKqClUnjQ0DJr23Zi7ALHqtsN1b2o
t2O5iy9oEMwuJqtN3DzznVBBMlLIsprpCCt23gGVEzMEtc377b7pik8BJUqilNQo
heVyjD///JwnvbwygoT72QJcIkp4o3OoSlWaGsPo3y1LCzoPxnxCr82rh3YH+i5q
838LBlFufd2kx24PslhNnnzEjPh+HO5OK+vDDMp+alUvEdc7tP/HBEj7CQKkNMBX
Kfq0QhB5teEcaKITwtuVLVvI4+42v/NlVCdOKADGEFqfwtC9k6uJkqpwwqCbO4ob
+2j1NZAWJwHGGFMxisR9+GWLNuvTTLrYJUUYCi/EFKTIgKGP7iFqjQP8hkYoqaSK
vv78S/JF4I+cQcSlqHXBBy+V9LzE94r/NdiqJ2++cl+qtmdQfhN2XE2Y1y42Wbzd
CFUNO8KwMiWvpB2A4lFZW0SLPzbGH8woKtbRiJHAEGB7JOWiaGwcI392Gyvxqg3l
Ani7j4AZ4ArHBpbAEjNhNoNAywI31P7kUogpMkUilQp5WsLPWaJ+viYibK1kqlGe
JEQCN0hfEm4KCjEVsBqZzt7STGKUyGFYDVedLiDGmmB48ulnWeLFSsy/cRGT9v6X
1qPwgIEvKdnex04GhaRu6vWd0VN1oKwdHhzvAqqUoXzBpGyxQqcI9dw9RGr0jAh6
z1cqhrCGMqWLnl9SBr3J83S9+iFUOq4QbAU4TBGuhCKk/vN9CcLpOHaKGbt1FJUa
KIThdBaeuTvUB/zTc+9sAtin8Xl6Np2vUzNHwB2DGEXIsXcvWVQ7Bf8sGGRDoE/f
BU24uNx4GTmlN6bec51MpLAcQXtue+vqdasqliMTEQIZP7FrlbAPH+mn0fuL34fU
Y/KyaQAtUAiXhsRzmz41KscX+Dmzc2fJguWpVpgttsjjyWw1PVmliaCoasGnFPRX
3Nra9CewcGO93Q319v5SAQAVxycXLyiQ+9vuWJgDo2Bc61cVWmAipk+PeNWCbqw5
GTqUqgdIUpzEFDHP5XqkrKwzr/lIIy/+Yg9z7oeUPZsJYDidcJR+UQ2hDOEw24qp
1tMRtYZA8wzHrGv0v7n2Lf6l0j6owkE7HRL74JBsbgZlKmv1/3jDEyPwSvC93jUR
TOqm7msFlnprHlGNRQhM+ISlHGjsp8BrmJAToNy3iC988RRcRr/VPUKXJSlIrO7e
YrUjXdqzLYYgb4i9SzI4mNH6bVyUwajkOIp5p39VZIzZbJYsehjpwSh0xtAIcgCD
YTbS9YA/3Uom/WpsvNcwEa6XEn58H2fOakdKMmLoI5IzaRPFQQyw5PT9+htzjLLL
MlgDMQ5qcPgkfCfaI23aL0GtEZ7bVjI+l9/7oHcqDlsXKhTU3+5zQBjTgmwPe5sU
6iRjhyXasVTbyhTEtm2B9tNGJ1obnciNnWycfVXQ1tPncoQnz06+7ThnQ2SwiGEL
YnPUR405GMGPgNAM+SXLg3vnmVYdw4ht+lltetp6kBqlBik/Msz7vqjYtN81Fupa
Az+w9fzgnizjK5hvnBGgU+I4MgYkqazgDKZBt0XsY/OH9duffHLgO/lZG578ujoj
RIspok7u995Ys5si8BBQ6cirFvwVq1iVzy6kZXVj9/sx7gvzOQBKRnCnahr+A6R9
h9fMkkszyiBp9bQKj7mGGpfLgXJ8Yx8Orym8iF61hO1snr5X9CCwdvceddFrpFMN
vS49maPKZe400koPn+9GGe2BuMtZjn2EliA1vqYdD4IhPrRGZgKVPQCMGQNMmP2C
VJp+7DK9299ZtVNgGGjoJISDcVY50r9pQyqWZRQgfekR7tpVaTjIDQZU7bP8s+xr
gYW08hslVvBn5gAsppfWiGTpvXCJIKXUmUGttEl7lZveBimORHnRJwg99Nx/o0fI
rm/yZvQ+Xr6TrYr+59bmiPSkFyRVBcZEopVJMe0HUQ3aHCpVn1F4xa4Hi9I/pz/K
mGfwUxyWzGCLDKgu4ShQ4hEvU/6TQXr/IT3KppgpySLeKSRNXARkDUFwS8Zwnej5
PsahwVxQZ/0gIcdc9hFrBJ+xlAnWgdC3nMp2iIQB0gpPyKzD910nAgD/5wvXXpTg
I4NQDcKa9YcwCSeH+HdBlVYPxiHSO+8JJZFpXoIvwJex4ogi0jHcw8PJoauxp3g8
R6AG9Q/C6TFzi1v2zPJ0XBLRVqaBE67mgLITRFqCwOscCzvZZAaIHhZEhKQhLrPy
/ze9ro20wie4CYcuFecMN85Pk33MD5WrC9MSSQF0eVKQJdujo2Ub/S4rb34MFQNp
CCXz4IQnjp6PPi7JNlCK3t4MUbKUOC7p21pMQdAApM0vz/UCW+oo2sAyHZqTWnQl
nvQicxd4UGCNCQfupqXvJ9GPv0WcIYUMPPRJWRnbaEIrLhO6giK5rk+xBnbjCcAk
37Ec5mSBUMolD2t6kSuUOugwqyq2XABTD1Swtoa1Xg/qb4Vey4FTtVrVC0eeT9vH
9QIrgtQqH/jRT5jccyOJIxMe680UZ8iJ7Q5vZ2wsS8gY8fU/OGggRdM9qfMN6c4k
VapaWJzpuOT9S0dg4x6ZoYTiSQc7J60RwPQUjP35iDviG8lbrfD9dsWGnozPIhsD
GtwLlkN9fXp6/N58IVs+GMDA1Q9cj/syVdhlzwvh+5963eRs088JatGe4k0Z9h3n
18xCzxqELIehGSUi5ucIIciuAwOt4HA/h4Urs38YxsYVIbAKgNc4q4p3052lemYm
tPb8CbcUYZ9Cu9C8ZwpA+zt+70eJaoIalqMeZ0hWQ3Y4othf1GoVRv7RbQtS43ZU
PwP2/eVmyVehDFg09rBNErEnWsc+KEV4USw/WB8w5EqBMnZTSvfSYvv0mJNZCVnQ
WPnTcCbTQzvl63gvMKObg161EgNTzvOJ3qsyUFSHZvpUe0He4GwTGmhPZiq0OgmW
JRB6etAVLre2WzhrmjKvjLtDkWygiDxDUotCb0Yt/pjL6AZcIjcJVYCpwbQzmzOB
h09StenG33DH/OHhFyTR6BICtHGt0EJZNgf0mbOIg7DP1LqrRQm/eeQWIqxq82zC
IzojUKxWzvVpb+2Av/Dh+XZKJi/ZpuNrIzGvW/rIEwE+P7ioGwnCx/Yp3Y2Z2JxE
QZXRssYlo0q+SYmpfz2rhLHoCKn5/pP4oaunjH9GlFiRBYBlKqDNkr9PfkqbfR7B
ndzsG7WRTayBgjuXa1Fzuc/VSVgumv9+pojE/nX57DgjknQspDw9FipTQ+JTSKkw
uAWDSJjwS8+KFtpGKTg66/bDVNa3NaPG239b8Zz3Buhak1Az30Qv1e5XQTbQ5njm
4FCQw+3r/VQlrNQRNXyN63Evx75aOj6SuadwLQWG7RNjpXC6CEf1LJoySOXJPtvE
6y4SwxDGdifP+ljWlHYiAZWZ/EcBzwDi4pRiOm2aqdvuUG/sjtByQUTTJsRIIOYU
5cfEIz0O0H2QYSfQikAswL92seEP21U8LiEyhmIQiqRT4yFhVdPbaJihc9g27L/7
zcjPD9s3upSR3JfXgmr9UNElr4+LU6ASZddMPthitYUlZ1+ha1+WIEg/J2zLuMsG
WpRtRuJ2eZzyXlDAena+0Iyl0KsDzhhIlS3vl9gZ9I/+cvRwrW/QU+hCenoWLQ70
uGvvvdKm4hGUGbRcP8RF3PMAUpL6TebDgEs9bj/7Qsi1cUE10CB1Yf2XJqW1nJDd
rVAEqv5OYEOsVZlrXVpdI1gOg70KpCPaj+kZlAjxut+1WXlD504hMk4BZySXmU1B
Z7v+nz6TSalCy6d7vU09eY6EPzs/8dLXsUGGQIfoowgLa90WYYWAEyFGzlvldmQM
s9pQdayKHhTMxwRfYyZeYqzo4np2pvQ1SN84T1NMVB6CJOrjwoendMMbtId5/Lew
xBYttSLRKfqlMBKn5WO8Ca+hgyHXHutq+CgCSMIW3JGOuFumUURTSdTxb9j28uRq
t7RSXX+VXluSO8VoKzsj1R26Sn5CNRi93gE59bT+u7PShvELpRpuP1O7zIxsc0qq
d8/iI3JMQ5nU0DsuSpNEgVnmkwmhre6aN2onFeZ9DGks08eQygFICgm/8xiMaJT9
JqjoXY/5CEVhy4/lqtywk7Cd6clxT56GKQjapC47BTbl/7VRZvFs0HZDbhhsTplP
wmCfGQAvP2uDWWzEK5GlsePT13DtJ2LbTxYPIfV2JzYS10mNt3taEPksfPrRsNoP
/rX3110F49fWw+75zJO04lklYMpBWUrn2NegTlDzo00gabX6HMRoVrVQmxnsA8j4
QJOpIvk5xYJBFCICwIRJtgzfjKXeEMSE9zHT8goOhvS2Qypa8w7FL96N6unSSZCk
eZOC0as9GfOuyYiYeTsO36rKV/zYFAGA23LuHiNItdQDrIkomRQ7rDGl+GXqIPxC
AXuwzws7ksXQ/sokfH8gCdYTjemZolyIfmkzzaaNjkCut2YHEprBYlBINVElRL7m
h9zxSp76rr8nv8Vh2qOkWwtGS23brO/rtB5FkiU0f1UI7ArP9Ud1cKyGVBJEJCoW
T88omEFJ8nJx8NFGfPgXVvMU5KFzRrCDqFajXEkiHHHP4P4z1dxTMjQWL7MYq7PF
tM2puaG488AROyY4sdu6gZuWUK1AVJuHNt90c59SOfn3z/JNHEVpcLzuNSvP+cyk
Lf7Tx9AYHk774R+SqbGtfPCSdeQMnYx0pOvY2KQgmZ6VaQJ9akZ6O073YEbych3R
USxcEecM6W8qUX+ecxfF1SRtt+ibAT4S8dhlpa35b9aK51jcL1/6i3gYGeLr8R3R
s/xbHMXCTyP5LY45A392vANCmmi5Ng7AoH4jbunL+E+5jHs6zokleFrDeuKL+qX+
yA7ZuSNIPDlPXmy3BPngbgMF/dNRnJJDzuRlYoj7nHZyTwqU51ioFxHAqkJi9vAm
jK0ickgc8a30Lkh5hmAOkNX4TcLlLLyBqsIZUIhVuTfVi8OXMITgNOVTIBeWT+cI
ZcIJV35mh13Oz0uepr0oNXp6+gJlx1ZQMiGOvJFxf1w9drQDsGwAcNIQP/hLSKa2
zb/gCEhI9hTuvYGK3yVUUTlXiMX5ICHHuwFa7se/0WKvUwuuVRtbjcVrx6dDtRBP
TPNhj6Mnz/ppwykO0JR4TMjg+M+WG5dXTJeF6hS4HIgNaCmmQv2j+ZsIStxQNrBz
FCOXWZGCkjjXV0Qodp4R1dv82AQBo15+2/BEfzgxaUXxtDYC3P3SMow1sCKD86Zj
MBEpI8gRttJYkxLcrtUTXYKljAl577KhtKClPmx0sv3clWmxcs0lDFz8qQFLLAkY
pmXSPYnI3MQSazHFUI0IM5M7oDyncgb/MEDiJIfjBq9/cjbHADw95SBN/7LEpANr
Ih+XKPh8zUVSBg+jKKn6+sZvSvxeJAkAQscJy0w9UIaWC0sKJRLEqVVOrbXe27+R
LXbGFHSuRJLnfmBXoeJ/V3ZG8DR8v/ar16PFfwejsrp+6HXE0QGnbdZTtvpxuFLX
Tn/9Fd02bAeCDlsjhCRJmf75xmXoIcrYjEjOZeD1G37WVWtvN/qRJ/gds0Nc4/4z
X+JspQ2mjxr+9zui/pzEPmjRaKaM5CHMxwgX+nF6W/OfgUwyMa6HWmoEZFtp1rbR
Yt9Amc6ceon3zZSaunTY4isJGBQdUPm78VOKILdIYeaTp+8QsKF0ORWvRq1EcfB+
8OgZZHCGg3rClLRxrUO6gjyBMvCwOIWG0K+LsWEoGA2e1hUAVgD7ncRTsu4Q+QJk
e83cjq8s8bfx43uE1U59ffRSs+qdMs4Qw58zMLttlwubN0lJ4k7GCHDNUmjON76/
LRJLVGXXthO+i2ZxQrKJiLzgFrVrfG4x9vZVHZri5ty8FFDbExwxIU8NzVwl0stw
z3gATleIxcH8THUvyOaFWrmub7r2aeM0MNSgHzSmWwmnDj4klCKc8XPy/Z/AeGzm
oT00TKi8c7S1ADorhv4WpbnWdjnrSKA4Cp9RmBbwAUAGA9riMzZ8OhUPi7vn7/0M
9aqbQP4j/ma8JtB1HwTAe98fNA32KFkZS1Dx1+HC8ZYiXPI7OXisDuBs/opMMh1+
wR5Hy3o5efpQtZqE+1Ih4uk9PVtLCSPYuiwkWqpQiZJM2SXfXrPFS1kHg4w0Fxlt
Tt4ItTBp14jTXu+ZfqE1VlcnkEx6SGrieye4uftjStdFPtdLgVl9DG/nO/ARJYud
Eyxg7TNanbtRRMaZ0GSHRkx9USfOFDF2Tk2GmaxrwmAhSUs/Y32XoqJvQnSTDBbu
O7yvu9EbYSLfIXVbQilqyJqYAZowSnu6w7Q+CPkeaDoMAVvElVH7Y4j17edRYbHt
1h/YWncDk6pOX3a6cOi8KH/Shyjqz0K8w7Hhu7Kh2ZPU/C+F2ZSYQMBi7A7/wIb6
nWtBhoLk0LQekHW8EilU8N/kD2x5FRlV3Q91A0ylcx6f7H2z/RmyPJghKAKVr8cJ
/AFVutgEC7gX9MUE4M3/9SX3FGQmSdZFLTjWxeyQzMrV0tHM6+yGchqLhhKGg+sV
nhXgJbYijrg6YqSA93+x1OknLLjusyCYl6l2qPsG9QZnu6J/URhefo04YrdpOXFy
Kg8yyC6wXHSFYcR10oGICGpG6Ig9mRx6JVODq3d0ng3y2S5TnP+CTquHVAe8KzNd
uKT6P8W8Ta0cwc9bNPbE6nmJBEsjp4L0GZnujQ1SQcq1KRDISCZ2MIzlZ0+c90SG
Zc1ueS3RllYMowdjDxJsLdonfYY7FtB4feikTe6xyAOnH6uA/pcbhnXcEcPI2jh3
FTdh6iwLmU9h/cV+Onirn5J34qXiEoYli7Ekx4GTN6l9kfQhWDTDUqMisoYVs3Gq
UpjfFr45jzrUlkZRerg6kNAM0Gg7tRAn4gcafwt+dVfcHWF0z+FXzPC+6eo9RgrD
u3YhFIhIxfZMyoGBdyjtuA==
`protect end_protected