`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
ddtXksX2+yylW5zu6QL2Lhnb2d1sD00763mmSITNX595NcHTEkwn0zB1Dry37fOW
FufOhVzEJp80NC5qZ/+F0Vk7Ik02dIR0elf3clrjeJRK85K4e3Hoo4xn7YbFUIms
l/8VZSb14+JVGURjfswrIyCUotIzlzVYZ6gzoZwDXIi5gQIBf/gI+KxNXPaKV+PQ
Ufys/12rjO6aI/pPlqSm0hCvftmBcnezN2hk1UeXgOIuKZnogjOsf0iJVX2aOOWE
6pD/psybjbnsNB6kH5uFTA5frkzIzkzl5d9+YDm9OyC+k84E83I/7/j+rk4L2dah
QJOvksSIzN867/4Qt8qYTQ==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="MvBXkzurAa5VTw+1JJ70nePUfoQXBvZOku/SMmg4TwQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
oRtzZL4VJ4iwysPsC8SXYCzXS8Fw2gtZTOskLcDV+1B9Nzn1zTyNtlo6lNICRmmK
ZRVu2BmCc2G+fmzynYlNTnSa7C0Cuel6FYpxCBlOuk3OF2tzAmLAuDyOH3Z1Yjzk
a0aHuoCdIRKv7BrZCdALt03JeUmXKPdOmIlkVGFl8yw=
`protect rights_digest_method = "sha256"
`protect end_toolblock="Jn9CQpRhJt4rnzZPRk+dOpzAubz7omckX1MrFd4p81o="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 10288 )
`protect data_block
gD6l00tciPUa6pDNTk/+tzLxvdHE2s3DQL3/JqqujQBC/Ei+vcAB8wM3doqg5vTg
mdfn9XB1bLOis2CVSfu295W2DNwHfMSTc/8BhCDRnTlLIX0UCJs9Za0+LoM0rMrV
T7EjVWppbP+Em6PkVKCwlmIQ7JKaifJ+Y+kjw9HCGboYo5074hY+K/CBbfsBQY86
9TaaQBreoqF1XYO6tFmic/SElYQ0CC8XuikdkDzbSZEhCd+p4d8xCK5BkLSRrxYM
EqbSe5pomH8rrG8hMz8dxxw7CdemhJh0WIJEa/xA4DM+fodK81WOO4083k93gEOr
AXFtaqckP6cDLywbzBC8gVPnsf+WiNhg4BzxiR6v/bBY0EVKvjwNXywEuV6/aaTC
wULj9kJmj1DTfrnAaV58+ivUE7csknUIxWis+NM0hqeZBu99SpRRPN45YeTUZMPf
rKz4bmO7jEOfWwijhg7muTjnHOwB9ESettYdhTNkvW7Q4837JOzUdD2sRWuJY4X+
MQdbSpUDqHIw1+bJ2qpcl7jxN6zWki8Fvj0hRXUoBeVWec8UR7FK4x4lxuKAFoeu
eFzxkojED1Zl8V0ZSpMebZwB7TnPxcgtfbF8SFFnvNeJAWCTkoq/RJT+VhkUVkgi
bPvzDSAimPoZlB6usxYSLOugfOnfjmrJCOcezPi7Wtk7AskCME3CQJS6urCdyQTk
FOEaLY8m/HboyyXIsYbS0tbvH/5y17z0ar+gIV5NHHyeCXk65Xz1OUh46jbOEtHs
sDkVoFKpX6f/3ukxlVnXtAAicZ+dSWruBW1wkTYEN6gdYOqvyqVRGXN4lymsGrOw
funonMgLIwb/7E1kUeSO8FrrLKxrxoefS2ZIkvaigNn/RBJxuiN/Pkfd012CrhB4
WKfH4ilChJAPmU+bWHOTKIR4GYDvReMQnV1ZtITZoBW7b4i241suCPwo9o3QsxsP
z1/j1r0xwKIreDZzFbY4bUktqEoABLoHEb7hY6W5I6nBdXg05hG52jcsuOfxBLz5
HLXXcW9Sx+VaUZs8PGF1anG0Mc11ucTNx2l9tyLCzVRIDzB6oH6/7aOXQWwR23iy
Hol22ENwY78OWXG+6Gjz2rEi7QvtzsQzxkMAOzmB7aj2SwO4QokxRK2WDLRsmzKS
Y75UlOAGhuxois9ZPzciUtq/E1GEMENQq6kMXcTJA3psaeE66u6NPHqxHOE0lZqn
GSS5EtjFBp9T49ogqwL3LeuSUV/E3T51rtCkce5Sb6SZDYElAvrg9zJQC4s8PJ0p
7NEJWzYq6PurL1RcghdMlG5mk9UtPvymFWRkofQ26WRtSQynfg6T1U4ZJnOK2JxF
KYLtFzNwvNmOUnBNANKo6+yhjJ+PmPscJ84gpVo1oYJkrzMyfMk72mAdP/Dp7Abh
rdXbG3Qzkq2L9aQagJypl6NOFIM0FVFLTBV7evZDjUOxgGHTpaSs2nLFUrY5KbdC
vktzl+1dZPgznuwKvNyQ5rg0bqKO9yRHh+3IHhlufn3sQn4FVkBBxXUuARCVqO7d
G4CM0oSUJQOloGP2mXBfMgIrYfFn95P1oj7LRuT8sN4aBsueWNxZqYSDcDSsN5HP
Ikfyh7NQyftmIyWeNazkNuO1erwenrntSO2qkGJtJiV3AmUa5aDu1pdRlONG6JCC
jiqmwfGh7ixdrzZQvNZBlgWsO/c+FRTpen1RKB3JQ/fzhj6MAwN9m+BWUy5bILP9
9UlEi1tbjNtqWMU/TUwbA7GE5rgSzqEv9+ph6Dat/Hj7wchOvJHRQeZHpk+qZEvQ
ubcNjBpvztEnAOKbvwW0VMZp5VwSWNzALOlarZYA0638bLiQJ/GpfT1tL3tvvRSV
hBId1lge/Z9sBS9Dj8Za4joT6n7ogb7k2pffdk+CQou/daBUA/5bpI3EptZWNBRK
/3nKnf6f0W0ZcsTPDYNMI11gcQAA18X0mu3Qc7Gz+TDfwj5CbaBlotGrsn4nv4LB
xsquIq/7jNlaTMisPqL58Z3RFOUXaVolZslAbB3e5BqoEZzIYR5Yzwjy2JejK6s7
KT2aLre55xzA0TDMFbSZdFlhJP+aAc2/dWgQM4sE1e1JjCImanuO5UXOP8mpuCY+
02vd9s9WFgVPY/ugWdWVS+/HNGzG0lBwOJQUn0EaovWI9S6PbnvbFW+7hbsLmK6J
SQoSmo95Tq6l5YatTC2LeV0V/U2G0kDf6GyiqxBnzck4PyuWhmQg9jiW4TamyDuT
NcBW8zKVcsbEJx4kLsuU6P/5GQTPqi3HB9VqHxNNWIC2r7ZsMhtoznBFZddufnhD
wZ68yX44AzkkmUFAkyXlr+OvaOcg9T81xdGYNXeYkvLHOFWrwtv5RPAZNYQouDd4
dhDmeOq/QUhviWIM7x9ML4GZO4zT6lf0zC3z1iAqieUilNG9XDdKhf/LwbeTRY8M
H3/LF8Do4hwIJt1NiIa+7UnHj6hjHqqW9TVCahQFWM/VByS8wmrxfl2ox3R1Iq47
S9e1XlOjOuYdenQFAeLNwUrMTSFpEzerMSQd9n8nUVMXjeQUBWv9bhjxrVuhbwGj
M0C38bPY4CbJVloNP7hXQhGvw4ny91QsXgr6xwjxBqXIcqjQHaJwGqYOGmR404c+
zh8nqG92WC/4KjFlFt+D8OwVn70D2FGiVZIv7t0LAAfAo7GMIK+NfkAJaNTcFHdW
Q5bPbos4x62HgnZ/3Avxuik374cP9T1ArTyRE1LnNbc2ZUV7ymFGJIAK/DsOBoyY
TqEkm0fNVIaIDaZ0S1HYnGzIAmyBDmNg4jEhWzMHsBbBdqUlaVS5wKIXG2AidhVf
pxnGuZLFIj5c8SWfUsm4ewx9lXXbBEurzmU1xjdDvSczZXvB1bB3wZb6N+Spldx3
IjiwpzEGLayv+dlB/wontacic34utfWh0sQooX7gWIJutzGp8S3uzQia8dKrYCHC
of2pOelyXN3cJVlNMKSM9pDRtovSRrT64PJHdG1DD0a85ElXFOdHpjctOgHRrPxR
W5uAaMKiCyduOaE3mrbqURqqcaNWXOQmw1x0c2/AAIs1hScWgmk/g6Ko/OqNMb4O
+whKIcR0EkriIyvclYlx/GufxT49Qud1MjDAMVSj+433v4XloQh3pmMRqqJzxn5h
VtQT2XkQYdNz1RGpMJ5ecpj+D/hD6XmE3xX9ti3EfRjL/+rsNer3MC+Nz8T72WfH
itDm7oUnEFVd6ALR95yHHemtvOIbUhNf7S96tz7jLFJeEG4GR2kiM7PC1sczEEgF
4kgGTRMw2FjibCXDYA9zDxHT6EVRRXyEyuM6BkBWoNMf4nlmzhPfKAS3c/2Ge6O/
Lh2x6nKt/ei9nMQh/6/U86YL2xg7BxLm7pq7EdKhsYQfM0lDY+tqnjGG0Xy0Hs/j
ywHUOQ5N74OtISD+Mw5JBntlL69IPqvhzWAvGMYctCyW0LTSbBq4+hNbf3co3fbI
oqhoaqS8n7argyzRNEs85hAXzIqJAHALhPofpLdZ5q9rNquDKEqTXsdIydKMtpXp
J2O1ILDfWqGZ+bDtY3yXiPfmx86i/7LukfWlPrcKC74ssrDn2oB4X/QO0H3Ivqtt
FszmGjvzw9uktMAGIJ46eoCVjSe4USvfTRFaK5CPne/PC5K5Dib9gnat8FJTaoDR
tU4vhbqjfHVyHGEWBnSANSk9Ru1UM3aXtCl9jovL0yif2WW7T/W2VzpXwk+JzGGI
0gOTuSRCn5tGTR8pojkg70s4pZ46wN2UKYOmrWaEDXiVjfsJWNRnjbFWk1+x4NVh
fd+qpLNEwqw/5sXj3z2DRtHzS9nQ1bb2RivDbtAF9LDyDUtnFV680Qi3f+NQ5XoG
0uIiBO12tGQqecOKF4W/jNAjDizNXR6wG4P43Iiw8eSCH1RbNR5Pg+1kmJlCDscv
QuMsEr5Zt7d9Ho+bh1of9l9LrG501J+hvhLAECS2kQLpUPKZhml7mK9jVA6Q3at4
kh2mSOo+xP4OZLMcHTH1aOJ9aGEwRq7ilGWrSZbk84P3el2BsJ61ybRK88fA0vuS
HmUMzvUrBcIQTFe3fmDkhVZMVLtE3GSEBvf9kKymt79rgkyIiWTZFL4NwmpZ9HDB
dkwoVQGZ3MB1diNIN7nnNpGWNKKQZAsZmI8SQ2Ac5M1QteDsWWCEC4FQNUOoKb2E
a+pkh4wcEuAsNf56nHaRZfPgKECGWsZNtY07ut+QzD+RO2HtIwiwEBZgqyv0hR0Y
9ysnKigXj7TqDz2fe7sY8Wh/CSiwU7gPSwtFBJ2whMnJQN7SDnMPQ6pfAN9AI1a8
Fr9xmY9m31D30l8lRILVpwnuGH51g5lJNbSw+wF3ozw9PhLhrQfEbFgMRWMDjdL6
UwuctsafL9QbGDzfgKhQqj0BGWHwbPBJJIGo9LiTPmdqzsCS0z8VTm38wvkLVAJc
sOvd5eFXlDWKI+CHYWzJO6rEXru7E9eIarKgocGdF+hu23UkiFxtd2BB1gmNTxFL
z98aWgrKQoxN6W7dY8LMknpAPXE26lcTf83tAYxvVMayPivJNZCbUhq3OLcbGctS
mQ23wiresPCvt8V2w32Rk6irvPDzmjMXFlmpma5gIisIDb1RHr+MS7kUWf80coNQ
JcewkTvSpjXRenGq/Y0kP/Zt35ZHrYH3OJGL2plLBIy0XOFYaVveGbm+Gs1W9pjo
SLEaVSvRoOKAftYOBHrhsxG/x87grjbUhSAzw19xkluoLXuBFGYRtt9A8A71tHdU
Iw8jbCqa1zgbWMaMsJUEUpD930bpKrCwOsXGvoK0laTnZzc5GFxNxVhG0TAiz1g6
ulaJh3KvyNyfUbDYnW3lkQEppO+EmLHTxGsjwygF+bni5cpztX3tBab8iANEFKeL
qMfdj9qIgCUMRbx3KQiNGjxGeFvKWVIiAZCH1smg9l96LW3Msj66K6HRsK6DPfo4
E+KDQU780AqN6ad98s4urSUQnX/EtSdIT41bI4+VYyskzUJwgCduTScXyz49jnn1
1UQHdMTVrZQs3/HyrFnoGdUSN/kZG8mZP20xddba8Fix1FVR/j8fVz+AIwD7CZ4M
qG+DiXDO2rg4eOZ6WrYhLyeQy2e2I1yZFzXcriBlJxQdrQAFk0IUK8YVGOIZ1RM3
feN6PcDxRvx8cOpkDXR2QaftzPo1RlFTrA4id/RC7Utf1i4xMTtIR7bAQdPWyqkM
EFraQ7yv1HnSDxtZKgv2v7cL7kc/+y7IeCl9Ly87xdDxG0WZG9dbceL9DyqsVUmS
SacLOq0tKcXKVXKpmWqnxv9gDnyeY3lZnKEPWwAEe6BxJhWUxR83AnhJiA3G/Ush
PBr00xrgujU9/VP+yun5+vw7Jr2FbPWDQOEWU8KiuwqoGVwGPWFQ954X0OXhlOnE
6FaFb8+zrE/h2yyVXnx/Xeuw0zmFnwKuFVp9cibG/fEtVf/NvwtwpFvSE8gbx6GC
aABwk5IAfcoENMFx+ek99WT8a6Nyy6i6Pe0m0JeyMiCGdCw1Z+vJ3Fy9P6iFo4ua
Y/+xNRw6RsAHHL6e55ep89Pe8C4qL8IUmTtd29ZUme5sJBO5pRrSeEEyyWL5gDyt
L+GuGXVV9LyeI4sEAb0hwMfg0h9jQintVxJCyc6GMU3gjQPJ3KjZkwp+LFcwx7Fg
5fvCi7zqtuddGgaTImKBExfhCfK2N4FeOD3L18cFKhzgK245PljSW1c96E1/Opaj
V0WtKijbE2d8bv5lp5m5ysM0so7zeA1ZhMCP4v4L2wyd9bXbnR+0vP1RZz6sB0FN
q1OQYIMVFcErXGjSAHd98em2BV05wgGpg+c2bvUEiZ8qFEsFT0NrxfOFhQoXyEEX
P5zXEaEGsKlQReTGdDx9qHIDvTrG3UjJLHdNMxViGGR+YmGgXvK2uHrKBK+0rYQm
wxmo2WVe3GKNR8rSraa3NY8nj8OvM0t21xgG74DreHckoPFZ8xL2wXka5In99Uo2
ejglEAxGA9jmHXzlS2HE2SYywpojCfUHF3zPpB3RSTBa3GEAZ6RI4H0M5HHPWAOZ
bomVeJ6OYz4emvgcMch1hHxamP3GwT+p39z/sVIQhquuPgAPE0wts3aaIB7LtJPe
A3SXW9sOHIyqcSxHHMow4KkkhZRBJCFdYYvvcsabx9oXjZWHpnEdK7jKrcdf0SX3
3pOvEIjbdCtJfZM77kFMRjL4bY7Uh06CGm471PNDgX6BY1dpNTiHNc9WZUJ6wL2+
XDhoFlGTITilG1j2gslfDOkCpB6aPmVEVepIxujbahL/yMegrLOle3NSgEqkrhwa
IyeifzyoYGk9bC+p+/53d0AxpWfkmz9VBDay8xG+uyS2xuW5mBgkEOAbrheGfGwS
k2P1NMo8YVbTt1IiAJ7IjwrnnHSKskW2sI6qZxQTMKGwgBeTRWTj1NKWDv/8mmMP
ldCMosxZgv6X/AV3Nh8BRhh5hVWlMtvp3R/3cq8nTNAvyLF5q1pNssD9xGQ7qvVX
6F7mNLh5q3BFFs4R1USnIisRiNEbsnY1KM4kQfzomuGl/Ve72BagXB9q2KlbOz17
FlO8acRCyiGP/xvxTPTUVZynutzOJjQXOjuJJ6wB3vvMDYg8BPoG+qUudXTOJCkE
UYdP03W2GDZutWy9smAoH+URVb4qAOb/9eR33eyd+RNSod4++af9Lx3pUM5SsgUP
xjDKaEJubeChYDVVZ3zhoVIaB61OPbmjqe++BEuutLkGKOFkDIbSlBCevFjzNcQN
HHn7LlmszNstlUS7sKMHem7yxs10JneUpTqvC0o5Tku20RrCodwRlQr94XJbjxf/
nHRwlgRil9vsvC/dDeIY4NpHJEqM8QeOaFkf80U2fKbCjilRLswBYqyaN2N0bEuD
ICQHsjh5zDU1j7VfSjUcP7HX1LUoSMHK5lh3ms/s1tnF+BsAI3XJlrMUPwOfY9wE
EdrTCKpRpOeGPJL7cRB0Jz9uD1y7JRVEucJetNvF6dhmnt05cszzNzrh2ICrW4kw
pc/WGFsZBaXcRuxRC0ISjUWDND8HbhYzPZvWGf30mYIvcE+2ngzhHq/eQYUlypal
gEtDqYizAWX6VnNWtXG+AbXs6CxtWzzeuZuQsQl1HibwNT01/mckLV/B73g/SYC8
mn1Ma3qGORea+cC59tS4x40FtAWhaKbYu90zpJ8JhkWqLdFf49JDTcZL6FfcurJi
57NHq4MaMLD/+THGZM0t5wK6oTcb/zYhxLUZV3LJUSjkMwYA11SVJ1YcBUTb8iky
NsGLV53f0h86Hx4Ce4DHdEqV41HPVDolXAcXYrWmmR8Yo+C+NtkbV56eEGoyc4NH
MU7U0+akEWle4R6Wq/a/PWgabDQIR291RCwXkDCoeqJHAijFfpR/+LAR85X9pjBZ
vW/d5FPbhv4proOyb6pCTBFii4KfkSJXY1lJeeuMZCi9TH7tv3xOTSmTGdImk+Nt
/B8cFNmj4cusbztukQWvlAqBcdc0si829tR2U14unmDgBGtY498cxEZvTVnWkm60
1BSYh2imkYb8VQYsQUB8a/BqtRS4Xmqn9UXV+XmYCFWQRnaveTiwAxtRMHpB9ITA
ricjBQx51WHp6aNQFWHU3+MWiDU6eJjiCLWOICR8qLsSnpam6wdrjuMN6xefctnR
9KLmkEYeamm83QoHSl+jxJPuOCIor0L8AcL+aQ8qiDNue2HPnHXQf1N/T3WcAXbG
th+2pOmKR+qb13XaGhLErZ0hq3hEgzeaGtVsC9wJOfPTyWRdI3Jy3EdDlRLYIW0U
bQVq/x2mDPxfgeE1Oj/5EVemwfd/dyxD2yaoeKO+oacQhy6yXDD/fjtmhVHCIXIH
KG0sNVHzR6Z3Au7jYttmgezqQIVXRJKZ8Xlu4nbCNaX2ZtIQjOKk6xZEPfnlm1la
N6pgn5i/RGyiDaYVIDRSu+szdeqc2kbtjpZFkZ2HRoZpRXgBNFV3zZTDLrxXkKza
hbw164Xc6lPTz8eYf7ycgphyQwOLJNzGjeVUnNYu7u2YF/LiRBg0HHyTHBplD+We
2F/vOHzQjTCoF2tfc3hdFMNLeU3/YxHoYO59toplBSTV6150tVwyGAVJd1+GD5uL
1PibW/nevNddnAa2IvaLwqPR5FUcKMh0BNe8qNj8jnHf/4U7Evr1f1jvMe1PyuiO
Pe1OkbTvnamwSjBrT36ihMB2t+vU92MZc7rXDPmxWRgehKUIfe977s/vwGKT8RvQ
SbpO9sTLZdMAUr3Mdoqa2NABGvfLE5qXjxxMWTWSA/R3quHRZR5NGMAxYyMhfPn4
7qDelz/lGx4zY4a26YfBW4GsiAdjPlC2J8tXD0fEc9TEGGHoq+eTSk5aZrmMSZQJ
vlPHnkUEFSapYkb7YHHyWvaIdVUpCLojdGzn67AwMmWud9CvHoQwnbPPDQM3OmVX
3VbgYESaRS2zJ2gZJIiVt9ZfVmbzZsDuh4AIqV1nWFBWdfkOrERS0iAwk178vkGA
rNu36r8HgwUaNfriAJODNf3cFfM71sSQG3SGulrQipQlf/onNYREYodM6zUiS1OT
6BWPOrrkdpvuQap+djv5Iu5PB+I1jqRwQ21RHW5cUPHoQ9ep31OWPfhkj0bcXyKM
bSNF0u9TPhNiTGb4KT2nSVV+48i3AjGYyUvERT+Gao/Bw8014oWz8C/TDZYgGhBk
XQ+OFhMkFIPg3H/pxSQZEC7CGhadIHfiRBoB8eTem9mXt/OgnzGBNMV5D5zT7Rvc
1K5tCyViLuR/XosR1PmK69GuyoQdKC9D5PvU4iq2csqTH4/pyYAHcNcx8fUct3aR
nFVmJnnw1r4iZ3JUinHUeM55kR+tA9rVA7kAMEZWAEFNkJHT4rXVC059Dknygana
0t7wYGdY+26Dty6zP1jBYBj50ctcZdJdDWBOVz/UQgx2aJVaFLJQ5g1OA3K2nJEh
W9Lh8FA+42vAuqcrLe5J4ygnXbs4mZi1yyPGm23qHpGOMpmR1wttBKakjGaX+0WO
fDTxlfyecglrT+O6bFRLCqmNPZI10rHPN6dLWYfdSx6sm5k8pq02XTJgFfQpZbIH
lbXBoR3VjdmJwlhMuBDgVdOZyPTt9jRKAszRTXmJ+IOeaeJ9JLvka9CnqMJ/BjVd
kIrpAvueBYV7XICCOvckxdujcOntr713tnjpLMrUh4DJCG+sGSM9Wb8pmW5yLXTW
8hXnqtbHLkZBcNwmdfPqV6HdUMV2yuj8rhm7XEqxiF3aGY2l0cUIGKe3rqTka68N
vmLcE5uyN+0ickzaQ2ut1q4XW8VpHuZwp183eBar26mNZvlKoTEIKQ06dvl9C6uy
WIJjyGVKBnPbGOlevNoWkw4zXHNuE+utQzhHQm/KFeHDTR99EJ+IKhTrunI1DQgI
ESEqrleqBTaqn8Stj3J9s/r0Zx2yvCuA7m7GWxBEOI6La/Wja1zIANGxQuIFUymB
QadFcf0yhp+s2Y71yjFR+s4XV7lxEfLt8ro0cWYl5/TYJSqnGrhLyumngHe1y+Zc
m4U1VkCX812RK6/HMIFtUlScJpURwuAxo3flH2Zy9ok9ntXrP0U1N9pmy0aEQ/0/
Sudr/5t5ZwACF6GpKF5gW/il0StgeAL/Y4NwPsx040yDSzN3CMQJrzFuFYFMN6XT
Kh8aHjJuyE2XaghakiktScNoj9UvEKoC/DXC6CJ6RKPSHTSFEWuEt8ZNnstLdzNi
XR/myRbnF4s1SOhM4bCF3EHGD2sOJe1RdaI+In8/HJyWIrI9IlA2qkUZ32RLjkgK
3OlliM8ysR3geDWuQ5BDRYd3fqHWDBbyi2M3f7y5PJuFAlk/JxLtP32s9kHrR+ye
p5CS5fmPdwbVy/WZYPr0zCljSXKM4CqnOgwDasqDemOs/4LxD23tCCyXSr+eWLVV
BTWihjvOUigjOyhhBWXiDeRB3WQs1yXb0x//cEMmYQqq/vfGGQwQidWIKX6ZMfMk
b8iKPFdyn4/oc/V3rGhDABuqszJFmxBn5gX0PJnW/As0guV66Brkvduy5GKlNJGe
1EJzKGAVMHw24KXFZsL3u5J875Cf2b3tRmbt7v1pffSEGnKjRU9zcSRbY+F86xif
37iZPVmFASr5utfl9M8AU+efkZ1bSouGlZk9DzIYQgx2Wb0LAjnNPMaMNqodZBTG
r8MqTsl9alWUWv3PV7/oOlIAObMCNlapheHdjI76SWvr9Se2Exeu4HPoKGtJ1X9q
w8UW6HwAOASuiBf4fzIymJKXv2e8QVOKgrmI8f4Cb/doBIhI+dDmFPthS6gxGMLP
/by/lkq91qLEXAIBV69nLDRSPmN/OLLjaY9xTQkNOMYMfqxbYwk/dQegmWDzMG4d
PixhOeG1G0zDxQ62OLx9NRRo+QUvjXwnx2HzIrNkbZ5hUVz7lnUamDIlL7tVbd1M
SR5AeXlRBs9mtcFmqrSuF1/Ev+Swj04Y6zLuFagGlf5x9sRzOOomqpDdQUnlgq5m
YVhSbwhleJX9pXS09L5yKCmvzqx/YBElBA/8ZhWrW1C1diJJep6IhTeJpW6fMSU+
HbU5++9DkPTP90AjbsERkgeYkMjBpqnlHqgjJZUvTW9ERBu/ojWFRo8hNegjrepe
mmn9UjFlmCUDhP+1IVfE9jt7rjpZ3wx3W5jo/k9a887Bv0BKxzVZQ6A9VWRdVz0B
6hlsOn3ap+U0u3aqW3BUXlBadog0iEFGI6iPRmKadHK2NJkBhKbF2z7kjGF3DUeu
FFZ3/FSZACJTb+8uAnwijsso38TAbgOrlKr8EN+SxWV5hG0N5jNL8CiL8RazBST+
Fujks7GtoQeUTwZTixNKJSLWIW6URZKk/ffxLm8jgJkqblzQsrfkLYkBiCo60nsV
cllY7k5+lf7quPRTjRcafgjBlXaiKOcLC+W6QmuqsPW5fDAim2dLITUWAbUciFa6
vUyYAjj921mtE5zZesxz22a6kz4pPs59gdiVhWmKANB8ZDrVqePBln2j+REGDoLo
nZaRwBYs0ZFO0cLqcTHOwtwq7e+hSvsAKn7vBvNxNK9WffIA7eN6tYQ+sLlhUv2c
kkxhAwSFJRYVAvxPlXSZVGkXbs2pvkRIUVeBvfiMj1ZBvAsnvsnadNhtRUabQnDq
J1pWkbE655WsOQLWq0jOGlleXBCghjE1NrY2DraSWUHl1btfMqUHlOzagf/MDjBE
n7W4v1JqyOWzJHkBaKKhrqKyjvoJ7NrpkhtSvifFz4k7wcna1aw7eUAoro3Gf6mx
nTvHXcLb0NnovmgVBey95F3EtKB3roJok0r2oms+OI8c1wa0v6pOmGAZ9ABnTzTP
kzaUSuOwlBgJB79bEKJzG/C9QULySuWq7nptq91J1bgAvx7jyvAM8muyjW+I4aHP
/T/jPvdqQyfYoGqbeCnLv4+0Ys4G842MPwPQWDyi6HgYzcAiWuieHhMqrVivyHbH
cEd1c+nLzLIntUaTr4u8Tooj7vZqI45qKhyuvIuntooNmfqAqNHAVaInlp2hzutt
BJ14Uo7ij2VKfkplrpWnqjbOK41VpzAm7kZAipoOdI9pyONzatrwDqx9Kwrj9GVm
83/scGAkPJLoRz47dxqJFRfzvnvYAv2jHhiJbFxqBvvNgv4gNGhB0pCHYUYTDsBd
mY+L7/SVS+e9b1rscqpCLqyBhFu0NNvu5v7qLf4HllsntS3PlcAFQtqVumhw989n
BshP1kwNytTs1bzT6snZLpvEtWUcFNI/N6o85ADO3Bs9PLG9mSx4c9XaaiHIk43A
U0qRJ9XQzHQ5ufqkfXLqsbW0GTe1NA4psHjltcL9ed/x8vXs6ZcG1+KoZT/Zw0TF
wtn4bg/UrlRnKjSpGbDbmCvBMXcInpz3iFbcRuHv6kzZze+NLbAClPlNbHXe72z/
Ccet7nKYnRQIm7J4B6AF+SLKGGSR/aCcAIFU0EDOOn17OUjPWekOzIrEd+S1IK87
/4+ARDyFG0FNeGkebdLNJ6yj0NpmIoNX02/W7pAy4CrKEh0DG8vsv5QbFyu9ga6c
OyQErc0qwemrHt+029rn4zvtnufdpIi7+gMPpPIQjOU/4GPXuB3FXnoXHP91Q6yt
Hi83DnUKLywdoai3dQN04qdQiHiBcI4xFH3HoE+7UAXL/T7koKIi4yA8pWbpuWKf
XQE2Mm7fVLiuGIbM+zmXiJMwB+70q6FYdnZjSD5zD67cFcGF3MVebagmDHwNB0lB
JCIA1n/4i3Y/9MmIH59TGEsCcyguKlfo3XP9Qbsmfb7icoh7rW9epY1iwlXZ1tZR
W293ft2o5q31+Ibjyb43dgDkSsM/pl3GWDrsDMpUreWfAruLPwXvB1mAYzHeyCQh
fr1hSFduSegnAtDwQWzjFK4TK6PbiW3mC+aUVZ03WoawXtdAuUB2HEq02p6eqpOZ
KwlrCN6sw1u3VGOCkQTNcivxq5VoNwASIQhgNvlsHjUxjsc6Q5yJwBBIEctQjbvA
9EqKfyWPT9XNWCBu9ancek3zZ9WMZM1f8rIzPw3FUrtA1vlC840fyaa9p2vgAeUG
uqpTWg5EtW8+AqlOS6hSQEU2e9VygWu42df1V4YvcLxlFMeoowl/kwSdLZQJEjSq
vndCEUEIrhDyjSsoziI8J/FexRflA5g/m/49V4EAaPzfBnwL2mrhHDR8cIKYES+j
f19JpnUMFUioHdy+NfXDsnMdiYNHkJxOj+ecXgVdDd/YtPY4cED1DQUS+pW9jLzR
5HzjseMl2RmgYoGIRH4i/I2nZod/kJCYPNHurUB3GNUoYRviHnBLo03tCDPLIokF
QuvE8uIM/b9VWA5llOPBJ8spAu5rYP4YXUlJxn0LD8eQbahgAnnEPTuyFC84HstB
YrnIOYIMzOs2E9Kba39OVi2XLuGoZyyQoTJ/11ejYVjo9QDXNSaYuwfKOEcifAL6
a48Lme0M9Je9Z8iQr4Y3yJ3X8a9x/vg+/GamljER/bNFjCtsaRKGMIUMdn2OTJhD
6FmZKv2ng4I3P4a16H+1RK2l05BYjYjtdVI4i1uUA3b/FgLcqFxSfJSrccJMUrAX
m9NqsrJqiGrd9nOAiuzeX0WElPKs8qAFiJuX0hERjydDRCQ3bRxuk6nWOVqwWXks
JDhj7TasJ5Uyvy9SwifAp6u7elOXkyZXWthbLKsXIP99WA4GUu3N6BSH1dVwbSWV
iQBuDWSqhEuzH4eJEG1z9+OtQUjj7tzv7suAqM/6Mxa7BIDefBqOrLh5QmW+dhM+
jRyHHm1Ht2svo6cHK6ZxVToDgvgufU2R0CwpCbLEpQ0YboPNyLzib1hL0UqNewV6
t4BXr7IEUJMXadhtS7d51RDKISNhHEo5ry0sUovYSaJrx40IHj8NFS/JMWMXyeyw
JfM7PR5evLGYLF3tJ/GrGUnIbIpdlTt4VLNQBDruOlQPzvQ13oDOH9BejQw+dAzg
azls/8dorjtPtUPI1EjUaTmI7K/jIUnoNjqLTLQExVsDv2m7pkQXNbUVe9UIrS2A
ReEjXdsBTjKumA3I84tSHV22+uPvWLX5+dMpl0vcsZklX0uzSkhHaPAHH4nN8Gnv
iAlcW7QFfngV5xIwd/jne2oRFJHIUewmXXS4wbZQGXMZSPdMBP1qPUhsi05GGYel
nKlZCZ5QbI4AvJRbiPVpSy4Xa22cec1NEGWH+UXXeqUEpYpzwhESDL3lXrPtI5r0
7Wb/44C5xRGjvz+cU2y9AMn6nJIMUmN+B5o2XjeZp1cnU2MeDe03UwvPBQ31Ybd8
kR1IihXSx95hDOxwD+2GJg==
`protect end_protected