`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
ddtXksX2+yylW5zu6QL2Lhnb2d1sD00763mmSITNX595NcHTEkwn0zB1Dry37fOW
FufOhVzEJp80NC5qZ/+F0Vk7Ik02dIR0elf3clrjeJRK85K4e3Hoo4xn7YbFUIms
l/8VZSb14+JVGURjfswrIyCUotIzlzVYZ6gzoZwDXIi5gQIBf/gI+KxNXPaKV+PQ
Ufys/12rjO6aI/pPlqSm0hCvftmBcnezN2hk1UeXgOIuKZnogjOsf0iJVX2aOOWE
6pD/psybjbnsNB6kH5uFTA5frkzIzkzl5d9+YDm9OyC+k84E83I/7/j+rk4L2dah
QJOvksSIzN867/4Qt8qYTQ==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="MvBXkzurAa5VTw+1JJ70nePUfoQXBvZOku/SMmg4TwQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
oRtzZL4VJ4iwysPsC8SXYCzXS8Fw2gtZTOskLcDV+1B9Nzn1zTyNtlo6lNICRmmK
ZRVu2BmCc2G+fmzynYlNTnSa7C0Cuel6FYpxCBlOuk3OF2tzAmLAuDyOH3Z1Yjzk
a0aHuoCdIRKv7BrZCdALt03JeUmXKPdOmIlkVGFl8yw=
`protect rights_digest_method = "sha256"
`protect end_toolblock="Jn9CQpRhJt4rnzZPRk+dOpzAubz7omckX1MrFd4p81o="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 83360 )
`protect data_block
gD6l00tciPUa6pDNTk/+t0OO0nC/UTtBwLB41d4inuAUA3i/ALrNyoJVcBnAmEQW
ptbcNp5fxEUJjnOxnedyZEuEBxWRieZFQnkRdF269oNDrATGT50FqUNlwEx5ZZnb
zi9cuRBiHSx5HJ5tT9OTLFnTHdPO8z/MpaCCURqTBbu7rAoNup3c+j6yW9zW+gth
PAHXOe93jFZxfG7is/AvblvRIPRUgO2tRUy/1gRXgtR/xHqjR7pQan2xiUdx3roJ
iU65zqFpB+zo2vm/Qv4LtkpvfCslF1/OkLjwMp2DbMfF8ch3iRY5P4T11J2mAYyC
/KsQXMMy4N8Maw/riYxqDUUZa05agED9CT2fGyLlsdl+khDkzMpQ03sSz2zMTCoH
qhajmqgXnkVvhZsG+kg638jw6/0UHzeJ8rUUhP71kwMinu4c6oYoZ+8J4WA9izmX
Mc4omfI0GKf5GukWHqm/UkieS56JuJO6Jx2B9qdgZrom083onAVKe5magtqnzCZx
ME1nj6TYMMaGM6WOcG/l1sv9Ml3Xe2nmvOC2sI40RYuF8GyayXVzhn0tPgAAxPEc
0DTHurvgyopiHZVLeFWYYtvL6Prslp5nu+eQmpTJgsx+UwaOH87lo8mVIoczDP7O
pxL21SDj96h95rQbdVQHbMzRHQpX4ydNyeS6TsJqY6aJKLlDqoZ7JfrfxY+5oXvm
CNRxNoUxoRDtZHmDCK6OO+xRyVPenmth5640ZEUCJX2gwur3Vxkgq4Hr4P7aKk8U
NZaEx4DHccgTN6sCKj/P25Tfricc5JcGlsZNSZf752Nkj7pGFR51GQ/3dSBoTT+M
LSgg4b+0zXpzgiL9mtbDj5/PrYKFd+0MSN2bi2vL5Fftzir4EcZs3PM1VMGaWG+g
nKJS6S/wCxEdNZzYV4SeQExpF478yygTyOl7MeQZEGjoMKEmqAIp8iEfK9MJPycQ
uUF31UkOZxnNqGrmKHIDWchiahWCjOVtnaOvC9Xw7umSGeFP81N/GOdI9zCo4vxA
mLi7bAgLTlZqCxnUgyKjuf4ViwCLn+rGkLeoj2efqYfFrJ6zgdPeo8cIgbR7+0g+
kTeWHPJCOIpGZ2Zm2bGimI96AzbMuwXAoa0XimSiwlFgiYNzp/45mPPiAWGI1xtW
Sg0z9sXdWyHaIgCJUrWI0I6L6Wjr1Fg6NEDKclNfrs//MsCHtlmB0g3AeSp1X5Cn
t10BnLY95Iz3kSXm1QNQSjdEgRfUt0VSTnA90PmLfqn3a6ZW0csET1EW+Sdh6qMJ
kXQ4Ad4YxprySdS0KvbrIlUW7OQNad9dei9nKyfXJMFFGT6NaL2n+eTFIpmvjdtM
I6nv17ateicrSeELtkBTtlCz1VWawDxm2RJ7xotJ0pX4C6+EaN/HdBCnv4kGM4+O
3fIbNNgK6Iyx0uairbNQ4GJCluDU6unumh3EvthJM5p55OJJ5t/9GeOjzEWIyguo
VIHbiqmcxprcfOhzgkfCmkGibcNk8gteMCpQM0dU9BNiQCf4Jj9jv+fc5TmsXBz2
G6Wu5JHPsCNal48hcAZiYt9AOmXt8zWuy2IUeqoMRlHRCjB9IXbhWq8741uAPmfg
v52qMGbLRWA5tFroM4+en0mNlb7DMlwy1C+yMguCHHMY1ooq5lTKLqAQcBush5Wj
YxecCh/jf6qca9FUpFVkkg7smRw0We/FZgBqUhjdDPfXmwo99Uyz7rSurCzsELRV
EFZXvLZ+1fFX1m7XaZoByKYhql3zhxMbbdVScZlfSl7Q39cW3xJzbQ6es/TDnyOb
1ozxsRgVeUA5W3xfGmBM6JdgwS67OrKZ+7NzcApgfixoIdo4rCbxNYa7P2axvupU
VqK7cfW97NnmeKn8QHAEgbSqxKoh8pLMz1na1Lkma7xkZqJ/gom9s3ez3x01S/sj
UjX0K4skLf9/ePgaU7oSnHtpBXGq/DSYHzbm9ugLptfNEI5FXkzm5Yc5ZudcmD+6
VQ/uxyuA309BsxUxAtHbFS7xyuAUlMHE+ttC7AJtE/CXvWdOa8+r9lQaqiTCvSsG
s8yDwpY9NrqPj59mM83GbzNa0u1zVN65iVZLAwVk3BAOjdBAQY1Z+h6QmX/0up6I
yJKu4UWv5bEzZnNDilJ3dpg/n+AVjBm74MLsS/M9cMydgzm2jF3NtMy49iHLOnLl
/UTj7LxqOERzO2Uzfu97CCCF72ewKs5se7toXWR9Ip3BRRNPBZ9gBs9GoJWGFUuz
J/KMAug36UzVHwefzU4Qq1fF/e3WHRN8qSQAB8Tvxf7Yhvjt2HXwf1oJ7HCg+ARP
hD4o0Ud34x0LKX6PfWzFjg/5mqvN3Ce/YE/NOipiXWhbtZJM8S0Y2MSThldl5j0/
iqBs+HEDjjHG7fU8QHDYHJMljgPX9FDEskrGGHVZfJwq4wC8Nh83ITK+hQ+icZcL
YE7fybXozgXZt/IfpynNf7K9rgqoJOqPcj/9NCaMAI2WKHs7LxSK0GbhlPI343dG
fMkAas3ezHvceJuxxnVrRRApFQRLkq5YqObUq2kAaIlmSt6lZD6idficopta16Pf
wXAPXF+phW7KD/pbgfgcv87Cp6XyykyL73w6yNP3gclPSjUvF2S2KDftyMilJuZ0
8tBPk+gE6nUBMINLGvCns3dKpdmit6KvdOkExiLi7mvRUDYJhve8CEJL5HkHuVcm
art9p5yk1Kps9n0rF8NuGEKBcDoEvPBExN1UH5BPmlEqjBLqJ5ukbXG6O0qYKna1
HC7mRyeiK4JnTejHVJL/gA/CbYIGNS2fSd5nb5R5se5vE11hIvjHtA3bph0+/nO4
2xMAJvYgDYMjpJkJWzAoCeenGQDsCRmdhilNSb/I8a9fzYBY/0ZdZrYRFY6+E1xQ
G5piXh6ekR86Fni9WcgTCTvInJRSBLyLYVq2VZF7vGva9KRHNgnRK8JwIVCbtm1N
E5a45yDl3OAH82gO9MXtQ3ufvnTRHAP0tHPNg+v5jC9TM2jQ3rfdts3RGe7U1azg
+eIH+cGDKXIJPj8XTmNxf3XoBKHWHfZNyQHdzL0pUVzYVYUn+hVlbbotyvb9bP7P
zo7NJqR2vFu+OfI5vUkxtrcj7mIevbCXapP4VZRd69JBaAFJiOA5fpr3MXu+H37Q
GEijX2+X+UqN7dzeewfB81pqA7f7q29Hqsoc4qMpb1WgKHXLaSdOHqM33lV3SFZw
fP1hp56QcMpS4WR4g3PL/ri7MVMcAF2+Jlled+0IxLJFO2bJ0njWYHu9OKd3rZL3
09Fy8Ja+fBT1U/ZNS/Y8FTYbETXEhS46n/xbqVPODtUUAn1tdTJLUEz+iw+b4xoX
KcSyQ4hzt39jBkN9CGcKQ66zySDAnRmriwpa6t5ieRMTKAeVDYz1tZR6n4jqwWaq
t9x6Ll5esrZVDXKTIUDr/9Qm1ZnxFS/LjP6Ld6/moEHuJgvDi7MWkDLEWpYlAFLh
VjAwAgadq/cFOtY1KG2sTYPKcZu85rmtWj1jX0QQItrwtOx4IiGuESW/Yjorpjib
Rt5iPK+sQxaBJzVVr2ioZlD1YRxrHzOuPvDGZVcoRDUPWytmCjwl0K0HcsyoybrP
eLkvdnaSFaldCZX6hv6TCww6mk7foPVEg1lj2Uj4qKbrCMhqW5y/bYFe0wcqLnXV
r6x26ZsvU12b7IRkIbZvFo3+vTnmvSlPPrX9mGedWqTJc96+byj1FL88vqjMVUAi
RQKrSTjTBvtIbZ9nH0DYUYxX2wvhkcZtHqoIt/aXQjb1mmYFxhgA5PFbZ2LB19AU
TC+HQh7louCILMFxCx1PVLsQAEUXsK/HJBPda+7Vb0XJS0X5jq+oP4ccIgbDbOiS
r8+oSlzD6uy4LZOLRLI6hkfA29MNemUj+kVRCD3HQkUAXwLk4qogT53+9jCZCMCW
sebFm4I/xr9x6MLCj0aP7aboo8Kt6LESUA6AA/lfWZHy5x52PoKzYsi3i3jsTLAa
1Vx3qZ0pa2iNUkNHKbxj6mCsc5nBDaTQwwczp0qEh9D1Hde9M2tnZHBMyOUCeAP+
UiXlQOvae8badCYpeOBtUfGfG++p4e8JJdmdLiLjsY7y+TzTy1KSLIEccJ680GJx
UFp2DqLra4wtJevPzrqzTKj3XkYoFt8zsTLNTS7KM264zAUKQX/yHb7efK1HGqV7
tvPaLqiw4AwHwGw2LiUWIzIC0AYIUMaNFBzQXjBvCZBnaTaxq+YXvTfYhJMIP5mC
tb/07Dp4+dBee6diTOJQiTQXF5uD2VnpNlgZTn91F+YpmRMcy2NtL427SfFrjgvI
kALBkp0f9xxo7wPVCjzU8g9zLTQ1PB3yogqF0U0nMWXgMLpgQcWmyhCsZbqTmZ5N
xDDL+JHaRmH3Rbq2MUvqVTo9b9gW9qidQXf8zU1/mfk6dcLIlWr+kHsDXanRNtR1
+jD8+PMoCsJW7kSkV12EuUbKHIRY1IuJwpDhtoYH6AaHEEaAJ06h8TfhL2ULSdsd
9HSTxmsE7WZJLP4udKCN/C44NeZspIomshFscJTxdidBsQBG/PtTySrXyocUm6fb
hs5KGIrS+jtT/zJ5gJYxr4zH1M0sHtqFKvUKDbW1QbCInYOFUHaS0Hc/wxjq6J+S
DIFAbTTash4LQ+q/BrSpFFNuU4U8mOJ6s7J+SSrR66yKjAAwzfCqv70rETu6CW7f
xrZG0zWMkuOUGLeYYl/om3lq9gQ8uC/A5npQV+OU+tKhLzq+ma3tHJLapoQKNTLp
72WWRQ4FSyOf+jw/NBWkzwRpFB4VaCmxXGGSFSiT7k+mrRXMfYAUSkloxdXB2P/Y
2vctJyZz0h998SsBiGpxm75FMQeVN5u+TvOTFlE/hiOdF4I2rKt2Ou+m48fs6qU8
zgCTlLkeKimAmZCvh0kJ57BX94DC8akAlCxyjGa6YB9O/DZMFRx5Ga7Xki014Fcy
ivWuddSuQZBjqX2oY7nEvCXVRpWhZxXkSBqhn+N8bjsHkJ+8Hh1eBEneMT++kziA
F/3uj5PGb0sj1TK6pZK/mQqYq6c4F6dfAoDpZgACGQHC5M80LqLxqE+8kapvKUv3
1RbYGxGr+wwI558JIQ2UM5V/E6hwZMy+7WfM1xhFK/DG9Mk/9m8LxtojnKB3HBj7
fT1Nfg+KvfBF+zlqZPHYOJcNtnm/Ul9SHXtiRbRrRamEsVbFiJZ0rhsLlbkvgVwz
rQK3psLBVTkZrta01gJ+F0tolMMOLEeV/cYDY90j+B/tovHG+eC+qVNIpmIv6HEx
XqyNIbtbmYxdvIhhAU2G3I2IljW2zUXPT9ZTGUzwaqcIV7CTvso8kkNbDtFunjHr
f3ce423k3d0RZmk7yGZlM3n67ZKNkitAzwxBldpQJlxvXn9sZ1rty+eiVvlbjsNF
AM+HK3NggakA4bL+TKj3aFXvYceMi9MitlKZCuO7ApsYCQgkvruw4JAQCa27jPCo
7b85bREdFttw01oGzfvNlyKsrY6fOvTgvN1dbGbCOSt+3EJczwovwHKoV1VkRKRC
KnyG1PIqU1tIkRYHCCqcOGx4ajAcDsBo2SlyIinIIKuzPzjVgBdCbaA3KYRwPCBR
kyS3E+IseQh1epFTAX6p1hqqfyStCOnTfaiMxbym/LhU0+bU4MafVtcGspEe4qEv
QsOO80N67ZnYDohx+CXQZDf3HzEhM6iiLWyjDZgUvvwmjxtSKsY9ox+WbZRhXwcE
QKY095AOarqwQ6mSp2TdRC8CHwt0J4uh9Iu1GwOrMeFOhe4ZyTP5sTn2PbzB88TA
4tdtsoN8Aj4o2wQ51nVYuD3LzZSPTSmPiYzy02eY9DyzWH/QbqVLB6+jwWPAIFWn
53hLdr0wDVBpRS/eV/0TqNP8KMhZsIg05PKQY9Aw/GV62GUhPrxZ2E/ocsSqesdT
CQ+SYZ+9VzSLuC/24kuBxVF0TGQZwvWb0Ai9qsGcVI/nhXggEJomsgfFINAT9A74
vtUsL5d8PQX9mWc5hto0Uw592NJiTGcIKdfqiLWY2MsAw3789J3DZKWj7vBei4VY
aUum0zfvFLHQfIx2rWlx785GRRUKV7+Tfv6IGzTQA7ycaRnaevR3/MERx6TGvZsI
Kt3S0tcWMjX5tMETO8rIMWku1vG+CfJzkhs0Jp/YUOylCUghGzxp5a5ON+nVo/+i
yNovpvN46HfxpczmP9bSZLphYSeRYsoHHEI0Navc6qyEEsaoGh+37qPTmYtwiz68
Eq7IrDFDsrtquCxF1dCfzrpufFYOwu2/CIq+FbZMpDuYoLya2fN22nwwIBPHkzom
zXlr6HklXJtRHAFohFWXPibLuu2LBhxnUSTNUWy/LQyP5diSvxsjJrBI6JhLc0/s
J5Q1WBr1HrYvcFPJpdogquZITV5rN7uhARvZ/vFWeEyVl7Wy825kaxYyJ5OKj23H
4AvbhLLC2g5kx1R4SQ1K1B2EfbS8uajy9gh2Z2lEhVJD9u7vJOJZaub9DWdak3I4
8hOjVmw2Y9ZZBn+v1X6Bk6f4YOhQcLzQeJGSi7V1uEOCmX2U5viEtPgkCN3lJvQQ
NnrsPJt6rOa0roN2HFZLcqN8DLrC0ZexfpolKto1x1pvsawpm/GsnGkb5xPALjTC
+icpd9hSb7mzQWJdX+Tnk7aGUzG/w1TDmaht6611gUhBtlOpgWllRD87Aloc880Y
/eVgHKoS9xvroIscH7msEdtbNNTW2NXZ3K8zg1gt/TUvbCXPlhFaH2nBw4ob7T4C
Emb1/7smRfOI8pr2uYX6Xi0uYXboRK4Rdex7fh4hAR0L+yYsfUF8IaNw/YOn9eaj
usZwNGDhbolYbBfpZ2pL7Qdkg4lMNQxD9+hwj0ZTxQWRkgUA0mh+XR8F08HuXCec
XmAPtzFW+lTfx9c6eT1G8SqQ2iMLF+I0VYTdq9quwO4eF3k/4uSkXmT8WlyfiLGL
Z+HM0x+8HqRSfE+krQpIEl8Jy6ZYcYQfMRhW9TvTnbiRyXzz+8TqlsmIWcj5IHqK
jhJV8ZWv+N/TkcjwRms57+6RsCuqCgikWrMtlLQiOqYPddUlFZNsfGgqqQjnBUa4
1LpQDouS45zHDzx4ZHxSl69xDahJSm5ooa+2/5Fzqx7NdD79p/qFGFOJ0+wyvTPq
LYnxkEfMz6Mx9fdkxXCjqdq09V7DyO1jqw6T0ziFVKGBrzDgLa51WYGf5Uk+mvII
8+wRtDldjiiE4okmQA2MIe+z3ifd8iY8LjigX0NMV/w9ysG+DLUWIiFEZZF0y2X4
zixR1VK2hBwIt+JgB7RxvtItMbgJLAbD9W2Q5aWszAR5VCzt/Tkf6+BYX7niIDwN
AsdeqJovWRw4gUz1GhtS273dk5Xlxmv1Oc/wOr5jp1uK3NgqZ1R7+aBqMDeXqlbg
g6iMf4ufRcnxrH2f4tL64qbaBZ5gV0VmNSltvPnGRvF5SsJWL9DzGva7llKe/OIw
PL6iG85Nqj0FGEBoXGy+zIkI9oDPQ1nYDCrLpAPgfidkD5PYPbHB7RrTCEUaa2TS
JXT2jZtVsUFb1ksb7Ztf9Oyg6K/pLtyL4JLKG+dTDlQH88KcuTKaEU5ZSBPnVBOv
VLR2qwJLNvDYN/GPYOumeyowl1pyqxMZ/y8gTLMbKm1IzbYsm9lSziw8t2WBpJJV
RgqXsWQLBGKxXNFABXAB4vWxsaNz+0uhx8ZqjgMo0azAsGhpy+CAvya6gLx8I3jA
J/j/IWGVuabTH+hJ7gKbkmyOuxAAvCPdHnfci2KslBoIz/jQrJT2frTEjexRBcds
d8hrnC9uwKbuveizxT4MdcMlhhY/6b9Sib/X7WP6NwYlflBRTANd3hSLNj9PariO
ilUUAo2ZtxTPv/XBfSSPPUOmIBonRc4XFlc/NUHtSdpE2T871GY6osOaxqPehvkM
krCw1AP+amHj6pxhdLKzDSrc32SV34/MbPjwSll/G8IjUarygdVyLx+ldXvu6vBT
3j5kPwK22QN4Mxi1h6AxBR0Sv3zOaATfd3iQVvyqs79LOpu2kOZD28pbLkiwlEfw
x5eC2WA747JXP6oZgbURjqNdz3iurz2nVup46/rQzcn82QYiWKpFaSGwsOHNcMdg
j/VuegygrvcEiPaHqk2tjqV2i+Wn1aC9uNQI9os1+HGhKVibxZlt8832RPTQBzLi
lqCZBLfpCkgTH79E0WuPc/1BJQ98y++9uwRmdk3/HTMFS8g0vn1rvb2/yR0+7EVp
eOxWi0DwpqJAEPtgwym886sszMKyyphZ0PMvCHCF/+Y4grEvR03CZ7GjvubOwlcH
WzXui441XzDYLY1zp45ttDckijLMF03gcbP/Bve07tJajuCPOr7U5u3olri1PUoG
mmUvQYS1/jykQGnrxw1YRZk6vNyGJ/Gw0tWPXVxSTZsYTOQS8RchpOsI0tawlNOx
U1w80X0h7tlAHZgHDFimvQHH/WngCA2jqmu7NzFXpao5NhQWikaC7wH9wrORC/f1
adV69IYxOvaC++ugCzAxHChh92Vx/xoWuXgo6YOk15t13IbtYAuj0x5QRNihJ0lL
qUkIhDjL8a2bXY7Ew3kCLxzI1XSjxTHRAAaFsjqkS45taPfcTdf4qMf0AgrMd3GV
6jKocS4OIKCDWaKs1qSCb5sZZzBrF8RQAIOdOBzasjAoz4VFS4uejmTZxyfpB5VJ
g1Nfkta9aOvam4wW5AM+kqQnf10K+XqXIFTOwgGe8J7VsDIR2eFlxkkXKaNMFuJd
uMWeavCflZs4V7Yw89Mf+rA9a6QAZ6lW1aurZZ7aD4tviDuAsmbqkmWNFsFierMe
0zchDysTCPM0vd+yEpZlnfSIAnc/tHIyrfQf6cKWuc2uhcYJAaOx/UHNG0E4Hv1s
/KMnFzDrhcVCsRtAyMs8QSD8WRh0GZllT/wictyFX3nPaqZIvs8VzzlMiHjQwWSv
kGkQK2WrQv6R9+XVC+gDw10RAzZF6xkphH4C73XQhl8qebhosUFIsCLpD4zYDak4
przHmq/X3hxDijAmaf9mPTjKJlwQztIp8i2Hyl/4oHTRNXHLXKOpWOSwHlIukYV7
x6oEvzHdRx1YX/zUyQeVX8F+41c68HrK5aU3Dx+AIIeGkwA+y2WLqC5W6mDfdEk6
SjrqWvLVA4Umi3pyJBf9MvbFVvobCbtMMo9lxZpwi+gv8RycXU1jZRpTSIEmkgj9
Zi1i+zMPQRP4SfCgNn4gQfA/OOy3CZov2BaUSEGIhgs1x1FgcfvP+QRVmON3zItG
IzhK3AWbS+w7FbnTXI2gC+u/WDbEU//kwYnJY8CM8IHmsxib9F2dJ1cl2fn74nj0
PglaQfKQ9622T8vVj7WSN3K322kKGnPncLJhSGW8fG6med6f2IXrmyIfGmOAGGQP
t2uNvKkJFyVMdqs6RImTkP26e9zPDtTahm6ss8gKYeR2QwhieiMFr3IR3ZTRjUfM
L0e+4x8XbeEYXbWDD50GMiakaX860e+G46Taum1+BEzmytHtw9bDpDez1kXdubi1
XfhPVfcTvN4CrDU47/e+4tGegC136ntCFvPVunEvXgN4iFky9l8dWb8U4ytJ/931
PPsoEi/Z0RUp60IYJjPuw+me4Bw8OCcntS3I4/w25pYwJIHSowRLVvRZnG6gbnsX
RD8cNiJcAq9PUbnAbVbioMSz5XMKaw/WtARR9y7P3b75irjrPDLjqLFcx8sNLJ5U
K98YYfAb1bi0tGB8H1VgjVoECpPAtGCm+9EbHAWK5WJhPjGtHG7Mi4mIwnhr97Dh
AYpQsSbSG+ep5AXKofByvG7RgRpk/1YvsJIE10GEnXh8jcGXYEjkKsmp0jXub8C1
vxTFCoZdr26d97zqdmDu1Z0OtMAE92FlS6rMTNbPgKYEycFIEp1XPNf1Rr1cYYVA
TPTaCdGLoXe4gkD7woAOLh9sEDFQRnAftMCArBphmdt2HO1vNqb52QhKqDXzqNqh
caed7MDyyIPQVRUaUlqLqH8YLW5oOIaeXJ/E+E4bac/QQQvj/Q2pYF4x15YpHEAB
FThp2BEtLwIq8kJ9D4renE68YVmaueKccErRupldzvNPtW44AXodkpcZU4TBWG/P
uc0eHwJGWZhOpg4ZT/mINBSbhqHa7rXrwRH0J4gRJ5a9zBofQz2HsoOno07XorJ1
PLXK81KYmCREaYu+v04UykOgbNQ8z8tbkR8uOkO9GdOJAO6BIu+AX4QmUjHyldQL
FR+k7vZ13EpNQsaUQcHc3OtBMcFEIgFkB9UFcbVIfEOOtCJ/emXGz/IXkbDtA6DH
viV34jtASRog3JpJad+qFEBU271BeXald0TZFrq6POpgrGNkkdSqt8mTBgY00pEE
Lg1vwRyuamkGzEZmLLb3icfub/Nz2B2SBJp8h8iqtvNyqeHzw7K+4WJZz9DYqHIk
oleSXEr0t/K50XAhsSFo4jYvhM4Uz1VtITe4MvCr/ymVJD+D5DRs2JHas62bx1bY
pvfP5RnlTAnKoLxJvSE87hU2y4EHSCDHsH0tukbR32CvcbCK9H+1ejFwXnPzj8ql
6Qw80PZqIRLXlgFahhR+mg7+HZAo6z8+2FK/ypeoNQmplto5fHhz5QEwlsASW3NK
4V0tw7W4r0Akzf78Ua7ueBh7+Vgy4dPqfitP7jBI/XopyEkE/DY0uOYlrqop+B+t
TbULHAlcGYQohtv0IvJZXuZMkpVnZD4jriYHPC58pCgRzdlwZ+mtU4+prFh11uHT
auoMSBQr6ggDBrH9nb0UGEi94rIxnma7nNunqpcUG05l9zO48iopxkidLtFHEbuU
tndFw42BA9mNxF0SIIXlzWCxHtFbsk2f5bC6vCKrU/4g8oVnrN6e3A2MMhJqdyTF
cvDTnfStYKIjxqThkc+H7JtMNkdf+w4GSTb69yfsfUSdM82UwJehdQMpQgdBc/Tp
ROI+yVkZtEQuyQk5ZTs2oPhUylsTWo5TnC22x+DIfuIXPM0lc9Q/a9vKI4k/qqX2
CnmgQpXG/IN7roC0MaPLUvqs9cxXO8vZkzcZhudPoD9yf5pebxQXsJpFd+RI65wS
YixVux8QEkPzvIKvL/aAlruplQ3J8vJeSHzrXpIbc7Gw1fXBOitB+Kcexiiame52
QLXXQIQDzEpy6shMjiYzN26CIn8geVYLlhHRSmo9YsvBOz1h0G8AQf6MniQ1WdCa
sGliWmuSdlxkMjzAlgWZs2OhLPwXz3gJegAtHcC4uOdKL2BtiA70CMxVhvZ1yw9+
33epY+lR5knoUy8YSeiqYZIlG5lOOm3x7lD60nUHBTK3Vp/nRj0UBz8nn1HCHsg3
vyZNxes/ZyHo4PZcN14Onao/E+V+MKatV+d4F1rt8sSq6iv+u/EZO92ti1Ezzdrh
X2B5TUhiTGRUFGLVrjmJmR/d922QHwRr0IUArzcOVfQ0yfaFLHOpCYjoqc+d8WWx
A+zfvKP+KrAGD/zYqa286ab3w7SPHOaGxN9HhTC+LfhmRbPPwi34VrBCplNZd/uR
GJCbE+ghz1zbaQa9mgcBP5g/ACpwNR+qkxVv/SskWclX1wmsMT1hn8nvcWQ5MC0D
iONTl+B0rlaFQOL49lwn2+8+ZWJQ8v0dbcfxz+z1PfW9U52qrnRD+5IVQgFPv/gS
5BrUT/nye3oChhrOHcBN1Z74p8fN//G4d6BhZ655iK8rpiBSNXbwA++gZNhIpAJF
hP0tVEj0zkE5kBwQqHlQUjwFCiMITWxK9qfew8mIwVSwL2cqZ9GosO3PTFbdU2WP
cbNqH3JFpkPik+/gP4mEoGCQK3mpAZptBZSBQh4ra4Ff04UAlvCEpzF0PhNiJUuj
27DM4vuAKdcPUs4blhKiz+pPpKIm+5s3aPizaRVE/u68XQEhm8SljFf8rPgsPj0Q
0KbdhKoeucLqWdQFnjyvj6edvizBwHORKAg3f0ljYN7FzNq85JyPv//mWBMA2f2R
OEHFjAEdttZTwjekHTZjG0ffnYZDvQyuGfCXQl6fxE7D5mwFEXOeRs//3o0cRg/Y
FXQZcScCgadXGTZIN8QdV3A2tyo5GhhwHJdopglDSy/JDoVUW8VnTLR/duiiRF3d
imX9T1FWOWGNAcwILSE6gmbqwiR/Wp1Tfy2Q8B+fj81FZSOEWATNfp/if2ypdLSs
AQJP9JQ5FGQ51YnnRwVXC77ZVIW2bfjd7rym+T6KwE+5H2DxzK6XP+/EalrKj4F6
bMlh+8Jnhk+z/sHrVfvkU3mGppA8MiU3b+uSkKwZxUNaej15dbfUjgURx843kfAp
0oaSBmmkqo4c6ccNuC8Mby1fbm0N4Du2YH9JJE6TIS0PKJk8a/ZRvl6PG8Ln5UpN
Z5APYQlviN/d1nDrSo2OIqzbHpfbjRs9Fl4kz9xJtqzZSzZa4RTCzDbpcr5LwuoZ
pJZPboYfZnGnlabiDJhD/HQZNAQbFwV/gx/ftVJa6L2JSE/UZ6Ufg00oydTzcHSa
PX8W7kCyttUkwAWOdMC5QWsAOD/pZVusMXVyXyh1VDaJ0cJ6O1txiPNQv8URA3Zx
uKM22e/7RC9EXF+Sp+4ioL8BmfxUO9h3fYGaXqVTf8ET3qRfpVeVDPr0b1K6Aykr
z7NmHqPHN24vuAZfBGWy0MtlE7EMPZKP8VUs3VTQIFVWATaH7bB9iTtaWT8vgen+
u7ffyxJhjBJ6vUBdXO97Glzfi8wbgzU0NHPagD10c+FZ9tbhhH31mLcGJq7Vky21
P0Pr/o3TnrX4pJ7pk9Qy1h7bReL3HyUDH7iV67RvkMxcUV2TiycGGAQURvOk2Sz5
Vk5npnNdwKqfYK8NShOYBwXYV8foLDAG25sjqmbrKoPR/L/yRnvKhpMvoKXy4u2r
O1MazvhrBZpgILgUHM/vHNokeWYI0CL1XFbrFSOudldS/Fw24BfCwZnIsyg/vimL
QGPAAplOlko8XkbLfuT3kjBlJgKcUJx4mzCRUpAZ39o10StxRMEG0eUvR7wALTU8
jOCPkr32Heeq3n/r5YP7XndVbffw5zmuOPhQJEPH4ZWnJCJdTGCyCdWmprIITYx8
cHkq9YCBel7enMhWMY7/gNIdYlFuns0Dadpl6UBiPPPtW+GyYKmxdJUGjxlZ6WMJ
JKQNXOL9Y7KpBbf07qFAxr7jOhsdK1eSalW34wNs3dm6qrIqUALDfCrJnPurP3wf
wKnbbUXnnvYj2P5VawSFY3h5BJkLP2PlZJampyAkfmi96T30+zSzdrS9CG+0/vaj
DmUUTkemk3vae9EMUpFPE3krV1NA8bgCU5d0PWsbVdOHCDZAc2kSOTVGO8wWITaI
I2ZQ+bMaCnHxtOl6V4QTtKiqUGDCGD+JGYeO1lf1DP298oPkGGB54FWGpw1QQ3eC
3N0woqD7mByRRxr8FqsUjA/uQtXkoZ2oQhpXZ6FaNzUosLT3FwzXNkRTvw23plea
dJwotTqlsgRfqZD2Bn0bBCFyopNJRQjg1W2+zErGzPjLNWq93nDMkKNJf14MLx6t
Dw4k78a3H0b1Ifn5FkxdW+cRcGdyZhXugTaxbjM7wklg+RutnON2heMrRMc15KI6
eYvQzRpD0xEI1SZTznMbRmeOj50RLLIvbFryzDP2aX/Hu+AUcO+bntR/4YYm34GP
t7c8KmthskaC4vmKEg+EJQd7hZzGLcrXZVeqLkW3xSLvNc8V8rIbRBv/qfjXauul
w/oJpuxkbZuODom/mwXJqU9S+TwvzyFrXOItw+BDgct71NN+JE2ShgxlZGm6wr/T
eAdhvN6iO9uDxdWiUW3DzWXCQcQFXZQ9KBPB9UFHhNhtJByfcqiPty7CWS8gKt7U
/IOrQz0GM4e5WoVjRdETGCaQdjDlVEzAKM3XN0YbGJsJYeyjlPNPMtztCOV7wtHF
GjGOq20eKNYYJctpomKRTyhL8Avvk9q1Id0Qe+mKkPYk+cxcY1W5CgsVHMRnmWIs
y0wlHQ8tbTh3pkNvhaagodGVB0IPQJNmUzJZanoQDKVDJfjzJvydVe9AFr5s749y
OvJ4H7mazVTUOXe9+agYSL8XUKJJddcN8IiU5C7nsleK4LMERh8U/YITSRKIAr/x
MQBmio8HDfhQejNlu7HbQsJrkVoEDpG8MQ1TqCrfiope9LXfYlpt0yMcka7AXjMm
cR6ApBK2OHqLil6Urcbix0TMKeSplpwhLS825/bLg6A0MwE4gGf1NE8aqvIBFnhl
TZZR9DGIytk0Z7YAUaj8gnA0j68irBMHjnGghs3ifyc8gqVDOjrFhgd07EBKDPcI
YNgEZ3rxGoe95CnU7lkv+ZJddHI+VvKPxfqv5cevJPd8VCkl1hsNmqPtmImvMsyZ
MQhA2X4dmUrDCI39i/L2o0dwOGAMeig0iHAnzn5UbKPeVBd5Hsv6ZEGquFrhQY7e
DfHgAIUbgViRjJ70lFtnMR3vaAgAE3hoy32HES9frAA37qOOO2ROmHmjOJ+T587M
riPxO9X32AEEhkg/lUy6EnDjztcAoZuuXwxaVd9p996tC0Zc9Ik/ybWy3qGJNl+z
PYEihEHcYVU4n41DcZolz+U2dUwplsN0ZAl8/fe7FezvOd8cCphddV/Je4A79aCY
9myF9lRyXmTisRhYO+WRYt8H1c9/jDIuEkpNLYS7fN/bKG6/DFQNzgTywUgr4UdG
oxSClXqtfafu8aXovlNSci7rnhlscvMOtyWitS48wtVY+CW18g6XtryVYPlwDMe5
fCFlGdiv2E9T76qTdz7O3DKHUs2RqZlPT3nQ553kpeJ33D+jNkAYBK41Qc01J/az
In4OYKb1zhTicAq9RuHsQGVQp60l6U3CVqKJdkQ/ZkWVxWiR7MDx/fkwy/Yy7d+n
PD+KOXb0GtzYgybLnIPGw2aaDXq0LoAGCnWe56uNxoZnhk6rJ1TJbduaRG9+iFbW
sCo4a52tCLaLe5U5gjUhady/kXHGuHhfEVTw+8L+DuG+LcI31XlNcOlwlXVF0VaY
KAfy2FnJ0wKUrkVIRzyyR5OQ7UwHGx1Gge11VleX1TQMEd0fXoUPltDHwPJJgKSl
jS7XDxoFr9aApqs+s4gJJG9vMwKzsUmNb0GuvWtujiKLTubirza/hO2W8U9X9QHX
b7HFKLcMkwoE/V28AewLg7Vi0khBPw0SUHJS8zH7A5NdGmqQaosCw89z/XBbwqBw
4cEM5LhEWg8c7c5ODmdiEizeBRGDi4BZTDALSo4WMaPp1bcyRkMcDnZEv6fAWFBv
rtg9m65HVvuOaSkuMEE04vfCRoV6tlRuTp1WP199vrdUJ2e52lihknzrJzYCvSTR
LnL4+Opab14q220VzooXp4Cgs7bOUcft0WHfwme1sdjxF0JiINhffpobx/3Pz2Po
iC+4pWzr7M7I+VY1/f+yso4o3Vlx32DGBPWoP0DMqw5iWRHPGDUD6D/GVagdNlQk
9IJSY6OiZnnjJo9tFilYiAvwWGnTmNYdlyYxi9dIRvMOXaden4DWhekD7gpVk9na
A1Sr0UBYuXf0EIrVYZUIsH+vmVN1P3L4I2NNtscrnULO93PXsbV1Ur/ZqtNk/v9H
nZ7E2IXfJnpLkPt/dM1SO7IpDVRNp4d2pEiwNckJqlpd7tE6uyUBpDVbDC+lYkZR
ZPCd9sC3X8S0FlAP/rdb1RHic/VNyu/xa7GiOi13bLKJBojOJGQxs/m+69938bMm
v1jppCDjftz4Sohdv/r3gwJw7wiKWZjy+7VJ2y25g+iO776BhnAwKndUECaTGnhp
i7vhxEXTEs4+lrUBngGKcnomIefwt3422N6pYcSHrvgXpJ9xiVdJvKUY2csar9of
3k84KNddHRbwmxSVaAr2Avq6E4u9p8T6Ao0PglpdH7oJQS2LgwX+NsHrjSfTvlIX
cfvO/60mdhlsAn0VCQ4m7WMVEVvT6nDKkHMg9VnmE3QjF8IXroIGVdIGyP5p8e17
CP+UqVd//lEAmMMedWqcfSmc8/f+w6ZRKDGpAP5qMQaqqB/hU0jZYbO9EXjt+p+2
NIaa6OVwgmUdWLuiiaQEh2hKeiqPyA57LpR9Qw/bON98W3E55UL5yaW9/qhKHPUB
Ape7g1VMEp9WqMugH46qIIaJN/O/WxMvJozmKW6niPQWwbXrDaUvth2qJmIFQp39
pGNuEw/S1HQt/flBpkQfmqKjul/YTOCgzB88Sn/VbEPjIKL+wDjs10dIndSbmB+T
BwTVA3b3G81n+uOGTB+cAw7xg6oGBwOrIx98RonUFq9wde+RSOgLSpQXDpO0sg8K
Qru0bI+o1H/8OMTki3iZqr09tfQ6h31Q7Cn8PqSpnmIJKwDZD/gMAZDCFYOyUQrc
cm3AK5TtWWU/cU68kNfHcA045Wi9jU99yW1W6Ilh5dvQvH+QpgxwFVF3Aibqz1GU
Sg4w+W3bwOTJrpaGWZHMDH5CC41LVkkz+THWL9TFrSFSMNKQ+bBpxY6qMuFm7po6
EMcceCCcCssgCt6QEZ8LT7E6ACbb1vjZFGpAx/p6q5NMGBYQLc0vgLkEv3ltwia6
6ZLWBy27upmMXBKFsEUthwpcao1qUHQjHqaT4AUfJvGeT5z8/G3GIeOSDWo5WuU1
XhXJQ9Hr2NYlbP/Iw6Q7/DKVbY1BmrIITKbysG2SM/tdplnjdXxv9lUgPlUsjcrr
iZmPKr2kYxIa5d0cPYMtG7i9b7uPfSeQfyov3tkz/kbhBRqR/W68gS5yYq2jEcC9
iLOzYqvK512O5NK2Inn+JPU0MPJyiRNpPZgLJaqW9RU6PKAgUlemwpggPzSV8sIS
kPDyEAg8JIXfRvYn/zhQkrkRVXmYCL6vXHX/Rwka7Ft9QaH8VNxe8F4VfXaJJaiQ
LYQBBPNX1BeEzcayfL56XXPA8b1hKESF+lns13Ih54xIhx2+X6WWf+B63sooUSEk
1epcL4+9nybGA8WAW7//iXNFKm6YM8fDlcq+B7uCMCT8+nFycXXemM6tyx2hJrCS
Sq6HuGKOupoLxv1YVkeS5dgZ4sQIv569HiPlbzbmPtz+OG+/IU+g0/LKxAMNRaX3
KZjePDLGFJIvDB1OXx+owcmBhdu1gd+dgG6gYKF695mQYHh3FMxUf/oKA1OoqQSL
DpbHtz2+YwMa2vOxEWXAsYpAF6ihEyJE6KQpWzGWUqbfzbhvtec6IvsWcqVeCV4C
lWnJ2bVbxUi+51tNghwMj1hcvBuMgCrXgr6EEqtKtCh5VmcF5GSVAQOolzoUMER8
qgemuur5KPmhmHoeZ26b+ETNZKQ1qk3JSXPiwdRgqInUbL4NbLQOh+QQQxGErPGz
gV4rNOE+o59+M/prI3/Q+sfgQdOUdIRDBNngf1PUwAZkiR3lgwZyucF1aVk+kRf4
9CVZbHF0m59KidnPZaHlaa+GE1/Ki9HkTPRvxPbbv91spP/snf3rKhhAZ2zTyhRM
V5b5b2/T+bA601cciudg0moUb6EX21ypplve/Lv5KNjrYKuQs0j+Uizg8ou84H1K
P5OCcq69abzNTZGqOHA4fQnIbrxVY1Q92putwv4gyPyVvSpet8oGoI4vhLDzGMzb
T8xvP1f2Eq6QPfNjL8svRxOfwHnOhJNtri2liQOk1bvKNY3AUGG37x7yFv3tMRn/
8hmIHveJeLuOsMw1Kv3IZAWdaADeFrfYk3uelnfaMsy+sTvAbob+b6NBtoKIYOja
aT5+PD4k6Lb7ZyZA31Q0oNyTYYgSop2csXCnwuQO6+nKYmfvcnu6itJk/Vs0Nz8P
i7t9K1jvzAHLsjOvo4sLGp+KXgVEOr8k6GdeA6vZGSC8RBqA4LfDatXvpagxX9PT
4o2svRTWzx8ubj7vQHPTn57V1C30Wb9wEHr5V7k8BbmTk2LTmC36j+iZxUZbE8U4
LwaaSE/Bo5Wr+IzJbx/q54gedkdfM++xF0eRMi32I08UmRPJVoUT3mnizBIF2jDz
xfS0WuMd0jP+4XUgxLbt3FEQrYzhwo9A9rRJz/NAws64xJPrMTPWUTMzSRNCGkT8
f0ugfEoRuzxXtNJ7n/8lc+URx5uQ4YCjJdQKWQE+85OdBovXGJxiu9qH3NKEkCTV
TO/W4++QDx/OG9fcOwDnb0065VtjbjFib8tT0cNKav/wimKLaanMm9nPAingqUDJ
QGk855X/0hJf4wppWg3465knegbdetQCLiwFf2izbycOND/Pr0O8my6VIEcCKHu9
BHTkQVh6hjuXRn+2QarjpMFjMRSQ3o519p210n/badmU4NRLMSAAO1CsFkFOKcV/
TmeQQQwzOeq0guVxowLtOQ58DgDNGtV3Qunuu2c0aJX+WXREAAnQcgbcJbp2FAm0
2r67r0DndoUeJa8S1Hq/biZrP7kZ2mOfA/u/Yg75NN0MwtegXIrNSIrIRgmv8FhC
FCWaGLFCb8Yn8pxE2/7nxtLdrcdfpTuBIGBl2doHV19V6v+Sro+aU8EI5/gVY2iY
w/IkjVLqiOMR/sxL31dJ/duhmsPTTx5xNTzrivSpLa/e+vc3clKf4wcrwllLx0On
vROAr2uajc3ZIejtDiHYRXihkbWLwiNbrAug7lM6e47e1tM10xBH9oQMwNCihSFN
GDVdFQXa6KCswHtGfxIrl7mEpuDPi17P/o6MrusJ+TTZC6rjyR0ti+AItbNDL9Ok
R8RSP9NtAaSiodRYHntDzZC2QkVIPASyyT56jERx1odJ85BdCJlJKo08apslXgTf
NAqYl7DJ+RJ8SisZ+MYiGLCn6MzUSLfHGQQvO2ynj0ivtRYmOOlwDd4C7cBpY37j
sxZAq21OEgxLHUM98Tsg5lOHvY20ogQzvTaT4Pdo52zGX7qvsylxK9jExmS92QuC
OatHppss8shjX97L8X70zBF/1WMBRIJJBsP7LZ+0WkXDlRCVjJKFQBp/7pQSWNuc
X7eWTB/dVF06HyZMp/PxJyDAekhTCbEuB1J6n9BmrBnoGiB32wDTVDnjZJ1AEsn+
TrMRU9/Fybk/A+ythb/6oPE4RKWq4OKmrpJvRFbThDqQehyNvuFmQJI0jdPeP4ZL
xClZ2SRWj6S/neSaUevEgBz7ZuvC6UHNwfkB97n8yOQtOFg+dMNSo70efBIMnGoV
Di9rgX5P99AEQShEqp7RWOiMi4TGcdeIt87oM/wShdFL9nTuUrA/tkvLuI0Hp88e
6lBu7z5sslAakZzvAncvH/IKfdmWM6wCfpTAvKGP3/tyQ2rHHQMpV0GR67HKTvKV
4NePjKfE/TAjEkpT96uBIUJisWfpeYB2PC0XZtAvKdiIu/F79OHdZwMMTZUm7gOD
gUNa55T57uxHf3lhV9EoSxrHtzHD4Uuwo4Gv7tfQ56trEiLH2D1wzs0u2vDd6grH
B4lSVY3k5jVTUSu/KmAIiDLXACQXuGQRTwODrFR1CVG7hukjWAraL2pozy5XHuNp
+h1IUznSP1V6EZKZ8nBAyZfYYUsrxuUJBHFC7aTg5LdqRaI3RtqgRbgO6BiDPBT3
w+wvVbOPB0o/SL9ixKPn8/Ih7su//5aj70OtXYB+oSsIojWXXyD2RUeF9vQKACSo
Fe44PJdXhB4VJKgrjixAK5i5Ycudw5oxLAC8NK6FIYqx8mkTtXtFT/F06UIWsUP0
0VInT3to1MzSNw2POP+o8u73BU/wWvAHIdhF8ljXdYxZyt+gLjb95tctKaihXOub
UiHXpHsrLSo083OAJp/hoILn/l5BKzdod8CE63nJXUV166xOaTfIYha9JuMbqglR
HFCkQZES/crtbJ3bmoz/KjlBDEW7u8VAYKZeoVb9YOLJILXuXKoBLngu1/pRic6f
0j+6pyGHy+dCTzyeFSDsi4xuaBwUqvvV1aanb6d1SG4lEXMvlMe0v7HXIhf5jhQJ
azPDyvJgT5e/Cpni5c5mhJZBtzJBnI90DN5oBpKZzzvnIl2A3g83Zys1Bk+SQLzf
+4w9p+PnmYhRwUosQxPkEPItSDr9T/9pordBoRDvJqTPtuO5+q/LARYL/df72GyA
Xik26igLs7TjwSG6BlWy/uLS2dtpi4pdykCUTJm8CR8N/jFiUMaCnc0ITG4KZYxD
upapatMYBWWRD8vzd2q0cprx+I77IZnavYRhLUiBLIY7/PtsaQVWFsT1KcOW7vMg
GZGo/l62BTk1dKapIeluZGO1yjrcmuhNjpu2NmS+SAXQL7E33J6vr9vFAWnVwwUJ
HPhZQvljzg3thYTZvJJwEEmWu3MVBeuhwH/2dXTdbXzQg9RNY57mSBoNS4RezEon
mt0m2eBqX0lUoCJAoGi65ahrnshXZH6PkxGkNahZJO4/tZI5tPjA4mFYGLZCed6R
vKcQu1YJnu2iD/Kcahk+cxJQb96BuxIjZFcmVyuKDvrG0neMKl2yAZ5tbgymkl0G
7MeYNaWeUFDLj9vdQ1TvSFWX9jCGvEiyDqnw9MQzRUDsGJV6sT5yF6OpkGw/r/vN
j6VRna/KddKXN3on50pWDXU0ijsg8nIBHmnrYFaAYMStGElF50aBWzZQ10ssNIZ+
D8DbSqD8CzYQOCornxj1jWQSNckr2eyHsbJ/kCw2NsqNkeI2PZed8rTpyyQvt7pr
tqH3puYBbh35cfMgPeJQwqQqwfcM5aPS/R+LE2aqypJKfVWoZceG6lY8tRdwOQqn
sXA572ZG0ESXokMrnUGM8i4E9urC6wCH63bzPTkq/rjSgMJuYBo5pHwhkds/fnXQ
/nwb0qiVUgCt7PD6moBR04OGCwSizgxSVLV40RJDK1z+mQmqhcKbwyH3CDAyaod2
7xLbBXnHp2x///HBoCosGWmzbY10gUE63ZASeQXfXKZDGSHtPL/1iu9ROxD/x9MF
WDYJhGS1QNOIQKB3WjleVlUvuZedwEwI2fmbB4Z/VDUaJw9cm/I7Fynh41MBj55F
2OcL8pjnXbo3IV4fbQNHVpea+hbpD39iZpVzb/bWmIfltJgw/pnGlm8gmc41RIpk
zFFrR/srkETAR/nkfSDCFU1+mn3gUExl3YywrzsuW4MMp4L3f8ET680+BVx+XMgA
tdKak26vv5CCNvzS85ghMnOHFmyjJNsA8uBJD1tnZANNA8rmuJdFBIV/xUDUjs/6
pAcIOxaeiUAk8l231Mgw9DQmyWJWUQwDWT2qs8dN+MIjgfgtL5+lu8EH79fnKUWU
5EEjrafaGTRYGEqba0+Cnv/LZfa3AbTfT48rsBvaqIE1Vsthj0O1LWvsuQYTwYpZ
Xgh8m+K8mY/I0bZhgUXTkKuLnmP3+McigARPCIzU+4uqUBvMabvyJX0g3f9fncyB
YV+f3Wrabuno5JWAY76wGRxPMLMv/qjdI6lGrBr9VN4exrbnvKiNr35ZeZp5Oio8
+2gagVsyo8QDdPOcWUn5BqmosTnJEifZbuW1fOD0ZB97AUc9r9A6Dsb4GPjQyIcI
hPsFk2WIeELIaESOYGefy/D+qf5VUnzN35HU5sXGSSpjNrJHbb3PPeV9oLy2ZLbf
7pxt4l4lOlZkt1GEL8p9hb7+kreNHWQLD0Eq9iytwwgBtSCi6TJ31oYdRvZbHds1
BCskifEnkDIOpCQe7lbjIE5eO6yS08O9xZnvUs/dWxF3HpUE9w4MibYtFv4g57Aj
ZwIGsNu8S4zBbRaQ8GEnLm2dHt1NT5FeMkC93AO9G2uM84NrQBwziJHekoOFKg/5
nvUzkcMjqIlA8CsXRxP5Bl78CHAo4VFTHRQU7u90WyNEpJZFmkZcXAfe8uNy+0aX
GKhO9M+niS2UIZEaZqhzepDgCRUTcbYOKIX4Lts2DlZ6/pIA7AnZzPd/esCLDDII
VojAUWGnflukBQ/7/H5r6VWuTdCBj8362bmoiUF0t2HM5EsblPbf/c1ZHbnf2KyB
DafCQRncMMiV+jUf/XLibIuR9xSMIMkWi0m+W0ZaXKcJVs+q51KLwxlZ0lkUKxRT
i2JyEFCockh/OGxhnrGF8zLzo+gFcXjPAdoRkvKDwzyBqWrWcAalyESNMMt/8Fma
kiz6SyNJBCkxXc+z/OLR3Zpph7E+8CGUjjauEiaa3rp4C19RbgkrVk4+TvTPLoun
BN7xr21s5aqjSc2wTSqMcunut8Z7ftGxp6rLFktZChZfOij89m3cRfhS/+gYpty/
dGs8YcAECaB2Z1wwUvsgQqNr/YFR/cMBzE+CCY58Q4nOsz0jKH9ZyO1MNZhp4Ebp
7BPxpEd16RgoO79NtJYJo9EOg+v3FH9xWTPp10sZNX4rayy+Q9qMrJ9dtnCD0A4d
ZSV9wfHiplQx5V7HsrnK62rymZO1NjvCaK0zS03z9VJbkIND5PhFCtEdVTW4xTvi
i+UdB+vL9K9zEdxqEVwyx9n/VRpv8kFpLCG0xCSkQ7pX7jDV7ej3/Sgb+R0HlztE
jtnUX3ccluLOuHNdaSQw3UJfuRTN97JYT4ztJIhcLZTeuEqViIqZFSDJ4urPHBqX
KRZLQYxKQf9zoFsqmMxE28wWWPfBSCBmHP/sV9SNVC1d2TcR3hTHmghB1BRdYOti
pgWfzs0PntYsP/XhGdWN4K58JbzFsHeuVjwJpOLe58MIzUUzrRKJwfP95U71rEuI
T6CgGKCrUvI8vdbR0YT7ncidpSsEG5O5mSJVD3GnTpKD6KyZ8gIIXb3TPXS7yAnw
T3aW0rTJsZOajU6Yg5Aj3YMj0sxhxHE97bLVleUppnhC1mpbS2A768a9ZSOvQVRx
G9O656Z56F/eQnAVeIS2NbsRUHQ2aPJyaNiUsBX9QnH6dmaSthQHHJHUj73ES7OH
qhOLvAlPDs3gIbL9ZSF4Xxl7ZESei86exKHNKP2Gmr6WI35gY/e5ehnpYCY/M1e7
I4weyKuAmmUMsw/43KW7O2OebkWDheeTcVqYrANywM88YQMelF3+Pf+heDeOAfy/
53C5J2n5bG27VyO0Mh0JdKEaZTky17gXpgRYU0yTi7aQq3bUpDrlFFbXmBEPr5W0
esWtoZ8+mLuev63a2B4ib7RbasApqMPQ8kTWi1YPYEgc7ivCLQEeMD1r3JCwfCqx
uRzBSuXDJNuIO4qIMkt4hNd9Yv0DU19triKRSorYqIfsQfcGdKy/pMll6IltcKmE
AdHnLVBenw98hhA0VgLsGpBmuskICmXOw9U4jTC6FDltV/JN8eMyF+AF+Pt8qASr
9NulalP525u8P5GWuG06oYzwsmgyYzEeocr7bKlmB0s52vPNJmQV3bnh5kQuBF1c
KmnR3ERkt1OVUpyMCzIqh8kQDS+jAFOb3yoWsVsbjAWOF4+btg6vqvgWi+6SAGp+
XX9UAxLEABlHDs1gHSt93eluozCdTtQi6l81CQBlvnrOUxuQak076/RZJIKWa5jn
bBNUYaTLIiZL/m5vPNu8I2iNpfBG8OwfjFga6hNSpSSbmjUP0yqeejUVCeQ5RQoJ
MN6XWEzz6C4J+11pNc33ooIerqS3VwgevtmgbQdI97+7+Uz4tTVeaOG/Bo+jnsa/
kqly82PaZDjZedkv+h0o0Wi5/DX9DP6p4HdzXy3namUSd1L65XCVs3rcBPp7XRfs
ahSh8MR01+VV0GVhEnzsbXeLO8JSRIDOmwFoua2nAqiPPJ+J5EK/tWwx/16RS815
zdXcxG4GGrPhZwKo9khjzduDJQRj/moT+OM34vm8hBlWQZj/sMtUxzgUUC+zBKtq
oMKEdXrVMpHfzEe6rc9RqJIbhP8KEwEPvjI8mKAOjBkuKr9ogrS5k2Uv3fxzIc4Q
1Fw4BSdN4NId6hGeLEqZe8Z6J2UxwzZkWQj7uIYZ9ZG03hjkEJtsiThXCKNs7kGy
Rw8moEW5FFcK4p/c2CsT8QKJc+RLagzJiCXeBRBW5pVSx6XCMkPdZtsUOCcazl9s
HdmQN2rpXtdFyymGlesO1h2VVisrSzWND9AuGZrqU7qSAFd/LDSByJyCxZoNza9x
jBBR5XF4uPnWTGwZTLJXVcXZe6mJQVsITcbKPheepwCxAjxSbJ1QNcLOchcJdI8i
YEmuFcJVDYX21GfGTFf0dhmZ/Sjg5rZVJ3usW5qYhSlUEW5MejWkAfTBazGgKSeA
mYsq3O7n6xRyALAx2Orik5ONvy8Edqn6Kw+UMm+xRLLItOC6nI17Rmw3PH+u6WXl
mn5oLCRUCfh5EC91QfAs6N2pIcKHho11fHGWohWSVTjw/60/Ng4qD7/YcQ/naMhr
6tX2sKEe/tUOgy+W+9NpFpDWZVIxFuxw9qiKyneKkZP8wKzJHk+tQwEzdTNauazO
yEmKgVw4u+ZhGZ9InTUKC2ln50oemF4p3V6zhTFOjWrFZXpiyiAy4HghRUzRf3Cz
0dWUb6bO4clYRzBWNBXrxQnvtc/G5Ss3nef35oNQWI72/qlulkjH6pSi+23e8FMi
n8pWXiZbxqA+7/gSUw+KiFMPRvZO2eftsK2Ot/+ngLNpzRGxT1OjYrEKBVBa/oa6
BlW1sPOliZqwC9FAabS9vBUvd/2jVS406TNmTOk56E6zUBxsvibE3Jr3Juwd1mXF
9VhUge4LCZIkIx0odrgGbRxXVYPQuECzR5rJO99Dv1LZqMcGpY3nhVirQIFn522o
ygqTdJe+xBkV/Y7iRmiPKxkayVUffDVgQ6QnvlA0HwWZ+9/mSc/ITzWiuiYJ3Wu7
UZUps7uuxZhifI4wdpQtKRLc6zE/pfW2lUUARSy1nm6BcXOj4hhVgJa7P5I+sMTY
V1OHYjL5TM8YC775vpMNFdXCaZovIr6AxgA0cU0RdYr/M2InJHpJqP05i63pEshz
nlSv+Ah90eBha01SUa3K1HKwIkawqKohgo/15+/Rx80DVclQ3LEBD2RXvROfOLWv
iP6zKw8gRbnJBZ22X/ZwZVjt87Bhx8AgN9zWxgdDbPuF8tsGVurhKS8kQOuG3mhQ
i1gc5zO0fRUX6PSNtAJdyteIHwD/hMdfeg+ddCBXXQwUXd6X4bW8/HE5D6HAnqOc
musF+jDWDnP8Dx/SrF76Vo7yMk5qJxKpNX//yIMDm9hjDWP0cPgu6auS1LV8BHgh
7I5BlkiEqCVwUJTe4rmt/GQnwwOldx8fJzYoyTEqfgzaiAHR+CHa8ENjj1ROcWF4
TgAVMYFnwoWcKDOQPqgIzKkBMLHsNhXumlT9DU9vdUW6xRN26EQpAIq9mjUAItRq
pHA0Y1cMAtXfIx5G5qu/MLJDOGGGoNj12fXf93eN31PgixhQ9veV9FuI0i4xW8gu
Q5TTZduul9UKxCv+gMmmoXo8vrUnr2XGevVMEHs5UZOzksAqs77aHXNcgpVt2mBE
HVYbLiPgrCofx/86jf2anlC993U9gamR8/K4R+6ftavcdKfKfCJtlcCmHRqd+z2M
QZkYfi+MuL7w1GEnZ0f7DvEDt2uGWFQ9Sl9kbauzrwQaLV4Syl5cUAdjOLcG4+nA
PtG4iWzWc2aeOn+4+PbUSWP1g37Z/4mw3r8X+rhXJsaSrUat18LSwBFBFQtnX2tV
/UCbh4+ENH9FzfgbdAXEjikKdepmHxKgWRWisH9IG6nuLPn7CA6ApgFFRTpIg/jC
EobOPyR/YtkpG3nz6y3CRTnU/VPIWbX4ATUgwfAihA6HlV1GQ2tG27fFCNscXsIa
zVLgf6VmHL7siKuqB3kSF4HIpD9TJxYRFkddF8DqL/3MZuKi5CV6ijA7jgsruxKS
/usycTZb7ykum+WCv10PvRvOReSp+rpv6iquCqrLB5F23nAAZ8DkYTLAriSZ61uH
32yJ/EdBD3XexVfwYSXsJSeuFLkbIsfrbQTrP8HI8OIkku7djCrYzfRjqHkMbi/9
Or2ra/PRQRU+pNGxFfcW2veEtGuC7IhuKdR+8M2iIgXenMcY/rnskrLGgzQPzizG
8hiLyza9hv1cQmlz/h+L2GhGed7P5vuUAN+49+iMgxT0Ta2vIWv1LHKqnlcYYsb0
HAo7XPOZ75RYuXVTs5o3K4syRHQ2TsHI/enZHbDF2QML3sGZvWpf/bY1w08js72N
LSRcs/e6i+TQs0Ofbqn934Y0QRPOkoWKNiWt3tOqGIZ0ZM1k0pGLFBSwAyU/LM5Z
3OEEkLer4ldoQSGiDSMoWbgVWzVP+kKcxlznj/KK8xdi7b2VWMU6urDggpJdGbrA
wTEtsyIpBzNGbUbCaLnDumZwW2XabezwcyGXdaWZ78+nlK5X9ShvXQ8EEfiDMLJ4
Znzeg/AuSEeLc7lAea5Dfj0oZUxljJxdacxSeZedcJHhOxr1FSo0S2BD2+hnv5u3
JzwkLPNVRuBlaHZrvwviAaeSIJJLNXx4bdH1iTATGKkrJqlMXLNBjJOvRhaCWf1p
iBhUiqSzRGr+qN72gXuIBVJcnRkd5DkV8JKOJeyn/nAp2d5tA9oxbPGo1LtqgdH8
ldvJmb6IAVbLfyaHNi5uZ+u0F39d2WZNKNwiadgG5eQlnsk0bMgdFXuy2lWmDrCN
sl8IFg8agUQNf8qDRcg6WfILTuY8JIAJV/llDnES5aaT9rvWKZ9ADGCFlIuXFy0m
HBFu0h8IWZhULe3Ci795P4MQOXiLJRnjffOQRFGUyOQ0NPonKEnSSuscqn9upPk0
e4GhN5IvG5z9IZ+HisPcV+MaJSn6nsj+mfla+BSF5cCxBogiTFh4zNzJNegIJcWv
7IXmEYrUOvMzm0HMkYWveCmChL0qKLESieTIwTo2wp4X8F9+xjwn332T/ndc1FB4
fEEUy6+g03vHB/aR9cUvTI8KhoY3U2FGkYRVoLC/XPEK0ELLkn83BTu2uj5WmLEP
qFQUx9MiqVHZ2/sT5UD0KGeSmBSyVfJyo4rPvrmLadGrxJdieBTSW6yqv8NVvonc
Aszyz00VfsoRwMHvFAPiNTgUid1evNQbWW3y3HWc15SV9XlcLjXxQteZw7s5bAXR
CcQB+M+fxY+NtqMXvoc8PVA8PICdQDsxv7the1Baz9wnVlo5O+Zd2ThSO8AvWHvD
d9qSv2n52mQffs/7Vp30cTss0VAMzOiKJyVA4U7FKnxorECgB4srn5ioCWjbOZ1i
whbkDWOpY0ncsT6DEaEGHGCYZCUjZJG+JIGDi/FnyrvQRUZWrrU6nucrVezxM6ay
i5o/a+i9FOCBFjANN+QmbzNATlcQTYE8Y2dvAimylVaUvrsr47bpiJL8kufQQU+C
CMh9oQse1nQxJdki4F7JC6ghnuNWKZP83zKuCIum145/IxTmU5KNeFRkWg9QzKZm
WfeH8sqC5xtUby2Ae0SVYaXf98NfeBNLpuyCgu7ucPPkzU5ZEQpHDwuUTyp3fZsn
iisML2yYmxd6l9Niz6UYxNF3T+7qeCue0dD94R5Z5X7DWaXaty7nqRLex/pgZvI1
a/hkprIndWVc+tiqHkaNH10BpUjetW2V4f7XtYTI6kg9R6JYTtJFnTaf82t76V56
AZqDDHy+dVqDiiZ55CjBgovrmypO/suFYVq3TupfMvOcIwj66Eq4qZfGK6If4kec
hzQOm0hdiE4hToKYe4tC7FfmesJCDTX6X5RYNjBGXNkQ/Y1KZsO+MWtrC9VEFDxx
tlUO0huiYPSlNKbki1tjuRQgBbn5O/YpcIskT4AUivfOu2yOklO2ZiOpgcMxTzeC
Y5qwvZjHjD56UbyUhy6DQrMtzGcxhnQ3ypz2cF89ofU5nTqOJzwUegZ+M67FJmKe
KPm+Qahm+YKkINCUd4HgM4PyB5Lza1pd3Ot7soU0DTYmCowoSIUl3EP+wcqDT3Ik
c8ioqMPKW8R8Tz6HpCN6qyaSZbGXMaGWhRuxIrzcqSalKE/6U0vF2CqJo0oLkXud
gZeQNawOLiX5vG04wir3fAFQc7s3qd9MAzIJ3qu9pQrgUeYJ2cTo8IGugI9SNDlZ
EMGsaW/TaZjGW3zpgcXMR95b6+JL1AevjVN/FXYsKX+VRmL5rx2Hmo8cmY0uUZwi
dDJ2cBFN170jhlKiPT2rezRhVVIyRi3Ix69fAvDsFx5me8mcl5RRDFdArtafLXo+
UWkU5d6b7CNG5Y1ubR4dEI10udUX+kC/n2gopsmiN8SaSNJESQ7QGuMIl/Ez+1fx
80+kJthJdGMaiRBexrMc+qGtnV9XuJw5UbWN/d/GKegA7Wtem2dd0m6lHaSv7650
OG5SRhEwD6BJcOTqaW4KbJJu7bYDZva5zs9MgbVacaAH1k1ZYpLxXMBRXxyI7kCo
ubUSOy8Dt7H5yNjovhmAMTEHEvszlq/MT27i49uTKDpt9IgbKOZRH4P6F53s8fgX
Ujproj21jHTtAR9/o7SFVPPftvHVKm/Tb4sBDdvdSQW7o6JzLq4wU2AgCtrA1Ik2
VkOmBuR8E+mMbistepsDaQOqi+GcvhLcMTW1Zz/LRSIwFG+zzaMWbPuAAmfYEcVp
g3+bSQa5aydhSqmam1vSkzvVeaJ5gNppO+2TG4axHWB9Qcddtf5E06cghnsgtXTd
WRERj6oegZMnXUJdP+hlD47lfQhtYXbGLzz8RZn4HOQtP0e4y0ajXy36wD7VZd9f
GIwLqJG1yDRC/uDUtG71uhjnB1iUS7keJrcRDDh2oJoB7H1fD1X0yzswbfXZ/g2O
hAhe1alTW7KzCSx57QRjJGkk4XUJta0m7HLg5DZSbtjyGBt/BoyRGCJS/WhtOGil
IIbQ8bVqJt8fZ6li+i2C3UYJ5rhOyDlJezC8a7DEC5k+z+glB3MqHyO/h6qNvUob
1Gco6fEC4xU3LJbJvg5uho/fJSCTvvlebeGO63WEVmEejbRX1+5nmqtK4rtHm7ha
wmw72PbnxwGgMlQ2Ouc2QXfpawp4u08yFllm10NaKOvBRE/S80xuPMTzmPVgB1i/
XYibNzwDbcvRyDbMuNc3ITkm/OQDkIT6BpC3a8a0Cxl+IC/xJrWwtTd2YRjjdsIj
NCv5tF1ChAtHHMoJIKxuvluvhnKeRdHtO0XIMP/89dJWn+W8aC6khMvqJX+P9r0U
W2OwEajZEqd3zBVXMciXktahNK/t5nipJ7KVcMdPTOPjCKOT4h4J1k/07xl7QPki
ob//W8fhXLdaeyi2ZZA9TiBhk2wW7t/bSDmaKY+Jyt6Q5hSAyp0RWfqMnhLos3Aw
bEtiLq2es8EoK4ivwqNz32CAtatWNkwgv9v055D514lZ02/RRSHFTwCdAxwCGV1S
mrZue2tUZTBMKW3qbeSJFpsfp+ZGWyU8/QLcujwknoK3fm6GJ+JzB8BiS9/u7luW
ZFidSDfajWITZ+4VaAly4bjg3cFv+mgts/00eeE8tgI+/O6AZV5fz7/P5bwpegHI
JDMIFpkbjAnI0DvjnKIBKhyxYcIBjL9Uq0xQ6joFTGjdPbSu9xrbqjihppy5NKG4
+5Kwpoyu7gjziRMVZNvnaHdrFrb1pD0SLiT6ZMBkDKQtr0S/7uHmu7xwOIghpuXU
ebcb76z4sjVMVhqwYI/lxl6yAA3Uz6tfESLqXawC/r/YO1YYajm8PIrsOKJiWGOh
Z54b4o/vK7cWssSwDRSLhfLtwhDvpmePCnrstZ4+NlEkieNlgaGYfk3jJk/G14Vo
yPfHoU1c3V42BYKO6bw3ci0moM3AzqVaI3n8XeB9D7hZZQ3hYfF9ml/elRn4+RUH
izVuxxpI2QrWdJYSxFQGZ2qFKQMf2MY/Z36IBSAL+Y2WgJARl3mgIO4+LAfMjwlf
UWw5KZXO3emkCo9KVK4zCR5iga7v5o8CLns2zOeory0GBk/Jn39mIfslN1gA/81E
OrRxcllXxZYCSazeOj938nXjBl9v1PfB5gn+xOuAFzxd/haSgDOkEVUNHzKLTlR4
IhVRzFhHBunT7c63EDkw7HfrEbo5oWB6g+xusLr3cuw4avi5i7ut83b84UXHzBYS
NHDuFE4MYUz86Je0cBC63DRBGDbWG3Wb4RW6ADsqYgV4CyhLJrgpqdkELiuKXknw
ZWC88X7x0RbN2wTdMgtum4dz1k35Y1jHj7fQvBvQutNA7Q1U5HnHHOsAA910E/SC
SHDu9FJ9JRxgZUMmhM6Mw4KnxLbB6EriWXtezs+FxK2cUH3FEoF8r8110B2MbyXw
74a+fzfdxvcOlE3Kx/Iggv8AyLTQ69FFjcmoXUBqUs1lgdwuL3bTV1BnRmuAI13n
8Vvs3ONLtLZHdmwRpgvvYB5pO0W78sD1a/i2upGtIe5G7qdWQjpw6pyt4b5YtEnR
N1d5pwY8tMybrZ+NNl4LDWIMfkcBKvEdObL2kv8aJIyQP+5WPYP023PW/EW9twQf
Wfwpfi6zi8j++ZlZGYbDadq3xn84YJPr6mCO8KcKxbi1alc3lyYCrYzZ/z0Nxx4J
Rh+ch1dPI0LkRwXN3BhDfuXzMoeOR04+1l3jLXwfvR2/lzL/xEC9mEFkvAvOlSXh
M1bY1I3wzimDq+9TCxpYvyvCcJBo1ePQjQiNPb2y8tq6ELwE4F7Rns4MRHD/7mO5
/OwSAgmvolSjjS7/ntiNtP3z2K/tn0KqhISvT3mK58gvjHFJkbsx6USigZspWXyX
ASGcZXGEPhYd/Pck+lW/prgzPAOOvMpJEgNqCuWkJnPEZMhD1aCH6vAV0f+yBtLO
O2XKDs3PhLf/qypUYEHD7ewiX4/Ahke0ZI5a9gCeh2eaxTYGxVZrWmApc4CVUbcT
YrFFBlLBU/Bz2dRUNZvXcA8Mcbh1eqmTAw396CYN6lz/SI6zAAvvdnsYDv50cxxa
ND7Qm1vpLCmqlBK6XE0SsnQxvz6j8Vs4pyCVPLiefybgPciCt2xjI+q0GsLcJY0O
5tpNdSl4h3wUodgFu3GJRQmc7yNPByRWdXqZavHj2k/BIXnVs+TBWa+dJQboqW1c
m9HgulRxnUWb76ua8FtLGOE+KKd+eFVhkNZwdyilculBHPKmFKgSjmqdO9rrO6CB
C2ZK4VNfkv6xMlrdrJwSd76YWkbX3X7ojnYZv5hiLz22hosdNtHBqc039uNqDRZY
lkaw6YDs24Cc9ItgCEjDOJZTAtR6y9i6a6I6DDUfB3ufkZaMbzJlnGl0AsNC+6zT
UiKK2bD6/hKLuq/yaOT3axCHthIi5QffH3K2d3yAvYZnPwqt+9ajsZqqr5QEhfOp
aAiZFAguWZfUEW87NjtF9GzkUpfEdhiYOx8jbf8MBlXQFAJTCnAn25H7ocf6z2Md
yGG35Z+kNsmUIdCsO9IqA+ukfov/fh+VwnKtx8iHInMl7RrZgNg3Zr5z68IQqWl1
ykcVl19P1fJ+NKbT8rMgdzKcKpQT9u4MiMWKDqqVirEuhcXyOp0vjloyHxA/9eSY
aNj2AaalHmw6sc+V3T0wgO5W1U/naYSVfKh/fCyZ47sCYSM/Gowm0jXLcMKKSLgc
SGle1RdDx2I1FdWk8xCQBxkwbSzipMTuy7QyeVztq7LcYEixtKRuRls+Uf+teVyp
YUw9ZnvECBtAQ3MImehUSdk79BP7z59AN590QX/vXmUKmq4WP0BTzikJ6ChLeYjf
t72wT6I+VDAm7cV3Egf5BoC/ulyZzsUZJClNGyFqsuXX8+wXbrgvC/WZjYLNHMX3
I0CfTRHf2orvsqlLU1g1etgHLGGJN4hPUq2o9ylUaNIEKBt+fPmUxvskK+y+yT0i
UwWsKBp88fwNHqNyygEIJSBoBdW2hqIpOuUOedxgJVOwC0HLKf6P/eKTzI6hsRsR
r+w4zA93XHXDoT5pEOVHcVdg3ktuIm/2hGea4BC23kzz34vyvHXS9swxdU6OBfcg
2kCAQvFwJi8JTY9gA52FAr4vaVWCwJOyNC5444/IlrxHcon7uvIkh5gg1ltB8/1l
8MV4vT3qnFsOxfzrdatsnTnsS+iItQC5eD0QI8X7f+wj9N9yagRLs/pvxkvls3El
NwmKZI5PFE5ym9dmdkjZJ+/igwsGe00WNDmIVI0hsMrbD25hZja4mnuQR4I0Vp2Q
5tb8ABYl72MYhkWNBM7bvhUqrSx7AWUjF4Jo8M9GhRVV2FsvXSCMeTi7d194PIEx
aI6WP2n8lpgY2l3VvuZIqsyBSGHohEQ+8UhOKlLS/c8uIBODLRJEoGmQqSOU6Zo3
/Nt3NmyfmUX8+cCY3WVY29xUGfWAwUyQ/LsHg92tb5W1ZNrAlQPeQyMu9YpTnn2G
06yyoZuG/ZaUbFE0/WxKEgONcXxeFJz1eBI2UA3TPsu5rITP93jB5RKBhzAUJGiD
y0STC6gpoarpN4BeQ3s7nbhQAE3TCZousE+9TUXhZ/x+UVb/OVhA4qqGbMCkI/im
ye/kc4V8zw3wojLKW4GyCCiAtHrqR/d0SVczWIo6L6PTuMGdNc5MBVA3MS7wR8X8
inSiQTqUwKUbGfhEI6asOvwjs2+7ClztFtmBdYXz4gDf7r28uuV3WGWCZeESKsws
aZqv1IVj8hiw8N7KzQVdsyAk0Od08H2/soxb5+bKJ4I8kQKe4TJaJHa5NaPnvmzl
BTm5jr+QoLHQP+k4EpglRXuGyHxQ7maSr1t3srt83b42gPBuI/35cMdn6V6IsJWk
3arqjsfE5khEAiMb+3JHX/yEjySP5z3KNv3fooItY4bvbM0lRfwaJVo79U/n81We
MvXrKICe0lA9h0409R50Mo2fZDQt6jQVqsAAccCH3kXwl3gq/tn766VnbfOzP0gH
usqJ9MpXOoG4OhbZJGwSUe5or+aYg00nKWvIp838V/2YJfCCOMEfkjJ/diii+ZNp
iIQ3ruZRuiTW21a62lYDrBJNztv4GBqbSwOxwHYdfrhejvAzjmUX8QgvdjbOemJf
yzxMPs/f4LM1tTVruvGQeufJJCmyibGSmPmOWpP8dyEYJ794q3ZYltj+Z/6UGBBj
FhKFxfuNUVxrKVCvaLTM/gaf5PTRIcJuzKLP18pl67UYXetDhM7wmRZnRpBw47kV
yweWV4AG2xk6uzt/ctciHpM2ZIpOqQL2VzO9FwrzaJddTVFvRU6t/MLD8YshcFG6
qBL5sXsUokd5CWG/mIrOL7jcFrXMR3RO407ZZPMS9B7RXm5IQ0etETjMaJQWd7jw
HbN4mEx5oczyYymQ5uCugvWhB8MP61RlHFdWy9oTrSDs8icueyk8k9vTlLGgb50+
PShQrtEObmxYWXGTAWGrwrCx7EFQBjGIn2PjCCxjLEVdK6K2qdZQABmwx7TfX5A9
ysxG6CMtpqRTnv/k1KgMy1J5Mxl2a/uJVcVeYXyAOv7RhYDXN+MEh4W6hUoOkp52
HJ1XcC9zHDNWDwE+DhRm2ybB0JLzB61riMOFtR7yP6Md7NBDggN/Ralqg1dbmw5G
QjMShy0yey8nBjPH7fBCkranG4taXMhSnO43TzShVgDZ7CWyS4XgBylXQNguLjzD
ErUCVAfrGgRslg/+gLaRS6KqE3NX3FChFgSeIF4pA8EsxrHbnS3mZRIpilkxHqUY
Gwfivphmf/I9k2Zx7Y7TFFsdupvM0WnuQwK7pAc91JUwNcpRm1ZRK8rXGXuLsKcD
+PeKmGRy6W/kCCDQxbc4IUy99IP9kgwjOYmNhOPTp7MJf1lOtC57W8QL09MXqQ5n
1h6LXL42M97cabUqSfrlb5oknK7AfPwQnVt2brUknGEnD8SnnPRQN127cnePLQnl
34+QiZ32uUdNWHIKGXPavxTrcm96suatJz9oTB9UXW6GDDVJqOQPw7qs0V7J2OtM
2ExMHstOKd6LGanN22MMc99oqx57X30ffDqNm5bYxaM8B0klqvUXGzRPoOnxvS0p
+FcpzGWf60zOsYlEaWJZvxGU5bbDrOUJCIumbVQ81rJ9OhGSxDOxKEAFjCueGE8I
vZcFKmsNlrmAQNyyjeRE0HQfmLDjZEf78vSC/C2OKrw862mt1VzNdfHzV4HX8tFi
bUpo3djUM/MRKzW2mpKFSd3r/Au48Ey50zU1zWhKoDHpr/YcUd9scGVgauDzgiHf
kiRwFUdmHlzg+sPQnzVogqSEfUXg9wqSQQxxVXlyEyE+NP+KIqadDpLjSAbo61gF
cjl9/bTJRDMwCOLt3Ybvk32d/KcWW0UF1iX8W3zC1L7HJzAi6mKbt9AXXtTRiPL7
BVXWHlQIZbvg/pgIGKMtF04g17wq3TtMkTzeKx3czuK/vW57zZVidLmTBJy9xaGL
jCdHBNPp4sTjBaHCXHaRLQHqF84c7gYOVP57cOTpFHoi5ODrGKK5n9UcEaxW5ayl
bwwc4vxeIObJxe1JxQZCuP7BbAvLyKE1qQbcCfmVlEypf/vuzvDU7AfJUnUlLqAe
n5AYNLS0Phm2eHdpQrJwggtQS1nkBc8HC1wH+Cvm1Cb2+7trmeikoyuL/ElBqp+B
e+MHwMw5+BO7fmS0CaBuhZ/YTrzYacZA+Pl+X+we2A9jz9SObEmJqo/uIJu3eyT4
kbvVGiDBL83Z9ZmDZ5WAJU8mK2rUhd7YqaqjUPd/hbv/JH5/Y33IjquFX3mejg5a
Q4p9/5lIDHmINlIHg7ThmnVFmNv0XBu4XaIWgLNJn8i2xRcIaGln4wO1QfzxznWa
oafid5ddYLaDdQJHn2HC6fKkQzK6g0v2T1kVz7c68aWaN3Rj/4jiPQNyftnqyGyD
SWl4E9dEpE+Kn/jy5nIVJFhncIysraYC1tk68yeE5Tiv01ashZjRCgGzZnp8vDiG
kI4eJ9DxOvrf92dNg2RfzFyTjbfZ6PCNCyNqLaua7gkg3z79KgfN6Oyb3OAsCRaW
RTdXdGEEOjLWtwtN/nnvHHBZY3TNfKv7iIWmYivz65/qGIBvn54R+Xj0sSCKMolw
kAFO/TNe+RtoFNKMwzNJC+ZMG/uZ/DN9okBhOvZEpiOyyQ50f9B4rwzwN0+5dJmg
HuL7a0KVg2fJ1TD9yN8/qkpofFaecW2tpQ+ivUeqL3x665OCOULrMNFTlqdaVOEs
KgV1JO/HYzX4q96CAOGIeFlb/nAYFC4SU9H+kGYQQSw2yon8IKreXTKlHpiBA7hl
73aqoFOWSNsw0BTmmWMHsIX3IjXAs6TWvG9HNTEkKjQpj39fNIEe4RYuRFKRyknN
DHkGFRaGxkS327BYGAo17mijO5OUYeFQNq2tjw0MxNQRcpKbaHKH8OP9JBTt754D
HAR6eHSpNwNDbn2fJmZ3GhopdF1bEDGLhDEobyjGR1ah3Y70vVN8odUntfbUJlCm
S+PXAcrVmMx3hsmLgt3KCHw1hQp0Lod7Wq1qjKIfPYPv4rCL371Q6Dbl1q8WhPeD
gHGmwdZaqPJktWgUnT+1XzFtVulxKQplm8V62FVdlvNLh6D5cPEn8PcW1Ps2xP8V
dp1fZgZnWOnq3XL4fOhlpCiexFfW+HZ7upkUA2lmpZpgxSdlassCLf2U+xB8z3fZ
2ijzv6hJZU9GMM4zWF/FeuH1gUFIwtkoxy/CVUrkAUfM49xJZ6bfrF4PjQng98w7
1Pz59hEMN+ZGsaPfu0XSALKs1OnLvyIWtAplnltMmI6ixCH0uvSbXU4v01YctJgE
ZUhdpIRHhp0zbEv920gD3fI3enwFOrcDbAg7A/C72ia2YQADi4L0FzpwPLDzCNKv
mL7eQ6Tj0wXqJTO4lFtWDv8/fesm2NGgiRlSCiikYQfvnk36vBWs3hHx2HIH41Xs
jwZweMF3YFy+foNB+qpHXLGlSpRE7PFk8KUJJZfUf2RTt7jsRJArI674BHpuw/r9
1GXue/SY3wHzjh2CpEas0wWvu9xKZBlHcKWAbrBw2vWhV5sLNP4slKoE7+bl5zH8
DHMiSXH7EkXXkAL1qH1V8fuZDCxQALThK8ameNT7TZYy7Y3a922X2w0WeqCJvW1J
I0808pV2zO+xTvZXVMXWItsGfqA3xA0mVPdzQ6j2mtiSUFGOt/MuHWHJmaQaCJyJ
1ReIqpZF96uZMT4YepgOwJ34ICNCuY8Ol7HjYgfRWdEp9NmvuP8klMyy7a0//5r+
ddZP1+HY8XHaRcezjrA6TkI5wCPHqLEfKkGQiaxIMIA+zgyAhIw2xJ3t+mViFHwL
7NVz1E+su0M8t55avOt8La/cFnT4i5jsGjEtUwo603siyvICNssRGC/i1AtABjqh
oTRN8GNTcJfFMjVWvPXG0EEGVcNWMa2K2yzLZurtC9/odgkQDyBc+EhwWmPdw+Ni
JF3KxlM7U6fa+azhD7Nbcfs/P08F44BV9t0xmER/lof8SSqd/iqB/5oXxzVh7+ia
NN9QbYBw0hm/g6mOimm+gzVdEUAwUxk0kBWoy/r+JuyWrPu2AJLXbgpRcPjHD4+q
n/3tOFmbYTtJPumcu5r7NC+iVWenF9u9mgJcC7OggZvVMVOW8JOw5tiZeFuUOdFo
ojG8wfCHVJVdjHotGT0E8e4OLM/FG0siGo8z2Bdn4Dy6F/ht5yqR0ou04ivwmzj2
bmd1U4SXFaQCcUqM0UkktYekp0tsTy47nKvh4Fqn0MDWIwQxTT/eE7g9NlJ9EIg/
kydDiSVU3CNG+q9X3v73GXT1F1TeuVTJ+heLuRJtniPTe6A7OkOdsew1mU5434E3
OQHwAjs8KslwmXLiHpWoxB9oy8qn9HSYNC9y924Xq4Y1qRYLI7qcew+DQEgJMEC5
BQLmgTnCYC7yKt6gklSSPGo2cn7DjcUjsMPk3oOYmde+6DJEwjQQ1lkYJzEBmvc9
OEd0ku/l5rHRC/chT+WL29cHceSSSb+3oTioWMDrQ1pHRdSokjw/CC3NzFKosjSN
378hhIK+K3z79ohQEX0AQ3OhQ2RZ3NkG0BrsquE6J+RSe1CW36R/Aufbd/rL6b/3
4IHPvc7+ut09+RLW9htQBhKhOb0Mzhkb+LrZV4wE4jYxdzJKUkrPWtOMgUoO3XGT
zN4OQPIGo5kDbftG02y2ktEC85yUP+flI4X9uMDhxY8bODvxIUdnz/wyuOO9Y+qa
PgHEbhMefCSYKLHj9RRYnKpfG1bIpAluDQLXzVJm9Jigbkb6zb4u/tNpcJN+L+Ut
TQBbIkVRKP11mzQpq5At02eK37whE3Q80THw9SvCKMkxz0EEtsSOYqfnD/+hxB4N
7U07EM+Bn4WZOVySx0q0u91eejs4q5+SvAcDte9NYx+Jz4esJhMVflfask/1xy6F
nSuE1L9y2EAaa5zaQasktlB58S0IHNInUuq5csjDOH42vhoR7HHpNk8g67ddoaD0
rzYzmUsRaWaXRfP0aXreAAhCuV2cXrMsi0r20QT1zmsxJRyD2jpn09s5yVN6N1rS
Qj9wBQqdZE9cpZPZdLVe3JarJZDkXsGIKtjPGtmIPu59sgXylTEbAS1L2dCwNDsF
RKHIAPmThihQ93tS/5CjbnkT80oDElm3CZr4pRPkNxQ637nV+Mk093uDpqZ3mWX3
AvDj6/oZ3pRU0ZWnyn6dnDFEMeUYGMz2w05IzHoThmSx7vlRzZ2JXxcCpL0n4uOg
uQkChM9FPjhJSSffnrry1IvWYF9ILKTR46mjlzctzMJvzQRSqOeIIVYoJxDMa73E
5BZ8YihsSrVtdEAJCMfXmljlkR/hTGWuwAdwnCoawWue4j974kEIAYsqYvafDf44
VZRpq4I7MSLAdDvanZ0TJh1DF+DR1nb7bkbmx+V3httuBloms0kkc7CTeEWZsjId
iYHhspz6gQpPIsiPP1ggebM2Xpf+Pdnp54+5Q2vQgIevypa6D2H/+QgHkBpSsBFt
qpFeOwdyAsaQmsBq+D57qPtXfFnBsglLxNM8963FcdPXPcR4MaUf/WHd5G2XUdvR
vE5QVaFHlq4oq8WyQaAJ6l2TcNLpZZZ41lfAv2pPh9UgBpOya7OzMvdUB2V2WNlO
BWQ8m54tiRgURBhxlZEmqMyh1ECw+xsrfNhvTLEUZWzNnEOQ491MkRfFA2XhFL+7
ZBjgRxVzzXGW3T3crtVX3mfQ2rWtUj50YIx+vsFuwfzJIe0cN/c9JNh7SXJqJuRo
LiobC5fOu/6SoqA7j06iqHBkRXm7zrMsvbFJdik5XkPdUDcpVcKVAX++x+50HBNd
BFmxBsX9LcdroFXyIlL/oNdBBL5AwbzU7JbAbFu+G1Ju0ghNr/sWloJ4Rc1h/DUn
dV3MMnKRCF3DKu6GCD5tolPc97TH/eStUHlzYY8KNo9QYuHV98FSEiEhj29mwkaY
IjAgQF5eRzsft+m8FrJGHaBJ+6yKHDD7VqutlrIKvhMncaUUOAgDPudEPOC9PjEK
LACxqBw3hDxYbtVCvgm3RTbTaaJg0/+7EnydfQCkNMeXuTxf4HzGoJji3zA6lM4g
1AbyfBpZHCeI2A/8oossnqapYTSC09pG7KBOfGjtYWzu1iH6SVOZvmTcwRt8mEeG
UHLtJByhEL9QRLGGncpjNYzkv/S7+XZ4H0eRIB/wGifg09GzbGm64zvDTgO50dB3
jABNB+nl5o/zS6zp6LXGd/bezh2Gmpg0AyYzeel8Yfo3DguxuegozTRoH9q8wIpB
FcjNS1mXkPqRFI9O2FPV5z/yS3Ty79wjBWHFRdjiFrEmeAEf5a9D6pzIIGSOZm7s
r0SEebtU7rq9agaOqdPzH1Yc3EewNqrBAHk83CcA1pT5N4Z3Q0qS8nmkVsWEVJfp
EHdaI8IXb/rDe0d0p8sNYYnkk0WsBCUKjKYswOjNlUS7dcldsKlnJzFhMx1VUeSN
zpzKhdd3G3Z+Xu4pJO4pNFl1DGzwELqxKjZoWbhYVygnpcT9F8g3PjEjA0KA1VYX
l/MyOEuxVkwLTD5YFKF8UrtN5mogVavNI+J9GGrz1zzqQ42cmv9rZOX1+2N2EEyl
igRXccFhrWQRPZDRml9C0rtCgh/RreZFxuRItH9xDOi9OUQRlk5SDq9zWVyinext
URnz4/1NqjOD69m4NCyK1xz6opolk6x4EgvZATIaJvS0LdFTqSVuiuditJgxXi2U
9FKFytSmxnkS4Cp69wY7mpqSc1GYr5G20iCVhb0Jm2i9JgiVYSU9Kb+PGAioexVi
BubtF0f34A54LVBrRWsROLU1mr+rB6EahRytTaHav69BiCTpghq8+IE86O6LUVhz
RTxx1I3WD4ovnlcIshF9Qcz5H07rmjVibZ9l6OFIX5tLtxxJX+yOaHCkCouEDWoe
xFsva2LxgjqQt1lYGi73xliWeX4+xUfm/nCnGK82r7cr5SMXECTXcAhdBquy9eVN
vIK8HhVtZBfrfr5G6fKpBLFkgjl9bD0Eu+9nT2hyboPrI64H6Un3J03wrI05U8QH
+f3gaWsTghJBwyZlKvVDX5GZ1bEf/8TnKphZHUwXObWP06OoHLYyHkYKGqyPqLbb
JL/732RPBuHsqssSdmy8KQk86MvihVc7750u+HTpLQC65j+UqVazDsFB+5P+3v3c
RWXa6Yy3yyXIMghe/21Ui29R4zoIrcUt/mQxoYIiWCZ4TnA7nLbhxu3qfwBTSv59
hvVFibdrqdLB+blN3052OfBuOf3LP7uS82OUW9FBp6xQa/d4OpgyzZgVYLnOWDgH
da4a0PP5yEdkvekMJx5z0zFPLam2eJl9UxShGAJQl9pbEM0E0LnXCNXsqYDmJ9Zb
khPGqcpIVOTAdeQqD0AfPByQFTZXr2Ap6tfno4223JGbOglaIj3uflyWG3mOxEsi
wEOE4yFhKtlxGs21WHFbv1Ed+nSdWFK5qlx60QjW13KTFFsn+/WjypDxbSim0DfT
X8MIyQmF4ALw2vPvofAKcS/Qd5DUz23jMznK0w7BWH6kD8uaNTr1it92xvGwKlIt
vWoX4VI3CZT5qb6+7zBhxW43j+pJ1zv7y3IvqpAVzfGIz1o9ExTesJpKGmwUiFU1
x3lC/7B3TJxGaqQvtAA7D/9nXQp++95yV81UmGOnWG+ghcxuXvHk3QijKw261toT
NQGfFYfXlPHfVDCvQsiwnSQaLLG1uAv8MESMicPfF60okvyyUTL3oQ0KMX3IPZJt
AubEW5r+caVM7SndjTDrQkBar8MD81lwAtkM6Db++zD7TC33aPgDraWBi+M5K+7A
iIoGdQ6jH1jGLCvEXJqkxuGQDSJW884SyfEN1/1Y/XuhmkuwBEqyJ/UMwGIHMfXM
Csec21cH2DCCsrMe5nzBGRQaPMtECZgSh1WrpIzjPZKT6POgPy5XlJiBIHoxjiF/
ptzz0wxODwi7C62XpYLgacipw1gGuTpJpfhU/Nc41mcTER5QMtQuBhNxmnQOWTEK
pDGiZHb0bBJ/HZttbd8JJUzi2abs2uNTEjkroVjvjlX9eA2HFf9xZ73Q5Y2LcaOT
bO/BZcRJ3eM4PFqZdLGVuiR802A6snrxGusZuvr2Kt+7UkbVpEKabe+wylYl/6wd
1h1+Lk5plLDPTxIbC7btKTEtCSEh+Ocq+r4kC6nO5A//zmG70wxVeImpudEZ/Ui1
SPjsA4FxYdlhg7FKPJ+Lj/2J4KzV1/nZQX5wXwoA1SeqWUbGWd6wCnXRsaK+5S60
p4O1xfMEXdkWRbdwrFhEEbG2oOJ2Y6OKwl2L0WbWs00PV3KMvmCoCnGZgF4nsnP+
UEv9fVvlMoM5OdDsQvfvbHMJnN/ww1H/7YSJA1s1yGyESfoPCdvsyJvPvrom0Xso
gPE+VgF26MB9PMBE6NNSoNkyBFqE4zsPMA94un1Nlo3jGvBf++xT4UunkhUVb0Am
64jM3gBX4GwmHyuag+HsyN1hdrB9HXumcejgXA2asz0lGnnJpKxNsBLhEuuo3da/
QaEZfo+bHDtGUsTQcuSurUgpxoRgIe7Ug05KynmmBzRq7khajOyzTrj1UhT0xbJD
PlqfAqorAqhZTkp51BHPuB2Za+nqE1t2rbmgc3z6UtMHmnsUJzfqPX1kegTemxBV
vAPyZux/jM/hc6Xh6UmRwnR+J9gZefEdwmdzk20lfL37kysp7PM4Qzi26R0H4KkA
2tcnvjIPsCs2OkCEYKxCotsXjp5sTasVNXgN6DljQBCItnTMkjwuYBA3iqI+32dO
PSJ/9pccAfphaAPp71DbgRGqmxZA4YpaXuhibhsWfGqIAZy5Wr52Up3rWu/2tN8D
g7ME4METM9w4I/0c6PMcDvx/AoYWs7SyZYIDWc2uMQvN4jyJ4PEfJghW3uuKquwi
cVFuB9t74PHwO4Z2FVtw8EyWcyH6Cd6iwHo0XU/wtxjhUtOc6td00r0fQuI+0IoQ
bFFjCn/aaN5aeaC1HXLWvcNpbBV6dsjxm2RJzR+ZeBT+P5zc+NTUblwcEnmyicuM
OUDxcmbzS4MwZ/l+JzCWxngHNcC7QA1znNOuesFO7u3y9LoPAfOXQUZHXojTAdoH
Y07X7lHUtFb9usgwN5HphVZTMtUYHVMtVPcZuFsCFU5mEnnCoPiFbZjVnrfuwe81
FuOW/oO+k+lzIN/ijNlBKBRasKe4dHEf9ZgfdJaJHpueDBLFpUz0VejWQQnz+K1p
egkHLGN4NwEjGqTcv8ZKrGQwYxOdMxudgmTC69+JSQNrb2zt5BcSrrvh8lIhnSSr
mg44bzlaPqg1ckpX1Vra6vkXnpTnBT+zplSnTCptIrxnew05XScKgPqIS3FTB51a
NEXiTxxsbWS76MyRljg6FUF2sDZcB4Dnt5rI+nKiU2bTlilzJ87B/xm91XBRgsLq
zc2obh3vpXRUqNfOuMKeFiw9XXgvc/ht2D4+ORQVuB43j/j2URv12ytwUOgAy5g3
hoTchy0/7ylBnbFCpVmXPGvZVEZVdwh/ze5agDg4uDVhuQjwvBUaX6rdOM0caSN0
IYTaUPIGYR7yiwGMTdmcr1j2i48k3jKrqLoqe/TH2i97fO7XTyEHvkJ6eaSMiphN
7K7HYa27Pzx0dEDIrXCd0IgDXeFKt15/9IccjO3YPW2bDlxmxBYul2lBt1GwV3Iz
bRxydsmW2tgk8qWGMRn+YqZ9VpdtQAS6qWNaxxXafrU5wgSISdhZx+8c5GVdvRCH
oGsZMk/JpG5mvaDeQqPHXI45jNOESaLPAM9khvtCkqJAsqZLRfW3bpH6fZ6bD4z0
fyc5Gf+HnAvB0m4TUUf5DrWs/pYe3FtSIJ3cJD4JE1NkGBGZH02YCDizOHL7BWow
IjzcKWhYwSXKbmtk+SBkGYin/xpRedSilxYt9XBS+gQi+IHkelZZEvq5LNHc/VOk
RsaELtfkGpupgQdpP5u5bqCQvt1dZZXXJ2e5SUnm2X2nNFolHiGobXkKXqaeVSPV
qU52ei0+WTS24xrl8DPU11pBZLH9LIPG1xPDAftfoNStyeB5L7J2LUc4J0PEEFe9
7WvEOC5mkc/f5wcCqANOD5u4xt32lUj+0uGpb0sGHsgALEkYatBOqcZCVlff0FyU
PvHwxdYFJ8hZPytMmFANLFy9QbKGqMTxq02Jqwd8/SZOXJucWHe5muP7ciTUnI5d
68x7Bh5HmzNSoxEoGEfsz76WpvmL+eGcphNVemTt5QcXTZLejRfOA+OV03VAGDBo
CZwLbeRAp2Kg6YkCAkYhzV2az6ayuHnAyIoWlZAJAyg+ACTi7/Lja6+gCOpVenkx
3qHRpaqWM5SJwF0M24/8lZKxH5I4t3PF04zixex25Ja8XXAmt5FeD1KkURiTNH2v
lpFFkV6t+MRXWvBBCaSY0Nq9hPqglkYj97IhzNfLY1vgYJ+BacRz3qaEMzp7VEtb
SkGnJWcWx3rDGRKrTxSNl5lqswtpTlHIzm4bFznhQwkZZTaBeRDXxMEwbnq9pMKe
NuH5N83h+YFXqSQTIVgTCi/LaT/URgycYiajd6685FDe4SYlil/mE2hRulQRLYd1
v5eECGWsSzEYbIGtkwjt69deisvLSDp20OlAj8yWmWpZYK5Y6w2QBBPf3fSc+zLy
N8IvmlU4qwyhgYMr2KXRZh/eZfaXpypaxEsG6O5b8/zTeujElUKlz0SyoUDqigmG
PJyrw5ZfHKG9Bd03jMNUHhpFBtKoutx3hPlgqaJYuzQHvsXswvVa97uBFmt7UDmP
vb4qs5+DDzXWBibXGx439/qL7bM8qMF/2FyAxj65m3zPuCOfGNB5IzL5CBN+Z3OO
OvGTKp//F7jGd5MoNCzxHxOQ8eiBIhzLUT5vrwAfewcT83Y2qzpFxSrtV12iryfT
0Ukm6BySvy3Izo778QfKyb4Xmc498knjQZOT160Kt2BVHdB46YQ7bP9zDL5Lv7s2
QPNwbuQhuyERubElwAXl5PhDPI6imS9HkpGu62iFqbek2XmuRsLZwL/z2K1ZQNJB
gRc2nt0TKAbxCUZh1kzkLQpQWFSjVBbROg7qAyT0NqDnurdJOMXrSIX93KhpmdX+
pTEuG/7A9FMY/rgTSAixnAvbh8xAzSFq+QWRzP7fxvoABixrSHJNJt4KphV1IZ2t
AT6rPUKuvSKgCxuXh5Y8q1svgrRJ1LyRMx3FU61sJwy8/rWWQg9gi00VMk0xF5xG
jgvOfl5Hg2TVVPGvLRDPiAjU6PZMDvBdpbopEQ2PTiJc06Iy4VCAm6MadA/zAAJd
1K025qdKkxXhKY+CaFZjGN7jUwA4wzcThanW6Pi1zAsbIqmmSPRvux1Ox26UA26X
VSls7PxmZTYfNva76cE3k8AUK1ghbwyzZ0HWFh6Lf+c5MzPofD2QogWUDqpT1Suj
ByPiozXIYeG9VV9VsHOUXXb8vMRCrGvlZbahfZz9NyncNWqPmJLgcrHctjfY+z+H
xh8/9aU7Ga2qoFL1E88r+yW5jd4eSi0WN7sD0FeICbHQQ6t5qqjEY50Yv7xqKxIF
Om1yf8YWSg9Dc2HRMV+zhYykv0r/YsfED790/O07DkZVEDmiaNOClx5XuYvxilVu
BPqXAzI5lxfC+JGw/k9if7NZty2WFFx0pPvGQV/AyB71YuQxLbuqko3rzdV6UC6L
nmso8A4UR7f1eFDagQ+Gjlde/WOYh1yfBS1Sag34xzXK9CLivDFJ5oRIS2Fj+SH2
dVoFjtFi8NJgilCjHt7sMbouPADFXZTl58BkT3MnsBH+Z9v8+VTPwkRsAzIxkaOg
j3+/eMXUcnL9I0YYWvy3jvU3GVh7pq9DWdA2wy+TKmJt2NMGXRNeXPJ4IT8W776B
i4+WsyncHtQW0tCiwuqtmIkTOfXYroqlmYCC8uXQ90ko5NzXWmBv2sHUaqvBjVKX
J4GOgtF5dJACtVBSwsLGwJoP5215oGgFzxH3g54kfc96RTNU2JO4N1B3RccGmrwZ
V5M/JUgWLHO8X6j0S+W5tc0drbuK4O2BJXdpZlZvAsPC05XVcubnsLD2q82OFLfE
XX7SlKrSWq/7WLcuqZcHCtxtEQ8oY59oIKSMBmW43g0Xht2NFcE7a+r/SmSO/G3i
vH1OZEktifDjIOI/tE2msu8XdHJLdTON7VYg5JyImGkzDfEok9D1NdPh/6YcuZDZ
Y+N0+r+NUWy7rZfq6Nu6xxfX5NYlsBrTvVYLS1k+l6kiGUGR+Urdh9JBAPbePmk5
0La5vbTSA6gq5vZcW90xte09B8uOEpaR1scv+lci9eeMh1RgRY9VHITILmPRRGM0
yP0sndlTWV1RtlIjnYmdY0SpuzeIjPH1A0uK4NbQExb4oDw0VgPhjoWNbL+0bAKN
S7IdX2vS0eiflbNOHfNOUa6goXMll+0LE8W/e4BEc5CfG260aZ+MLHJjckNE9C23
XbMuilrHujK8h9vTxy6tdCHNXZ81ouGfGVGUvUF78ImQuQn1fQaPJ5owQStDFZMJ
olFcRzvpllYxSEcHrkxbFgo2YD9Ue3t4hr3XTkHkVkcvlSw7GW1w5ZRnyxRBo/+Y
eBgcVQpaPlsqyC+UuCnAqz+awz3Qft9KPedriAQpNY6bOnVJUzWxMf6LuJ6KjsF/
BQBbc1V5w0EhlTamdGO31Y1IYoZR+7d+b7wphi+tCrhKSqbGuOrjFvYQiOZkboAX
CYfvu6iadimoQbh/wyUG1xy+EvwAd4Qpp3grYe+6fP1nf9G/pkgrsClzK5mqD4c7
OeyM1T5qN6hJItJbpaD4KTNAiipiE9yayko7PAHkXCuTHF7i6X7ewK6tMm1S9YMK
k7ITitlqRqWLrUCEpL/ZDIEDt+FBsFvK1s2npHvzGFyL9zuPCaJ/4FP6zXvGaX1c
HDlN3spuy+FODdIJiPusY6W9XAEEM6dba735efroOuaMwILGW575URYGKyJ4ZI4Z
u08WwNpUf8OjGzXpa5OTm6BjFsPakFCFvpNnMnGsU3zyIXo6gY3TjbMDKEkEPqXX
iHVF3DNa1rOa/CCMVkkUPigz1u0h8Li4hS/yL42Ib6y80SMcScOuXSW6CuCYEHn3
akWWF1T3nOYmbuFLo3rAcSFXXj+64OQaTC39yed0vB7GpGENTLkDsQERzAryaQtU
vjbj0TnxiBz1mDjlDVFCkRqPCdwvLi2kiC1ZbobWMl+gq8hGzhuWY9WIR4W6LQLg
dU4GCgVi8xrqBtuDzXLxwn3AZ4ppJFcJ/fFuR7XH8jyMEBpcJJ7T8HQV1zFCqWfO
zpWqV38S0UfI0DJ46Wb8MKhjtOTchbgKuw6usTyCj14hIUto5so2HpJP4figVfaH
Lcv61/e1CuUvPB+3c8EfQS0/2ybrKD2O+O5CMPHee/DvlYKSCgxZUGTc5ENdAX49
5QuZiHYwRRdOeKDjlJQcU+aqQ+Cxd8+hMdfbrVng3fjMEWU0E6uerBEcsiRcClPX
vkhbYyiras6vaJQ7mqH3QWGnU7F0+3kxBXRJFy6lCaCxg2GBu90qssk9jZfl5YfC
2bHIkuD9faesniZEgFyQQgyEzF0IMZY6Wvfxg1GBa2/EvkADYnUavN/wU/iftdyi
m3C65RCqr2vSp6RX0qfkKF3JblYvtNPIubvwNynJTgXezMmdCy0zcIPt2jk99Jrr
vKVSWs8ysp6EPL156wqnxuurjBAlSCABSE3v4xY4YR7oTmPn3RkHEhdRchv5KT+K
eOlM44nB1Cf2bsiUtsP8mAgV4077d3FD6FH3+oBENK/mzXHthxF4aLVk7mbs4Bwo
kJp/xvZOVZDoe9foLKpzWD6rdlrO9FacYdlqJ9qLJzNoupHeH72OY9wAEWadpHbr
QYq58B4YQLQuGoMCMLOuGYbvVG916xJoQLAIzg/QgItTxYHX0tRzG4eGKW1K+KaF
NOaEGejugrIAtCb5JRNgL8YuToKn8k7pwNTlyM3BvTgIFfS0b5zrBZZIqEpZ3Zif
KYWOng3FbGJSnXEApMGDk18H1PyGmOQHGaKzyxXJUQ7IE33QnydFul+q8AsurTDZ
6koUpXT8CWsu0VZQi6aRL6u6e7LXQDnVwM/3RcPHHsY8ItRzcODxyLhrgvgSm4s8
X/oNLSuq3WFjKES00DKp5+T5Hf6egDH/UuBcqpgBJd4WssWzLfEFHSWT8Y8i6XeC
vk2XDEsVFCn3BGlGdZmocoEZ4O12/ajxGkLVuiDtVt0muAKFPWalHvmgVmgv/XBl
NC8bZqTJdFl6UesXPh3tZkfKnPD7bmudc5F5Ohwnw/0gRO159owljGtmVTGrRB/v
ICRJHvV4MZw7/HO1BxtOlMKtRzPrNLC1/YwNrs0/RWZsIqovmTPM+Y5HJ2b8STLE
jUBpFU1mmNcl0ZbcROkvYao3R3bS88wNLIHrnEKeKdZvIF8X5Wr3cI5xA3XTveqz
jXUtQ6kXhcwq1TOHzYXKyWBLpd7fMvOArsKAX0i9nHFy1qf0S1O395UI1LkIA+23
cB2MhGlHjvZemByNVHhY3LZuo3kjuYKKsd2NizSHoAFdDwXXHCd9f3aaQr9eUGtz
AFH+AVTacJhBQC9ee5kGy5v0xeqUqGH52Dvy9XGACmn6dXWIB3UL6Y2nJDBkHw/G
oVZQrh7lpU8Y7mw4TSF3TXkDoqe7hH/4Dsy0BJUJwjWKl5eVV2tqQycqy8KDDEj5
tRxGiSTLBlMRisnRUW1mI+rnfnl3sazlgL2mHhB2beVT/t9dc9BFlDKqpyTpoC4z
pP/JKWI6jGG5GO6QAeMtcbDZLGeka9qX2xZ20FVuEbXpioKBUPsM+SQhZivfDnYw
isYS2gUk3+ho4ueKKkZ/7yLIFabQ8ucS503xGNoxTuTLPxzuyG8XjfeS7Uv6v9xC
9AZ8Yk86NJF/WLX0DqQ+90kKUMRuHERTAdJpBjjY03asG1UQgqri/GhdtBaYy41R
eAy1TvRNAbw0OOQidItibI51l/+15ee0BpeUy3FfP+C9z+Zu+CszvfxhddNRDhfc
UxDdClGkTe5RGiov/xoD751on2Q3gH98Xcbfjb28UOGmAmRTbrRjc/IOPp0mFHgx
oiRWTJPR4jLRGqHrYFldlH2tMjeQFqF0DWFPeOOYFijQCtsvZpj650UG3OJoYhBi
Jzlz+vS4uWo7OEgfWC3IW3uSo/PKlp+2DTYuXu8dkIvVl/pWhl/VeorpEPeG3GCN
46ftgFIcuV+M6rwRzWb+cFEj4lHOUasUEKdp1yaXMnZWVOBknwQJO6BsJyK7evTk
gzdJHWsXGCVRpifa8SrK34znB9CDgsqYTL/JbHjgEDgkoU99uSPAxGBV0CWZusaG
zoicePNcjqlVgdXKYefTFMvxAmZtIlqc5WCmlN6Fr8wHhRwutV/6dQh7izmBMNrr
ixSH2XTCh0mYgH66kT0A8/DqmjFIPpnxjEb+R1IyNLtvB2/mvjIMS7TjJX6uch7r
qvNjSynVxebwgpHvtE6zDkMfpTcjDRk2pa+u4Pw+ZWN9Q3htC6Ig3je0tHQdxx9x
NAFIdPK8spIf1UfN47lEKZ0j8bpyBffI4RDAXJ/tlTZWLE/9iyjSNfYJo3dhxa/2
a5I+BkAbKMMht/QkkCL+PbP/6EOsbBtwuJhn8vLPuuSBVUf4HKsrT9CHAy44mwHc
+53+niCrNbSzwzYZX/5lTurcDC5dLeT1Mxp6tW1CBB4EHwz3k2pbwzkkIQZCApJF
mllMLVYSzoZZgaWw1RjmM1taX1VNjbTUVxDNV5kzh+Vaft3SI1C2DqBZhMFz8ypE
bI17MMrPDtWrtbAI+n6tbAHAyOvNKEXgQN3u3HjdDcAzEJJItXNsHG7YQOJ/m9ja
JUqv0t+Ze7M7cEQVmg7LUnYuKhXL0ZCQvXXrcCoIgiR9GeDN+XH7/t3KPUu0imc8
YXsQoikX1KZQugt4vU4cf91rxjWfPrCUKcZwSUUH4hUsNSYEEqwrSBm94cuGcyCU
UCCTUFAVShvZW3m68moPpY0opdPhIBh+xGen9qnKOUWqaN8qyyeVCfoyRHNew4U2
1f58KALvq41UzDNCEMhEyfiRoU0WaNS8GN1ZmbwbXiC6Tw5ZXC7TV4zzMG+Xf+yn
njmbeBsnI/1IM3ZiIaroisT4l+bSgEI9T9xMWqt6bbe4BCo2dDYiMgpN+o0jXqc1
JOjvbGut/XtUKKBPITztLweqVostiMHtxHqe10xviRZ+Pb4vECPspQO+r/u5i62g
NE3V6kqHBWejiU+endo92b0hsgPT/cBL0DP65h/Aw4iUbybSvZgA6MeT/Gib0cG+
+vL1K36aD2ITXwpl6Pn3nrHr25JoRvA72Vq3VgsfE9Voci4YiLodRynhN8UWQnIu
+9Y3bdxPc91AHZ3hv8qyMZEsVzD5znTX6TVrg/WdGjni04aAsZ6K3PVBgTlwwtZn
vjTbQsY+3w32L3vakS3V156Lxn8Amh8n9haBY0m4AJfWuPbPZVz4kHTtKZ/WHy7I
zuLNf0ySwVy8AItrVcan1GB3o9RqlRwKaRSgXXdEmOWGL0gKo1AVLxqjcW5Ecf7I
jr2gniyaj4L0+idEnfmtimmyZjpjXTh5a/oc5oHUy0nKa39XH8EEY5tRZrPKwe1J
vfmoT5v8mbfJvbYmPToAJSyqxvcr6+yVeMV0LYn71I0YNYUDU2tBfnxkRL5XnA6+
gkpNVtu0qyuthoWK7bs9K1w1gQBxWAQqzsj9Non88CfiHQL4yPqTvYTpGRVv+vu/
ujE+WGiATJEHYPGcxkN0cozpohUU5EbXlvItuAeTip/Plup32nwdkQqJ8kXJbi0Q
s78fF7eNfPSf7ju7gkzy3YWQ/tXJnN1aJw6CMY13vHcHHf+NN2l85c8m0u0JCiFj
v7K7VJmVVgn2+dpEQChjNcnBWnhEoqO8ITlBzD5W/1odJCIvKPuzmMb1nASGvPE/
uP3JM6dt509EM3I8aUn2E3o6uoGaKLdRswz5VxvhlCD1Tj9YnH53gHt/0Jrsp5Qh
EGySV+B8c5/lxxPNMhN5nxB6alr7Lp5ytTTy1H4fvy6+/DgUJkCpt7Y7Iin4T6hf
1EHsPUznpidZRnuaIZQNRUoskPQpKX5yO0HNQ6d/XhdYhzp7mMXRkol4Jbpr2PRy
1/WiqtnzEm2zYnAzxH88eFmPgq6H941dXxu7ehifOfurRL+r9vYxj7LYgG58YWp4
BrsrmPmRiH+/nbqKjGY6qjhYXxXQsBdc8WQ3lSEkXFXe/KHkts1gXA7mRmbpmO+T
q8TUCX8xq9XtaZ1OLG2Elq9Z+ZF6L3ainGmHGSWyiyMA1nMPjDYHKttsgiB7XjgA
ozUO5QqinzAvJi5RPAPuy4D0JjzkaCaXGFwDenfvjRi7nGfCyLF8kNzGUZTjDQm6
Iv8DL+jbA4T7hvrZUxI2esjGTwFqY+BUNEaogUp4i8TKn9NbYw0ukf+I+Pbo5n2F
/KhmK4W1gheDb8sGbHm2Rw6yQG/ISoFVLOS5QxSbdakyTIV0dYX+chcuBsDD71cV
+I+/e5YGCpf+6hYpwRLBEKmaMpOrn+FVuY+L6hn/zvx1Bj7VBOw9SndGtxKD8ZUY
yQm0kbsL/skPWbSFtd3j/ibnrotOV/Ehj6m41s7OiWLQKjrW0sl+9uP91OgWFQqa
HQs5ICWeec6qL4dk5l/z8izOAKWr30p7peyBTYgXGFHrGYZkGhX6M8W5guz/yLXx
kwQnYqQyKzyusrLV2G/t3fOuCklGX5f52UE/HVYA/5GOX7Po8sUdwY6YNqKdb3kD
P9nUvb56tSxxhM9fH9lxE02tTEe5kAmvO7Q7JleRPoKXDVSUMrnd13d55yGPoWnL
8lfNmap0seC26g1FrRXvDUlNiIYgtoRgfgq3BeyCboOOVU/kQsD0Fz7vU0asKsEE
kbgrvROgS9sneMXnSq2BQjKWZdu3vXmbDMdJqO93G5Z0yKS9c/W4PRWg7PqSnap4
T3QUCY9JC+dzFZNpQiNFQDW17a+Xb0cw3gTueqzvwXUTurar/aiUs8OssgEBli49
l/xdIy+aQIyKeEAB1asyC7rb25yyUjN1r/YTKWv4F4qIIqSvz7Semo5K54Ddsfig
kewgNNZDdaBtZ+gJf1GXOD2wdakApS3J0zQiM0AgR0Ajhuuwkrd0eT4cnbTVqQ5v
ZKkCMFkn9IS+0fGEt/GKCQT1cL9awkxxZLqFAyuvRTHC+fjU10boPFNxJviS8yL0
MbN3Oi45uyZ9VPZmWmmqrOHv8B0QZbbxhlvQL0EE+47IbeBnYsR0FSHP2etezH3k
UofBi5IjYS1bvp6W0ay9c4PoSNvRp9xIfFijAYm/AFYQkZnwpHEktIyq/+WA+zce
gK7vV5GUAktugDgIeP0rP06zV4JvYZlUnX0Jyx3Vrun+2+JPDIa6knnultGFPFA9
09jTBo2t5SWyZqoe9NEUz9gO6jL+cR9EP76BmZlAp+Thayx+E2FdqGqpan9VbkQn
Tdc48zHkm3MPjXsMP5BCx3Bup+q1y9jPyxpWz5R+fTfYGI65E3xJW/dnO/4kGVti
35GxDhbVYTMdK3apsmvegZPqlw0Mv9p3bSXWfNHxZbp9B6Lu1Qw2Y3QdDllF0mKA
meLubSv56QCKBIocM68N63P4D0nNFjiXCK/B+JOFlJhhOHLRPGV5FFGrl6fYnppp
AU37j0egiXmqJItZjxEEMBw/tw5rubM+2IwSLazjObDKW1mTpO5DA1qTjCXIVq2F
vtWlmWMz5cTz4QgrkHRaRmRX8Gul5U4ciuyjpeG1/kFOUaMwZ8IYf1k39kMyK3w+
4oXOoKE7XT8HlOu8iddhfm9fyYzetUascM9W6oFckIcrj43ZPGsCKvfGx3Ifj8dT
r6Yx3PaRt22zjqh6hR9FgK0E0JUCg/a4TYdRlNhZ79Q/f+QZh3knI2sMhSKAqZBY
i9OTO8HgkQFAvtBVjUXloC4kT0qY1FwhoqXdnSmttg/FBxIBn5atb8oBxzWGCxob
RpVyqLODOOM8kEl4+hyDu9pNzsjJCr3f/iR0WlqeerkpEyT5NltZHPdQdeEh5/AR
MW8FynDtuKDZDbR9BvPtBI7kXeu0PBjntktbwKpq4neES+EdGzkQF+imbHM0BUVv
Bd035wwGmWpIyPFheDA2WbQvYmKY8YuzkXh6ZcrY5i2gV+PdvqawYuWbvz4R0ql/
VT09NRy02ow7z0ucN0yRAex1tjS8d1TCiGd1p0KMt8iVi7tb1EHprM/HzlnIORRN
Qs5BtvbR63taGikFBXODWa//OVAc410pdh+L93ExJkjqwwkobxxDvexx+8fJI1Y/
qBquxUMnUSHJ7l//DugOp+sZaIvpwPOeOZSwZQVpAVc/db5vlwhE9xM1JBes+qc8
XsKrKTadaly6KPE7iwB5cIZeKrpQHBPAkQ9JTV3F9a6lOb8ve7z4QNhmYHn6/SSF
1VKqZVTciLQAnFbXCOkYHaxAx53qBeVSLb4dEeWjjqa1gqb/Kmc3vSH05k4mVK3h
P22MUPW/LBWFK98qH744SfE3zhiawDo2eOOySji71njWDF6cHXMjgXVaDCZOaRkg
RLcWl9nRrtnDS4vz6C1/VF2lmPILNYBClBgugD2iTxfuvDnSlErczH+dMBqRVUy2
uE/rfHDJShb2C9EaFFoic7bPelHgD268IoaP6CfVS6mFYzYZS2fwqYga0VEJnYuA
nqosqC2zCnYy6wXeSkYjGkgoh1aeDwa1owzJA+l50Db8Jr955bbuoVCFKn6KXDBU
wo2CVHPI5bAJlCrpXl1tFqjonWacGNanAKqmJVMeD7c7euSL2+YJUWNKYjOwtY/A
956prgrOhvTUXhUXBWCyjWIo0dDRC2uyxan2NluX3wt/mSjGETM7xbz7KpgkV8oN
xFX2hqfpfrNHmMWXsqO2CH/81kRcv09AnIds0lYIF2XTviSybKeJaQj8fafaSwER
5TYrkQ5av3aBulkr7wTxvKU03F16icQp7jlJw4wsEQRM2BTr5C3Q8Z3+huwvX4LC
dXmQecHjdZhtqM5CnEcTtLJ04HyG21vbKI3p9kkE6AwxJ7BrV5ld7296BZzJCL1v
wEjgKmtKQzuFhRM2riIVT5YXS46qL2kHabeYQc1/JJG47pxDAnma+qDEIM/VflVz
/1Ugu1CkH0BIplXhDOYETvn6Ot3r2fpYZ66EU04vVTm3f3mV1hnfeMsWAQAczMwx
pxGG5ZWSnPYEqJol6Vigi5KT5SOvfwAtuwyF5HmyIuhHrPbFB1lB9lDAwK4/pfFR
XZnq32TPbrZv+cLdeogZFjdpRvC1jG+rVYqdnoQcJIzlF4h2v95yp1FVmnNDKax1
lezU6Vk4Msk9Hb42o81hBiqFpCODbQax2Y9gNmsNK91cbNbOwdLyFRomncFaAL5c
H3u3bI0wlc9m/7WRc1Zr2x/PAOMoyvjWv3VR+JSoVZELbLO4JlsowFWox88hk7/J
qGEdiguFqZrxe8f6Xy1/g0xHuJu1sU7H34D3nGb8xrlsK1mCBuCSK5YIdxW3/GP/
Wun9Q2+CmHjM6MeMJhOR9Y3ZJ16cTBZNS+rCTXxTiPlZaPogSS1TxDinE/i8IQmg
YMXKczKc9ssV91aBgsub1ZNN8dpwtN4dTdDiFVqAqxtY2rWGvwG00qn5eRoK4T+U
5ecfkllKrxUoUpG6Vxzp/qHx+nY5Om3iPVfeRLHy4mT1lPaAUhjH3UE5sNeRZ3sV
dvCVyg+aGi2m1C+/AhFu+i8N7cGjpW+g5K0WKiws1DvqABN/ua+69ba0wFgcvl+E
fhamxmEZQOPepeehxKDyLcxg5M5ULKg/xLxfjWbv4OvV9ottKrQVHV+aJDoiONzP
gEZKNyRs5x2DEbZ14vMExzEi+c3mSEN0jzv0Tw45GimuanCodGOwaKVnAu9OB1kl
rduEYTaGR/6dpir8lV/sanWH/VW82KWxmgHKE4uJ6CRw2DcHWlW8o/xGoxYRyDBl
Iyvw3iOQzrTHaTz+P6Hr+QsXrDsAxla5Xd5MAx3Sh+TD4uqcpO+c4LlLVvH+XI5o
K23y5FlvcR+7wlbybRwVsorytea/KcbtGI74NsmomcUC3W9D9yoZiw/rT0IctXl4
zcT0STpPA0MwTk6KYEDvE2KvA+BhyhQfN4QlUncrO4c97BJGzuwy1kBPJzwB9A0+
zK2jUqQ96fFmGTS4JoEZVYWyR27wlGXzntY67/jpsI15bNpkRlQnRt4Bdh3Pz5GA
fsqhhOXkFXQxryScGd40mVYxtI/mbbalxtYO40kvVGefP+2Uwo+PxDnBn4CZL3aL
J2BAFqlR0/d6GpnCMe/6WliA7MCm/25Kf7xd4oIT1D5WkoAh4t5RWprkpVXhTdWZ
94YLVu8J8H5iFhIOwJh0H4iKUUWcyM0JPNusdJk0eFp8JY85tDrqOjc4TBg/fROY
7TphhS7U5/dopEqc13IcvcX5x+lS3GC4nXk8sJEJQv/teQzc//Qo6x7rXAEvvxjs
I/wzp5LRTlLUm3x3/7RmA0fwQDEbVZEkzHPClTeB77beVussoSRARwwBJL5BNLrt
MmhqWoekuG9nu3eQ73ra3d9L26lK2kJ0CWvUsE/QEkmvI55wMF53GwqURpRoyRVm
6XyxZjVOivpNPlfoYYY51X4N899x7wQSQXB4WZ1hV8hgLbeF3rtCdcw/fgwLexl8
fwL3lR/EP0ghGSFOZfaYw8++m9eS/9cnaVbKKjvEL7V59AyBOp6YwLosTy7dHpN2
qVUfwWi/fCy6jl4a9qcten0Auajml1x6Sv4DPnHQMJeUU4iOYTZFaxKPRszUGrpR
6VaQ5eVckeernchJ/juSx9FhWnTphRwsd+JiK55TQA0V4BOqgW2zi5VvZQYRs6AS
W2biEASePF2+S++cZzjuIcB3efeJXEIV4vBKaQoJTEj52tZ1Ycwo14EwNFu36dwf
GzAwm/NtI81pFE3ng0ZRjDonkGFONR2/LLYux8xO3AW2b0W5NM85PjKtXYgDKgdu
7Zbvy+fe3EYd2l2LI9Gk43phz6X3Qp31zO57HHTlCINgeF4cHEywhX2ttn29AAo2
4hg7HjSVijz/u0I0GsjhY1SqPQzQjyKnAhIAte8INwppt22Wz72H+LZyoISPcB/H
5KPyi50pDc7ubcrRDv6Dd44L351lDA1w1uqgSyF/HqlzH/3+crlWz8BgpzjM/RpJ
16sJ6o1e78Bkh+qRua/UxGksCV5wLrUphvFPg9EDyZN9q+j/rNiEnv5+eC9/zx1d
aubLE2EJ3t/SPJo3VF2T5O7Fg+FVpxKkDZYVHNDY3KxMkp8qUrY+VyTIdVRRjJ8u
jebC8N8zOhWdJo+4DzM1qkz+N/pjBWc1/aHsZw9Dftj5fBoQjf7YIO7WbrzZU7bl
f5wSqgH1t0CpRpviyHbQmB8xtA3gzQPUtMGrdPfgIQFB/MibPkwkS6IhpX56aRh9
ibzYv4W5J54iO/jD5UhE6txU3da/xtGbx0EhU6pZGJy5zWAAzTBx/sQ7+fyfvcW+
6T+GkmDvUo88bEh4RJMlHfXh2MT62jamY52KKskZ9Kuui7X+CU47cKLpghmBbsaX
sENExfSHjQkaFZvRJSLOfWCloFOcKuEIE98m3l4aQuVaMpo4a3r7J9Woo9vdBQmC
+Ec7Enr3vHwio4rDAVlkwAHO+Whdoqj2FEhPFZm4pSttYqWdBWt3GtyWo83oOMtl
UCk1i/+78Rdj3EdzvioaofOShvbPGPw0mqz/20dFw+fQrWI2O8gXQLTV7RY7E+ya
ZDfi98AtT/WQv/TFwRT5zE6Fp4hhCU60S9E2a6g0L1z1lFa7Bov21/t6kN9F8ETR
BOwTfWRIk2WktbPfsL9wg9keqQtvApd2xvx3fSIyyd7ZAC3siE7OGF5iFewtcgws
Uo9L530VYOGW2M2+bcc1LZGWSSHZ+pfmBA0remqLNRL+rHf8LwXv3840OnKUQan1
2j6B9lYh1HZ0PnZvEYN5+rQHEpg1nXILalTDA6L+whg6C22ud3BNZOnOgD6KG/Vp
ssVqS+w/MyH1X7WX/72e8TwD661gOUmfEdJs4OKDahdB2icikG9owGd4+AuejWT+
fI9ByQhOMzWt0dMm7AXkA2Uv41DFTiDF37qcinATi/zw9RAh8YDzKF+WWLikJHKK
lAY5gLUplb5AcRdPDPX5GQmGxlm/U1pUOWMffCNyOTn/3v1lHeabJYG0sYVE+HWv
KE7yIJcX0f6xrf8WACHaEMST1+QCG6ySoH/cI4fTHycnJ+r3+vokxngp9nx6n1ag
aVXPZqfkE19+N6L32OzX8k82+84o2/ZgE/YtxbB2LvH9WLs9We04WbWNIolwqCQO
/aqnaWFhpJiFkoE9yGGiwib72eQw6icodLZLS0e+o66nWxPU9galoIQ8G0Zw79aS
ziVYy/hPMmVJxJsUuQYJefNadF6eqf4c80Ka0INqgO53eOoepCwgj9YHyqb146zm
a/qrht5q86GmY/Ux0lYHCnJN2JqWlo71cpGFPn4Je20UqWcOdgl0cDZIRxyxYsmR
8gDB/nPFBQjB+UPIrag2ecYohzzO5BF/Wn1bDCOEfn0wqYWXg++t0qccql6S8O0a
763y3i8AqKG0MuD8TgfgkPZeGcK4f5DM69m8rywPzeLJgEHEChWEOsVDWAjrlRPt
10xTYlQjGAUHmEzfaYNEoNl7zgEhvOesD2h7ipkiE3YiaJMgAQ6EndypOmYMIS1x
qpV6YhHWaFKU5kBlzXR8y3ZlaTe/xO1r65RYQlMioWQu1I0Tvvhckbtj08yNDP3H
9BFKzs1ZY5tSq6DGHabpI6PHxjnb3uGp4MvOQdPKtBXVJpXc8p/siLP5hkc/gOVV
tnTmQXZwC4Gu7xqbdu6LAmJYyFg7NmY7GtdO6bUCmd7ov1ENiiGmu/3sYIy/bb46
1Dx6IFNrGUeUXju3wB8FJ6/250ygzWgvDGN5XklPUNctwDquFIXZIlbouSXm0IOZ
YqcrMWQpCoxZNDFYqxWxRcxIs8TivqWj6AsvWDiFZQOJ5Bcpt4ydGCvwpSiuj/hi
pxLPYxDEzjAcH3fqbJW7uFjf9I5u+BWxj7SL7jIoCOCd7GN3b7CrwSa4FHx493b0
6MmiFG5F6WqeIERKzNwycuaNRARqXKOcCV6+muookj3IA9Y4wumNnS6H2qz+lhvY
YtD73u+ei9p7zmHaJYapHbVfYlX2sP91mrbjre4cLkGFLbJjrKWfZRneXcClN31m
3nIyFvqk9eaME501mbXxxVuHU3i6CmDJaQXyJQPCQEzvxHcsfziRP47Rdlq/V5eI
5mnn07OVXRX/Lw1BSLXRtBN6EqP5yuCQYTcjVttdd4tVolYuuo2FgzfKhS3LMGzj
sPPptVFVR712vx9tNEJEznj7Zm9uHt9FOLoh+LqWuFQ1EHAXm1ZkKT69pm0uCQY7
JqaDq1egzerzFZMywuis+M4d0JDJLdIMfuWsPQArQj0d6U96kGbBNYkhazKWtbvz
JcoJb6peH7CPg5KRgJbHT1xZt5G1JEj3Xx54ORwrQvaInlvDymuRcle6yBEyhM7T
ewdTRKB8r4uhJdGEp8WN3/UekcY7QNDMkBZ0wX2Lm10lENb31lBeeFg9+mAkdfJi
oebToTIHdcUVEIBGW8dQedjax/MLGR0erf1+E3WKq8Wb0mCfkihhGBOWomV8ljYZ
wIfpYg3hKEbAomyasJJHcs1eQ3fco8khazxwTtI3Uj899mrMJAn3dfZaiqKpWp8C
/5Pg09ICJ/3V39/9B4y1723A0hmXc/yUE4PXpiki3NwPZ8yYn2TqkgNawZFycPo/
VL04LkYDNubxUCt1jl19Tvm7RNltvsRN5ZO13wGZiMSfFzYdDWt0y1yqkr1LQYm4
aHvdHzIm9851zU/YmBU4i2M9l+6o6350nVr6DCBMosfGKjbHSRN9hQgEXUGLmLuJ
2WDyPPZkaLJTayqqPI1SteUti9dzpv/gX2pWDghbUaqgi/Af8QAWik1ReEAna9vs
I2OJU5gfU7r4cXQl2cuFsvnaH3p9kUzd+HP62O5uRCSENuRds2m0SgP9McBbmlgk
qWYVSHwsbImCXJRuzjMpUEpdIGJiwzJnAbbLSZnif4Ryf3i0wmnjBAXGIo4wvsFC
TpUq4AQ1abGJLZPExoWbN1PYzUPJzPmSq/EcU0XEccxbFUaP0wjT9MDwFvgsT3p8
8ieZ0diJTqYKGlN9Zg1qK40n6Y+FsDdYR8Ew01RiMATtxRlEGmpb1sVzuI+ddQ5m
zx3KdXZF+Sq2sF+m3/BizzAp9yqkOLfnkp5cK2+6/j1TCSksipDr0istMGmEWn5k
tzoZ9fUIKbhYn3eV7t9mlOYjFkxl43jYt7kvUTy3LcV+vVzJTyrUlOYE3tcxcIv1
gzbehTlEzAvZs1YPU+i/u9qXE/jH7xVzaL6RL067/oazieQAlm35M2RaAFqQy2d0
+t9EauIcMlGRjnGU6MzdGvIGYNiU3McjsWyzA5zYI/0APRoDzB7IpGaVcBRKdwYy
hSixEj3Ty0IhOrMiaEIGxqyeE/r1BSYVxsSAU2EwTCn0eYU2S628rn9StHiYPmj5
BKZWlsRZQXnf80WLMR3djthMPncdaJNb2Yobs5eGtHeym/3arTWLGhGtx1MWF4H5
hnn6KBfvMTwY431/EVGk2rx4x2exGgsfvfn/QZub26eOOSwEzT3cMjNEp16Bl+CY
UDJsDlw0lhVUJCxVWFNF4F+ehbeE/03T0eUe1EOJvRhQ3NGg8MWEHR0gBq1/VQ2I
ftBsa/8vAABbheP6zWaJauGX1br8D4jD+XLSwCXtsISB4NoduwiQobRw8Jp/V8gd
5d+VYX0PUJhS/o8pQFZX0W2C97eXt7Q/wtc+kzmdnpu3tEPPWF7tePhWTo65Pt0n
Pw90rPiM+sn9g+kR8i+LiB2Wqgl07j0oMP+OJmneMuQaKIw4pTlYFkI4YfgqBijz
9aWogQQWq1RotFa7DkgV9It+HJYgEX1pFT9A9i1B+g0RvITvpX8kt9gLPupjSzsi
/9oiDJ3vgh6RHsFgHo649QS+j8Ud8Ba3fdw0WR+ETI0Sz2G/hYqCN7jiWPvnx7IX
/dEijpEssPfarZmBNmvYnXAXvYEU7lSgCoE/yEM6vjAcabaF6zJoDtdT+6WDD1UT
K5wDlRZWBW1oBId6v+mm58CqE6WIouQxH0p5pfCvrQ7cbXfzsuXQGNEsMt8dkYWy
vQIZuThiklfaOR6np3vbf+VjOhjHgpcpywXMyL06n7SlGLtLMzGbbHs1oooSCm1d
P/48MZTf/th4yE6e6RtApmjTbs75c+FErRlWArDCXQepqURx+zcbDN2GSLsMbWQx
ygoEdoFl04fi5Z25EXV1ifIX8VDk10LCLnFCzRrgOz5p7AkAAdU4NN74jIcOF1GX
GxRJClXllC7O8xbb3BEq/sfUUjh1bN3aoS2p+sSM1m6g5+e/BVROa18DjCclFm0i
LB/t3DCbSJfcIbNfSeVmOiyVZUbKDhl946nSU/i0LfSnclQGIHAbJiC0tiCQ7mDy
iFyRD/lcYzPPFTYpvSsqn6yD7IZGFBxg3GLCrgJOpCeV3V0OPmAOgD66Eqbb32pi
as93yBG6ePW1JfLBg8A3LZWgb5BqCj3C3H84DOKrHgMS2Pjoq9gbwxx/1fuMiZhB
U5r2KlQ03asTEyQnt5YVenfyo9FKyzOC5OVgENOsTET/613H36GwPVZ6alIHAmvp
6LUcKbgkwvRGFoV+vOBwABPHm9aVKa5wbZMfYmLtJT/IrscW/nFg/Mhhb7ysRo/E
JEgzze4+07b/Bdtd3fDRJzly4OJjFkDsT5IPMT9e4sCappY5u3XVa96hntw8hHWy
DSyvoXFMDjIUUUKFx086ELYNw4+7XnCOkE7TDe2Owlr/31m4cXIUCeE6hRUz3UKI
iDvzqsMXEkc9N08naLi90ijBntc/hw4UZ/Q1q7rYI3z/hIhRfXkQy0tn1Vadgn9p
8YFsVtObBlpX1MS8lgOsd4+msLLYqDkLm34kzxOU81mZ/7Hanipi+LiZ+mg3zEgO
0CDQLnxhIURKU26Wddr7tfkAhyg8DWNnz9ANqw78LA+FtWcRXoyI/9wbzetrjGTW
vmCYHQaq5xnlpXiftCJelXt4s2MPL0NdOxg/j3976dtkPxNbwAcErohvdiuXEtNy
VxIqRqPpihQZEsYdjrjYNpb79uMvMznFypDNM6QeeV4H9Be3TZUUfrTZPjsF3Spo
wqhomMzOl+S9ewM9b0XkK/k7MBikrG006jEbDhH8fkgVNFbt+QPEG3l8XBGJWo77
YFfH/qUM1yutuZQwzJF70NaIqtyL+Ox9X4rFzlnqtWKJWhZKfh4eaJ4GHVU+3dpI
8fODoewjnETmO4SqXFlnsFe1eHcqOuhRVKPxB/+/EnvZ3YJirv1V+rcOU4feA4F+
X6spZE5LA3hcSfAkYthi5RJTeBPaRPJAAHtMduogmcDvfXclDtDj/WVr6Ch7dmtl
816tudVyUz4S9epFAWy+GP1aosQDTQ1oyygKaPlAoOeCBHhgyVagrUSYoFtOQr3j
05z96tJiFOx0M7/NwjQ/2lMaFh3nziMjpw5sS+DeR38QqftPNHNiuGT+4XT946Dp
nzBRT//1ErB+wrE1oFMbHwvkv2kQe8k7b9S7w6X1bCdT4bGVDUlb8OU+s85WAuPh
lsKYhamgwDrAaYMadaoMjiS3du7ruzxeSkiRhAPnTKMzu5j+dqVl6tlgcqxxQQz3
fZeRXx6drCdGYgBJDo5sKcglOQx0lmnMfqk73ugJc/4JVdchpzqb7DciGNZp+VBF
bLbVSzFAD7720cQIjpuN+H2hLk52TTfgKypN0kc7gaH6UkRAxlcGvmMdPu4z2QtD
S+Wdb7T/VLjeSak21AOP63J6rpB366rBMs4HpDxbLwROxGS/kveHWarExUpB6ijd
/EUMf3zfEW7hWPTxhC3DbxzrMcW+IpK52G3bHa50peSXzduT5t8qjQOL3ofx0hXs
jHdkucuiYHD+5G7XRC6fnL0+MpV7ibGwkEcVjpl4A86DzHUpn3SPtuKIGFDS85QD
UeKdY9TvpFw0MN/xeqh6KZ+w4U7GMXjm/zluuc3WovMYw9m+9aY7F+G4OUE+r7oH
3ae3wEUIoDWc/1uZtDRkTJdlSkoq5oCptioacWFiwpBob0toAyl8Ku/BIuxsAuJD
j0C/VuD0v0jcjebwbqtBHiLDqFSmGA9ytr4WIYNjh0CSGehVKpP7iCAJpEkKRgDQ
c5edHpSWbb42zytzN3T6PzsH55l4rnVWs/Nh5sPYRmfJsrhg3anrPa48gsuuBITl
ZCpMlFc8qIMgygOOy0xhOtl511Ksh6IiC2r/gUNJbUJEb3HyWeWGXW0031ALi92A
Go8iSM9DGmuamy3ULq1pk0HOl26jO+x9XoAJ9iwy6RMQbR5XOj7+z7ZiITep2ih8
yDgCRticjT0SMUL6aRx8zOQSGH1ly88ywItTxSa0FYiqPnM1BOdhN7BqnvX5kOTl
xlUPpfKc6oDf7w92ZOXxdF6ZH7tzexKKr4uh9ysOIwXghqwZGPoMnleQ7rhyBHP5
pnCdHIiBUd+TEtJoF/9HM1NFKYg64DKHgd5z7c0gfyYxQFv6LlT9mH06TGBrd+4g
9lwWJXABSTuQLe+b+dM1ymPEjWdCeqr5gzgZjRY7ZbYKZTd84EqmSBuX9oJMJvEI
XXHBIphUt+JWEQSYo+u6x578Pda28roxW+M+Eahtr5ZiSPazsYk3fTfUt325kAqn
nurhdmtgVx4/5wmH80phPyIGrsXXypLo3i9wy3Ue3pHpEeKc58tBJP7lPOqSHQL9
Crikpa9z1nyYu2K9Hk9Lxb13nFdV/zd6ZOTLkVMMcomfyJQVw5/kvRrFwAbgklA9
8S3h/2lTcx1KwV83bUxp8Xb8HMugDUKHJNHItO4exe/uJOUIcbwfdmTk/2WrtWFM
3oeMSx4gg0oXrAGUaujkl7rw8qDjePGntMDeYpxNal23xBdIpXejvPK/CIrgKeBI
aHaNcI2/aHfF1AekxV8myjfGu55N80QMARuU1nrBSrErYlJNSxTPbrBeOSUBpEID
xHcZL+fUsllIrn4lxb1MyfHV5jcJ3C0voOJnSGHzCN0oj7nkF/AiZVEeucMSvNoY
7wb+z5qKHVIph4YIeoIghRrQmBQRuskhZ7qqvGnO03b3jUO15RT9gTjJ1U/AGtKH
7qHKvZFkbD3jTcIil3oGKW6YppqHyqVaWONPyuP4fOVLLtW70hGKUjQRLv8Yodkp
JKLPZWKQ3Gv91htUVngMtiVAfO5hphNixsdywi4AVyHhGu5PgFFqbVD5/LeFcEIT
Vzx500L5zvypdwjCaxY3N20Uk04b12/6ufkZYiMvpwPRk4vptSfV/z9rA9XEXJJi
532SKTHqOSMC+UnBXWEFjIMlpcIXhG7ib7Tssg7Ab6oi3GfFvv71Jn3ct1HxGWcw
4kkLDh6zwPrbjwGVJKnptZyz60uWnFO8Y/Ngcs2C1Qr3cxFE3he+4CfTDvKMweBi
JLiEMF7j4QSEdsVNr5+ORBzu59q/wLkjmGvbd1wIgWJfPq9B7AZV4kl6oV9CLy9k
vu4N4YbshnaOcXFpxpfIqqYumhvGRB6IB6uz/SBT5WVdh3RrdCsneqoraR72jgdK
Cv/E01dnS6mJtbQYVQR9AbY2mqpEAYRr72rYv86OsMHjRybcML034oe0K+PCnPjr
oh7cYrOHIasX4/BhQfdsbYWm3Hi4FUsAHZRXHTW+1Xwycbf5IkPj8HkDfI3uNnmK
SUNEPxgA5aqCfaE2Hy/yFP6rIviOpM5Z1MN7aPqFWiV/FH+cRWoOOUxfur9CJjLp
4lzTJTzpR32iTe77Wm9sivDGZOHtK+kW+1AjxlsMUBLa6TyFTfM1EeOlDbTytKNC
P6cEmEp5/7E0kRzQufN1s1QJ4dmsuf0Pbg377wam9hPTW3fssGk81Zy2MsWNyKmN
PrNuTMCA7/o/bOd8Z31sZlyoqXsYKzk2d0v4DzTtCv/WxAapfUX/lg0C9bfqKylh
3OeExW+ofde8TrdusEwAkQDJDHmaJTFT2AjqBFSu8P2Ij1nX8bwWEt18uE5xXkJm
yvx/H+69pzCZpo6XhB3Lb+byIswN1Us7sa2Ech9awbFzM9Vi57SEhIawzlZW3eKo
EJYpZdHxJt1Sf793rlxWCW0gZJDnRk0FELk6x6Z2BSZM2oGKLR8mPLCGVJZGRYne
L7ZPQXhXNbddBLfPqZBLWay33uvARULUfRYTWsJ+hM8pSPjEQMFdEqV6f6tgigcZ
va92mpz2i8JcvzNrjMSr6SMVkN2LazwBMEl/8uy3DuVAQ9ij7eckalA2t1cqrdcD
8iwlbcWFCNZfSAdGXOjOFdiKOGoMrL8t6luU9GPIOuZqBFZd9N3vVSFYzj7HjtGu
UYBb0oNQ6XSNYMaYwgtLFSitWO3S0c8K3YRsuUXwwDGf91wnnaTokdoGZb3xUz7E
cwhSZ5vo3GT0dsPvHvqQQnzr2Gk/oZkyv6vncr7WWhrvCKMBZaRtWAnLHAWpmI/A
AXQ9QGQ/LWa/S5WKVCBXEe9iSrTdQjddVccvnqgiVCzpkMGxgyriFK/EtWoxIfI2
3/bw681UZ9Rbc86C+cB8aHwohtkeUHxJc0VLZwo+Sn/bW2aU1cp5OJap15w9irCP
+YBh5MjEO1K0xEgetj92gHeupOPRabiy9E/yF2LRXSpg8M3kORkXnSXF7rB5HlnH
4jMBM97cALwzXYpEFrz8TqAnhqxqdQxKziroZzCWDyOWAxm/g4qX8rugXEx9WD9N
bRhM2fbKJaxsePuu/NUmXbfgNe8MIEqMGRFTpAs8UVpMLC4EnwwariJh1/mLu/lF
wt3XxaJobtya70H7OC6GIzNeAmArDprCPoI09l2pygba7K5/J5uZpkzBZk5M8pjp
lTIZVc9ce5nj6ykgVqLFe5S5i4s27Wt08mmESK6gDalDNpHLTL9zh6+aXypDGJvd
2NGPE8l6E638xTUczZnelMBTn+Kk2A1TyOSlDNyGS5oPrcNblV2UTU3og/foDoBc
UOeditvx+YZjd8kg35I2wzc/Jnf0ucxHWUinoc3Iq8qG+ECC69XkaD4jn+bhxBJ7
qJWwrCmi0u3y57956iMnihjN1PTRnsAwjci32u/S+/fDOuZ5IyYV/VRxQJV5xtOS
CYlShQRxo8VKdwAxHF7dw7Y+86p0HfIrjomJkwfMLKwj1G+BKhFGIqTeQicvd3QM
CHdx57a8WrNztYfgSBssC/9YkIg91p88B3V17eJm1Vow5u7t9NhJ0qKm6SvSe4+B
l7sDMI1YTkzN7MT3zIjRwtHitW1Jq42LWj/KNw5mOjHGnZ1tzbCm81qGVW9W6wqS
a/DGEQyEZJgBr5ccoO4jRCg/m5TJg+7QEZ6UCqPBCv8h23WtXunu/Dkti8FBgkY8
egpgwhg8zTaQWllVBHf8Ho4MKCGrbrtEoHivG8mfLZwGVqk6DqJpztfy0MntWODv
UHwoTJmN4zbyx6HM9qUgzs9ze9jK5wm/GXL3AD3yxnpDLacryHIauvfsuNTClm1e
sot8ANuR6INO5ZtUNVBJ+8hLsGsxP3U8W2mwoEEjQZ28X0gmGuqymNhXOQ4YswEE
C7pYpi+T5RnkMCu2CeRiZvlgIe0YsWj0joR2CFMLs0RPlesA7LhQueHKhvwVtwEW
IcdgB2tmNxkCFHYORrj7KwXU4UHrhqaUv2kiBbMLx6zDiYwDrjKJgUAvEpAJ8eW0
F+/ZmDqgXiLCbVmc0Z+BxZYUI92uckD9Lw9+3DtIQSglZyb5AbCHFxodjxjHcvlP
aOiX1xoF0F4+LNwoImj+UmTgSozMsAqSEVWn50AKxrGAi6OCprdQjVATWJHHO+Yd
np8Pj4Q9R+occtbhxO2STsHMKQeEOVrzgQd3jcv+C7ipltlSmpZJoDqceOue1SjK
7eNuF9JH+HVRlhLdW5Dscl5StlAlV2B8MIkcSwRiUVUOXTlpzlvVjtXFhbLgb9VZ
XbsHZwQdYqobMVCLHu/XauyMLzg66M5ofBxMzluAeoj8zPKITYfGPPOr4d/QmwX7
v/PaG7tWO+CaRnLQhYxR5szJowIfMcKhDg5/Qh/4vZXh15xasU+81f7shZNeRqJM
Qd1CfZfVa0x3yX4skrjAnz6ofeqI71b4r18uKVgpDAVUl4F6L7Cws50FJSg1gSc8
f7qhoC+CgV6RKf/dmr7hVjm/z62FPKDdGR5a7/8fXZjApmPiQhmz/bLVg73hvIlC
0fVPZXb9yTu4G4ZuTFW4v0rp78HiN9LmgHqTImpzTStBBiJixUoZL9MawVfDKVf8
DmGgiEDvqnC0CAX8o4UqsojfoFYtI2aIu9tbFbiBPOgO/ULPMrg0J/gfUDnqDmR/
PXPKFHrP/RboiaOONHj3QnvuIVuVvEhdpg4r+vWWuyOkUjmBHsog/YoilWnIy1gM
5/JwXjYDife3kATYbIs7rf9wu4lABqkVTOx/OHKl5roAKHyGX/NwdW9CfLajY+1g
NrkAfBh14l2x2DSf3C3E3yUrC0wXs5DHvVEsdykNJxoRR8W0R8XvTQTNQzRmCM2y
A+31M8K6qhtLsBPfuJTyOS4oD+5OLCAIPYhYq08d6MB0sFh2j0J/n3CkcxsO6oPs
3OIdufJajxxxg3QHFMivXAyiwjBCTcpkGWAToFAQVSsEiSRhnRozUzHAtcaSwcbw
Rwj3WpZPBLmcu8EVpHecwPj07eAwioqFZkYayJDi1RgBpGaJ+H8xo/l0hOyO6vya
mZvmq3wrZCUc9RAI+0xcZUKLKntSPX+qSN+gVwEMtB8KOcrLeSAfPNXFJBk0ooay
S9B+/3dZcovLEx6P+A3s99KjYYw4/T2uW00BARH4worziW80KJAPEHWZEd5tVapC
mf4wScJHBjOHacvlfsI3XjRZJN6sVzTlto3/JmiGwaP/ga/hPM897ymTXIHOTnF5
DiW6OOw6bNiWVYdHrsHo1+Nv4aVeQyVeXuJsPLRWHpNLszrUgaZ/FbCrXdJOPudW
8UKRXoYKFnoeaP1zPsJqwnKT+uWtEKsMEY6kMrnkWFBVuoYwDlBWm1xujT3/JmeD
ZhPmyF4X8eqqGzWi7MT6f13x54Kn2y8vaUH+ddqF/8QzZMSXchPWTq4/AWJI1Sgr
uFZYAiXKl+aci/CA27LbVK8KW+80reZqfCvOGNNCGtRDK+BtjM+1Uvg6C4Qw6nNG
x8kzJ/cRD7Rv3PGwBqxv4MO7QrqOd9D2wl/Mgm2hKCodie99wLQJnWfAQWJoFz0b
00lKxkhaXJdPn/Eu/k+m2zvxKKtEBYFki3DYrMLJ69NrO5sld74gIU9Qg75gGqWk
ZUPX3uYzwncBkMXKcr0H9pDnqr8voaL8/6nIgV3eefy+x+98HzmGgUPNUWxltFTY
58cftlylJFsLz1lwGsKh+KQgba508T87Nc94TOJs9fEXWiF+9iHJjoDWV1kl1oyf
Xb+9Z7Bnr7w6gOP3iX0zMaDPwGwNQK48aDKI9dN19518O3g8otUAzwMJnDu9bvxL
Pe8I7lZXcrJZxPL/hORJARPQtx80FbOC271aJ1yiUe6PPihODdq357r/I0l9ahxo
ESieOqHqTvrCsoYoTduKa6dcEPFUsWomxEt/gMSTMLHBjUlurSIMtyldV0CiCtIj
iPCworYsOmBrabh9dS9t8hSG6t7aZ6YCmGT+Fhb6a6l4T0JeNqx/uWrviaNJDowk
ttiQY+9G2KwS0XTqkTxBkNgHmxQHa1sqNFU/nHFyQplBFYSxAEQsP486hzHydgHa
xlfuPtdDEdVdfxgMxo5+H+fG8/O+PcyiNLM6Ql6F4ko0X/TGYKfkImTNiWajv5ya
1bZ7S+UgLvKVxqQDofcEEGiqGCG3sGUr394WSLEpPePo/Sn/QOArIkUclju0y3ky
DYFi2Eq44GrwvnNxwjKbWUXP5byFXOP39XXrHm1tzq7epiBXTWKvU4Xi3r/HB3h3
8c8g7aanddMzLpenee5a6K/FkXbbzNNVXryHsq9yB4gV8AfssTgd5LI+0OPzcVWn
EmrcdYBXp2M0PJJV6HRmKu/i8F2bEezv6IuCGBPm4AU9fz7FXogolyd4ZV6ASf71
rtb+6MPG7SAlAeIRRLBOENdtvGGpJbwBplE+TyFm0oqKTcEgCY0YwEaNcLsuh2Vs
w7wmQ2VV/RpiC3mCIXFKw6GYJyoZwnAFGJICd10rmI9NBBc3MOHbTeF5oX6GBsDi
DzpTal/bI89K8lKLKq0FhzN6mgdiw+O8I9WWZ7Kz1bNM3nOvZbfiVr0r+NprtYee
HfmeMAa/RbeoEsKSO5A+iLCnahvo2xAX25tH8D6LVzAWpqrXdZ6ZJ/78ZmxBpgao
h8HUTn++vqZLMKhQgyldG29CkOTTet9F4wuyOldCSVeBnfob0PVN7nXeiQ5Gpo6u
pnq3dqXOqpE3bKGew6ObVgoM4sCtPIzdL61jXz8mS2tlewI3Q4apsxVAeXpUNcmW
budu6VbwYlDNqooXupNtSXFLD/iGaM5FhDKVGwNfJKjNjKZQ5fi++Euq+eEwQOvh
6sNzHNU+8EZBg048fGvzW5hhQKfs85az1lb6deuJqHz0wQ+o0MeJIebJGnjNct08
EYIpX+G5CuQpItELVNhQ+zHP2AR5rtQID4X2rlh+f+3icJXXfck2pXGQ0p3uW8hX
k32iTBpmrhW8Wl3KXP3GJ7wBzaWBh7YNFquiBLFE3v0lqw/alqkUlVZvgHRHfX3Q
/EsMRU+G2dge8RWgG8fhf8jeUHDtusjjDVxiosiVrfBtRP3nTPRDskc5SSrG1Uma
YtMVwqAtbVs7gGGg6e5coe/s6RRZUMn26j4UQMbefyyKeeJjjAchOA8oB+/pxNrN
mcJIP8t4VJbZQmdAB9rwwJgk5h15PHddEzvRFVPQlDrrZ5a3O8osMjlTV4qVjBtO
c3PmAiBuzQ8VL2Kyxcn4no9hvWFBPpQPze5XVcbFzx4U05Cp1ZgKyq+HZiVNMfvN
A1SrUtcqbDHtAdTb8Jlnc/7pCO5E2DJeOrFXYkoY/z2Mcrt7pRLUJHK1luOTvWbI
VD6aWHBjnBBzgsWzN5GqPXgrd0aOashelgm5TgSqQmrxN1iOqyEhJC6PCnkhTBXY
NuWeBWo1dWlFirQRHMyRe1nZTluf7AWDQb0cdFzwbrGWk4u0Il7vy0RpJx2HXDUe
F/O1zEFRg5JfUA/g1wU/Z5nGwdUdTeAjgG5IQG2qHOI4En2AanuDSy1/3Ttj2OTT
ll8G6Z7aGJkCdatoaAE5IdEwHuH0sL1LHvIScU6qSBryFfPp8hoWO/Qsp9eZ4j+R
dKUmZrWmPL2/tbHR6NcqGCPazmmwWofOX83T3eidDyA8MODO9PyjZzW1R/0TCFgF
C3ZC37CRsbQ0o5ARqP1Q9GfgYblqY2zdKihm4pYVanFJoZ07bjxo2Z5CcoyCjJmD
/mP6gA6np1RM1m6hv8IRD750UhbQtHwwIMSxA/lkhGH4Xh4kgLv2us+5ETonN97a
uQnuANiR5k3TJ8I9d/KnM3Ra3CDXx/QjMlgT5krCaTzi9ha6KyMnxibjxkl8IPdL
psURVVDDGL4UKAeT2ZE54VaXX+p/eU5mdHWbTCWcNDFntmX4sGxdP1DSLERTL+Tx
TYvXFhoo7TR+6acjnyNYRLb0Xp6qk6+cwB6lT9pwYACRN/9AY4+Kbi3ta/j+I7uD
DHL+fMUGjFpiB9GUxBQiUdo28P9664OphQmbdXkS1ZiVfPx27Ed8EwD60e8regPF
67eMW6QBxpaSzhAGOwCWoJH/BVN7pF10GzRfChYAdVfAgYBiEPQBROrjC4KG6hPJ
3YwysVH25PoD/A5CZwy2A6f8ROEFOhbhpFv9N5Uxru/8raGasSX4zfKSEbbWOSbT
+uCFi1mfJnIOlcR+SE2Bza4dB93rPuXig/D7vswDJtvDGSektoSqezc2Q2PCGyoF
lY/KBP7QsZ21g0KKlod9WwfRORi5f5qKONza4VThaJyFsr3G2pQUfkj6RTYM809G
pSzCvKIclXyKjR0Hk92oca/Y1zFBkkOm9U2G5vx7XYQ3nUwrM7wjkuZe/SHjYluB
lzVWhlSTiF+WCoDTXcgfMjKXYcqh78jzTa/VquNZ3TuyuaDkllWj7ApotVkD5zV0
dttgYCU818U4qJ3Dczwu5Pd92W4R6qfjalcldNenyEP7QVMWoEpLwpzmz3CL76bA
d3wNtIHK+++jbCnIULBdb5eOzKe44QREK3MPeQ6WKcmmsnkl9JNZfrCpX3Vdk2a/
GTDifunUcQDIaEjG4Y2VNuIpr+TvzQKOWfraYtlwIIgo1SiujORAJPnTDs8TB7lA
C8xm++dA7WEp+F1wdq+2sUTgL3NF6TK3eSb8RQ//eCgLsX0EaeZZBYZZMnuaLBjQ
mB+INKXo6xYWyhrJeu9fR9jW3T62tHvgqtSYZb8BqoeEFJUMLA3nXcYarVaZP2wo
5JCAQaArygledF4oqBGQA+Ssn+7dBk1cNktZCCs+ykrkHkp4ZIey3eQCRru9pFtb
DnVSyTeIGnqRWjjFZiDZapeDpKdKQYGRYoeoOWnCeWgMTfsbmdoyEAfykzuq8L5x
hJaNp+gr21pI71aX4cX5rs3rnsflBrTwZFVCNBKgY49w3qGY+pYdzj5vMn1G/ais
DrEuQv7lYBjT4aQcB1TJRIa9z6Z98uNRZCY9fDzKKA7vB4MBHTqJzAT+lTtQp9Xt
ubgeZz9JK5u0g0neiQVzD+JvzukRY8AXh62J20PKSxG0PGKRlNICg9sS1DE6GRzn
hapd7x44JuhJ018bj9uDMvhDH7sL3PqHg9ZZKQKdIYdRLm5ZfBXyXt9XX9gT0Sg5
g3IEJpJy8R42mmMrbheFgEAHt1v8Kgs5wmzzCPTZTcfmnKrEVPlIlp98wa3rAEom
ZF+uxPMu7CJHCKISGTCZoGB8P5JF7wqiO9ud1R9benDiygLB0lIl7+QEJnMGUynw
Z7d3+5O/bd7JD9IUSOoe9emdH6Oo/Nd90KbUjKFubTuRTAHMFggGdMDFWkXkR3ZD
EPkIdwsy6MWN/86RO+0Hl06PLBVqUuVxyG1n4Pl3g5wmjDJFGXOFgcMwHdH8Qu1C
rRsGlcFDE+ZWULee9XBZ2hg7hHdzS9553OrFUddSI+/2Dh3rIbnLXIDJ7CXXHo6p
Am1+l9xY5yEZy0lo2nk18iYZtJNao46erocs92pYSE1VEEQqQi4lsWysQehScrRb
Jw+MNuNrjfkQ+jsRS76a6fQZJivxbxX7i6umHV2zDF3a5/KCa2h+x/4nE3+ImYWl
R40q0UII+0XIUPWapKNml5oSxHhUbTrHK0sq3d8tU6wSyQnOnxfevGjcaD4S0tB0
i3wtV/HFngE0K3669OY028Ns4d+8pC9TgXyGiw8RHbBetIHo1J3tdzEWZn29r74Q
0PD+ahavPMOwWlClosaj33wGT5jman7OxKSgJe3+11aKTeilpFHtIG7PzESBhDjU
yraADmiLoPkXVOMtOEr/hv8pk4NeAODaYynCkiSqA63RC4AogfTRXku3MNUPJ8jV
UxVRWNo/sdDx5BGCK2ygFSZT7pCop901PAQePZ04gvV3M9hEleBl6ENUltuxHx+e
rlaBgqhjfbRWnn+5C5BO38QMlZgSlceLY/3VkSFWZz5psSXEjZOEjknVteST376m
RwGkjMSwF10Gpq9yuRQftuObtnm81BbhjPCpJdMAhh+QIH6dDrwhnNP2osa8q4oK
6VdgQcGwWhvUgyiX9xrNgVFj41FT1n9PgieB8NtCNGlsdFeV6cizgvyMkMQu3Jzk
PD8RYqCWgVFI5YxWT5oA2U+Z6Nev0617HjmSVJNnusRSiRnOjlaQfHSpmY4Tnc8W
QReBFZObSQXlSDSrHJGkElRFxbN5UisHq8X0OlpoAzTkOzxHnOJ7FCkqp2gv3WnC
1XDP+TGOA6EnKrZqZogXj2qUbblxadUoTobENKvk/CbggSYNa4wovPUKLTbBOEOw
5xWmjUMDw2if7fVw4r6Hb+DA1yGtr78QjwTLjTOUT2OHO+9+jOfWjbpTGunsnGXj
O3Xye8iK+V+f+tsj5jsTw2QPEhVTZLgWQuG5Q/hfOT6xfGllIELBo0aDQbDWXmQe
VmeZ88u+70HsKOYBpskakV+OKHK1tlJZTFBCcslmJ8wkfkYXf1J44T+EetcTxLRh
JMr13Rvhh6BQ+ft5IOQt5A5OuWnd8R2WfJD/eAADSWe5qWex30R9egKP+sz+hwI8
3D/bj/sUNdoD5oFERy5c/VwR4aQxbFBI3eygI/KotRWkbGJNWNqLzIsQ6v9j3Ek9
ho8cOQXENS4NE7JolzT6UPUUqX0H8F0N+9Xc56oeEp+BfMGJtTrW9fvxnHkAgRyg
dgIO9m+Jy1iuD34MQrAQb95XWsj4A6WmRXcq8H4PzPApW0cUQpIS9El+0b1LOXIh
9BO2Qcyf3HQW/Bdt7wpxqLgMAtJQ1+0qpv4otac9YjNrFr4vMORSALQnJO6EoG8x
/DtB8CL/OtQA6CZchpvOfVprHeWdeSGzhqkYnJS1+XQ0wk2xwnPobBn+Es5v0cZ1
5vpoWv6UrgsAxmkwcwtalM5ngjYP0MhToqw/fMEULaLvikTnx0dogDLKe7wAEuwu
lPcLwpcpToUFUtZWEy4BtECR9+L6hcRM+QcFI9suQLfe+gsWENLiVn35i2dzQjhg
XYwlJb+Msf3+Jej3UFcks3VIRs6TvOb25TQ69oswS1DsFZYtfXhOLkaiA1uDxRXn
RI1WKkbbHljatEbEUrduydeQA5vxAlk7ZwhHbLTotV9eQ9cJeipmD32RtB7FTKCH
Sm6/qBDpOHGbwkZmLL0xlW7Lbzv5+lBVA42LqQ0LPhq6XCXBYCmVMP75FlKtFijH
OKyHiG1/QHEN8+xON4cwzbqogXL24plV0CXv9gmostV4p0UMENc3B2qHv06BAP5B
w7A6GyTLJgSwXj54cWfdRRbJAs0OUJF4pEr6giitWM5eE3MXiiLf4k6kFuWIR4Hg
QvTjeyDqWJI1UigDDj5wrmsn9tpFiTcs7gQhUKQjclcsF03WYrwe50MMVxYFP7HH
U1JblHlW92izExNhJYe3kMySgu390qfF+TPuG8I1iibjsTFbr8EjqUmogBJMvxtn
1tBkr2qbHUvoUih6T95qC6myVqikMe4eFDDZzqaPh2gxQdvBsH2kUzXda5GXO6ux
oQE+knLjAr4x3EusJkEkJGpgPJwEOoPddH2EBDMrXnO40H0EdsB+BBcPHmmqaI9g
pi24HarBwqSrdsNDIwo0LoKnTI1e4blgklPFBPooNDB1fsir0ZRkixQF4WkR31zn
JsgNZ+qGghp0cnaEc+lIvX1QpyBhbg0z4RJw68pSq76aZWhOjB4MQTwS5NkOb+B5
0eUde39Rnft6WaD7yg8AvhVAi1BLRRy7Dc7yCzvzXg4SgZmCdWWTHquIgifkRAVP
9b0yEYVASQFmrsBgvCPqPi8TL3jgKxTyz1Cb4xir8hqIvjGLLuyLWEsi+xGAmJR/
rHO9X13a0hXCXVURLX2T4iGckMTN8kGWGRC8chEMy8Uv4rUWDRQeSNo/u6BhnqHf
/A8+7eB/G+vGefJlXTWpLgsUemjjc5noCxXzjh1coaIReSdCYu51dAzYqiFdvXp1
OQelaLMLQjar1ArgTzerUiLEiLD53nOsbmJeTOkOcjN3wv3Wb9jg0H5ewi+2L9BX
JICSChikmEC0PA+m1z5pm0gtgnMRjiufqLPVughItFirA3hTaZWkYEI3K+h3VlAs
m/mgNTm+QIo/Dl+maq6XBsOjNg2ilBe/PFnqXto+UPcIIe6OjTEurGK0M6aV5ozJ
J5itBVLEFeqKv2jzPdtAaGvHKDGs0oiNi3H2xzceiJY/GDEO/7Qava6xxKe4e9UN
TjXsTwgruHAjSIWmyN9aD2CdJaOaInuJb6ZnS0L3U1J2P8RiXzkknE/nTi30S5fn
JLUkONI1dlQcd+81CInyi+x14/SG1CJV9OtMypEQvYGezs5UbQ7ed0tg8nJKo89k
6AftpEb5adrSzHNBVnMQ7qvI6QfTnHQgbxiHTa1lULIiD/lAWBgjvuQTbK+YNjQe
kFopwiuUgqZ0lnWm2bUZl/IQ6a4Hnd/Cc9u4bR7lQmQu3sQpKFWTcA3IdGfROzV1
xbKW/d2YK5RyWZA1ZtZ7fjp5cXQhphQQiCskiBp4CwHD6y75kCZDvZJFDsBFbRMD
hCIg8pWgHikjUiq/IHOo5wikeUNYO4uU2C6tx2ZF7vLRFHtCD/I8Gh/5xRiSb1o7
3F6qwZWbBu6U3azlB7F34aSdK3ZJSHX/lNgo7/x3Fz51JpEn6bzZ55bTWvp/pzKZ
tPE42rqec8om33mblOSQ67+YDPZOtuNOBusxeoaobuw82V/AmwIsULrulWiL34KB
3eq4ljw+GlghgR8sKgFV5gzVMSmpYkhDSisKkl2Wd2EoNcRf/CwsvGFLyfNSxlli
cVp7YMN2bcX9oMna2onkyHfIYYxuK7Sgz6cCJunxNPfTSc3mCL6ilBE5brLxx1lp
OVdbRNZJbbj09K7oH6xDRpzV1CPOWfAVo2F0QV0pM+YrUWuTawLQabZEovlSQMQm
O6lBX9mbs3+BxZwi0m+9w8pEivfONnG5RxgsoxcsuQDq0i75vfY1S/1g9L09MkEu
WxAsFvionPZhNhPK9eoO/hpi6BNaIA7+iOzY2szfGeaiVP1082OZYUSXKdHso3SR
5fHA/ensSQ5WiOuAJTfPPRjmsv/VUdB6PnnSMwxWnkvU2AnImkRigWiUGRVXqjkF
20OaSBFuqSEAbT2njRZ5QKWK/15dXSRikjG7yLqbFPo7L/0NR5KWYdFjAbLHdL8R
F0jSY6HzSzRiZcD9CZG4fZqIatxU2yIc2JSWKUWjEgqJsuNCGciLL5DZsMXAEJV5
SEgLh8CEfcPaSKL9sdTf6AT/+HHWJisK/SkcALvKdDu3CheNo1gMkMh15px/1dAy
c2dfKkE3wL+YIX3yQEHij02OtMMji0aSZttTwgkwzIwCmf1hUCzVCB99pes1L1Nu
hCLB//ZfEj2/nI2ljDvCRuoKFCKUpp9286MHuafFOZOEEeng2tuDrHNJ6NdQye7b
xyLo0kMYMGyDWHD0d6jUYlZDFP/9qrKH7XSVWyjr1098e4I26b7KvA68WNXfEA+V
pw3qGEjRmz+df1/uiMn9f++dUZvGDR9Jtj9l/F53G4InVzlSMepSD/mUfhg75yBD
B4kKoIFbpMo5lhGPdMLOGUGqRUHnCnFWtAwXC0sMBibhtvHbp1UdDgqOLQSflfCX
OLnMfd4VsepggbW7XBtSOQL4D77OEDrWIP06MyuIosa1R296/XOMMuPhrC3DtZ3w
HK5PHao8EQnK6i0ieDmlWG4lMS5nqj+RpUBzW0L/I3naQEA95HPRWVyyV9UVO3aD
HFwFL4D3U0aFlA4qf2SAloSuJsW7S3762Epy45qT9bzWZ038zqro+x0/tWy5dqmf
zosSyiJDbV9BtzgnRCpmSJUwkv0elVIEZPvh4NZqMD1UwwKYxTbNYFj+T4mA4Yqa
snOV77wq9OtsRnT4Z1Cwu+izXC7tn44OkXlqwJDN1w8axK4KK2u4VNZMn5AzVqdg
Mh0hTbGGfDMJXPfAuPGSmSvd8XHgvxiKN0NAUt1g/ZPfW6oCJypkpLohF8EfMmUR
9V9etXc6/bttjpKa1D9dP6gA878o+cfgTG/eSWcJgQvlY+j48hNELV2C+FD1gles
1T+DpHB614cMmnelnmXdMHK2qT9bcwXkkKRrqKtXYCjUOOBf2I5XpTMqun+E1K80
IczLqtbnIO9R6zPaqmHif9n7hlMqgeU6Ut3+OgrUk/mukNuevc4yl0WvG/rYaCjC
VJKHzpH0QiVVXMpPuenNS9UQcEYcRU625QG1ZfRMjwsqZin5N/30u4NjPFZu6sq8
kInvytZ8wIkRXQBqho0FtiB89EiIIJVGKqgA3MQWRBwcty88pqHfoi6by4t2FkDu
DpJwBERGFOlhwjKcv7kK86EDDiVlf0+aXHNuhSpSxOyuLwQMsxCv4qyVQV7uQhrm
iRBWQGUVkG/zkss1y15fVM8oRWVqmG3vRdV++Kl+cTTQZMm7/7XBCC3rGk4x+3v3
1PakQw2/ekb43mpkGP9165LLQPBuayBH5Q9zTPC1KiSCKTc4AEIdTgAq9zKnAKbM
7GF8mc8kkFC9xpGszbPyQhrQG6+GDZcb+mfnyB8bdqIDeCEYD2FEb93IdZZaei/L
NvVRWe6SgPFdudlNsHSP6oC6r+a2n1JFlw0e8pO6kysf+Oto96xbNNqw2gHYxC/y
L0iv5YUGuQY/Pr6fSZK1/+WzwKDtegpo0dmn8xjE7aK3iMB6+MB9DgnOay8iS6Bn
zs2byLpF21nxdSs1Iu+mtmKqo3o0MsbFnGAsLY0wrZ8PnPHSLat51A5pDO4ceapF
Ow7bTxoJAkFn1W7et1xbWjPrBQVJBZyLWzoQCURE2/golQQhkkkSvSqonhU88dy+
my89sO1b3rSt31trek+1aRf6/GGeoVgcSdocn/Z5NItJkFx/fP4XEL7UJTRKkfP/
vmRX89QttgtNq2TFHHUWsyOew9+c59YFmXNaSRPJw3tnQeRRT2nCI+XSmOMxmUr1
PrIxMrhfxTKM9r+2HpULZV65VjeYVkGl5dr3dbw6tUxP2rGjWPi0p/LOWFsJfFx1
55xhBsVnkGFHEyVl+V52b5tyabiLjgB0l5pPjAK55wDMHIAq2WsV34RLK1Mbo6gX
CJxNGZITNd086N6fcCP2hp5GIgIYq/FgIfRxzGeVC9XwB8uAIdFeD22XA7R47H2f
Xx/8zKVPFa9xdGnwLCxmRcnICmOjgdhpCqOmD1QNKhZIN+DFwWdeMbjKjqHI8rD2
BWT7UjijT79qyPCWvsRZLpvMVijZ4h2tsB0KT/GvEp0RPsXnxEWO5jD15Jit/DkZ
dHleOMsutoHbIHvqxOAk4/6eqHQMhRBDRL0dnGkf0tGuwvY4+mujfOkEfWRmS+PD
p9vD51s5aQhm2sGVy4EVu5knbaoHIgNNNJFAWQpMmgjJQ+AGMofFLtFd2Ov9l9yS
yIFK2efDvPior0T/s9NbEZwy3OV2hASwgaKCTHM9UuFt14dRXWEUY//jzIxfHcKh
TAohVsXjJ2h8e/ucUxDmRLw3o0D4qNfzMnGj3F+voGtkRBpgCLKXXW7Z+A84uRPR
FpNdk9XzQ8obwlkIchR6QmuV45F74prBsAgEGiiAy3Suny8uBEfZVjH/XBe6tFA+
WFh8NrGDeMHXD2FkxoINZ32AvVeeBONMfLxwnnZVH7UEXveLoMPBrCQ3fRtK8sap
ATRqtwBAifezKFh8UzX+AqPAOPadS42jsryxlHyEQt7myms1BdPQoWlMpEpBwHxy
dbSaBSKv8a+eTlqzVrcV/zVHed6m88cRbIg3LpLvv4UorVA6gYMa35u0u4cSy/my
AJbkyAKu+f5XQnfNOPLJbi4VRg+mn8nw9ym9cdLjdlYNbamk1OnwfIDG6mvAlFJb
9/B/K5uP4n8MjcoQ5/34Pmm7KUmXfybeyJHtu8OLpJag/PJCkRnovlqyIQnBn1iA
c0nFAUlumgGhNhDfwRe4LAKYN7jQLQaeUBOc2NikAuGyX+7ZtytkVv/6yYt2whv6
B1RqLhLYbWzKKAGnIneDWRWZJOKn06f40Abonwh9oN2wO270RwTVLNwfef53mvP4
vknSKnqoVs8E0Z2wt89NQx+cx5lvUgihsQdRQT3YPWRpoSHVNOD893x6CuA5Mwrv
6E5NOQDFzbaCX5YrvA9enqg6E70TTZ9xzCdE4prqVYyJQLPOFBxYtRQX4Wpa6iBu
Sl7V9l4i9ddF6HuY0gsq5wyBuDHYoxvLPL5DBak3rXkFVTFJWZ1pGYsHTotT8vTE
PBKOVlKRsFIAPEMLp2XbTKaCfFHo7jNOPaFH01+Y8FYhsA2KJV2jcPWLRxz1Kj9l
yqZvwqN7I5r96dao3sEjlZvi5Z5GQmqvp+GkhkUCO1KoEme6emymypG3mV9o+S4N
wLAjr4REB2gvD8hIsqqlg8QXdwhgQyuPj+2wHDb4uynWMmZtmsgkk7xj7ATbS886
pV0cShG8+mtqiCcEIdKqlHLeB/XfNCmh+El/nAmbQ4CPYRaHSNbM4UP21s5zIYET
rwQjbENDb7MMbHKqFSNI99ceE8Wj/7kXEigyRnF2wP9+HauthR4LhS7x03lpRxYz
QbE/ZS2v6vRSBnYh3K7lQimwqnFsyMupWg9N304ZJTbrq61an7yJckFP3uI/soog
+oE6WmfpG5DOZAy+2LTjye90ufzVK3xL80US3NBTFJNubVf0vT7s1mytaqb8+KXx
kdIrWL1IS/NQakRyhMLETzLPoiFmx+N9ZPYLY8u1Sbk8cs1BFdTL46NGstlkgyyD
tR7Ds8Y4o4hrVksqH+s22Al1fa//0IVI8FlMprWdYIEhNp5S+VKGqiEMzyyQcram
L1FtvePvP7bgyTLH15N7G1efbFlC82XU/8mQrDzoin5N/ivv3InYsdxuqevuQ+RL
YIUa/TXne0Ybdc0mcXXzuNc0ZVCpGdQcLib1TCo7q6XZbnoubW8T8EwOOv0gBGqH
IS0Pbq/yYqSqpfNV238rXr8JFjL7dMJbQMZInN7tDHqA8+Le8nLtKteCfdzZWZ8t
v/1XKqcbCaHLkC0AfkLKm6avT6FJpncJDrpviSqQBUqGayGJD71EuWFs1tF1ytnP
7AJhc0e/HhY+DFjMSk3mHEXtRq6KizX0mkSz/oONBqXEJfbdmmqC8zkzpeCqK2WT
p97HdzwM5L6uxuhC38+NVIOdci29YFXKs/6oEeXGfXxlh129VTHRn6SVkue+QFhh
B++1x5KaD+h5VwclO8do40DfZtOAUkkV44Vmj2A2wxw9g16UvA6IaHtKXjn3934U
WI2Q0gZe614DKLKlCVs6SoQUS4IVD1maAhR6Vs0nb+924hr79XKOJzSgGm4Jp6G6
8CnViXWA/6OB5y9XllP03otVbnhfLrVkA/C8aQl2fYw6SIRY3u5+ABVRK6djLXkD
F3SAw7o3zdrrtNSJPrZFwhytynlnnineh0O0iIoRj7kpOTtV1pV7xrfTqCmIod9N
K9EnDb+4DrA75t8eQ8Wwv3JarAR3Dt/77ukmbTvAgm0QgIqgra4pMid3CJ1WyBk2
T3f8WpGou5NNjkV7thlQC+KK9Y7ZNGgu28usxlOrK0+WxcTqaASocs7xIwoFzg3d
8JXjy5rnR870q8T8PThUgUeY7ezON2Z17cxmBJ7yNEaUjIH6mSH91Oa/WjFI/w6x
mhXzrTNd4MCf9w3xBbBvmkxCz7Rrv9AohsK2aWgdn2lh8SyGNBIvMdyRVeong0/7
ZOKNGfCZogRSw3p+wE4cZH2uuatSh5vbaBriHTKZwTNrMwjCvk45yLYlrs7EqQTf
GqE6TdFx9EdTK6J7SBFOAUxuDwwG1vx3b1slK6x3EZh5lSvVjyOWF8cLRNHjorBC
d/46LhtRmfAIZaAbm+yNd/W0TSoDBwY+LTQhzJAxqa9+qXDcB4uKTeePqkx+xgeu
vPSUTqm4mdz/uY3YVe3LpqyzFBXdCLgEZDLgVR9h8YqaIozTJghoMJVbWgFU4U5v
zv7Py7NvOJ7eNb9X4w9PKcQE5lvkR9P7sRKpaExShb1nVm/1GYM+cslbYvOzY5L+
HzQ8/vEHjcjKgTWi+QEqELMHmudB10gMxqraL3n9zCureFqTfUqL6QmxzIH19FPo
cTsK8e7OYJQxI3GQCe3GyV1WFYO3LBRUkzo7e4EmCZNspldzxrm31jxO+PbeQnfh
LtatLtW4B0Cejx7MKz7d9UhBB0elxaBzI4l+Row8gBiRavWH92Dj3WpLHOz4K4tH
SX2QUx5P726dm4TCSspip7JUEkQpp2eathuIzp/+r16cNIj/KvpEe+wqy+piECE3
onW6Bf4/2xny/5TaSdqQ0w2lEDD6/JE27/gzWXjRuPYjiGDiE221vJ/u1Qbzi1lw
tsqGpYR7mEW5wbS8V5Tw5k8AH7RFKQnoOlZ9MP4E3dBbHjpMVcBwba8fp/jCA9Po
pLFcsep/aR/hIVqqXaUXZHhiIP3KcRVt3YAg7pRDHoZ974fg47/2mYJNrfjj0K5u
ZnPaq23En3mwU8y586LmRrhIucOnE/BNzBMndibWG5R5HmTDtTh0+dyQzk4jAj/V
z5MnlqalzZg9IlaSxAQizamNj7jXts4AIkvXkOEx86MSJKowmA1m6tvtasZOgSVk
9fb/Fl5UrQC8XxWMUOnqoc6CHcjpiiYTKXK5viomZutSqt52kQHVj+4ZtRfB+a4B
pcGMw5j55u58NsO0bnQ9BxYh36GN10B+IsWOMLpfB5fahkJmHNPsLa/FuhXLTx+s
0N0TuW05bJjMN/35SWzEDUUqquyDQp3YCEg0wSNB9jaApdL81z1CXAKVq38fF/QN
44e8ZS1pcg/tx1/dmypJ2oDA5t99WXi+pqaw+R9VargTl3/GiApFpvbvzdEJcmd4
OmORJeqECMODdQzeVcUNsZpKslQkn30WjH+U+SYmviZ+D8TzAfgBDtJNGf7PBMqA
CPOYkfQ/wpU+2vR0pXSaaZKqE/bICWP4nzIcFVXUd29J/RaD0dBAi1j99qjsOnzT
nrtg0OiWQszi1j4KosEvXgJdygkFaptuAImFzmxg5ggM2WmwyS7+Y2++oSeibfL/
sLz1wXfpnnVf6EhVCArT6me1wehPELM5Bl5D4UEn7SH1Ue46ALlq+bunwD37kiET
sZyLeOIrU9BX0F3fxh/lSvZ4t893z4QrCiYNU5xmwz+0RraT6F6iXNhzIRs0sGST
7522H9S71wBpfSVioDrxDybJCqN6wULzIL3Hpz2PB6/PrH9ajIYMicCpTLD4tI0L
xRzxTaY/GQgUEkEh9lZhTc7S+lmqgCtsP7XqUBYtgXkc9T5hTK0DT83IYbsPlHcq
t/X2ajqySpwsfEiN4RLWKEEMP31zE37bD8KBt8CiQeo8yyobakdFJsYp40bkBcHP
Gwo27p7ImSI6ihsekkY3kmn/BYpBdw3YV9KxTBpvcSbkheT8qc+iiisIBoC/PVZm
gU/cXg1FFPGEig9kvdprJ+yHpG8JE14JKePTLyFuXMJaMBK0TmOMm25WXpo3Mwgn
SZeYzQbGr2JBxx2QOBAc8WuORQfMzFEvmffBmkqTlEUJovBUeAVDv4UC7j6rODOd
yt3l1VMLFZJhobJONIUlDAL49hpsUNCcgwsKiyzYzMn0ITJtF4p8QRsScisJzM/p
NpS/V2gDNlsVGzdaAQhmMaHl7viuVAS0faVe22Pmr8n5WlPeD7XX/j2c3zbMCKDI
2HndwAN+09iPryMmixy7YxHIr1NXwNP3Hpy9jn5/yjN4w/zj8J31antDppBiwIVf
svvyOoR9+3AvdccLjXHZeE35X4osuSmGMMJO0kqzxyfNp9ad/Exj5sc/wvjmPwZX
rVbegYqHsAuxpyw9vzWSiwYJ0n1TTUr68FHBaQlz5iee4EIP1wMn36OL3USDVMQn
PhRWlP1ZE7uwmuWmV/91p2TI1hljdnYx7sf2nO9MlatI0ZC8BBgAX92jdXeruH0S
ifsdE+9LcSZFlUuraEkrVuspcKeE73uxTfu4j56U7vOQRFaDRjFhSF0TNWXZYRrJ
PM+o9nEk51CV63DNOrg8JaHFCp0rr8fa7GWn5jhUc/0hXsr49AZWB/4/zuzd6DyO
wJo8utCKTjdUtG/KXFaKGYEFIPGsIdBdTRrEB8pSiFBICFPWlVK4KsQWn+wIQMho
JSmBjkEHa/0TbG1TZeGlXQcvEKsot+nZAsM5jnXSqOLp2pANAOwusP2DWkbNdC5i
gLj/XhiEgNzVzSWB2Fjip6Q5DW7xa6q/TsPDB/42nwJNi7R5qlPEYQDBSwwnJNBH
4D5vmc9PfPb5ZenwC84wV51gjozRgdIuNTRCym/NHWQOXXJUw+7/n9bfFuuuxZdd
GqPAQXkZE68H5VElTTfoUMy48EByHGbI2ln/YveJzxjkeDxyfyTT75jB4GFjh7yL
Dx6Bp8l8HIRyeHC1iqWv5/W2YQhMsFC0HG+s6lN7pTWbDrB7h80emX7i0WvTUA8P
ShEcJNFYD0nRQPrsKkH9o0+W3YwgAsXBQ6AEBQMj2hoD48GCohShj1YVvwyzqsrf
/dCd0zNWd/FnFRuFBpWdaURQFTEYFkvF+3dUxOA3bRSOERiIdQbZTN9IK/GeieOh
x39h4d8M5nKj3Jsq6bFlAOy2G2XxfoEgAmRsh/urkEI+5NUhdJGt56d2f6xOgAmt
6LSIanZxy0vqtAbqmPtcBLZSywnZTN92XCEVGuanvI+AmA0bxVMuyCJsEs9XKnpx
+0WlOdTf49cyJNLKmfjp7gw9kahY0bGtPHE0gxX/neVsuAukhMCb++HFqKrEIJOl
E51GcTIZSkEPb/N3hMAjmbqzDY/kop1f+xhzRTEnEyeBzwz3DrSvhpsVSQiujX9Y
4LptAQDzAlYn35HG/xCDL8eXj7ciNTDRkG9garCSr9IkubgykrB1o7Cu6LolZ8T9
StWO2iRRqFBYlcr0Cp/e5VFhPkp1tcC2LPb15D96maOjlHHkaChedBMJrIieNLt+
FBqO+WVTsDxqJZv2AaxdU5EqR6FkzTYZwzPwNbADMUn4FgWGDagx4bxZUgP/+ZVV
z+RtkHqkiQD093OOqApskp4spRPZ+itVZgZG81e9NSgmkTqWo4YyI0EwgFqRplpM
e+AP0hqs/MffKDN9fwVstuDuJgOtyXDns100972dGCuW8tdLGRukxWe35t7q8XCV
38cmEFcu8weW46EcPPADxTXwTPW/U8gxNhd7gCf5Df5bgpCtmtiDSUluCiy/4Xpu
KcVcQLGrG8V9qR7PIo2qpsickQULLzs/64WGNEOcikRyzxA8vT+B7YU0lzAC93kn
dEAZgclEw7oHv04SqRsJS1qHkVWYFxnriO4fyOmlqPLgZcvc+ZKr1fMBAZvZE40O
CMQU0U5Eb9N90UXVnXt4hX58Bns/fOtdbaNUduU8jx0izEJ1qFXjpz9z3Oq5lFy6
G4oXcWF0zvGzzlE2eEoEF3lnDqivS/qmrfI+ywUKBhueeeaISa4xUfb/ooqew9av
zxAue85pL2zq50xUUnIKXIaoJHYwlgsH7eswVtQRqQb8Y133LsAk+hkGXuMVGLL+
STcwtCMRp5lgrtGDmX4RrLCtGdMEXlY+qoFNhg3UM0LKabU8EJ8VGx0EIqT/6aT7
JK+0t0gVhdhM0tg5VgY1D9ub5Of/4PxPdNI71yfI11d+l3htuekzgbuVXqexzxMD
EIGloCAnInvo3OHXPsZsLQDcPgH+UetsUQFuSFTirirCgdCxeIqVDBMOv2L6X5JN
D86/7p2GJvlCLdsBb2sPct9PalUZvkSRh2hCiwSkpOnLR2SjkPK9lqgjGeIipN5K
8LE6ouWcww54innerU6Z1RzOQQ5K/udorPYXBcAdcbrWtxbXAfHzN9AoJ8/aLxEV
JbHhzXMM7C2Hxys/2IQsqheRRsUyNceyqpJRSVObKr34P9Ve0VUa3NenTIHSG9l/
Ti55TmNh7fFseiN3L7U1cVAm89sL9uspCKDTN09EmwiXxE4PVVhuNqr+5lho6k1I
h4iD3cAGDUjE9Adpq1aGx+VvewDRKPtVpgcjIUn5ZmkhWJKn83RZuaokTSWj/gDd
xLHr5PDyEJwgmUBC94DVgbKlDyofX9sriyVGbHDZhlIN3H2FgTaeBESUw+UFxhcI
f/OnGmsnRdD6pbcKBCW4Qm9ymjQ7ed6jgaCMXRQJpA0vFpTvULUM+NqNUt+XH9nT
oIH/+JF3/id4kVpMqSKqPc755g5qEhV4YTwKk5ZyBq0KP38iGcIe5x5dradv+8PV
FO0Ref/2JK3NJ2mYAgB381jFly+kqBLlbM6pBYVBcGYH+1dsbE+DnrBlcF/PJ0wv
+pCdtB8UEHt4fkah0hN2BdJkh47av/qSuwe1ZWFwLw/XWDQymKUmeZOetHc1AVnr
MZVPqImaTb7e5T7qA9czazw16RujRDS0A2TGCLtK9rXFOkt0R4PMmAuIq+rdaEA1
f+fG3SWV8pzHJvhB7FYSwnT7cI6l6OMyEpn+KXgtRzwKpbFCnnfsO3p/Lq+Nz+NV
Uqg2P/I4hsGkC1SEpM3RlD8QzkdiTHJqqOOT4QHcrM2TKFb2E2eY/XjeoiIazHDV
jf4hcSSXuKblA/Irsc1m60/Tml/hCd4UhH5bcSB5/DPZBX5jObGVKe/69KCKn8sA
HlOrlscdEotzavfyVwgs6JudnJPALDOf6kESA/ZLVKJTIK7Q1kiLF2Y9bdy0JcmC
UZwTlncfdoCGAPXPzajdTobQ7E3zMDfxdv2oGVOpHHWqFlBsWPwdIvu2oVzQIEkE
/648YuX2F4BppV1HAhoG4SCMN/HUxRFgOWfJTd/09YRC1YP4P2ngQXdaNLBzoM+0
kEtH2cqNvO5olAjYT+58tnZwpyTG2T/ZeAhlg3iSTdM2DEb/nQjjwvTYnVdtG9Uj
uQEa6u/Ut89b6Kxt1IOWOPaO6eDhiIAGBe8tI9wDlhtGr9KWFTMHwa08l/0BMT4W
i7Q3x7cUpkwN8Ps3EBH5Qr1O7KyxxgVfxEM+X9veprRrMXeeNM843DzcQyV2O21+
+IqS2pAmQ9flski5abVwpR9OBu1lX5Agz1eYCJ1vvvNqacjl+qYraUqEqGu1mzz2
ZKIxZ9NevQx7ZTkqAycE9iQQQWP6uZkwcvjfK/bDd/g0bE6g8gqliGLbPJJO3J+F
Towl0z/B2QanmwBbZb+6j3gF3K6N5Id+i7P1KppBDFo8YXk5CcR8xZW8uX4fHPBO
YgnWAGLDljC5+C2cSW1RUHGwmsqlRmp/5yZSIDfQlMKf65KFtVE3oNbBV+rQSPFB
I1ePgEoDD6BcxF/MPz2oslZNIf1foKsH9oY+qeIN7+dqjodQDmLHp4lNWqBRFzlD
TlCYLCDM2LduMBf8u9JJG7qfCtjqT004WKLuQ5ArkzKWQzI0gsasnK5nDt0DzyZW
u7QNqfKHw3qF4sx1PNKI1a0SIOXW9gzp4h3zOIksgxgcEMYqHlaH7ym6sYkQKpxw
kHtQ+FgsdxXYAau63FH1IpfCo3og4ypJSWS9QZJZxLCjZ9joB08c5zN5B35cT3zW
MGZtduuXjTbeuUsLwdS30RC7NUICbqvBwNb3w4Rvzf984wp771cQU2+iodiFgoRK
ZCwfeIQpNX0/t4OjX+5dmXcAlDVuOsXOP1f01xgiYjwppz85UnvV6cE0WKct/N3y
GLHZUJ4buPEHDEE7bOQEYvSsuRtvAfe4sT1qTE+WwoFryOl7Pe1hpmbqvchC73r/
jof4k9dFT22uOFVnQFizG3Cj9l264iluyDjmaZszXldT4f6pXsT+Ja6QFlBqE6Et
HVhEqB1BnKI/baG+Rw6FBGQu7glOAEB3lAtJd3+Ff28FjmmVj2giCq8eB+b0XnNX
G7eycNLRngkv1HDzyl9yaY5HFQ8CqkNa73Lj3gMdUEoIeezpXNqeUC9wlJqV0dfT
bsvlLU316LFJBPGuoUvDFth9ydI6+vdHr3bWWxVGp0hT+/fqq9jKz7kRCNELUVjl
6xOTNhkWMWrcZruXQ2CZNymXxL8p4aIqA+i0XQt8ojOWXnn5BfoLIhxMYv2INcgQ
ThkwcoJIQdCasTnLJ0hWwPx0dgWGZaPHRlX+Q+Bnfv9t00TAG6KdW3u+grupKtp8
1fB8zoPujdoYyYlahLI06565jRHLdpscUbebwLIK3VBEoZ7YzfR5Y/T1FUfF3YCY
LfiAwBCvZhK/s2Z26AAjunEDodOt4HJW+pW4XLklwECxbNLdeohTvu7ydXp06ylh
K7gN73v9J4WZCEw2nSef4yxb4YOXfjPhrdm2eDeh1hefUsw6fznrl7lir9VwN35N
WwFiN97DxgzsRGJu9SlqPUdFsol9Wk4Uxcf2KIQlSA7L/FEj2jS+Sf3Ma6a/+tro
qJEZUaK8ZaxYC14PF51wYufvL17fbUAMPYR1DRk8C+pDekWs1TU8e7nULGpsYmJY
ib9GDdaJ8+PqhnuxgC7UV0v9WykqpW1uqFcklfxeuSCS7lllGyFKrRMx/ub6xmVT
oTIyf2U6fB727S1hF22ok7qJ6q+6uwe4y52sbNbojgt6zAK8s2bcTMcOuIAlQvV9
3crEOrVLyzWtIMrp66oP/ylN8SOgaqLiu1rmFf2ILXdSkuk/Jj2hqv3kgmh/gLxc
ARTEAJcnDPJIXfN9eagbVjCnZq1QHEyI0ip6ZjpNvMtQTL1Gv18wc8A8+t1y2sqo
U+vfLaiCs7HxSE9XopN3I+5ezXNnf4v11U8ad8cfSWj4y7deL8iz0PpOpeotk6Cy
5DRIAOkCjkD68MRI8mUjQArtqigrOPL2WNqsUe4bihW9B+6NcKS/R6aoEXkqgD9d
pYSlIT4Jf/iKVfUQjT0K2emIJlNUsHK8SAt3h+Ccu8DW2PFs2Sh2HMtosNQ+pbeC
qLYAvYlPqIOTCtoexrajQ4HZ+2iK7d4BmNiClWtFq5wEzGvgPJHhP69HyFtYQFhB
0X0wfeXQ4vpfD21MhE0BXS+8oYSwaECJ1DFWU02t7KadAB/ghfiS5WeVTblXUbiE
VWKCVtHngpdi8R4sWPoTcdJSL7aQkCpjNlEndZlvcVa0agsKiuyEBAW3zqK62dkS
Yi1ua9/ZKPA58Sp776w0jeF6nt5nPc/r2iguiNWe8ovNMU/th5+gMUKONrqmCEYl
FtJiog+GGzwVMnoDKkaycpX91d/RLHnwzOHXwEUj+NKQ9ck0WBFLiJ+URH1bHtDm
rk+KzTiu8It5AI73iC3IvtE0z1VS4foS83xQ4d/8BR1bX66qxdOagqG9kcBbGR+p
oFL7wc/LWzyZVLG3f2xtrBX0NcqIoMKn5KEuokMU8i0yrTF6Gjspz7D9KVDsGpx4
1Yo7WouPD4gee6/luYqPhDG7oTqRavjguusUPltwQeqSaGsFvybqibz0WhTCoHg+
VQUBqglrpIB8EptRIpkjgPutaYHOQ2zodB16k/3v1xIH4aCrWRn7cPNyCQwJEQEH
s6Yghzajtd7UyZAQVgAmuiJJdYW7eBWm0agUo4eqcDY6JKnMDiFCnMMBiacD0eqB
BK8kRHIlkSurG3AiQlYP5J0ExnqIRDrSQkR8f7r5nUbIOtTo4FJj0dtqr4OHRkNs
CIDwTMpKrmz6zdHn/0hOMzkWWijqNoJw8Dvv5kncB32Eup1Eo3yTr+R7rQetjS2k
X6rWdN5NifunDMMeIIbkempWqGJtAorNqg8ubBqCI1MxPpLeJ8jOOPfp5mcQmWnI
AQ8aNZZY5afhu45KHUJFZatM4ZOEJUwBRvKKJPjTpQ2xh92Aot/svmx4s9Yj4xeC
cabfw23N/JEF1egRumtvDXmQyRSSAej1Djrt4cz89tbZOlklbia04OZCExy/qVex
w0Wl6FurXjopyWFzM6ntuR6bUu2QMbSslQ6gKfcn/I++P1rlhPriKCBppgNLpYjW
VhMaQdygq2TPy6DA66iH1WdWsgGA4NT7dX21YZcl5UzUYCekgL/qj9J50RUNz1rj
i5S2dSW4nh0F1R9lZh6wSwFadsY4xvk4xovOsFxXPN66UVxrxeSYvxES7iCszyD7
HpC6Jk3bjoVfV/BFCFo1yhsEZQEqNSIHoW0olt0rf/1OMjkyJOAYt7w4YglupKww
N5JsQVTEJYqW5rK/oSMq/kYmZwKF94c+CxNmB11rUB0YrbKXYY0lkRJFlbsqNUVH
D+TKJXySKqGujnyscGrR9DI0R6dG0acTuzccZHrF0n9yPI9UsiRJyzPCSsQYMtUd
HAxYGMGfEpP7Ekmn2AQ1cab2IffpsbqfoHwFvjQ0jyo8uZzNMrJosHR9EC8x7PyO
HBxbJKjLxvbAZOtU1RkNyMRRH41amRezrvV9WtFgw9uuUTDXI74C6kzHEXJ8msyQ
96jYAnpulk6S8wV/HAudJkzPODwR3Fr4yV2rZz+BLIuUpbIQinbXGjo0hEoxwdhE
tAqZezOzY0PWuFJMyv5Yqt/PtbS5I8PVX42cvZZ8YPOsfNw1uRc3DWRpeh/r77Mh
xPEiKV37+DCtmUEkUySH4XW9Gf0jC2n94etcPp05/tpjxN66bIts2nrROc4doPia
c6hjCaflrsIx4yl+LAKEXN8OGjbUsdoLoptf1jQLvsttfEq+L7JJ+6PLXieL3Rao
1874MExfFJaS1Jih0O+0bVyubjaFnAs+o69pbZl0ny02ITi0arHWkLpdFxEQVaX1
kSq2DdcKu1KhNyNSsatN7rLV+qLloeJ+/cNQYE6VIOH9kwxRQLKNWo4rXCi4B7YN
V7267Rn1paQe2JeeHhqMCf5plhEmkXgd8WPt8tufrbIVHvR8pOkcIFdEmeI0wG6W
sLYCo6v0ngecV8N8tPnBWYSpce2RElCxVemOhLIBGeS1dICTze09ncoFPfdfOGw5
1eTcrqQupJjN9u9lZXDfk20yMtV9zeVFY2DROoICU2Wd5g4tNwcMcF7uB//fQlRW
bVk291FJYWBIxwWQUfyLCwJf0jgH2hiIICrfWU3N3htJhtVRrAbKuto02/6N1jjH
T1oKBK20GLpQ4OaEFVsq76+HWyz1tyZ3zCePlnqVoeblin/M6kKFsMy0eSaByRHT
ix41heEf3/3gp526xTADXBvx/liwlZZ2Vt40bM+EDgt1Nmeu0pegQZ7RwWbLHsg6
5DKMv0+8dwdClooTHRca17w3FPDijvekojp14BAeDjJIlApQQSEm5PvyTXfnVAOw
okJ38o+sD5mAaI/CyOTobjLVFd8A7sLve8lfwXUsFf2ZHE4dy5gHp06ZQlP+BOBZ
hreJR/graWrlTO8AgLiZo28rL3sraS6iQp60WSOFlH12SHE1vpwF1siBSEjfOdy7
bzJYSaKw7QCFJH0Dc+XuK0WTKELy3iVw8qPtfquISki1/tZ3xcUvmB+KrDCq1nuZ
XapZDy+VOSWQ09XH/OBV+vSYTiVqqezpDNp4r/Tdx4Zmp5cGQck5GKmdRaNt44/w
O+eRcv6ZffTrSaQXl0nQRFg6GQgMYQg4XPBalhORdFojAmJ9RsirG/Xphhemy9nE
hYqp3/kufXFLZ887R8dco8Erbi8iOfaEWIYiM8JdUjNiYsn5jiOsrLDq+RKaMqrC
Hcd2Wk8CNzyBp6p6zJnlUzpI03pEzm5eeR9sp7tl/1IOUrq+/QV0UYlPY10v0dw7
mvB73l3nqzgc0jhSGDxU+tuGa/ap317ESaehSv/RmwX0+nEZuC/QOzvAmiXcEHTr
zIbeG0ZFTpqiTNOOtB48KnOgMB0xzOnTkaIbBwP8C/fcK+lzFrxmY0hWedqHPzZJ
CNhBE9/Qyg1oWvaAG90Er8kWqD9lmO/o1sa93TyF8CFBqv6dj5LByd3TIKMcSD+w
/tAe/Lb7wIQ9gk39YrR4iSTCUk7C0Ehj80IO63LIeLYM/GMfji6WWAfa8Jfb9yZl
4qDZD048oAIVZ+gJfgnv9o2bVpng7Vde2IVajdGRZY2yO3wZ9GuvfOIpH3puM55Y
Eamo/w1eKgiqcipTIKJFLbc2r8vq8zDGaY7ezzLuF6I3B6JMAiFhqMY6HCyDfa60
CWdslLZZfOKWQ37Zso0bbaQ7x5qUNqkxjCoRgipas3rbJobXXR6Pu9c8uMwFjIGj
3SmyjnaHipapFVKSRlybqmDrdChpQZMcpLvaNunsd6A2F9AcGJXeSCsAsUzLDHsB
Lldi7Lz4W8NotRli0eNvaGeDlh/TA7t70aS/+7FpjWYWa4VL7KuNUsadgS6lYYd/
7xnz5HM0Fr1+j9m/fPZmz890bPS3tG+Nrhu8ypFmpdJWa4VAlg+PnHBQO1vrsH3k
tgSYZm1NPDDxl5t/FgaxJ9g3P8BDedMFLL6sV7n465dTAzBoC1eOaD16MfoZJkmQ
ogc1Besz3o/wQunurONinZJ5QkWFHoxoC0B2goyyKBxXmAEnivqmppYG8chRLGeP
gaLipNSejOdZ6qdUAQmh6I4HEDukL0EeIgCgHjq3wGrMRRQQp+0iG9MRZRQy0CAh
Ruq5ZwLpI6Dlt4jmv7GaA7e25y4AS/iIO2ybTc55D5OJ0/QvS5Cl72HsqtuqM4mq
6e6cWXOx2vSrlPvSfEg1y5FGSLj1C2ilBJ+YCN8PgHz5r48IbNieDcxfHbqVqDzG
9PWE0EH9fSYDeai2ErLhhN92+RthdcxEnyb5FS5ImzP57ijZy8yrK7Krg6MzvtFx
DLoGj48Q5VdTslQpboVC/EdCWkX90+gUzCGKlFPPIzwA8A3616jX4jpIPkeA/rIX
y5eRcR42u9qCXW95bZNCA3M6Iad2IkghzU+sMgAXxNSsqxb03kC9tUNtjG3MO256
/vxWxeHdx3itfAap/IEehr6NtXt3zJpKgLUvkqensQqldFBMuoJHq1wc4BtBKsWh
Hlvaebe7epB1QsxDrGFB4EeXOUwy+iY04fLfviPwIlrbHSey6KvwYNSoMEk8UEXm
C0tm/tStzyNJxVcqXV5Sk0UW2511cTaMqCwr83reZgu1o85f2+AoKGyW9ef9HuBP
YFgKp0Cm/ruCmIzVQ8gZGrEYFQkm6XByOqs2efYgyOqrjP84uJn4vb10RCthfQXm
1dzQ3qZtX2XoVJJEGY9Urst3ri8Oei3e4xfsgiKC/hm0iMKkZBhSqoCna+a71UdX
uhUwj4MXh/pcCfdlZqg+HeibbDKE0wwBhwuytW22/4CHmGq/rT99GM0NXOgo7LDp
A7LFIWdxcaO5OHwjxW40DmRgVS8Gl1RktZZZEQz6SDGzt4+26BqQoUVTSHO8Lp81
hHokemLL+P0x+DO6KD2cmKuf379JMr3C9TfYRisws4ZSj+pIdJZH0oheuh1u5o1c
A3OoPEvxmNKYMUgO11zkxJgfT2dKFRmpjb648v1V0wAEEPfstO9Kn6Yw3ntT7MTS
AgDD2df5Y3ddf23JBMTB0PWssp+gtHoEGp+oiA5rMrpkwHekOPYa78LMD3q17EEy
oW8BDlnEgZEoS4Z74e3Vn5sfsEnMz1YMlYLxhtNBZrG1GpBbeH1e05/cFcQvDaIR
ZmtbPl3dkxcIcz1+dtx7jumqCALGTvGJoGPbwSVhQGFSzuL9Y9ERNgNNAUpgqlha
SpT9zHwatVI2cLmMDqqWY4e8LuVCVdfULWHCxHN4PkIZEz8QGGSPSPvp87uJfU3f
oKJJKzVfU/F+4+gumOgcQimZxGh9xhF0NfI+hre086DCxrRYJEtlAtB0HJwdJrKX
JYtYPvpCSQFSfc477e/w+3/tQWoqRByASFzM4I7L9s593lzS5ahzQ7SO5PHYbRLc
hWTWL9b2bgQ441XTqg4sRzQZi6mhXZnXWDXDVKS0MF2JaLRDW5TAzFi3j26TfuxR
nElZUr8B9tpyckHM+UqN5ee33qJYiRIWUS3Wae3fmndpvIELFlizDmUxmcFVQiiD
zbfHy9/S9mF0HlSqZMP2KZFV8t+2YDPjoN5y3bNDepHxB0DDMv79jRNtGHXU9NxS
is+qiQafxt9mBH9cEENWHPC9ThnKm3X+yE9IVthuDZ0rdLqhCAPjY11DSTRybfEN
eGvoEIy6dPaUfEWeLZ260e+2WH0JzXh0JdFFKJaI/fj7vM4t5xUYyHYnHtexORVk
fT2R1Ah6Xqf21ezk1ZH41c8oPeI6dfXvO9zl1GWGyw+6udoHzftmVAHhOM8d17FI
bKb0DwbdTrBGnY0vfcT44zqQCXoVzY0JX5M7YdiTWdjFx5BEWzCcF4BHqhwrxxN+
Iieqs0cXefoMGsSb4xa3SvE5Kq1KESJZpf3mRt7C6YWcm91TF1JgmoK5v00m++RM
19qWnp/exzhgLPnonCtX8rtZOAUdKv6n0k1OkHvQGeptBqi0JGYLVB/tB6yeLehW
1K31Z4oVb1/bT7Ez8UuA4HoNKo8EfPKZCP3n4v7puYBYLYsf3lCN+k+ZsMYsMnR1
COfBtL0gvpigF9XFUZie1Aijb3zE+L1h+DgIOqMEmUvaXQfiitwnaWm02StqcRYG
lP/kj9FeNgrr20DEnRzgcoyw+ygTPTVD0vtKWww74V/pokwxArDjPYKcOR5AaVcV
d21uC+rcrXtbSd5xsGnW5AQ9XpDj6y2IypljA2DJLIckMQmH+DjmnTkvIkZCh+7/
uvQeIJl43C4dndolh0sT/nu1nwBtV4yGy8ibqpMLdAHNp2mQREpaKKLQJCwXud7f
otA5SZwnO7LHpUWEk0UkHNLQQuHhLIsMVcL7oK83dRpxLTy6CMHDW26/yLONt5uH
T9jD+54he7STFLaAD35jzwGFC9jH0yhFj7m3jasDo7iLRd7dQuY2blYMlHk9XxiW
szDl+0xfiM3nqp9Y/7G4IxH5YQRDFy00N6i17LvTGxJD6goDUfSt8Z/Bzrg4PltA
PT4avowToF4XGx9iRaS5f8FPuETSaNW1I8o8hQM63qloS+ts3aXol+NZb1dM2JN5
jbfYRIEnhPae44ciIcGB7zOlOsn0W0nml+G//1BaG47zftaxXFEw0tGZgBIrKafE
5/gkAZaMiCdQjOOdbmuwUcgYoCHjDEm/ujNGle/Csyk4hRbUelmjr/RoyUdF/n8B
N5UYJB7ubkwpUj05ek7gLagV2Y2Xn0kBUqESGFxILJDtRKBAh3OFXPJsJnD5YUPZ
LOIISfLKlGEWyl2LGuZRJviMmsbmCI7y/eGomxw+g2ruBkqMllT/si97RJaPgN/Z
X3K/fN8aermiE1YkXIojbaeV4zA6+YP6kJh2KC76oxYZ+2PNEgDpmlUPjji34FVJ
OQ3s4KvkOzqByGowqTgQZeOdDoYHh2x/gSwvXwJDLiIOuXUMq/kdRYImVqUmwsZa
giXb7+dnyR1jgD8bap0df2yGPiDwv1QP2eksT2xsPvCE1beA17dtECM4PWcqS7M9
yN+foSTRMe6gyZALTWlDyNSSeAZev4bYxaVs9Tg9XXoX5DQvwuf0gy8zBHNygb8y
9dcVG8QfPn4lJfYZQBn/yGNV/NebMyMRuUKzfbApchUtsR9IE//IbwhaTJO/cXuk
GvFiyd0d+1pOJtUGPFQs6ax0Jai+n/bP6a2e5A01qxCB9fCDkvubakUmk3ddnRyh
8xV6TqMKvL5gkO6MAJ6Z7pPm9kW2JhCj8QTkdt3v2TBG5/KCMCyF1CwaKuGXL/8c
0VwaTTS2pe8tErM2pTqJj0U9f2sAhLwKTuogusN6VAhemqtIhCA9ZvLwArixLjAo
PmEWO6cfft6ZjHWgy/PhE1oYjQ6Fd9HRYUlS/gkscDLx0tNheZNpStfuFS6jpO80
8unAxQLbRDADe8nW3KcOMxkWTrqjTUejiTmgRC5EkCK2wFdaws1Fwbh8dDXgzxKq
RjMMU3eK8rDs/U4HlZ8ekObxBxFj+33oiO3t126allzQdaahdZhEXt35snm8nwqY
OWXfts+T+Rz1OtNoIqxJzKI/o0nYGhVDR3Bxpa3cF6aVLyYVE5LUzdKchxviMg4r
Jt9mjcaeuJq280O1tjUwBsNeeupcOrVcDcSKQDHUAhDj069BWkvaet1kukkZNlBq
WkHF9LIIVhtaDPddTo43U06CauhLjynRPISwnN0rrVjWPamritPFOEp8rMKlZckR
8dVxT/I1HRYYyk4i2NnhLCVWW6npAeuww1fqUvdtPMIKFvQN9n62cxvY8AlfxdR5
sAOXtq0WJd3e7pwFUdpkQmBoY8KNhlt9RY+/pqNCFIO3n5C1Yyh0aNgctlCGKOFj
7LvC+meQKB8e8M+20f92lpqL927s4FZXfwFE3+OJAvRXLYQG5ds0M4R2HEKlADXy
+3CMkYFBTTVIZKMtRxbRmu5PHpqAAeR4UvgK+x1q1yeIm+dlA26S78ldpb8A4co1
Huz11yun9/7v2bYDL7/Ay9/pYlH2j8NjmbPNRRE94O5XykZrVoRIONLzsuat9yJ3
pIc2w2brLtxUOuoeByYsmynDYDnk/m8Hnqo0L4IQTYU9QkgdemW9VzpFDaMaF21A
W/Tu+VMbyJ76v/GEmfHossN2c1iFaT8ItixiGCtLjYWsId+JY3DBbxJVTPItlSu5
0EhHF1qRIaYwrlvQZg1f64KxV6HZdDYhaPKyLbLziQEhZAqc28LsAva00g2bY2VK
SoJH7T1zarKD+sAkJbtvx4OC60y1fmjFYrC0K+KAdOPSn87d3H9qFsdg+VDA3bxq
UNib7X0bzrjkpDFDpJ7FvF1WoyyoAusvyePg60hES8OiXnC3fCy2Zvg+toosTC7n
zojwMN1TOR5Ft5YVTE16osCsLgJQ+54Uc0LaMQwjYLQ1ewLwZYlBcwz+bGEARsuU
U2WTMEnlB3aYPkXSaQaVzKYFJEXmY0CXsxMxsKas7RFtOO5/uKSB4qwywqOq9VQg
c6y8qjQVPWY9X/uG5LqtYQjGFnj8D7oKkyJox4H5k4pm+uqfrBwfQ/Z1MNaXAX7G
oSfOdiiEC7Dl8/lviVatIF2AaCwxE79Bbuqym7zgQ17oyjzx1Gl7Hfgx2ei5OU7V
7ndCMljOIU8X6IPbPPbQJrY0Q/mgBr9FOJYldxAXkxYTF0L7bt/eDGsm2/FRzN7a
Wble9riQgAfKEIXloTN+j/ytSzJBAwXjt3ORLiokJZ5zQ2Kl9MGDOsY1A/+avdoE
Hstu6Zx8Ox8CXEKKc6eofmbyc4+eohryoB5l01Y/2cvK/canH41kucCZ67KR+TTR
ELz/2XyupiMU5V0Dw3AHQSYoPgGsDLcHmQpXzUFbPZPwrtIfTZ9oF7xfpQFZhPS2
drnhmaHSmdiG1g5O4uWe/8xxTKe9SEMWJBnpT6SEnyEU2hPoOGsLfygTIEKdvd/Y
w+dqhXPB0iJBviGiu/tOtF+l1hUz9EX1G+XiWXJeef60sJSAZWZpE3St54Pv2FVs
x9xdL715CCBHxlJS7QR4tpUlBZ1+SDco8wvbiiiisEdQabUmzw48BjYwEisMMRY9
wxWlxSBDcbsYBPsXiE4DPV1mM+dncmZ0xnrs+py8BjM2nZ8wRDzv5vOdX8nGoUle
4hLxtlWBenIs+bI/PPql89wHsFQ+S3nGku2fwBQJyIZf/NA5joUJnwW4OG1TBXIv
TAASAld3X78ZlY2CfJQPjzz6aPaO+FnNcKnzyPQ92T8j3YeMGbOVmsVP1cQu9F22
/lJ8bIdd8V0ONgbNL4ISC4kQnrWlu6tjjsvVAG1T10U8YZbhPk0kDdH+Pg4YRHZ8
3Udxbw3kgc1CaRA8Yw5mZTvWfT5WNc563R5tKNc3J6nvsMaNF6Gr9KPpmDWF5qJj
I7qD7yLxxidv80zoskfSVwwETADC2F2fL/cUIFpWIYaXQy16JFOyf2WyGtuDQf5W
eJluKAW9qFv2AGcf+sA1Q++6O+vhhbYRXVPs9U+b4xAFHpQBZ7qpIVsrP9imSany
2pYa3syIXuLVuLUBXoHvXXngVdHObVDwV0ZexU9qpFP0NROqbBPThGjGFdiGQGIg
dmeNkRvO/jJe3o5mGQ4WQIpSlmpdiaTrzBw6zPUnaWgS5LLNatsVojVSbfsT6x70
d2UdNEXxWjepoZq+NDgamrXIo4IqEaCROKo9yt4Pg6d4yMrSNXt4r7I5aW4mnG/Z
EWWqHnhJKxzsdZ3i4eHImBVAyUW0I8syPlzF+O/a2DwEV7fmFnaOFMYomYlbzjNS
SWlOoj2ypeFa+g5vcz2V03ucMa/uxTVxHtOnjslD5JN+WEgqvSkYwgnj5mc7itf+
Z4n19IQqRUNnBedAEUS9oxknP9g6ZgGS1FpGZhgBpwVUbaD1XsDc/Hb2FX+bRfF6
Rxf1E61Uj825FZ4LoLlosZcSdurmT1qnqvxSy4GJp1gy1gBu4Li/g/SRr3DgRx5P
+JcnWx1yxTjH6veIoroq7QGHUL0B6ilAL+WLCQxHu183ZZ5GgdJefx7uUlkKWttu
s3qcxhMY6yhbiGS8qgycGgMXeylPp+wI72tr1qkWPb92avYAg/TwGvEAEUswdM/m
QxjNksKp02Q6cEBqHffc2PKeFyst6mDNJePDGy/qNXebKDasRf9alzDUrjfxf+IB
OHVB5dDAb+peKQ840WaBPYKHQw+n0Vy3BlZRsQs4D2nd5/gOCYoW5HLFoLa/PcQb
9V5CkR+9ovjx7a9eGioClBmV6VYklhvzvFSw8tzjDxTYB5VEUgxIThAqjvhlO4u0
au8JNmZpgKGwDXExQwqduMJI77XIyHQewGNBk4DKz72hVpS5DfL8f/yzbpfxAglM
UHjPH+KJVXKjy6Vk6mFY0ND/g3QKMCZz/kgZbZ4QI3rjS4/dDRzULtWqRRJDfFV9
KHoDHTllW9AIrKLwgS7n9+xoxL1aSSFcyjhY1pRkbO7Cmcmr/pDELc8k7wLCpCG2
e8PyP+blZivFJqWMnYf5o5Fv+avETRLCo3vKJyHvbs7Y1P2i3PhyOW+ZCxvH+Z2o
iGSxgdha03b7lCLwuEEnBR6PyeeL5HKsacJ0Sn9ZQZcQOCJw8y8biyZS2tGc5SMB
WjeIV1C5gUQdOeiLG67hj+ERUmEYGj8gsjoIuewMak1BfdL+Mj2y4zPOntY0zq30
Iy13gZxztfquu8iH+xuR4kbhyvoC4SG1E8ZZTeUAdzv2IjdJ9SKSCs2VukJGLRfo
iZSG+FofM9dREgKDKpLJe2pPMKeQDi2CAE0XRWbZkgVvqWDTN2hlr6EAQlnyrg6F
HX8B10mgJ3QWYCnUYYqLyNEI3b1cOuusmHjwZacN5KAqE1ALgrhAujQtLtyJ+1QJ
myLfeXf5OFV58V9UnmLrE8lDLekcAB5oz3hN/Dmtnysq/Zvy2HGXu94QzeoEJu1u
p4UC1NTK0Om1Q0byWKISrW9VNtwOGC63hCtNFEFo5JzQw1ZuZkLuoK1ufWCRzlKZ
injGdRWhwgs92xUl4T5DNfCjgE7A1DXe2vrvafz5oCFkQEcvIKYX+xkRLUO+KEvq
ZZzDC5YKHLD+x6FXNqVkg9n0k7ykOewEYBz1a3m8EUbA3VfySLw0IEz790yRm+2B
P2mmOe3l1RneuL1coRUw5QaLe88sC4FInAZr8FIlHjmwxe0CT5XEU/Gpwj/nNrms
BzbFsRdk7/wHZfI7TK6m8Gh8rusblbYOzLmAnMd/C/HzWpOUHKkjExzTs2A2nWrJ
XjQYrSuP99l8Izl6Vtk3GeDjAKrUyzWdDb2tzIgNHPfOGuZ7vvuR3KsGUClx1kBy
zRAuCAyCwFNNVbdwcrMHeCfSluWDaINst3zoJB4W3BdSKoaZwrQt8HrjUjpfrIFa
2SrQHRpi5p3q4jJcVPboCeMag0Y+UkrGgdWEUtqulcADn/WLVPNnMe1RP54YQ5La
5l9vyG7o+DYa7AO7QrE5jKQv3qViB7x9VxhlPfegHMU6LEplTS3bja3KEX8CuuKg
GgjMQBhMAHLAuYNoEWf60ocVuKArpHlY6e5E8mr9vM8QaY47Q+XTtpVciykvQsWN
KitxshRIebTe5raz5LsuPKHfKqgwQK8N23JA5fnaQDbOrEC6uogAHno/WB3+9cjQ
1bz/a0XIJfEoSINg1L3cEVvvPibpKNdkFpTW4n+jVHRAbK0vCOT+7yb27vjVz25x
nm63tjp+efjrqrBpbVVQdXojiunVpfhFJO/DcEQ+BZGg1R0/8dyKDt7EU2z8qgfy
+cSVuCn1DQXfCE992ydXSQKZnDFpYOO8yxFHyq2m4s0IfLo5+Ar5+vgnM3hEeo95
s9ejroWiVh1nu4dqwhDy/cFk6IUnkbqxPbdlUMd0a2CDnNHIAVnCRpjvI3Gh9tlx
UhvIlW1W3B8AXGO6hVbNZXNgzvVeNt3tg8OzEAuxNIgkJL23v77vpQhpRcAJlvht
tiZcyTkybZG9NPCDG/1GS1zR/hRb9mea2z/4gVuOTPFttAHdVEEMEnexqMpSsv6F
3JhgmqtigCdRz7v34YXajNLjErknqGtnpeVLqY0pdLfQ+vlwk0Xqke3CAdTNlnz2
WVNTRICtTPHwZr3cQ9X0da6fWAi6Eua/VbcGGu98zpai4DR33WrmPqYpcw7Q4bH3
nW4/F8BDKATMnI9jEURLr2cYCqKDNutVQemsJFbFafcYVMU7RQ8NB0+hIR8bmwRi
T1v4PqRb0+oyTAK6uFz6VCiFbRhnMqsyisA8W/BuJoPxwTDl+0mpp/PyuahvmAz7
1KC43IUQQPIpL1cxYb+0Fc4V51yXV+JQnZ3QhNdPKipWec5O7Omrn9a6OV3IxmUC
vZSxSQnkSR6YpBDVnmVJXh8pm2vNHd/UWp9AfmrF5AvOqUapzQrWqVKgAALA7DEO
juDTT1L5aRlbZS1DWrwEFc0m5LlMvxu8evY4ntEwkfpKArOxijqdb/Yd/DWdrvkz
HlxRROK+dBcpecTWB0oewGjFNgwtRiT6Jps1KMF4FcsHP/79lWCy5IkCwre/bqwZ
DRxVyqJf3PSUKu8UNLW0bn0P8F/sCpMWwCSEXlwECsYdFPnPb6vq8UXZmbHnAud6
Q/wXSvu6/fPGv7D0jWMUpV73ynct8inrBCFsASnNPH9ALXMbwggLJ3ARqhBPwTk8
FMc3mieT5lnETz/byaifXzg4rYR9MLTs0iQlH2QS7jHEvkfJvBjpaEvqZ2IjgC+U
OIhAfL3UFOOAJRDBYoDi3o+5aYzrWSeM++S6RN5uFAlcWis8zsXZCb0MJwkvI7fS
UFryGUtqk9b1g81IBDI6s7ivIyg38kQmj5PqZ3V01/NzjXt6E/WvgjAHUyR4q/9k
M3cTn2R4DF0leMNunNw2d5wrgwrdYFFHrZyvoovdZcDRgkXThR0fUXW3L0gIwZe1
h11J5+RoL4rJINPv7BJ/F4CeZQuF/cQQOCSmjbNjk6p1uQz08g88JGKVvOQvCW9n
PTvtrnhe9ga7/vHGMpWxERha19KcEg+TJWI9PqIzWeaE9p0T4/fkjTxtvEiNGRJ2
CelDx2ykfaxx2VceHj9yOuCKJqG0dykvu20GAn+QxtHwiDh6kQ7nAswrIAQZPAfp
2AT36ks/CjNgAZzobBMxX4lRH1lwLWYYSH3fKFLrOq/FheBDN5quYto1OCHTAoYa
K/YFVUWsOV9OUfFukIS/9P7hvO0S6eUa5WjvFPF11D7axVRoEvcQfVQpXiyeAy2p
NzpdbTocHj9RLM5/lFt4tR2slPL/nG/N0n+3VFzfLFLzVROPuU9tAJo+XwWacuDd
biAjf33IHhyjG61Zj0EGGNuTIlyzE+GuWPg/d3MPw9Oan/E+xRZbvpdVZuv5btdT
M0bz/F4R0vdPKtlYsjbu9yoBeQM6Rs1h2X5eMfRprjoaHwRGGNhgz/rDJtRcnCM5
1L3fR6/JLpVESvO7KE2vyKgTz0aBZNDmLinUci8YjYeWrWUAKGI5XSMfgjHzyW4R
ZtB5HmWkWsw99arZiGeLzi9w+OW/v5YeFcAKhdtBo5O1P2N0P6ITz5lm4tHxeWC8
8dPWhlKUnobnxInDaPEPqX/HBoq2jZpZ/TTA+cw0URIOLz2J+pYM9lcbYRxL7hR2
9irdUg2zbLKHRdxnQHKz8110MJXbe/4wm/qklWl3ZlvANg55gknVB9qgzj/9giwi
QnxpCsWzF45eCZjQKC6YRNJZ6Ka/JpQCUgXcfw6Lyn5++fHd5agIAr4/3OuFhleU
p4HSuQnd/W8pLgLsH1DpuP818dywnXNG1dCtiCFMelBytjNucdPvYn6gXEI7lLzK
DDdOv2pI0pjZ2skX+V/jy1WKU8h7RIMAgaid7hI6icl2UKFxWSwi9+X3jyn13d/T
as/5kK8ThNfg2d/tZZA1BHova1H6iezCydqc9Z9OwWdmh2XJzwqCBH8ZOHGj9luY
zncG2d+IHYe76N6WvEE90zMqStJKJtie54P87SIh9HEaVdTtkF4GNL62W6iNmX/p
ei0iPeWJq+QfLSA+8Kv7BuXMCms+F1v/3KKEjx3OLBpjmByF8CeCYksd7MC+UHMj
iVKFxXY7uwx1BoLdgpgtOg97+6BxIF/Tx/0rP+6ch08oalONAatJyhBL/ikwVf23
F7aHDK1D6tuaynuBWl9jRfoqN4wocapaT2Z5GVOEHIRYFkxJkE8yb6q2o7I/0bI8
+RXdZxtpx1+UyRVPbibVpEYdliHQ86ReQC30zzR4j8PPrX2HPblIVlzLHqVUBHAt
HauWA5y5cB6DF31LkY9GkaqUJSwYdCON+hZmArea9Ua7vaHhyNQFj2OXqlvgohqk
yVgNF4NWVY2zfwJwYatifnZRLqR9BYtgRMXQVEoHK7ejTGhESnhZThWh3uXV+907
MSYYhG0RuW21TjMVXHiiHk+2C58kmTYy5IulY0R8dpAwig0hJNOPq9stRqM8vwiR
01km/rlzUzUCmVpLvaUjAi7gKBo4v1kZlLqFa8v6z4o7icgubXQS8zaolajOE5kX
fOEZKItSMsZhsYr0uo6iHMNpmgGqhR3ZT7VJAHmaLBzqJRfBCzBn85zesS4OzkMq
o82l5W1ZBdu1pMUWTDue7m4fKEAvBnNGZQskMarqNPgWL520WB4KX/iUllF5bbeE
5FD9MuI7uiT0AKvxjHZAI1UyM2F1TNG5PeilPife8Om4hqingoRsTAduBiLloN6+
fLBOZhaXSw4b3A12LeplkhIjnbtMT0ekFgC8BeMiDzja+H4UuAxFlMF5QQJKivz1
6ASEcOFq0KUSxNElcbUpZlOWoKnxFCPdLE4aUvIsZ8AzwQMLu2vCaAcseGUwsHtn
xyeAoVG8Ovlp1ZWp99GbFLXEw/1OoLVuw5BzPpI3Y1u4qsfXPMoJES1tIC7uXELS
w2HIJKrS4P/hYoOI1ovYNpmbOx10xFf9T8YrWyk4AJ5ocMu9hcZekT6y6Ic53J4f
CgcOA/OMLIZE6bnnK+gFvIUmlmX86mSEZpD+2Hhu82Y7iQL1fw87ev9mrGDhyCXk
skgRZvgbG5es831Gnraj2tgkOgqtfUJWZMjFYiL0Urj/sVldB7MDIxawhXSzF6+0
EDi/yzBYurAHwHQRJPTmWKG6FXz/1wZ3t7gN7hwSKiiq1FpLo8/Y7SxzFngG7iAz
ZcvHEl+QgWgKTWScR3EfBNCR/Y6DYKGB6OVuFvJMPVzvRLAdQBbAOxc2nWQIdFrm
TW1X8atEei03YnVWE3STvM6PfAgjUzP99mpzWAwnBuQe1KjgR3jfhSqsRUPNT6JS
am+yR9DKCSWAh11AWQlGSn5VctJQhXp17r7/Dxql7b/yhiM0TnMU/CkI4+lXI+/6
nvJ3DkyC+9V0XM8DDfR+05stNMp2lraMk2fzP0cM1bugVTWIuq6tpgaQ49umfZz1
mI6xIowmnPMmarEK82idey6kHV7aV9y6VW/i9XfxQlXEUkgM8XnCF24X+9tJ6c3v
snmAgGVefVMpQCgLInCshTny8/t/pZjh5zgdDXfAr8flmpiDGII//ZcDKaJM3oFY
NquWtaLqhPRGGYxcWE8JNLY8bD7fRVEBg9c9VaVNENfSHJUDKkXcrhTXDscAKB5w
nFXiJKvjagGCuA9aA0ekQIxdXyKI5xrEBKQgTr5fC+wTYzct6rw9YN1qJnUMaUhZ
NvbU+aAdT0UgcXVQhobfVc7xNK2590WqH/J4Gx/W557l6XOPOsVwulpVn9Yv/bq0
bjS7tHymf4b3pWPR+Y0azZAIGGwiz8xfvMNYW5H8ZwSmIoMFT6fQIQ3QwV1kbRUL
lcDq+Zyz8cDE4IAS3lbhqZnsCAQmcdwHu63QP9IZ6gL8X5zCHwho1wpqV4yW5FXA
8OnWziVkoOsoJithb60L+IZpVBzhhyHUnCV67neKB4wIVY2QQRz8UxQ2mr67nYgq
gozKTBIZngaX72+F/hj3zkPhYlBoDo7E3rsCcJMMeoWOa467WZnyrzqjZRDl4pl9
yiFU8KLMzLlrgR44JdXYjSr7qwt+QHdDXs1ab9Csvybr02f1PuFg6rOOS688kCAM
LQoHNk2GEhreShgmINNwH2LTbx1f56h6VNMbr2AtWn1WjkMAI/wSCsVttwCy+Elt
1g2X2d+0mk8R5oCMKZsAPzbTPCSKz3wE8rJ8++lnI5+kmxB2fXps/M/XF9h+zVhk
KgzUdCe9SyEsqQws40Y4eHWCghZDisTwlE56CVZ5WWNCy0/wEn5Rt30LKpoJELfv
i4Op2f6rx8iZqDn40MM1NDwDuFzrNF+EBEJJ2yuPfV9hpZGRW8JtG0lR2qqDj0gn
1PiKF2Iu3DND16STJsLdcLDLWtrl5xCKFFqml/BlcNNe4i7j6nhrGKLvRMYgj1XU
51JlL7q1AVLTyE7R/pshmRTlk0PEihwSWKSxVOiW2dHUaiFWVkLluAhlyB7Br6cH
bL7MhKsERJiTMQkOcYOFByLFpysBuNU9o2zO/N5cDC/meT66ygRaB3ZxvLlN+r2+
S062GCDBTaEn41/bktd20b2KUlLAn7bzYU423DdTjczA6O6Q7XaEH9TjwR+5FsJw
qnjRHZCiNSexyjTRvBYEm/3UqnjbJsDkjhybPnUYdfVbKlVnIIueshCmCKAuZcKQ
nzOt/ydxAjCbC4er7rFn7CIdV1lJBtYLkjjZmrqkwEbzMhdjXTaYlUP2FS/45Wlw
2di6mIikKFDjDb2+WV9NE285NNv7sR6aCMSHQCZ7awdWJn6zxO8mPMRrk6RTIY3i
LBSPisYolK46logU2Lu+n3cnQTIwLeQit57LmowDwy3RFshLoDjqnpMGKLmLM9fK
+q0nhrFYRs80bbQLpBsX1ETzyy7urzMfrZLku8ohbcHb3ry8FpjoZ20RJgDinlfl
dpERj80ZKCddM+yxzF3JaA7uHQdPsLw8f0tI8TfDwcvIkaA3MuteUpSgMcQNwnEz
TQ5ioCQvoupMTH7hSTf52k5SjTHfhRtvLykT89znaLWGurUceuFoP1xQmunCvhEp
IBniEJ959gXkIsRs+z6rn6LWoRarj9Qm0PEH7q9IhoFKjCStBnj1kYA3ZOta1epr
6KnXqAZ1Xk91Qm0wT7dY4qOIB6S+yIukw/Nxf3qUWD59bYCVcA6v7Ia/bqMIviO5
v9l6VipyIm9t0hT2VNaxUQAmWCvtePoCB2O1YEZuRMsaZIPmZf+9xCYUQfLRcSrq
BVxhCACzXtM2qwuUsFvpekeSRnKXb8sijqG6FGieIACjE0KsSWSMkE9VZztCyJRI
1WpMQiZ5Gopv3EhNeWcmzkJk1r0uWmuvm21CGKA0i3TfQOPkz+I9ko7W6N/F0dKE
rvHtujqNs1hO/OnTRV7UZEqrso4UI72LKBkCvmNcH/bFO7t7+/FULNuCyQWdtpvD
qlgubcSbyOywT7Glpm35qVqpkMpNn6fBrxNq+vUwrKP8mka8vZM3EeXlGFNQaeun
hDWU2yrEn7GnQoKCq+hgh45ajGFA377qW70WzEjnob6c5Qa6nsgmG0cpeEQz30gS
shfoPEed8ilp0ae1FRFSfAi0oI1NTXgHWU4fXT2aV19ppTm4nFm2VObO4xgBOZhK
SXl0J5Ns0o5Fg5OMiAk+8Rrh1supfNycOLbDibnwxbr2Msyapx2qGPM21CjsLJB1
CZ88CSiCqZmPMOa07KTtESSnn6fIZV3VmgRydhaSFlxrBF/4bfmpTsA8199qqSBq
PgD2LcZqP9UshoYE/ZEiqPuTDStoxREHQFPXVuyLYTrwILiXqxGpihQB1zvPu8aT
/1OpFV2iTim46215G/bNaddrIJ7J6LQ//p5ATmk0PvYCBtnG+s7cUl+5idE5jfzC
rXRco0uPDwjr94ymbv8rff68dmnMFgsDIkhG0sLbTVV7gEVdK/CUct8wfeDoanW2
KRYB/3UR0DI6ZJ7/UxE2j5bNbQ92+KDwysKNpIcLR4V411vqXilqkVCq1yzlPvIK
G2RfAik+gHaT64pmS0RZRen6p6qMFCmQZ84YcEFYeZC/vHvivKQMxVu9xJKdjJ5e
exRteuRf9FZ8TXp0H2J8UEzejJvHZ1GA6wpl/aFmJsc1ndJgcazjoge7SDpzGQIK
CoIpOrClceP/I03cNxtrjOYrJ4+53RtKoJxRzvbYuRFCW4K3Ubg44OZMzAGPzjj+
+BJ0YYgqnWwi9Me5CfwE68Ig5tK/VC4fEluG8WNjZsjpc/hQXC4fDKZLVD3W1mP8
/ZlijNUa7YS+DWwSgh1nQsQrMp6tAjn1MTgafn5XA8HjbCjQzmaLpuYPAoxTJwxr
Ewf/tukOccMv6ZE/aY7AvT1sn0h4sBYkqGAzh52Fw/ovXxCdYAGcnrLtbJ43XeNt
6LxgkiLfI20SKFqGynlg68g/7xJS3JSSYLBUW/dSG7T8XsSR42/7dZGN/HPmaiE7
oUmuMXdmQ6a6wmrIoBEJeJLeQr3A8+74oC4OCMjOCyrlcETrTAVHE95cgQx6JZ4X
IhXg+a0gi6M+xUfEAk8n1B51TIC1s/NPQt7F1ZZZuFCBV3S+ULjXVBquQPPgZN7N
acRnsFKRlKiawniFaNB/p+cEsM/G9ncMruV1yCWGsxx7Axlf3m/P74am2tyncXOG
/OiaIamirF7oOtw4u7ZMjfCVSKgcM6fopD+2jNfOHkkzrHsMPIt6cSFVU+Px6cFD
uNPyu5ZIt/QpTl5xnE7ZPTcdGC7LLamDWCUE+D5FERb1eLahK20Ffzc0vAJ3xGw7
NKmYexC9t0h5Gbwdv3FM5FOKBeWijTw7XW7iD0UXrmpmVQl4VJLElBabSXVMYSGu
y4OlZd/6Lh8sCCl47vrk0D00qkc+8KziFLG0o4Z8AbLg9ia7D2hBCK1x76Tez34L
i/maZnCP8fnAqCL/Of4UBduS9eP3wkDveEZMZ8wXSZHmOlmEeB4Y2oHcBYJ4M+Gf
mXwVIQjAD948wvJdGXsatqgFuP0rhntAMNyW4RMJ+OWGYYTyVhH/xAK2bFwZiaRk
DH0sXPJi9W47JASwlGQio7BtPDpWaCHHJHajW2ZbQOPHAAyHriD9A6fjwvRyuEMq
onxoHx1IBQYMmBeIJzOQP5AYZb78QSEsguwAmc6qmJrg1m6nvUZ8yOAYd9k+Ko+4
FqAO5q1TxN9jX+Gmz05JnfTfXDsOGD0FHkJ620ttymYLVI5T+aWVo6sloee2H/Er
+B/B1lQCU3pu4R8cIoZ/Qob+hVqE2sx3zqLRONFXtyB4cI6rOjD+GyUTQzWcZac7
xfdUbIoPbERY6Z9zhukHEoAaFgmoQoxDxnWcZzqW/pEwKtaHjw5/Sq6zUDjkwqCR
2J0v+P6HFNc3/K30THcWLxYgAd3l2bEIdryKW60R+ObaR2NwWPW1O07hhynnKpcK
izo7tXaxIs7NcCwutWFyazdF66iUASiI3Uxr+zbY43bKOdBx03hAyZRofkmzKaRm
mylLb4VN1rv2PluGjdrse+x8hG6uzRsUgoP1SEyDWOKegDWt+fWsTNX1aCTHob4B
k1LmSvIZguSk3Eg3o+xS2sf7KeGpl3mMQFXlZSF+L7xHcBHMgGccjisiRv3wZp67
whRnipHVZY3jd1Rl9Xe6lLroIHlT7OECBa6HnPwKyBM90a0KEFLVXaimy3AfOvA3
3QCSfajdhtnY/OsvwbL66Ke8L2sWGUYDf8aZTU5j18lSHctNofa9iCxok+U1YvXS
eWSRb4H3+udbicxHMVn3+ggR7GXpi9U1KKM/O3BjATKCThAv1kqhgvmJTSBI5rTo
J081RMBy91Is6T5rjPMmQUSsQlUrjdxTnVBDHZzU7HcjXEWh82JLekfzSXUzKYJs
H+lBR7ASV2njXta+xrY9otL7dUFBiZ3ZubC7b88d5Fht0XYAoPUkjej6Iwlj8D/2
VcMLUJKPY+3vU9MqzK9l3Tv1Fd1c45OgFWxYea4VLxANnaS1sw92pV+n4U9ZfHWq
MaujJY1X2kNZ6gMFl9Zrf6oJ8wmTdd+Qdbe8ofYBU0bYNFB37BJg22FCIFYnylGj
DLtvlvb7EQaGDC/pqZ12OSXlk0pPAuJT9TGo4r8MDGb6OEZGINbsA6A04DaPcx0J
uh1jbzHP5vd0btw1Zl6NBn1fxWnc9c2SIbdfSwW6Ne8b+mrKjnDIwMkFMR8E3T//
lSJl5OoW21g/DOI1ZAU+8ttqyXy/TzqaxZnJew+/En1w8/gt542sICp+gRIgOoD9
6QvRsK6+HcWBbaxET1KWC5Xo9M6k82MeE9hXSo20BqdvAwiYHVT3NB1W4IenUxHw
UANYwNROBmIrbhcSltTOCv1o+iS9bzMpL4z5H9GRdsxpfprpj8q7igjZTCcqongj
ga5XZLAMzCMWWShknu/hJljsAhdc/0uT9rXNo8qxADXgqO4WPAARyQi2YqBCELlD
CvjxxHmzzdr+Wvpsyg0rWB+qmrczwiESAeN28X1724OQ56C410MCIXsATsewC+JA
yJYhZXrhdsAGZHMI4kztx6lLy4qW76rMg3e0S74OrPj1ZnTzcdqw0APB23JxqKiw
xpdBM+B+hFKdjKoBho6FyD/x7wiUR5+MGTRdrPF/hZdOk0wyDwvis9cOMJlHGt9W
i0qfPKbQUPbaPXIlBfE/z50BVASyydSwp9qLCOO+70FO4TPxuKrhePxwnncSz4zJ
fVCo6zdXNp+M32igQTKzRpVtT5TFi8oLoyugC57fc4L2sAmib0p9HbtUlGQt4PVX
5N3A/48BSIxsibIsriniVam8V69Y11qmPzY1ikfcESc73A6qoTp7kAIOE3QQFhv4
LunVtzWENu0KsjT1pNwwY0d3xyE7nO4tC7TDTBNs80aQd8G3CHsFCejN8Ajag6JG
dGb9LP3dcfsXKdB1vF+gXmKWJbJLjrrc4XaKMXkFxL88kXqGpbrkjcurZoenoTEb
m3TiOwvL7DsgrXOu+iRBD+mK+bUu6X8xH6Vupm7Ft88XvYno2unC6/BcmtHO6ToL
dqJdHxFh+yqRydG9M0Ndsik/0RYQn2mKZDMYlGwVn+HHtYAaDW71jjrpqVSavva9
WywqcN32fJXn1g6VIHGEpxbB87JpFs+eBtJHfroVAMoPnLMBUCj8J4S1StdkMtAx
d3Vjz8YZ5j8JISImsGEcKhPVWqW2Nfn8iWO+CUfNUOTICZSuPES5v5TYGS3ASeHC
l1E7iTv9R/rIxnMjkTLaNbt6Ln8jMelrIM4NvQy7m7srYS8ijVT3GtA8TBEKrK9d
m203daYOaTqAF/Kdo6yLT19birDpGvSJ8CMv5XzjKQzuqhl7+n1KImEYXL64Ly2C
/yfgE+OfgrYsypozYErULCc7YKnZgv9KdNmpRCXy2ARwhOhH++x4VgOnMJ18Wjie
dSTp8lJHI+sXB95b3/UpVqvMDCcA+YWG+WwQ+dZ6ggJ43/8149FO5+UTk4W5NO7o
XZXa9jTfX9K26TgtVWXnsKIE1rEjmzUowl3M0+JFAsMHue+VfpP/pJGGaaskXJdi
4D0qiAilyllpeQp7TTkuNcXpL35LlIY9nP9gLNEq3Vj51zS1IWYvlXPFlx+oCu0V
6GHZZFKo3Q54rvNh/mSdRCpkpmQ4XS7FDVDE0uJdWG9yHR4M/eg9Wq/ZFwj0dvmf
yTEkaZB+gaByc1HPdDDYndXrePxBLcR9pKfIR86FNNSxb2tYsWldXdMX7dbvTztd
i1Mm97euvV5H3VaAcYKWGwQfsRCzzKOBAVnJP539XsJR3P2qcfnMGZ2ySwPJ7jM4
gyz5X9NwbOZLD1aTg0Rwkuy1AH53YlDS0pW88LpBR3ObBaqWbdFZftnt4DrhsddG
fkve9rnRkAZrMaP6Tw6SqsqyLs9ryVEaZPHEhDMvOzjVCP4WhzePics9s2VadpoM
4YY/Mbw+CXe9UJsXcwT7tS7o7ac/8+3bzdBkHQj/NUW0i1vuZVKRbQQOktk2yVg2
50GStWOsdvmCbQNtoZrKTfZs+tlKGmvkE8sECnny6wG1OgbLSPkitHLzadIyNEth
8vHCOJPKc9Qj1XxhGZZW7LorGsRlqnpTqdBwEOrZqdyL5A7cwS97eWZAgPrFUU0o
vo631tCXRyfJfuudMN7liZXD4hUPz7FdvH8Do3/vldrMVNGBYot+Ji6OAuqMJs80
HMZyT3Z7qClqLNvned5Frqi6RDrPKaImisqsWXb75/16OkIvbs1oATV0Mnfaqc1Q
HfSY0qVDLAAYTgVf+NeN7bEiGu/mn1sLVDEIWN5UuJ7uOo33TjRiMysowFipxG4a
ZnIE3yvqqvVIYi6t6sknrmvbtwKZIdcksw2jCwxovqVYFRiX5yF8b9+DKAjOisY6
VNxKynW0iiRU5EHqVZWuQTnz74T9+LTVYtAsF3+FQgciQ+4z6Sd+IUq5RIluKy3v
GnlknlXE20M8Eaj5UQz+2dXURsOteeVLGG82f1JFvxIPWLTY7MwecAk9c3E6CXCT
hN+yrcSy7Dv0xEFX0qhIDmGa1+Lclm4vN7/JYXYdwGDjBCgv5XQq0Y8Es4sX3MMk
WqL3CCCR13uKakLzal9OV/sBKlRqgpxsv+KI4PUVF67RkRF6YwNPfrgP2XVm34o0
G4wQR89wlMKdl6VKCDqQh1Aj7Q2QN44/3kB4j6+En5vQVySjoK7B3OhbD0DEiv+n
Nnf+jzEhxieIhFTcGxvWt2fCkc0PsBeU/1rMqEMIsL2UOrZJmnmz1o7b19dVTzG/
Dm1JT8eniI2yGCoHGRqHrDcywIrCs0gHUL2sYljFj+8/1sLk2tbaibfm7RDkUvUE
pODTzgNKUb8Oa26RhK4Hd57Fi9PoPnPjInf0Ql+NSpOZ/6IS8RzF+zftQT+zcoXH
id/mxjTk+S4xC3G091XlgEPVuFCGKc0iUQfacF9tteO7PUmuYFVGYVSVtEMJ7FPw
sevJYl6Sdw0ihjHpT/z32QMTPl7euv34QICVZr2mc4JHHNP8HWy9yvL5LS9qoVuo
sy9FW+ixWvYiPnQIjhBl3xHDstkATcQTFi2Q2WvibJkP6tCldpaH9cxUkhBzPPwo
xLTjyJuSlKQTkMT2yK6mZAFzCCEGrKmmxJdt2QqqKXlya8U9oEXmxCeNPG65kpDq
VYxenyzUm5CmXReKY1kOydjOPsVUTuC24iKRcGxO4MoWJCSCAvb2eVKv5JKSqk3t
l8UxhedaLlK72OrlOnTvQCGLl14D9Pgx+L0nJdw75SO6ruS4HAZnQ1p++r7KqPpq
zspmzPloZkaCIyiFp87rErvC6drVmNIx5g95Dk5ATpQFsAIWdajwHel3LWrnh39A
aMf7BJx3W7upM0Hi/2jNCQQkI8DIY6iAgUcgSSyd/W/GqZKptpXGNMuHWnZ/+D0i
STma9pZ8k/f7sKSwYPUjR/SVxcEqtDG13VmHU0y7DEV4S5Fkd2UgTNdCicmyuQGT
+KuX08cdOA2RivkBruiyXD7/zUa2JBBorp3VzVY/46inxlf7D5kQTdFvmmooPXbf
qX2ZfmxNRu/Irjct0fPCAeeM+FEHY0T69uyQojkiTNdA8xYd7jk7yqGuFrLHyZMB
cuhRxfDvlhc1Fr4U8KzQKmNgbGNqi8y8h3P1AvMxGsWp7OOvxNHPLzyXv/wSS0iP
E1XrJRXw1Zw8Mo1l3QgrLHhBpBTih1yVWvqhF0g3vmNGc6iSKQQaqnqiabkitsqL
unpnobTg6Wj680RN8bP3DYY+3ZAI1iEIrrMpUctRPP7DaH+8aP7vA7uw3GN7GOVY
8L4nJfGKho9LdvAG7Zi4S5BOK9doMzp5sZqb9OZkRE4Ty48SR2TlivrYXndL/3ib
rYtTQ0cWBL087UiDbXWrgfCRUJwrhOf2Uk+nPnNCLEbXYlYn/BtGBss38cMTGFz/
G95TIppTxdddFlesqSyBYqSzIQBBn2tm3n6RiQs4o1NSXZFKeTc9YzkatuoV6lPE
2oTNnzt1Y25fGxPdeIGMzzQPP7c+uWG77N3CSpkrzY0M/lSYDPXKXH2uoZ5ugMcN
YSF5DKGoWL0o3lMgreCXd1Zfifr81NhnVTUmnxbIrsMZZRixAj+bsf07i4RPgGRw
dWeTIRlQOJ4EBmImFcjYV7weWfS8hn9Arxg9I2XjDncWRf4zevGynW+jxpS2t65S
Sqey33NoKvkL+ybjtaUoDi7bkbzd3XyfA2Nq77FTnH53s4PXs7SBo1YvpZjSNP0y
kc20YE4CHmSmFz1btOAWe29XjQ88QvHDO6TZpTRbyUt/xlcxYOdVQaNKMuzqA8mm
gQ2ekrnJw1Z/T3G3XTFoSSLxvwCM4pYZ6nLKcmRfQ7p0iT11yzqj15aVjgmlOI20
vwwmmxxSRg2PaKJcDLK/f4P2dSA1lbpEnaQQ/5VsOHGD1J2imbSBNopQ+90lhMCt
zyGViSPnwKVayt/7UeN6w2xxjf8R+2T4Q8bKpvNLlhBNqcCTGbhrQwjvZbJelC+l
a8hHLoe21l2FIBuPPd89xbwmy9rjAskzRMp5K6oRho2W2JH4yQ2+jCFPJwSov2kr
6ytHwy1Y2k9IWNQYZa9hHGRk20P55ngGmKnX6nefo0Op52RHceVTM1fCxt4BHYDz
OUrFTttaEvyRv/U6NgBozGp0NkdxTk6ltvZl+LLAVA+NZiBDNGwCWdjS7ujZt5QF
r0r3TZCCWB1ZO43Pjj+SAVm6b7KQDv1K2Mw0nyldUNx+wi/c3maViWSuIApYfhXp
WpoOTOSLSj99s/8GfIu8h0EgetZ6wTlJ1MuPegGtQec+UYu3XxkN5qEjDl+4lpOM
qv+unKhhzcnoOwjlPEY2T/38cYeVprEnLg3VZGKAHD9APLWU9ZX8o7DKBo1NlV5O
g/TkOKEUZbTyYgC5REJXzRl+aT8sgyOtaEgjTYci3FmCcGlpZWBajCQgFjCo/sSG
3x0Na9/07WCLPsfYuhoNfT5z6b8tqHS3whUlxRio92+EuCXBfzcJbJlk5/9oaWzA
Q4rqr4+wErMgyMoAq+hvuikQTinIpF0oVOaRc3L7QQ51sebxbg3J7GfiFeGKeJUM
RCnDFyZ7bH6Qnv3J5MatlRfYD5uXYQlp1RAtUoiUZJzME/zI7LViYzTx9HK1/5XF
6eTBW2qDB7JRs/9p7kcqIzYRqG63VAuieBV0qCerTl4lyL3UNi/eaKzdl4javcoA
WeGzr0aHyhtyL+p9GSw1Rpm8fRspcPiWxmHzSJQRzDH6NAGjb7GDpyZSdUOzrDRY
2IryOR+8fnJinU6JrxKh6qSO156wvFnY8nrbfGRqpW91Ir0B9Z2NQE5H2ZJXOeXW
mczo6YT1GkV8ITyecH4GFj6kK7ZG3qxDRgK5vEnMhVkXWfidB3O2AJm3PgRt1edj
l9XhOO4S2FMEegwfjGOrr3MUazYC1Em4b+EjbzRpL7ALrK9fW/A2uUSI5dNUeAFn
dTrhLld9rE4g53pKwnpC4MGaWmE4N7jAp8IR2PwkdzbMEITzl+57uq5eneh4fdaC
HBkuqYaukbCe5XR8PcHhL1s9IOHAtQQwSfc2Cuwrvh+TH4pyW9H7+6qLaLpI7itj
AJWkoOa2iDFFnVbIfLqSQpQ5E3++h5WRMUW9XuHvvjfDe42u4dk2bKBXHwAVK2oe
+b6s8t/M2gYriXk/2DMlhGw+TPXRtLtcXC3a/JTp58qOCKsZ6XCJ27eAZiTc4FSe
Cnf3QlUx8VcKIQ7U9PLJQWQdKV+nSkwlLP56InShw+uZ3xP+92PVjByKWIhbcPCX
HJEoT6EXqp0BKdLWtWF4TZZcwWzj5MXRQTcBbGTjZ0xp/BoZfE9s4+slskTmy+nn
fcum0ibO+I0o/eDeWcCN4AJAnIt8viU70j/PFsdSEmMjPKFr/1aiRKWt3z4mRHCQ
YqNbeOa94kq8HgIjjEKEgxQ25G6eOS+KTXke1R4krws2goQc559zhFx9vQozXIbL
igSpwJ2s3CGbFD10w4IBfmiw+p5s3LijxA/ausLwn+OWsMokN+wM7ajM0u2LH5SS
NtYexHUGPD6iftAsT2vhiO49/rbTdHWll3IFGhPjvObOtAGbHVPEuVp0XaOFjQxc
Z9pnRGTJtjQtX1XoItAodjBPhLFwUk3404YlUGjHC2FqQEn+WHxeC8nw7px2A+Ux
Nhx79gRbkhQrvWPR8d9p+vtE6WYmh0Wc6arJqCa8BZyUJAhJQS8Um8qaYw9oilJg
R08QVxkWC2YRzCToEoDIi97iXZDsaPeuJnCX/OCQafeOHY3cOuJS1vc1Q0RGALpP
/4x4QqwA3D43e9A+rQhAhSaVF1bxwRVqaSDvM2XVzOQ6mokm1pwBrEOzkiWwPC5n
zrTKsj60QKp0Dde3TS+Hg2b0tw/PPTu2JTWVwMaNamj3u/WbSjZJhJ8co0LoejLl
NS9ugvnYg/5SuX51w5M/QzwPftW+73avDxaWV8Yy/3fYQXvm46lHBaVPj7yXE1Ku
bHHfOMCx9MFc44DSap7OFtZVXVhW+w9KFaOPjgMx/3HeW84i28qJtKfqxe6VYhub
luFD+0C8sHtcef9O7l3vJYZgDOvd0tVucPLjCc033WlLCThrJkjIIxn5XQRiG99Q
kGa+QggrHhl71hm+biAR6EYP0WN24kaUlmj0f55w1eSdnRfcUG9Uz8zPCaHh77ba
JkMS/ZwlPep8L30fGWa/dkrvV7CHuMvlJiUNNiWlzKeHt50drvA9aFhn2fqM+gZV
jp2PHa+G+RtXPRU4IhE7vHSbVOI9pgZp73Z7GrFh56+6u2RAhy3miIIXDSiYQLky
rwtAk0jC1erphraY5J87alDn0w66nxRodDhcn5+2TU6lTCDwrOQxbdKHrNaghmR8
XMTlib1kAjKiSYEBIHh9HY6mC55VfzMYXGxPvhFbMJUHLsUCwWgj4RCSC4qW/MN5
H69VYPnXMSOaTD8UHxU8bDGACWOdO/TtIkFuI1Th7YKwDzwycCU662PXFPzQP6I/
KYbn1vgZjpVmkyJZFjZUEAY/lKu7zpPiatmYCGBaSJ0oRl58SxTeaoju0pAgic+q
/rSuh7QnankiWW2QrX5cBONbOK1CpXrb85SWI3xRg/K0OLMSgv8oBNvQjktXOMFo
Lxss5MxITIluHxa+jCBHsUeA1dj76m3bRP7lSxIXVLa3bD8W5GepPQF7IRAwmxrJ
RHPbPj3hOx2OswWTx6jY/a1Wunr5r/Vr9AvLln4GnpE=
`protect end_protected