`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
ddtXksX2+yylW5zu6QL2Lhnb2d1sD00763mmSITNX595NcHTEkwn0zB1Dry37fOW
FufOhVzEJp80NC5qZ/+F0Vk7Ik02dIR0elf3clrjeJRK85K4e3Hoo4xn7YbFUIms
l/8VZSb14+JVGURjfswrIyCUotIzlzVYZ6gzoZwDXIi5gQIBf/gI+KxNXPaKV+PQ
Ufys/12rjO6aI/pPlqSm0hCvftmBcnezN2hk1UeXgOIuKZnogjOsf0iJVX2aOOWE
6pD/psybjbnsNB6kH5uFTA5frkzIzkzl5d9+YDm9OyC+k84E83I/7/j+rk4L2dah
QJOvksSIzN867/4Qt8qYTQ==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="MvBXkzurAa5VTw+1JJ70nePUfoQXBvZOku/SMmg4TwQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
oRtzZL4VJ4iwysPsC8SXYCzXS8Fw2gtZTOskLcDV+1B9Nzn1zTyNtlo6lNICRmmK
ZRVu2BmCc2G+fmzynYlNTnSa7C0Cuel6FYpxCBlOuk3OF2tzAmLAuDyOH3Z1Yjzk
a0aHuoCdIRKv7BrZCdALt03JeUmXKPdOmIlkVGFl8yw=
`protect rights_digest_method = "sha256"
`protect end_toolblock="Jn9CQpRhJt4rnzZPRk+dOpzAubz7omckX1MrFd4p81o="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 3376 )
`protect data_block
gD6l00tciPUa6pDNTk/+t0OO0nC/UTtBwLB41d4inuAUA3i/ALrNyoJVcBnAmEQW
ptbcNp5fxEUJjnOxnedyZEuEBxWRieZFQnkRdF269oOv6LblK32wBMhUdx70BP5a
+mCYfghX7zPnkAXOhWHs45cKJLfTBHT9Pw77ohAUUQkD8TjNSO+Dvb8sY22jMgvK
LyV0AmEW4lQV1HSezrEZSFUO3SFeyk5F3zZGgR0wSwMWdWr9TmbjWLKZwRQCjts5
4Vjmffb60GC8Re/SjrMTQLFCe5Mx6hH9TZriwyCj5zajmy673o/DusG+p04VLD9t
Gn0YI3tykfISfxEDuwjYNE11iW3o2iY8EImP3lEBF4v5jTyx0DwE2Zem7lQ/JVW4
45aE62g0cKcLzbGoPSGZ0Hj9sdgR+Q/IzJs26OxUZOJabGZzZA7ILi0PoVskHxrk
okqfQ5K8GZGXS9TFh01bExvnrwU4zuXPMTNj+zPIwmHHaSb7jEy/fL6SGg/q8g5e
mg3VyOw7WaYgOMRRYwUVPXSnd/TQNOJkeNU8Z+n9Vy5N6gXEPESU2p9HCLxdfgZf
L7AUMNWwX2MsqY75/KHP2+XIjswEbWkbSSeeorZq+HWdhXxHpKf1AnY2hB0kiFP2
iqHRyIGqKk5RKVVJAK4yC0tc4PYIKK3E2lm9kH9bodbMps/iSIsekqCuDIgekNb0
TjAt66mxyBMpWvxtegLQJj7PbKDf4RCSjNGShWpXn2c60oUah745vo/ABh1RwDKL
Aqtt90UxMAF61InIEjPnKEQJ3Fb45Zmul1hsR3Qmf4ar8Ip+HDdkD6p3+3OW//8D
zPkIOXgUrYrRDMWFGlD9U7rJLLY6Ltw7llTkYaBJG/gemM7Q6iHvU45vlRZnP63p
/qrUCSYff37s+sTdvH5MV0qImCGAL1y8bjXkO7FfXJhc8x5PJU0NEZ8i1MSdPFCI
RmEn5RSSNTaeFekFSvGx0Fr5JNqJ7GZVTXXGOMHZLgFn4fFFLs7edKLD9uaM/9vg
MJ4TTaskxquefQ/HS4YSXFtHzkcbzKnN+0sLrkjJsvmrzjRuxwYRI/BNJ3b3qaZc
f+9J3HeskWYFJRvgZ//HuGfDBhF6IH6oDt8yB58eSmB5rr+xtgJHyzktC5FgF8A0
jx6xDfmf4UP6fVz2QRaDaJh5G9kwsG9MrdXdoSSlcwSbiKsccELFqrfF4lVOqk4w
Qsbh6S1GIdA+Hch3AzhRAdwcT2GTscUGSyp/4KxwhuzCXCGabUERthj/cb7QvGcM
5uOsds90sotSbfpgxLimwNu7uezSL8KFmd2K5w8HSg2kj79DdwceTzjanEDR7h0o
Gc3tPNBWeGwm1V5eXmyE7rkIAIMNSLJYCvQjucRMs2H5HQVOml0P5+aJHaebcPGT
rX0Vr+SmQVDsodxyMI96WcxEwQug5DDTeChCeV4+4WjJVs240YaLUi002DcZW/pb
gAwi4Ll5aCExTG6MfTPtDJ94xkn0d6cwnadGvcEyZ6+30hRZ4wfUXUG3tmniFUqz
a8Mxttj7o/BUGU01zcQAg+XCF2oWEcQG3dnWszSssRKWJcu5J1zsP9bMIaBDMoRh
MZM9wptQCVhbOP2WPkQzKAftwUWHKRG90a8lhT7qCbv1HGGnrhA8+bpcxb4ZUcFz
kvOv1sUuz7yozZqQbLWxxd7RpRKRTIaon4K61I6A560YJhxNhuTd5NTH4jVKCriU
JCZ2bivlvuIkCRgqq74JLRH4zzm6cr3kXkeESerEGZ5asVP2fzh6apVcgiR+mmYN
qMpktxGnVVngyrjhm727vYMdPxFWXyRqz7Wj9sB7tC1TvARqax6aEeqY+WyBzxH2
9xXppEVsqTSE7bkL2aar4lwh47SZ0sPkT85WZs+Q4WD9wt9X7/KGnWAuxGMQjiNz
tSmyAOVgMrRBRx0GmYuX7eiWrhIYZXX94Ys93ejA/59Fn6iEuA9OoyJ9psXCwUW/
kCrV/9Pr82lbAssdVlwKgwXwKj5if4y7GIGkwFPjSxjMoqUd0aGeDBlpMNVVlGyE
i9HPGTuZjFu22Zz1vYp/H9psWHxqJ5HisYH8/NqIogXyT2wQVyQTwauzKP9cH9Bx
SBERFfdcytqvLKlwfbrX3hDScRDRVnU9nN7Ef7jA6sT/SIVJfPbSTWOQGMFkHO4Z
DtGKve/BNOsguPe8ZZNKXpoyoz9BTfFsKSJrj+Bd9q2GJ9ZPmtp3OSMnjv0Ex99S
jrg7rdf3W/t1baXnPB8dynNLsaW1eJxPtWx8/v2vJND4QFmKPRw8W+Km4HTyOkeh
5qWG7T2N3lHu4BInxMOBrnCjzUivmZh3XB1mBLzHChW8ydWFQxe+u20WDqkRx4MG
c+ZJCqnISO9n179cYtACNaryHsnlPPcoSxNnOe4URX6nr02c0GtJZcjk4mPCTU1w
+tgwHMd4MxiUY6hPJgs0mtgBhUR2xeGg0XV/gfBWV7ThZHocUyeSTNCdHx98I6jQ
U4hFNl3lUjuSVwytwS4PyPZzTnScrP4Tz4MCdSIDKHcsegCfAZRCOAYYpn5Dx/sW
4Y/oz/pcXQUny81f0A5/oX8hFeAbA9jOGoopaeKGUHUaY0AC6wOgIoiHbfz870d4
zqo7iTojEBBSWmrx6tim65qm/mOjB6A3DLRDvhEdtHXC8USyse6yudl0/f0Hm1aT
D9yrDSyiJS6QICp7Xw0VSRCJmqDLl/U7FDVPwxnuGtnDvWSNkJW49SFXHZNFKzVP
VVdYDOHHMOd0rSBtch506NSgBkp0ZNPLSk0vKYOv6hWHngA5lAqvr3rYyhnwdQcv
iOhtW+PCjGdfZsuowLbk20TSmeU/BXj3qD9ljbDkU2kcg7usLWa+dsAW3J5JRXQd
9XxfovHijyRLkvY9UXVGyBBOoHh7SJ0QWGgri0QjXd9P0eSKQbmiDOvNhD4nKTMW
1lgmEbKQGXZ3ADp5Xxe0PlSyMiWLLQxmjWSDeUZ4uGZlWVWumL7ghvyodemHqUPq
mQ6oZvvla4ia9KjZzQQrnSAVb7afNh90nDlSDOWBodtWjfdmq3e4puQbhJ5/r3hD
if69z5FjDDlfoWJYZEhcgdYL8mEvSVtfN1ytUdkBaIaqen+ZB9+kfNcXjjpSKH5k
85RyHI5riZoyei0baOirKT3QNbvu43ImffMtkH/cnqiCpyZwwGZhXDWdbwb2Ms7d
B2tl6bexUl1h7XjUe8t1lePfRah0bKy7WeWXAIdHR/buaYJjakP9fdThIzICTOAf
Ftwo/C+V1Ya/6dP005/jjMa5aQs+j2HV3mk4HuGidjD6HztvtUtS2i5cs40vvckG
StodIGIZiAt4mwPQmZxmbFOqyKYUfYB7POo9SKW5jw72aojbnoOJjNjDSRUU/Ta1
Jw0QPTABkwvuoetGqInEA2UMCmZB+xB+4pmEFYmwoUy3yZZk2xZkiVl74fdvfMpc
yvwF44+5jMcTk+RtA7s+Rpu4y4ufwTH8WMJIKjdYXUd7FEPjdW8yrAuQr2gUm4xO
YTrSNj4rjpdHSV5EqckiPIGkGiwIFm7hshyuzRjtyGyBgPkxLXUX5iBJsSgpW09e
+mWlkhXSv6QgO7IztEg+hkLjwhXe9QykG/9snPnpKoncA1rLhCxKZsLTxzGmR7h9
4Td62dppUzP7MfEej43T1i43dcqZmJcVOHO9wUdUsfO0VFtAJjdBLizxvjMN6+6Y
Tfus6lFMieTrapp8I9J4XgjznYFgR4AWCB5sskkh0OWD8Pj0SJX5eCFIl3ubW4Y+
YyuqyEwzp6XjMhvn2+8lWyzzAiqkeGB31QNIdhlJypEdXCWMtF2AQQgjUD7rvEBx
YMlIxYz78lEdxzjUXigAGCpBII19HybMPxrk9kQItsBdVPMT8lP1Q+tdcgjRm6MB
TLZmMm8ASr8q0slmHaSsH+V5HlBKMObpCAqOVVSeovWCWDHUt3TmIMZS24cDSZA2
6xg6F7Ga3VaCZSEOUYzFr2exyjUOma+X98Qg2IFfJOSlrYk95zbqgPmIHoRd+tHT
+c67QjEBGpY5MJ0vfDZSdIvTHvtCRMH1t9C7Le4gjywCV2iuvSkjMq00mirrc9yk
hZM+oz2OnGm7pWudskPOdEaGkiLcSvyznMRAWh7jU4/lSWIDScExXPGTy21OFKGC
RWNLH7DA2FCpHPHw0jQjstMHx+enSx8nVrRqzA+Js26lRYRZttoh8DfESdknQwMF
hRiJN945twxTp/6V2rQuiYhfXlAYNhO8cp1Z/ln1t/Y5IIa6CVEK50UDmwp9AaFc
iVB/LACyFCvPFDGLf8ZZJ/+I7owPUXmJlbwxhgv7kMyO+jxrBnr4IuSKN9BGnUWM
pclK0rLOisTEpSHOb0UhTeBXrBNQcIbWPyhk93W41T5B7oWdir8qJiNq8PQXps1c
zBOGKHOqFOKKqXOOq68ibfyuLJZzdSwMSbxyHS9J4IsKsA9dVDlhmOABjsCAct7q
e9wuADJvz0Qd/o0YyJloeQ==
`protect end_protected