`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
ddtXksX2+yylW5zu6QL2Lhnb2d1sD00763mmSITNX595NcHTEkwn0zB1Dry37fOW
FufOhVzEJp80NC5qZ/+F0Vk7Ik02dIR0elf3clrjeJRK85K4e3Hoo4xn7YbFUIms
l/8VZSb14+JVGURjfswrIyCUotIzlzVYZ6gzoZwDXIi5gQIBf/gI+KxNXPaKV+PQ
Ufys/12rjO6aI/pPlqSm0hCvftmBcnezN2hk1UeXgOIuKZnogjOsf0iJVX2aOOWE
6pD/psybjbnsNB6kH5uFTA5frkzIzkzl5d9+YDm9OyC+k84E83I/7/j+rk4L2dah
QJOvksSIzN867/4Qt8qYTQ==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="MvBXkzurAa5VTw+1JJ70nePUfoQXBvZOku/SMmg4TwQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
oRtzZL4VJ4iwysPsC8SXYCzXS8Fw2gtZTOskLcDV+1B9Nzn1zTyNtlo6lNICRmmK
ZRVu2BmCc2G+fmzynYlNTnSa7C0Cuel6FYpxCBlOuk3OF2tzAmLAuDyOH3Z1Yjzk
a0aHuoCdIRKv7BrZCdALt03JeUmXKPdOmIlkVGFl8yw=
`protect rights_digest_method = "sha256"
`protect end_toolblock="Jn9CQpRhJt4rnzZPRk+dOpzAubz7omckX1MrFd4p81o="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 18768 )
`protect data_block
gD6l00tciPUa6pDNTk/+t0OO0nC/UTtBwLB41d4inuAUA3i/ALrNyoJVcBnAmEQW
ptbcNp5fxEUJjnOxnedyZEuEBxWRieZFQnkRdF269oMmKf2kFSxRwb7nyv8SXM1T
+Aold1sw+20bAVHRRTiBdHj3S1hGLLzlNceoFeCxFsb6r++CXm6tn0Aeoi/yErb6
yEbUD6TC1uViXhIEB6313xyGZ7/QiuM9H9N6khTSZaMcqYp9cIFeQFjIJcr63c8E
e6ELffRstUDANlA+tRJnYwGV0KcImTlHcbka0LpHjK8CZTW0V/hBpueSpGeWIjt0
6rVfUpf1rSdJbHyEjawSJX8RIIFfryP0M2gkSUctf5Ze/rAiECNqZGHIYtE15Eqr
dG+1bjaghq3QC+woXaZymVj6fCYSyoprl5Mw8EF3IvHCkh/QBhgKLdPQ79MbLOZF
p4jPsJTzSzjuk4yGB06HHzUN5F4DmaZwP3J0TNPuJwtHjoV5ALtSO0DCkl4F5Z63
mG2pJVnyvzow2lHKhdY6uC3O9gCpRLEJVyQM9E7hAEM0abkDQRi1aigN/QTTfQTv
tf44gVKrC+ZlRPgWw2UA9VfcJ/SwsPd0GOs99HGq/idDDDdSOQM2kCF8ssELldJh
qjEnDSq2mV7dBJmu1YSJlS1WcFnr2yvLRXLxPL3PxvqCPBk3iapyzdQwt6CPviBr
YAlAqVCMYB7x4+FZTqleLngQcOWV2Civ3Eag1QtCgn6XC8TeauIqccHiatEwyo2Y
NPTdsfHoNFF5ZMLSMqbyK+4R0mpvPplrKFP/Qn21s+eg9/RavY0+BkSuY0YoJ3O5
mFlkcjFJrX9762OAgRLMnOVKTjQkf15ekxNlmC4dhQFyfBtXnuw4mbrvWYxBNqo2
9WH5PnDNtg6CMSK7U8bQ/VDT5vY2NR/aRR+1yy96OpBAbZjgNtzOVzVEV7UQbeoG
zDCp5cLifkbRuFgdYNZTxrFFs1+QUEG3w0sp3fBggeFEBRRt4nr7E3ImW+pBMMn3
nrD5Pd8Gz0bM8S7cFEXcdRvPPYy7evVOitvR4UBAotiOkLxSNqK8nM/ZdrYneIWS
tfR6GM7BSMaLx1JB/CA3V3INK6odOv91AMETppClVf/uqYFn++MzUvNDH+JbgtVR
Xsvl8uyAfptv0YdQ0Z7jl21TSJLqv3eO5NqtghyGd6ozrTayQc1VOAqxGzbuXafI
2yNUH/Z/wNuku/lyXRVRjHJBemlum7eW0brwKrVsDI8ZpL+toEtxaZHP0/WgN7lK
8OEbbHKRi2w0IU59vnJRx6n+B1nd+pnHwQ5B7OW10P3XAZQLIKXwdtipECZsDrXQ
fdFf1ekcIilqNLcopStS8x64F/JPhgsdam1Un7nipI06EHA/OEFjuRNBz06Pn6YJ
ne4CJUDY5jl876jDL6jtln4x/eTbq/IJfj6zsL06Ylu5Yruf/2ryk3SZowRQMJQl
IHQ7326RWwOFrlw+ZYKaleMzWcjzYH5PyccISg8EmXvfVdZWKklTz/Y3+Wy4ZARH
0EDqtQctCoMlB20wdCua6rk48e68HQEHQbVVY4gXJjObMZsF++b9i01F9aff9se/
Hgrcg+BS7Ecna6hDQ9yFwopvb6xZwImAN/2ep0LuWZIYBiZf3ncze1YaTiZLSElL
C6bXUOgrguyjWgfHkfBBdUiwkfHQyb1XBgArcl2o9umXMBl8hDcHm7L3iau1RqeJ
SjGkqpz1oREAXE4UbMmI2JMOYRfjFMZAe1svtPuXtPKFuN3DBpcScl46xAo6gRdZ
CtNhtN/gvqF50SdVGIhyGKkV1byICd9FdkLmx2szyzOFvJWXChD0yxOgMOfZ+Aw2
h2LH1u8vFz+6aZrbwPVZ2SJxqmvWYMK1DNPsXb1rukbCfL2CUsmJ7yWCrnKlhiBg
hyHO7SCegJJHKDrZwmMwjQy55hpo+axXl/QkZSI+ME5qW8hxDh7bCSbKtugueDlu
l04K6289tVE14pxa8xWtFZjw8NREatp29B1xIWnWlVl7Lt7QPzQbXrl5cJirU69O
hIypznKcgSpKODtVlWi7TX7vTxhmN0e601ZA4BuVOEINOcipn8yOGeFXVjgxKpnW
86XlQg31lEllrUPH/0OCmunPBG3sPqumWavrzjWhIUIKX5qUSNzdnn0LzWnq2B4j
8Kc9w+A3mxw3oHajM1nP7m8WRmO0lln0SLg0D5H++ytoNhgnc/nOHX85B1Jkj3E+
KyuwAGcH8VJq0lNOzahoZCkDXHCWv1XTr3JmdxRKaJOiWBkkfG4D576iutLOJ2if
2N0VFwCez4O8YsMTFIg7/sU6L0oKJIldaYSSxd3YH0yEKY0Xi65lYQa8c9nIxDT/
0NZCcVjuFpIt5MyREXR8aWPy+f8RknFO78ynVXFSEbvxw3N6SL6+fHk5FMurSNgf
OkI+9/SbJ5yJ9ljcGTByo9208UnGSzR2txLv1czPdvAuy3lhnRu/yeUfzXEj+8pv
Gx7Ec/ywbLk2WBbAl5QI+XClErfvRQl49QsDKUSI3LnBkTn0rNYnuMINh2ojrxAg
9UlLd5XQ8sBtjVv/0ETAsCKOW3O9mf9PrGSnGj7KwJM04bkcE7QIpH/zSiCAXSUS
IgmlbHnz/TXtkCKprFEmMahg/d50UmaFULzyy6mn9wilJV7JF434guPcLcVHbT0f
FDhrI5yBxIrvNfirkEwxhLWxt8uFdl4kEhRWCMfTnwtrUZXUcy25AtpWnLB7jK4K
mrUcjKA0rQZ5cvS6u5RRJctck5K6CfjeSGeOB7jJjDCaTWuJM+Stjow8E2nvv9EW
fQvISBF1Rx8JplTyfGQWO9X/rR3xmoBalYXRe84037BahcemlTn9y4jQivL/ZWzM
Q6eBbN3F/loU+g3NU1DH24kXy+oq7kieOdHLGMv+dNbyQvE/N319gme3VI8qZGz7
z7XCuFlyoYh1an2CAG4kV+3pO8U5E2pm4Ab3Q720gEv0mJJrgGhTHwFEEsbaBJLv
s/XyGKn7i8nLwl4lRtRKPQcC4h2ceen2qSIGYE9Dpuc9jsJ/G9Djp/58P5H6Y9Fw
xLTxQYvNJq31lvc63dRvOFZmz2FpYAKKaZgDYQPvoMoCZ0Bpgm42+xSN+CayO0kT
NUhFpm6FXx/+Z/tirAZUpRFjoA4PSyLoRsqebomaLkBsUw9NQjOgg/wdgDwh5C1J
JMvyQiGFaekh2wqTg1lgDifCuCkKS0b6CfS8djga0W2D422cfF0GZK/E4py4qAkn
Qi8Od4AphxhsrHDqTNM6CML7ZMCnzxDp+vnPs1SUqVoO0jQTC8AigBLq1BdrOszM
cYHI6QC6KHmFxD4/W1So0BdH6bD9mqjpKlLsUTOARfRWR9khOwxRgXxJ8hdfT2wu
HJmxUiIT908YAQ1I6lI+rO7Lipix1ztS2PLIQnCEdb1zx/ckgBzkL0QuoBR0KW1X
oVQvpIYCJ+zgLNlRnGt87hbp1eqemeN4IMoYRVaK/ssH5Oc6jqBgwFSnHQ67HdJS
14QZTL+4/6WWK6eqPdQOKdFyIb9l+z/cXWX8AYVrXbTWJmhHLHSZwyw0yUTshgBN
tkNRGZpkONSPNQCZ4GsLw6sg2pQM67CVfgj3eSlmTAh5rnMR7KL6JKmN0YuOUFoF
N7QZlXzOlxaYnF9gCPsyHSNxcAvCujq0eWe5W1jgMMbMOsxUhAMoZNvGmbhz4WC2
8FlD3vXlJ4flaXSIMqo5rMzu7ZpUEnmnidX+XFZM5JwEeh+/YHFMRWr4kan0N1SX
6Fq49lvr+nq73QVfX+uEP/oudGD3X8iJHRIw8l8TnMEHV/haiDdrKqqnbATta7bi
fdLiHNgiEWLSasS2xeJI7at4VXgkzZutlFRyT5oCHoi2IapQV08CxTwKs6ak5toU
s37joxG3L0VCd6v0mvsg/GyeUkX57puPvwM3l1cwxJRYWhQyTdbl8lv6fujFi2fU
RcEx1IkWHnY5mk4zwtCzDfeX95jhVrGWKASI6olktRqb2/22kcOsgmBpBFGe4uPH
EyFlnHFpH3+LvOsqwUo5bs/zOcwjFTYuvp8VzBFr0OP4Ywo+I92E1NpaABSlqvVz
E8ltWh1/COgAv5sactLIIuCtb3LVEb6Yn67RVXR9XqX94FNhfXBBP6W8uhyHWQX8
318f1qb/FJytNoJZsGLHTmcFzDJuzEQCZ7iiozgZ6l3KLTnNDKpNH4ZR279A38T9
Gqlxvp4jEe+B2uaCwTZF78Tb7qiXrwVsxu0pwVIgobSFRFUcOdlM++WdODQnDNzS
P9a0rivnXaE2Eou5BZPFvCOGk8XrggFg2pgsnKAy8aADf2B4PPKUd/6cZ/5jQlzu
+W+NRCRQpiK3vCCv+3UtnWH+MBmo4lqYzGWeI6jiXGgb9U9sc+qqGLNmtJjGyfSi
Nly1htSsG8i5aVwF/uz9XpGAXQH/MKk5rDhgcnT2fHB+q4EE82iS06gxo/FI6tes
ugVmW3T+dKa7Fxf40vr7kVMyvTLtQ+5RMf6lDaRl7grmB6v9Jb8tXTx3cx2Hz7QB
wMV2+zIFZe7wSjJM2mWl8t40UMJeI+vqVkh7umbuXun4qnlS+iRJtXPpYZnNSWE4
C8wdq8rq1YKi1efnkaM3UexXDq90jQhzZ+QKtOyfPkiMLSz07jXiq33z3tp7wFsz
Ty8jM0Zzo8B3zeScAdiqfYdxL2NxU0sNV1ZgZ2JcYxihWHi4JAK15kHWf/ADJpT8
Dzr8e4wmpte0xhPveCevsRUTLGwe5URZmKIzfkp+yXQswGVI/lnHcG/RpTFXMSkN
W5pyZyJvRrxkRRYiKyy1pc08OtAQ5uJkFDgsvjZio6lIQUW/NvT5eHBlDXrdwLu3
Txy8h+Va+HqcO1Bl6fG0CBDCxZVQU9onH5v1YSpe3QKpkBIiEmahY/d86vZGwAiY
1b4BxTux17isNxvtI6fhIY91MEsSb5UUUOcXK8hxB3YUjV0aDPTiw2wt7iXHP33d
dlCvNUt1Kn6pPYl2O0D1fKNDJJw5x/m0M9EMLD82XIsTb0L41U/eh/V3tkQHxExE
JPo74KsWrirgbIXGd9gfmG6NC1PB7K1Htn5TzgipCAxlZvLii/X2MZMV/peSCYlM
h4bagRf2e62eBUBy3DAM/Z3fuaDaCn1fTk85oH/sqTk0CCqEwygxlhUEJ4YtKSVN
Vw8GpxsgealrmboCJAnUirthA5sOSBEMEVVp1z/fdiKozz4j/moxdwcPogb+lYvN
NgQCBGLs83bnYiZEo6rNrPW5STxlWXPLRFBuR932VhMA4MvMsRVC1Y0eMXnO14yD
2dWWtI/JY0reYgFzz2NchJ+tqwE/aki1hxe2OZV9MD9MKLVhAOckpIwzSzfK5PtC
Ik56TA3j62flo+t9ncB3gWUcitx1Ug2wu15+YR+QB3ko+Aw6lSFaMk5MHhVzpBO9
g/nVearM2WzVrcBfAhLhhaGm4zTAYjVWjTB7nTCXtj2xG3sM8Z3jDM1uHS1NBe83
22NILG7KCaYHKkhYDzmpVymOZJ0kX7zQ0nMRmhHndEMCi9YYBedPbCcf2M5mq9YH
iaxehxzmg1IOZZymRiHvelvErszakTddKoKPKsq73PYYElHyu14U2U+javnPEOpg
x6qVKJRQ9FnG/BozTiGFa5GRtYbwi4PZ5bSMDbZYOe/BnKIVDNaHLn3ZjcpF9tMJ
VeGN6an+CguI92KYHBVlvp253mteZYDkfRVuy1WLo3dC5EHszYnrb9Jcx81eTBeN
jD/TOlPUnlDZFyg/Z009x7U3oLm17M1cOloi9EF59yGe2S7abyql8ym4M8i7n+E7
JJUHrvKAiOG1r/DIoMC3BrvLyyoS3dXnI9ezR+s21AvUqWRfEgJFATq8+qdbzcXc
1XMEz6Wf9Ug1z4jL4HsZmO7EkuWY2OfQ/UHMTc9Zzk6raUOvXPKRGtazt5zp03wh
bmQxP6KtuYtDD1c2VXCm/s0BHdbzsnFockaxpy08xfPNmeD/vVKW3evS2GYIoZcr
x1mgxrZWxDulmUdBr4MPZ5Z9Xcnit4opjSVwywTHBA/G1pqfh2PnlUsB4icRkHEj
DXL2Qyg0YROQ5C11+LRRlYeGF9vDCYMJm2bKCVHavLAcnL9xzchBpsJYKYff0Wxp
u3qOSvjPx6QVg48tPvmM8a1BJJuwEahCnM6Z7tv/Uvn32lOIGQ+0QVMI2SNqYI8S
0q0JrIbEC+O9jGZygx2IaYkMDLaaBrEw53QD0kOzGqKTqeEQyIyyDHXIlV7DCOV4
i/BGDJqCCo99mJGHWExVsCVFpqGCCpq0L+CZIMssrkmej0SzHuIVzXR1az1jBGL1
tbW0Xe1RgSS2FCouctnYXM0/lQQ8/5mfo6yZnkfISwKokNBVmmkKVyJpuDZYq/Wo
ZWn2WkJaaIF6bJZ2eXa5nGmBKFeymrp+1uURF7kMhEuby6brb5HzgRpbIzgpBe3/
NawaVFY/Hpfg5wOT6/MEURX4smA3KlOI9A6aa+x840fZzpqim9x6XGLvA0u58Ytl
rjoKHZkjRpUXy1BRzhAWBuZczdl141n9OCBPtbDaSgbVsKvFAsMprdSeFs1EOUjM
rCUCEISmcoyGBg/dRUpcYZqVqCQRG50Ttm/6dZ5fkCmgLI1xxH8jxU5+pwHhwVEd
oK3TKaL/Rih8TwD2vRpmyLd/hU/mNpHpU17eVW1qeudeI44MuK28V4/Aob8k7NjD
PLcg6kGL6l0m0GInYb6Lquz30JLbeR8AEEoSaGADSON0X2qYciPS/re+ZJDjGEr3
3p8jvyVcFGU4ETbA7cSAqLTR9C2In69cs9BHXVUnk5FPosO6BD0GpFUtzwjjf4NU
HE0AMZXdGekLiPkHFOWblb+jTeJhgXQVT/mI3QSjZFrF5BFcQuDDoiZLqB8qeMMS
CfV70hGZoSczV41ZLR67RWdnmUrsp2NnCTzWlMh9lWSSxNKJHXIjRqH07SNDHhIO
s/ltCJELbiAqNZuGkPCnvZ64ibuDQyO/DSZjAN0KWSJ9FJASfU77uaur+WRvf9qf
iydbDoQOtWl9X2aAeAiM4oXdu3gpJMd9DOX7bUnh5eKXxtyK/hylliF33KN/7bpU
gPiHwpa3StfxZy2buAMNuae3ZtfsasJU8HoIh21zFpKEy2xT1VI5M+Tvz2qO31tC
InQNMGsagMf9pq+KSuebAxWZaDbrxLk/mr4Fgf1pmErKqjMjU0vHdavt1C8WoOhR
fK5S+F4F2ZRO6Jnxrh7PCX3Pi6+FPSY1JYpMm92xsN+jbhlZhm+1XQdpY1Sz1IeI
AjFEAb1Ku85oqK23g72Wbrr8ViRHkCvPw9Rukz9n3YxHsA9n+dX1DjdbP2nZ2ikw
ZEyP/0usywKGYwn+HPVfWH9BfHRs3FXvJeYFJhDy6pCXSNyZTaWDciMAEI99BjoG
kh4cy3CLeq/hmgXRoGJGEGCQpZ2axWk7DHBeqFkszKn/Ao0rtEHPe1XIDgzyQ4Be
KDYkdWM6xzd2Wfed1la86jtjOd8BXADh06vXv9sm5TvGsWPcfbSt9DypmZNXbSFa
gvVuxydZfPy3FkcrP4oGZePJIfNG9tYBwc4E3g66UDDju/ynRpXkyWcU1VoNnDTs
lGwOazey5c9fzI6JsEQ6ZsI/FHZJRuwxJ/RF3kbA8gHnTPl5yRVjDoGZ1fEObouX
TqZaCCAi6w8fsv8I5N5aTejUK1DzbgNahh+hIvo6OnV17zrTaPzvrh+fTL5SfDjg
Px/aF8hF2fzNMRSzCzoyL6FoqSFfXhFeB4f9gnntqSRZwp1S7AAU01oAuzxr+v5v
fZzszd2IiGK186kU4jTOa12RFDZYAgESwMym9nXk3rYN8DlmTDJRzump3OgOiObS
0jVYVER5ai2InpHLbmrS+a41O/iEQLrI/SJIU8TBi8fG7DGXdEIAl7+BgYfcF5BQ
c4P3OEp8JADZVm4hgUUiwpgEHBBTWL4/C9CG28pTOtSIbWm5JFWILPxZ70p2yrlD
Xl2aiZhlS/00iqVXXgpKE/kxhAaiBPr8bnkMygSW4XP4a/4m35vv6n5Vt8gqBfgO
xWMctQujMQDZajZNRBolRXj4hI9qUnj4uJXaM8c35NInYha+Q52gCSFdZm2R4V7F
pJZtg9BWAKg7a8Wxt0zz01vORboahO100u8TYu4JBx6AFQ0mg21CU26kVNA5jRbD
mU31HktEOAO+8IKnVoHS5VYIcLeZzTnDe7fD8luiyLsrGZSs8Wc+x5m0QZrQXEAT
Ys/+GTADq+MqickR8lqQKad55+lTCItwD9Fa8hnOGRBFab8mHnVQxBnEHYue6FD9
gOEnj21TmlzQd5XDkCWEVb5mHxXg+f9u5GdP1zaCpWy2gK/UQGK2ULnxE95yCH17
B6n9Bo15GMFf4e7/vmG/8KEFpL498u4Qq/+4owY10B3hHMCKhQ8FL2mQJN8GyDoj
eKcL5+P/STgdPOolIlt+8MBTNswQCimc950BFz0LXoZqQMHs0ZViQY8tlG0CMaUz
ywxRFlNkohzJuKBCh34RFqXVNHcILFbmJsgzbwF5rUXim5hW1Y1xPCZzi0Sy2Rwy
umWjGFLcRYbR5gbv9/lCEMUfaIWvN2Vq8VVVu3+jz0+L1TztiezbOu0SeOM0MrU4
ApljxfCQpfFigtcLKC8pEbxGib7r++/qNtEYbhG6oNw0sAfHMTw2/8A3uLbLSTHw
PG9nmJIjTVat1PuW0VWuxJ6jMx2vTa7XUgjah1f3CpxYrpXoWBdPTDQ1nwoqmsp+
prS+WMnO6GLvWT5ZcfIN5ilHRVkEG4uqm/S1NwLAABzxaHq6SRAKun4W7cMAtWcX
SNPiSYDJKLUJj/LGs7YlbpjJ0HZeoN+Bq1wRixhJpPHjrKmyRgKkGDC3BzLMuTat
ZRLkjO8TFCqkBBbbJUs5yUSJ1/XA6wBDgnrvbSDf12+Jy/1o7V3655mXaIiflFnB
G0sHcoai+GCMYVkmITRB4eYhzHKDbffmlKcyp/m7dl1xtGYYWARmN3Snn2cMUHtl
/6ahbVywnX4wlJRatihTLucshxFIlSRoowCjK7LsN0fwbe2OfqOxbFUVj1QjdBu2
8hRqCI6ABZsFpp1GkUmeodbINEjzK9b9GXFWfmwl4u5BIk76Ik9WMTXlYWD6iK9L
6N0h5IRY1Vbg8EygOMS9LWzO4NqNqTw7eyduyckF6e4ekVC1KODub5SWEih2P7ov
WoGxCkkwuYzZstE7oockhzYqXXqRe6PzVBFrWykYOWcLTqWvSjXc7ugZytTj7JQY
9Cvw0QOjfV7b7dDm3rPmL6MsnBDu7IHDyU61Kg038Sx8t1Mjzr0nwvj4IibaL0e1
jHhBCnrFoEetT4LQ5CIndtGZlbU0Q49ESlVzmjTCQYT0ZPAf1wsOZtCVMCrnCZVA
OWvg3BwZvJza2e5IcUcf7y0iUhaozeo9kqC0Q2vs+YZYFg31+TVLX5Tb074gQAN1
qHDNW+UnocB+GWZAtSjraK23Hw/theZeqMIbwpnZDIT+EoA8md5V0rqkR8nu43jP
rdyEq5ROJWJXRz7Mafe6/eBNlH8fXV/Reulowapk7AhonfoRFODjnC8H7Wc5qLt3
wc+Lc9CDdwY9pb5OtZnHnnRJ4V/NL+/WQB+Gt+YJEkhFI88xYEI+78pb4L+TUXvG
hbvfq+ZSAdlVMMEA6LLK2dnIQYiXj/HttcjR/ESL2b/BWuqlhdmpKC+RH5mNV98/
i3rwtSLaINo5u8pvYYi4rlbaQu834XN4Fm0+Wg+JKWoDS/39zOFee3T7DG73HkDt
F4q/xpF18J1gbZOfuqPW3UrOlOUX3KinycFWtjEMYSn/mQNzD0HwZmNksF/Bd8a8
BOo1+6TSsKwjdz2+v/5QnPUMhn7qRDJFB1Z4xneP1BW8C7lFuGPHfNVsbZ+2qO0N
39fVqQ2qLD9/FT3X7NCn7cUIfnjiRLDizZHwNS6lGrg7dlOIGjsdSVM2Pux5ZUeV
W1CSEOvWe7isunmodWWsCAYdBFLulTkZE5O5FILjCqvaAQT9FzJV650CGrc/pD44
bZ/A6RtIsjiEGE5Rd1AP0bdOvZyjnl2XApnOV+Go+Q82r/o05T8tiR7D/nAE3y6p
L4efbaW5xE1CtE0bbhz7x4o5uEZzTjN4lOnkLmfx55UvEsBM8lg7R638XqzAk+ix
MR8ST8sAZVb5P/nXnXZBL39fbX76lWdsP0LAGzrsmxpypKL8BjIXHPDARhjDTTA7
sixp8dtlbaUZcdNV96U7AvmK+0Vr9iw/6bNFCQZJ+AVE9wrGz4eNgAJqBL5LIGgj
9FGM3urXoMY0TXSGZCzLxXnsWC/TIGzEwFRvKNIsm/CbX1bNE15VQbz5xmHuXLc0
XXzUS5+Apg2YXmL3SFsLvmSyNR6N10KAn93prKfwzRu2rEWyFlNq0knzJ9ch3QGE
cqvgN5xn9a7zBpLL0HT8+x+PqnsTgQjNtHaQgqJLXzt7eawfS2qGJCoB+SYraoX4
ZYSVI4FM539uWmxOaJ6GeNNVPK86inQE+UZRxfoY7WX7bmgPyef5exbaA6klHjtc
/t61g0tCp7XHEAljfAGvON1Qr+2lWZngynLjgO92ii+or5m2ehICA7Ilmym/6vTm
RUyWQZbq0vuo0nRvLCsvlhOFaQs7/9MRVErH6/HvDx9Sy+nYu0KHFV2kyPTPoKAU
cni8R+gwSr6K/g8ScEcOUPLmTwo8GYoHugY5kimFdFdistCNGj+cXIKNOHOUx7F6
FAfMZcCQCgwu3k5mEMTKrrHLuJTymHTpkCjcBH2JJRyBIRzxBsAm5uMy09RtDt+7
biCIjWKRL29b5CAWIezJDzz5OXF/VOscwTyFjIq2hJQjRG2n61TJcDdx+Wdvn6FT
ePGOF8DfTe4tdRhpgwj80wvlxsolH/u+x6uWS9duSCzqgLzDrGLQdbIKUHIQZACT
5HILonAE6QVdUM9YSKpeR2DVY8/lULgbeZTM+4ujiYY1wnP4anz9X4n0YXEeJWr1
chCincdHuGx9S4TyNFu1OGUeTOXFGK6fmYoY0wsMrABckIcN8ILIEzHHEPVvT60T
suMMvGn/J2jBWVYSXDA7mElJxFqoHoT2klRMr3qbjjKjy+muyWD81/hMkj3s7M+R
RjC0ETSDSPwTmpK8l973NHcKzM91UNs8HmDOKsc+vHdBtLyWfQtFLSw7P9/Ej/YD
25T+qUIE/9LF4j6/3OtHU5Wws3ajiCpjJjakBWxEV8d1BKagdM+SQCOoaezcPtV3
Ub3ygVQ9mgbgGjV/f2egI3/Ozc/FmxHXM9LCcB97pXVoJ8Tz7HGnTMhBcappCvnx
0VeBPWxOXP6zAcc/f9dC0iIxLrENHfq7+nhAovsIsp3vUsHFMCEDNDIqt7OimX59
+CV0hzv8zAhfXOqsstZ4ZhuQFS03y1FGAG72gmsyLJpCnnmK4lJSDrO0wxVvNcv1
Kd/nwVCP7I3Ad1sDL1dcvxXH1S8DXWxW3xkEb/KAdZPS6Iq4QzULsCVgZZSnbPJU
svUUDy8XumMsx98g85Rulha6+pOH1rHpEUmgWkDecuB6EZ2HY/gbHcq+oJ/BtPBA
VPXE8VHg6P3Wcpc/W8yHu1DqVIWsVPMn/wCq+uOa89tqOyW61e3Kdxt1B0QEMXOR
ZE3uzs25c/QmcNv4fECqgehHWP4kbml43/CU4dMLT5Icm0r9uHejY+abTiVFG1AW
JEulxtYaac1PqwzN4ge/wS/o/iYS4T8ojB0EI5wKrcG9QU0hFznizoWs7LrTieJw
c6gTaTWBRMB7jQMoIIepuNShS3cCEn7OczMVB2Vk6A9q6eB6U1j4OtFxQgxPH0j6
GltV8tVEtFUrAMhfr5Fticd6X5hwR0YlENbNKfNqmxgETU8EiRPm/aVirwyJb4B6
ljHsjbc+IPHvAfb6MuMH0+5ad34Vw77CZHxT5asbii4CO5Y1/TWLmkRfBkbp+cM9
KbWAYTrplwQJZLchm86BXOvHywGqjhlxkpVozLCS462U4wnQ63KFuwbJ+I0sdt7/
PRsRpKC5l7sDntNfrh8Td71OYDUUo2ZYmkzGT4zcZGmrXQgccsaXblLoTBN5zreF
w3MG2ytDKc1OKh0W42v6peNzZmc2Le6r7BVM3TbmXwYyKAUmb6Bs8SNN0JEXs3OS
eTUSBSPd+EXE55Ya2uYS4AGB/9j7nFDSs9GNZQYUOdQNN0PXCOaTAgw/UPczh+YA
CRdSK9ps3NOa+ZRa6Neba4Nyut6DzO12+ILFjy9+MYynLg4uI6MOQoUKjFjyr3Ag
qrrGcRKKFO/6zHK0f6DN3UQAiqlnbHO+6jv0QUfPBKlf1DdDl6B3VD/dqrSOzKwt
SAs/ziqN5FQCPO0Cv00h0EKn5eRfxq+Cvt2JJD2EIC594S4j/c8iCmvfwFmEx9CO
8SygnO0RKQNnSTuE5e8w1apWHJMpzKmodPbt6J2u+PmYCoY/6LdX+Bx8r2Gr/aZj
4H/Z2JfoKcbx8duIwCzb0NB05GoLrLMGqVNAnP7XuSbPlJT1I0agF9DynFvzI6Zy
YUJCGst3nn7f50Qg+Dvj067VBrSjb6uQJ0cB9+cts0uBQShYhH6CB0Z1VU5OA+Ni
Hrd4+G0QeNPYbpCZvTyRV2ooPcMGDDqPS05ZUGRIBqiTGZbN8J7W3h+0/hRiebjO
y3kV2GE+Q4GFh5CN2/WPNwoxR20q3LCjth7WyCzEBZJNYZ5WpLKfmVhdv46FQXxC
4up4n+1R5af53uhgoNttwrWXo9Yah8KPJWAJT5/ZewOKhCcHxArcGjZFFFaiE/Ct
wXsmQvY+UO8tmfoSa1SfG2PSqk5B76+T0w40x0+hguY7UaM6IKmkbBrAsb6AZhhX
bYNHFH6O8P0+DdUDGc5Kta8rmJKOg82o+rDSiq2i1c9XUeaIMH9gJDwe5AYxozdJ
WE0fx9Kf4QU/z5bEPWgiOLEt1+YUmwu7WL/SUjNMfgFrrk55fYtC6FqIS8Vcc0OZ
mAl46FEP/BXLSM/OGhBi4upFcn2LpR8rXiR819rEe25BUGJhbqh+vT0dP5Cp4U5s
XUFYfqFDk7vd4tv69ue17p3TPxX5JIf7Zdkq914aRdjp4bBrw/pwAVb8/vky70yL
snLAF+R2lBqoo45Hv6ZugOLD9WT/Q52cYgKPSRBeMMTmKupgIYpEFaluM/OoGvSq
kZM3i1kMEj/DHjZWDn8GxUMUJIRPYYktsXKSEblbR4et4N9GeCNJH0XWFltgbz6G
e8mQwIq67OfD6XueFT1KSrHVWZKYPiYka09dBuXx4/aA9QBHeQ2KcrtZDjxtc+zn
eV9P2jWvYpzQ3P+PHpPL7neZ6DB0qld6aPXg+rdabVp3aomx5dE0fH5r9KZEJQuY
tK6ROMYSvElpXbbvxb9t74f2y8WNH5yPFUpPCTzhIST5y4v7CMZ2nOlRWL4TC5E2
wEhS7ahAmHSYStcXsUcW6+uEwVs9W96xjCHgthulHhWOY/fmj/wySh9ynPnih/Iv
dLjSJalYXodd8Sspd9rkb3ftsV7H68UrR3iqJwC5sLJa7rU+PiIQ20uYSGalsGFG
t0pMo/CqQusXTrALer0nwfLMlxVdvJ5wZ99AAeg6jOXzHmISOzFKhMZmVqZdJRXk
UWxF97KPqz1p1c4MQNjXuFqbkQDjTRcVldNE9WPU5+oKin5NHyOo70kbJPboK36E
+ku4dwBs5nSGP8ntESpztJnp+kQpE6FAxZBeivv0ZfM4hEfRYYkZrpFtWfRVVae4
hMGSxXmff0JGcfO4FjLyqpIxxZ9FnlYdUc2A82FOpdXPEd9GT6YqOdViuGqlnI3u
zVGMmj1hQb+PFHRjOHSpwD/XsAKx/V+9imMqVAgZwaVK5IGQrHqRgcTKkR2Sp00c
0XmyqDn63FXltAfd6oxXN2CbAAaxBftk89PQsAXFjDOOAaaEYW1n/T1nqKWewDbA
sSbPP1Rg24l5EAyEjv/K4Pqpdytwzb2J8z3ufNql+CQ59MHfcp5YTZKBW67Qr0gf
kEA8fYIvaSsAZtgr7h+BE1MCQ/OCmcPdIB+i5opNw/PdgReNoWrFsCsiYB0ZUaW0
i73b55o0HrPO9VJDUy3BOj4N1lOlNHoyYPbL23FYEIAVnXYHsWsSS88Aafftmjbt
LVDDrKmSNSi8DJJGwfTeaWDUBCX81CjuuYS1DSXD/vXFLF6KcGRiJkRDD6ksw8k8
Gafzl2rvkWyZQ0xPq92vY1QrH6Mjw1vt8EuNnElnejQeU6zacf6nJJBfWvXnSeqh
tKgI/yxyTMUHDBQkT2b4860S2vD8v+N/4PjFFOyguT6f81uVhK54DPJJ5ODu0Ams
9zLxPwf866EeOT0DqfFdYVWM9rvW2tQ5TtJIusjy/5+ztxO5SzVx05IbXPhA3jeR
C5MoW8ylKDtb9c6msur/xSmvD61kdL4cuq9boz1nDtDPWD0kwtxTfqrgRnfKEBvN
EuBrm8eoPMsZopKlQqeqJkpff4YLwwIDN0V9Zua11Ay9yIQNRI1hJU8g1HirUxdk
8DMrD+Yazt+ogw5iUsFVg9niAAiG9ypg4E1BAGmVVlMyM32/O3X5Y4KV3Fg1GqLL
2nF14iYfn9U2/20J6vKZ2OVRY3d8F+LcLgMSB+qFxdncsOcoRAtiZ9JPLhlLFJAj
jIvrr6GGiS5DqmQzsNPryGFloNldpQP8p+COgVQFlr2drUeIyrZJvgYbLv72FA1E
wyWvOmX89F5SuLZ6FM7p815v7c5JvxoH2B+9i5SmOq050p9czPRTbJxzg/3cK49N
mns2N5fZ5q2csjpNizV+21nzGJZS6kE44lL16bIUMiEbJRqE2XcFSc9vfATzeMYd
inQmS/44VibxhF0vXz5b56NZk1GoIpdKPC9EkLq2hi6/DXCRI41j+F96Z9z8znEu
kUYfYGR5lOVSvXnsB1FEh2ZPCTeUL3Q5k/612Jt3wA4xHE2y7JN0PhUU4xwVshms
hxKp63wa1q3h5qj4n/THXty5Ogqbqq1Nh0PzygmZa8Ekvqg2Wj+hiQ/+RorM56pI
tv+UxuA8xkv8OSE4tE/R9G2FaoSKwYeYesXMDfqszRtWDGEQwnbp3iyxMVhetoMR
bqaKJjcC3AnDnfyJBdMWygh3y5g3PWLZI94tvJXL9o+9aIuoSD5KipOmG7Z7ALYa
FvyDURsAWAR+ehRySnWZw+2FdgXJtk+EGpXgUqZ1w/gRAr6F8Im4dKRrwi4fYZhu
fbBC9OiWjtrkQfG8clP1s+MxnyjBcZifew2hT8TQPMVaO3zQppJQO8vCJJvRXUWe
6wqFIFP7x+F6mKT+WRj/UJI36VTKaBCWQxV7haydEwlsnXNkiLtf2z+AmGn80Etf
PMcGGhtQbjvlf40ic9rCuE6M83zbdNJ9YgKmIaUDglm6mfQYHbtnLvN8ci1WLzVY
/KZ9hl9/QB81pbslxGN9kb1Smeu/X26sQ/0Zw2yb7g+SujWWh9u7V8BB1G8JOIkx
QWF9Dv8ab2TTG+vb/pG8avGBYFbaMH7iLXoTZmK2Rcvzy5F2XYG+d4AxGGK6x95L
507EyxzGGoQWwPgeltnsuaCZ+c07vlbLZNmgD5Q3MmxuVqsALWQF3pyx0z1xqAgw
KU/ewtmxUb2AF8jln2hSTZ1cVKJoVC9orioscmu3f1kol3DMjv+VvMR5cGyyD0q3
Tu2DIpr5yb/TO6NSQHyp+C5KCHzPhB9cB1gYfSgJaDp9al5kaPRsp/Fq2uknxIOp
PeaYV8DURQIyCaEJIAiJOGL49NEf5mKbX8H5HaHmdCv/L5RPQe8shClZBDJkMKEp
lmVfP0jG36rtbqkrV9TgaiIiyIY6N/47ikHBfFkLX42QBcuRPdAOaeFlgJQo9RQ3
jZF1Cs7uvsML9fKSc8eNUY7V+xU66oXDCif+ALJOZQuyjF5jTqMk/cxH8ihbtIgO
E+wMrV6WKueTiUlyuOqgKLuT1ySARfWecfXHdUzhfZzKYSrO01I10ozoqH9NRC9i
wYH7y6jeR2AEIjcTRsnpIwruCuu5gXbNxn7N+UWwVWFGVJLe3rOcU2IKwGzUu7/H
E//q7RqFn+I1obIe9KphsauX0WfhVC8J/VUabAYza9SIBOpm3vxonrp6JSN3FDlC
HJqAiglnM1wUcehTItFU4InBq6AM85OeS7mtXnsGZ8yYNgSAmsyUgG8+H8bHIK5+
j+XbViVKrDBdvcBisHlKKeiEwcFoIbRWK3sGEe9ZFT0gt7tINjKKkQ7CrW/e96Lq
LU9Ml/MIuSo5aNcfkGuyI28WuxhGYoc/ywBbwd2EysJzpFkLwBp1a1JK3M3bVmpK
P5FfZ5h6OMlset3UcKmj9Zeh1ejRjXt70PVwtKTqB4ahu30r7s7G6/mAJfnTQ5iQ
F2gsSkBJxDZ9eRy8qhP3q3V8CSY/vCUz0/VdV8xkj2GUxAG5w8UaZ+bm8i1U4ZIb
rMFe/N8n0eJnMlq3G4X3vFynPwU8s4xd1juX/OpGdNkwtKlOUqNvcUBgWRzcdlTZ
MVsZVL/PKQqZKZTYFH76gIQh1s12FRsCPwg8VTkMh0gIwqThJ95Z36lnDcrTXlir
yq3oF3VEmmd5ZUee9RL2/U85FVvcoHMwJ/gt8LGyNFJJjqCicQHJmxvJh3+0MgDC
3yFCGyheozJC0n8IX2UEW4eCxDWxdPqXMZhwQwY0XgjwdMDCz2EqWwzB7nrn916c
AUvwwkFdTUY7AbcRj2frqR87dUjM5EqUhHB9mJDDQP58YXPuo5gbSnYVXDZc5Nit
C5ColXoUcnQsEQvpKZ+rnS+lWusnuBoYQc+2yDAh9+0KVuGVK0HcPsnDPEArm6Ho
c8WpJ8MyJXUO3Zj9So79WjYHs4bFdHIxB3d8JEpfCJ+viMmvHEfGgjEQsBuqdxkr
GFBatwTUrdhWRnWCyJTNPeio8PJb9cQq1wBE6zzNRKeu8XKycm+0rCsSmgx68U6w
RES++7VYgenBXZGU99NG1bId8oF+SEW3N/TLCXMz4oO8y0Rtn5/y2jAIR2HRLoh5
rhlaSKQWp7gHOwxMHS79NA5XOGwEMLD5PA5dfY0O9bN0R/B/kzDTaz5aN44hCPdX
usp93WINZAMI3GNP4GKhgFjB3Ql3VBfxSveiJUZ9cL3+kJjcitYeDibIwR3GNFAr
DWt3LQ6h9bN+kv4YpdXX8s/VYDTkwbJuKZ8EGu/qiJJfy/sjzzoN5cgAL7oUY2oN
gHWIpVPpaHXV4La9uldNnZHl7TUhFttlbEauwrHGxxJTDfdi51QGFfQ2/VPr033K
Nssdrkls4+vSWvPSAzDs6bC67nCz8/yRu+NqU/nSkO9RIMXT/awlns9MSu8bA8gw
yK2fzAMni8Hjwr7ZbHI/RZYDBI6aH5BKA18JehF7mkEDA7MhRYdJrgWfJ6OOWLgg
qaj8Tb0tCrsUPg/u/ndT7Za04CwQJtiK8gQO3+4q2d6I+3VVzF3GDuq9/DHubjtG
GPqTbEt6xHbBzmVtOJ3O6w+HzieBd+x40f0YBYkQ7Ho9Urc6Xl8v2sHYj8cRnVOg
nHX6flZH4o9ODToXSA9brx1WAmMEhtXDV9RXVUrlLIPRxfRZGmdvQu69MYeVCmDy
maCKvLxod4i3Jq4Ewx4yq8eVcJWseTJPDeYxSVrwsj8huE/WcFaploDY1FciEmz0
lMy8s7g6l2caH6Iwt6AdnIvtfSW5AL0e/Ky5JDnFJirC+gD9tuSk5vUBRD8ahb91
IijYFGeqBxR585d5V8zMT+rm4Xfittcis7bDfSDUhKNASyWiyFHHJP52LNQ/P5+v
slNma9JRkmZ8SbFSeoatHhOWk6OfHYntX6xGjBLEDkgtGOBFJcH1flOW0VXul7Bk
qpMfVjVdSMGq0NBwr7dLY9bulJCiPLa5r/UHrJa79xfMJ8K4z+2HLSjoZ7KmfmZX
eQQ85/cVYIHO18iY6X6rqbCG1VNZuFiDTZWceXuDFpdYWRmQIY4jxw4EATZuImd5
hwZI+pnUwPL/AIkJRIjsOMBgOevQQPYQ+QXo1QkYHecHitZywh/1OZuENAguNmtb
yWmrGFgcYdc42MMVOhcBme5U1RxCPPcGgMiXc62MJl5cN8tQOBeGdGppJzYZfzDa
M8MiDlQjXKgXL0Gj19gcj4sVrKQf4GPZiFJbmjzn5xpxxWP2cUu40SfDLNsS0YCU
ETat7LZdx3rb/5XJa/NSDaA7Kz2hk+InH3yotc6nNcx500T6kU0p9eT6nHuMbunn
ik3vRPHvm9JsjSa5Z78FkyjIXcGbYou2FoGxmUQJT5/xvkO9BWuyBU7YdFCsSZqk
J7lEKVRqjKcweINhZFR1PJE9OjQcCqOQNv6Y/vMmCzZCYbRFE+vDI/lhZfi/fPaR
95nCKfiOIJL4GaGNujTIu9JGWj811xZHFuSJPhyaDVaZ2P66fvkfjq4+uIePTsyY
iv2LIfqA7sIjb4Hk2qEOMqW66CyKJ8tKJmc4p1jn/VmhWKsZFzZAC/LfyoeIIYaA
T+Kj+orB7ADvb44hMS3kei6N/vPFUOmZRBC6b/fn8ox+fTCFX+iRAf5DM4Gr72ob
0OSvy4Di09SAbw9/AwMPMT0tGnZyuv25H4muql3t7FFpYikUSi5m2hTGqc9EHLSr
cdGaqbYelLXNz6AUulNjitBGbzs9qNbSuFVpydZyx3DYYnywu/9IcQ2ITKHXMNc0
BrR1df6ueuKeWb/TSlJAXRcMoHm5XpVgLchbefsCLbwgp+Y6k0MpJNTjVk4ruACJ
eVBzRenp1tDKFeKCSRZWe8LoruWfPXjPgsvcfDLuD3Z5vlbyjMLU3jl4Iqsitzfx
ZfvjOHK2qFsVHvqFxv1OrY/3tT+dWf2ye4H88TXEI6WZ8YvfYOR7M/VQHyk57VG3
2XIC9KZHbLEwjOlHhVFSzpuJOGbQfNP8hPMdwXmmedSa3GK5lzKxw9RHlsF/dIcK
pRowhH+fGHhS1XpEJabeOraTBcUEGtznzBqgz+ZHIp9ndqOu9DgXfzwfdmcXohV6
lkQnv3TvyeMqtJG6CTafh0+WOpDc5x7bQ/9sWDVTSOrP5KwQac1NfOESx706l1Gy
+89X7scrfHF7bLa9RsHwO2Wo0GqimISS6qaIhK9idy3HkEfW42aPwmhEJKxfwMof
8pIkv+/tTybppn/2RYKL1c+T71twAOPj6GbqbREYyt89RdyNgc92CfuqxqBVPCMd
WsLhocqaiklWwvei1/PG9arp2SHa3hf1vcYhZwF+g+AlTLHR/hsh3MU3PDTST1r3
UipRAoFA3KL7vTc7GVzlnd8j2lxzGArAMk5RnFay47T/j7NnHQUw9gDp3X1wANii
ahye6VVKEVm92SIH0U+KbPEQqi/PGkMsxUpJdcWiG/qhnUM7DPPKMOR/lvNEyd9T
PPzo19Lk4KEpb1yAXWGcaLwE7iiOijsg1vRN1qwhb7qAm3dSMzbIbWMvFXI3053I
m1ZEiaADFwCyQFUxRhRGQP8HFRCYpO7MYxRq3I5Nzr03WIRAK7QfwOhz8+rqU4Fw
EzRxTL+MfKLlS+ZH842TdVof1mEzyMfQgeJKg0V4cdcm9UzbFMoAGzKMRRdqZ8Yw
JWszVBEQaa0zrhODB6pjQzTXUJdOTgNMqT0QQ5v0hxgOLiGvUXWbMBtxWTxxbjSW
6hN/6ymnwBK1MtWxpI+33TCgCjFJn59f/0tSZU6hsHpbaVXF+PD3vesGFVFODqOu
ayoFfRrYlV8PFhD03SRxu04hpgP9FpFwP2t6QebzqrrIZiiDs8geDcfPjD5m9o2k
mbJcEZHvA3gdzgIok/3JwwN0P5MPzrlsYMXkmPLn7cdJUjuyXWtUjBpPyPVVRzd+
nJoZ1Va38z5zfGxHJs6UINsTNRxle3agE0KTOkhX751+bWQl23L4kJr3sSYA7z/Q
D8ifmSRtlkp6cztdW46LRf0Vlbd1AafYFJhZ4ppZR6nZ1z4vt/S6KDgBLxWElbXO
z0Pq7shb/GqSJDzNgxRta9I8ETN9/NcHRdWuW65NuOdZNznYxkNbS6uv+kl4cMRW
YAvhwgaD5cj2MerKxP9Mg9W483h3sG7qIs7usaN77ygk3VOc2lydWoKpk6iRFK5R
C/JHSFNNR0aAXs55pEv5aRwtiMoawRWrOehWWt1XCm0lke94wqtaMsifWuR8RVyd
8xFpV1BFm2s7pHyvKKKNxQzBSVXDspNLYdrLAQ7dmP/bf12Avho7NGfyvRQw4eG+
6Q55js7h8dam2gXmIs2J0wjjjlEboq2usCepJaOxzGOQPu8E/ew9YykNjqSIBYeC
3zynxeKA6uhGOo7r81DHpl9kZ+4JgFwjOHCq3PSsNGBTAX/mqg7Z8aZdfsMQW7Vo
yAZZh6OKgU7h2j2sWwDIZ8okIBCKpR6Mbt0wvufFEEmnGf9K48oW+hTZl7tCKX9J
4C0lG8t3F+Ey4Zullx2WlVwOxfjkkDBLsFub/+7wNG9jesnum2lo4qXY3ekUg82M
worzs1VtoNrZfowIUNpkIhUlGvxPbm9/aGOBlZdPkTVEUPHtFgNiqcAqTmUrd7w4
pCN1zganW2xEYMFqcyE4PH/sqA3AKh4suSMpdAs5WWB5olXNxMvJV0F8e8lB5Vy4
jDrh/pyLs0G1Y9R7jjdJ8w+LCuYaA3kZ7WYiSbUXGQ6xRDtBk/zprtfdX1th7L5+
zSIi0DTKl3A5hIkSKMkGtZuc21UDjBYO72WcE/0QzHw7UkA/hWVXxMmg4IthZ92Q
05x+MS39w8zaH8yvIeHphf0E/b4zMC8Cn7d49AmvH0TooMjUxEzu5Sf/zTViAxfw
nSUBy07GN3deSStK7xdoQT1hYKnWnQRRFgPGAdG5Js4VJzi5GuTxZtNcUrdIqCTV
1T86nAd31Thy94Ron5DQiRlZ9M8lUuuIZi4xIx9CowXaz4CFGXjZ/z+/LN7ec2J/
TkraqHGYfdc6bkgCuOG+pjJo1Sp91D4bXLhcr5pyKUk+Dmlzwu+JGBSptNrDJcy7
RP5VotNpzjx5xA0MrJ2PlGJJ7UJvgL52miN2cwG8Tdn4s/S9tWX090ReGGA9Hz11
O2LFQoiBOZP4yCn4+9Ouektq6Efb4V551GuRlWLordVLldkmhF2xF0Yj1edY/Kqm
JREb6FuVmBKPqYmWbGbuI7utP142vdfGI6l/vlJ8dFwAA77vtXvIy1J1GdP9YVsk
wLEL8OA7L2haRdqdUEmyw2cTh3r8TkT4RQnKsFfUaTVZTk8F7E5OHLtMVokLWv4/
winhWVFOsWLIL2EPjHiZnNAtz/MUhrwrXozBdtZKKyV8cRxKrvDBeC72utfOV0IK
Py0E25GwRRpMnOKz5+t6C+I8CDhhyID7cMgp+0/YiKcCanuqLbxT5N5xgO32E34A
R1qcQRvuZ1Wxpt+KAYuuq9oB5q2UclVGdh7lrY3K2o+GJpPqeMd/hDakcHIqE3ca
BKExvch80vgGcJqToepOA24Rsebg2wDdLepyrDvshJf8ZqoJO6DfmGo8glCgbJYR
yLIBoSDCDVgo0sqDGw/8fSWL32f5Ef/04kwgV1zKZC1Yg/2obDALwCag+weKqaGq
/j+4S0/sUDX8BwgKL7u9t46lqZo2QyHGVf6eOshzcx1UYvknQW8FhdjMTlnnlVAV
EMZsWQNwsEqlGHshalOB4Qd4UftU1/7xTnucGHbW6G+AaczE9tf8GntInvnl2l4h
P8IJOHmyAzzx2Lu3nRrh2kBPoilBZj8Ibgj1PrcMWbudt1OU3MtWCk8IbNzS7mgo
WxaFFJAZQ/4eqdvBwE+Ze7TXb3JqntbxRnz8rMAGIvvprOlM6A8FoBe+apGvBO3a
+taVJoXlKdhIhBnkoqe232VYurQC4aPjKsd38/sZ+K8O3rgmPO1TloxPqa58eUYT
xjbKKOsSAyghFDOUBx7Hq0/IPBjf/ypCcI9KkDSx8jNHBdx1XnAjZFs19hDtJ/kB
GaRQp9SC/2Rm6ZQB0tHrsjJR9BRSRcVWoAkBSVKzXY3naL8aCAgl72lLRN09g0E4
a3hyZblj8SPXlrpi56Bz3mDqSVe7RGux8dwK9JoddsCtQMUE9bvy6jGplOreCfjW
bfKnUs84p8GW8jWcINnQamoABDrsxoCDBna8KC43Elpc88TK29JAZtkew/YQcdCD
Df9E01O8EssqFBp33WeYCvquaN748xerZagxzTcSm7v1fLIA4pb6iCt/9OJtaexu
azo+pRx8yvYeqBvoHU2fIecVKO6iDh3JbCzzd/h2xFnZm7yGw1cfqdBLqzNCYIog
msmnJ4YPCZAKnnW/YWuFYnmdU/53nXbbMB2yEeblms1NZFhgyTgm5UonwvUuISy8
ygo1lWF9reVAo4G9hCvBXJwfg7TZhfhenAWXfbYMBCq0QRsprnPyqg54Uba/eR4S
j+zUbF3leJPkPvy1goP/jsQWjvDsxeIHz271gBsHWwVykNA0uJ1+Q2nXu4pPbWsi
6yIcXyWv3m0mTFoJOkjRKvmoJFHldY6Sqp6JHHNMloIc1Lm4CMI75dSoetZiVqqX
3rqcNQYKCjb6T14B9WXMkv+M692ednB5w29aXNnfckO1psh5/26vpFrULgUhXS8g
gx3k0CcbBsINFpM6JIbxo1rO6/KfWFgE19ZxNZPB5MdM9lPtc02k0fPHy/ViZMmJ
0F0lhAbu0+sPCQKf9sLSfmR445/eg0UBiakDfnfb+Annjxb4xacHFTL2OaBRbS89
C5wGjyz+hxbUXdm8Ttmnvs3XobZkzt8IT7Z2BXjmDlbyk0lGDYbFg3e3RmzD2Gik
0VKO2Jlkh+jb00nuCBoIsUKSBzSRAnW/fKbiY9ne94o3iq4aPie2qSXrgEokvLcn
UndZ481LFMWJ2NfWfQYf5QNvy23LU4oUP2uacfCHMtDsZjhJV2/PBkI3xVlfrOo3
XZVLdc7GW17UitEk3hxTvUAOzdH0wlK9Bs6dAeRRKqgFdTiTqJWGkEMACM5zG1qD
dozTxdG/HeC3JzuMWVdqnpAYscskf4L92UiiZyLVREKKECpYmZ23jVTux/0jBeEU
0ONEkjYjrjnivonTwoGOeGWZJK5igKhsUrF21ntMr43dPDjCjqr+5jiBJiRftZLQ
baf0/W2vtscVKtodTm9QQghnPakXBaIZ7pacqtfgnuQF2wMiNCgYDA5tEWq4ee53
dKgFX8t/ot7vHOse4ssgLFi85digLm0Hs6r7OApMNDdjcH7ujLdKyOIZHYiwwYek
44XaOLuoU9FLQaEMHavGSngH9phOOddsOSSfQT1qY6FUKC6vl9C36Fx7dtsokodC
y3dzCl5P+iv9ree7zDFS0YrOOb8x9760CehSsjjpGehU9f4PbXhDSYGdly8kgYM8
OHttViIrTYZwMip7L32XZmQ9pr3O9IR9bmqcEVojLcDEGN391qgYSzrqMzJxyq7e
JyvBawurBn2hTytCSpzK8EnhEevSbF+Fo15JCxi5zJT/4tPziz95aS3Spt0L63jK
BrQRkkXP3+7YOlYQIZuSf3Cnas2qcB+sw1apTFSot+you41NDOD8MrmDDmaJkNs2
er8LZDI8ePr8OEd0Km4hSE/c/05RGXJ48mCsdOvpaC6iivdntZ5Szt90f+67hOwl
vNQADTV6sy00J/G19Y0ItMnUKXbBdthJ2MJJu78CJX10tUDt4PK4zU5BWVBDqV19
mQ0UqZDts9oVjD+hV6Xx01YT3EAdZYb+98n2rkATwcNQ1eo5j72OJxcnKlwvUD2b
eeJa6B/bLlAaryJwHWVHNok/v+QBm3RMK+3pw33SboeW3Rx2Z9aDoa8hrb4r+2ul
3yfZnqWu1z5ErEszqMGdBruBKi1CHu/fsXQ/F6biDka06QkDNwaskD1cO/DIcXlx
M6ue4zI8AAKXoLraNl32lrodGEW8f8mySvOj9lFRgYONNn7ehV1CzbaqS7fIGf0D
9yBNO9RR/kjFu37iiJwl0cyBDo3UJ/FNYy4Tk0ORghONDIIlnIImuRCxW/qxbNIj
qZmX80Gs8oReieQBtlrNwvbi6nQribkrlCEYEOJvrORH1lKOYF+o6td6YMiV49mk
El7nEscC8rxMLdX6eO1fg+IntOW5eOWVMsN5BfG7OKL7VWTK4NVhjBURSXu66CjU
JQQFxZdkYPs5agL/W7Y6grMwA9owFUU1sScyHNaiNniJ6YAl/SNIuU7KTbuJz5cE
Fjk3jlgq8V/3uUNp5uZPyYKp8c/bU0//z7e/hNKcDTYzejtrv/MzjgdWCOxV/5l2
GhmSNCdc+5PFSS+ENkgZmbNPpI55GvNxEZC3H6Lp8DflH+sjHUDee3s5AkEE80fQ
jo5DPEjDeu36R/B23EyHClLMZOt8CyxFOJCPIgJRlxsEMpO38CEmlcX7UBSesl3s
w6UtGxHBQoah+voBHnHu/dFJAz9lTOuhoIdwLOzBDPNDrlMJLfDJriL8C+QO3umP
LO2zIgJ1z0qlsgLzaJHJ1iUB30Hsp4Npwh0YVrmwAx21oVutgkt5oNDDm5v62j6N
qILRoeos0o4QPlgOceuCStiiRHrrzU8aRa+K8HZmIFNKudy/B4wYGNfAelIoeYYX
Vk1HmFLQN5NgmM+XqsUx7EFg/w7BM0i708f5YM8rhpTjSOfrjjiYjXGWdZSWY93U
uL6lXIoiTIgDgoDinC+ZHJos4cPmUxj7pDdz8N7oWZt6MRBq5NqAqzgDEv8Iaf2C
uArjV4s6JnRy+Bfj+afm08sRUbi43UI8Z/nnniwuziH/QN/Vdo9wEWVNIMm6+XzZ
B3wAZeZJ02aC3Lm/XrB0Ol9pu+l8lSRMJFryaBkZ8GnGyC0v20eqV7+q5pl+0ux4
B0U142P64aPl8VcblGx+LHbPqdKzzjHvQU+f4bBQc4k9dIhK358Kis+nU2G7wZ7i
DWSKp+Xn50P486cWgLZVqK97aqAdTNKZ9XgD+oZCwEZylqZjwRig6V0pWnpOyH+D
Fv0fRZgWeFsiNlTzoZ65A6OXcXi4rnSYLWt8WfmAzp43rr1UJaKqU5PQSMGRL4D6
`protect end_protected