`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
ddtXksX2+yylW5zu6QL2Lhnb2d1sD00763mmSITNX595NcHTEkwn0zB1Dry37fOW
FufOhVzEJp80NC5qZ/+F0Vk7Ik02dIR0elf3clrjeJRK85K4e3Hoo4xn7YbFUIms
l/8VZSb14+JVGURjfswrIyCUotIzlzVYZ6gzoZwDXIi5gQIBf/gI+KxNXPaKV+PQ
Ufys/12rjO6aI/pPlqSm0hCvftmBcnezN2hk1UeXgOIuKZnogjOsf0iJVX2aOOWE
6pD/psybjbnsNB6kH5uFTA5frkzIzkzl5d9+YDm9OyC+k84E83I/7/j+rk4L2dah
QJOvksSIzN867/4Qt8qYTQ==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="MvBXkzurAa5VTw+1JJ70nePUfoQXBvZOku/SMmg4TwQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
oRtzZL4VJ4iwysPsC8SXYCzXS8Fw2gtZTOskLcDV+1B9Nzn1zTyNtlo6lNICRmmK
ZRVu2BmCc2G+fmzynYlNTnSa7C0Cuel6FYpxCBlOuk3OF2tzAmLAuDyOH3Z1Yjzk
a0aHuoCdIRKv7BrZCdALt03JeUmXKPdOmIlkVGFl8yw=
`protect rights_digest_method = "sha256"
`protect end_toolblock="Jn9CQpRhJt4rnzZPRk+dOpzAubz7omckX1MrFd4p81o="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 4160 )
`protect data_block
gD6l00tciPUa6pDNTk/+t0OO0nC/UTtBwLB41d4inuAUA3i/ALrNyoJVcBnAmEQW
ptbcNp5fxEUJjnOxnedyZEuEBxWRieZFQnkRdF269oNX52pJZj7FVsbTppwRhr71
ncQDYtLPvWDvUKItueijoT8NPSbdo65a+gW+cmzxK3FFsv4jHlolpprgO6JdWWl0
XzXPbY7D6hqr76ky+Ul6mk7R7aQkWenPOvpFagxCZM97IQravtR77pcFZbdOSL8f
Spjdg3rb+AkoT4UJC3NuW0iQD/hirZUviZn3GzVEWrB++dhds4OLMVN9qEbUQ9c9
Z3WNC8/hauBF3yyL9vC2/ClDypUhdP6/D4IiNAC91oLUtE8H3SpbrAuodaMSVs4W
ZqmvOGSHONKQq4i4dDTY3qNUQgQ6QHfe1o/IvK/Gtbkh+HK+asQ1jb/zer2rknp0
J2RmQghlfwkJa4jy+L9KX55f/az+07IDAs2AV2GyY4vNd0Bx61Q3zyIcbWlyjyOQ
YAsC1TdpuNCyfVrEbbA8MBCNkE7uBljmKtV9mUycGeH79S9kVAUYxN5MD406M8gu
0qGbd2opD0ixWH+thaI0XiKHFEbLQVTLr5+BoYSCcOdYdBqKGNZFgMlmEWUgokti
ovu6YbiGJ9/yFRdgYwrBRvxCVkNM/UXDWGgVS25cXZfCr09UqAuIi9B7AV1d5tm3
uzLhfLfjnN5tbRsDsmJBwfQDIQQbi8pRRbKjwKrYmJGMh/9aR44qk3yFPImS2zbs
RfM363tBp6WFkHSUdN0TLFTJYFhRrDGQmBpIcv0XWseA5YynXGL1PhFMOj2MT/Oq
3QbOlL/+6rkZPkbah/KFm79oYf36Zn5OzonhDUhT/r6hGDLHFmR8E+oh8jdtS1MB
GSqU8rMz5rYePMMXVHejIAEEnnxi/C9aUnaL53MATp41jXpwd2MvtbyB1ax8Lni+
v2BI1X8l9/ZxyxFyrtJKS+gHH0diF4rxNH51oRtNSWNDkvm/pzfJVa5POjC8oKrH
z+KRZKJ3Bb8aV11EAfvnBrNvGKFBUYUTFbr8gHy/DGJJ6CE2qEd4DjSC6qabE5Oc
0xHratgi++xp/cKV7PEy4oy6jWZ3yepnAzMJ5yHD+zTI3v/y7nF61md0xRc4dFek
witMNkr0KSVlxom6r3EII84U3ItdaRnH99JYPgkiVFdNuprGkMrjHfMeyjtlUFEr
YHGEnI0Qe4//6bXlzNXDXOmp8VLznKhLIsghmuCusKA9EsvnSSTTV1NwcjHc6vth
zU79RwGduxd8zIUIla2TKTYG6qoLJYAFFKqT3LzvSg2GRr27opLs1HrW7dF8U46l
JaQuFQ6KMnS+eodfoy6QJLN/3xAT0rMOOfVt7g4J8HjUjb3N5fZgQYzwjkTjaJNc
Li7iDE3+k5KuZNR3jdP6gGY5S9M++vjUUGCyRjEP9f5m6E90rp5HJVWh90CdnGBO
ISiuxkQNHfTCo56Xl/5aqzc9Af9IXnHmUyLduHpgm6jdknUCYW2yX9DKvmR4CfMI
mi4U4+za1jUukaMqNIHaLHR4N6W1vGqzNpweaeDxUjFDRQ4Bg9+BGCvJCi5oT7/p
PABZDwbPzkPKeCs1jGJH5m5vWcl+TyV0y7BkCbVX+gggCqsfyqBBxAN80WQ6TR5C
9VGPn+nFldW0qfYfQnGeyYIuL9R3V/0M7I3nmQ4qU0l6b2Pe+p9n8m1KczbPJMde
WyRzuDXbJhkz/HbW9kG4sJdwT1kcGpX4Jyt/rnUU+fbCnCEbpspU17iPdsXAHaFr
DaIHAZ56FDCD+zd+2QLhONcZEi93/sWeIwJwk5I5jBj829DQnIyYcYISy86TYHpM
+vOWNiiZi6cHTSl5begiMDJE6MgFvknL7XdnWBfwmCt+y4gqa2YrsEUifl49BYUj
qyk+8OT99q+JyKjQbQfegA2W268GnwSJ6B5vPVm/i6CzUaIQh16TNyCMApB4hIbr
0JJ73z43+OsD/iZOQRiMEuxEYCCCngQo5UUachtaYddrlK2PfLDsrMx3k0OG/Q6h
cdXVw8qdxJWX+KtxcIO91hX06J4UPXiOu1XeHkJFMJCMaYsGx8dlAht5ZrMVFbkd
uHGxGD0uGkvckPmcXjW9BJkQuelAAcukoMZy4YB0PxzAVynLFF+2fiL3zZ7fIcsx
5sVb0iN/oRMUutPUFosFAgMFbTrTqLYIzzUUZZwu2X8AYS5wdKZkVjUOc+Sax0Z/
/VopQGntrsOJgABVM7+UJQyPB7rZ16CBrynAUQ03Mv/Fhy53LGvZKfAph4U0WGL8
4O2CIm+RfEa/F4EKVfgfvXdNPVC8facP8tHEEeKw33B+w5QbWLJG91bIQMH7JKZ+
wP/WpbnKYxqJNmKAB1QB/9+vqsnumCyVYCJe0BcoTUKnI+UDdfgRqe/CgRkI9q9A
Zt8lkGVqjjujtC7WmLUWFlQZ1FA4z/KsTlhW9jRrSuKFF2KIsVuyitlEkqXZAO02
Ih2jFRp9wXasqzvEi4c1yQb2ZX+j47o+wvj3g3wF5Ancqt6Y064OY2xcht047YlG
LLNw7cMBdIBuDmn8IkLDMJxi+4uAgSdQ7crI+aHbCiSmudLHWEPrPCVf7Lwt2TQG
vkKdUogkX8txcmTQ/XbmSdA++027E8qihkBGjoSrAzlDU9pPB30h945XMvfHlhYv
o9DzXP/P2vIvw/7B+UlBG9kFxmrvFGfSvloARSD4aB7RNKmYyx/MI/Eqeh2XsCBj
DHYrBUaZmpILmxdINuV43erkV1uzpPTV/BplZNmFPrN9qzXbipi9OjX7UsQ5582p
Spt0jsdo1BP3Av9jKUI10cL8z4NWXp9p0C+6VmqpPE7knr2oYSGy23Q6InjLpYJX
tZNgqSDWBgFMZKUCChCR4JV7M9tZ9OK7aeyP4D1yHn/y/EcgMBBLB+Q0/2uCu2Ly
KlhBcO7AFrk6uzlPPVAAE18GV8cFsNSiAiICUn/b+esr/Z5r6JNuWdS0nsHQnYEt
SSJdXEjt6/mU45IhS7kqqr6oUFUaHABfRRNy8whv3ceeI3uxbQCBAH/hbrssLqhY
mTyg8RUyht1qV/BQhor+lBUL2s5DhZx9lZiyfKGDGBMUiQFf3MDNScHzL+dg3HMU
NPjmr8hIdjW6Yqc9Wf9hkE2mx/951hXA1jOUTcmz0hb4KvV1ROmM29geHtNopjPq
QUhgro9ycg1adHe9IDuI+WeQEdjfRiseVOELcwPOgxFwI4uk4shoOCPs++1OQXsQ
cdSkwn5yVzTx5bgKRKlsVt+CVpylk314+l5aFGcPhFeFo+MqEES4CpkAT+ZmzSkm
YGyqy2yHHUmXrKgnGywMPgjg/qgPtcoc1V1CxRCdwTrUuw8Q0nJSiIyIShaYx7eX
b3+OkOGE5AmbuF/vKruJLZJ8VDpXqUuxNDMeeb4aW/IgDS71rRlhs1L6bygkfYdN
yKff10dnz9zbZAIzCADRTOu05k0x49dWae6oLd/icYgOLFZ5dGlu8Tj671Z7NkCX
anrgO9lPnjTydjSbEWAZqZgdIqPGfdewKMSFGaZQgfTVLG9duwmsFPyzs03LP85E
fw2eWgt8Ytny3sGaZSCjnk9mSnmgxbsSUBtmgBmSnzu9/vSBo9hNKvqukU1ktou6
j7YXrQCzDA2kgevmpFI9i7ONppSrT8/b20ZmaERnodtdnI2k1cDaySs+WGlYCBoj
pE8YtzDkQx9HeiTFZnCVFkyHn7Lpvjhau7zBQLfLPpP30aa5p5GjhUefHn3jnngO
1TvdYFxVawpyrwCzcuVC89U9nqt3X/FWCOkVxZQzvzN3qsdE1oUqatQEjtH+ZRgC
9n8Wjiuj56yaNv1XqqVNcs/xO+F2+gMJpsriqzbV61M1fE9GykyRnnFjZy/q8cjD
Rs1bc3rsc/cMLalY0rqdDWVx3IhLpXLtQrVQIFL02noznKh7XOf4xKqHuuD8lqK6
EsURx3R8PzT9SI+AA/qgW8lFkDZm7pOapid1ez//K1uzibgoZD7HdT5sLm3sTvqu
fSHaDjP0aHQ+3oowyQNXRtFpSbG5QFAFzXx/mdZOYXXCiLsX+PCoRcdHiBY7hz5g
ifqy2u59Jg8HwDYjtbNags55meWbPBUClnu8HNtcKy08xe15HMkbMoBjl5q5Z1Rg
U5NvdYsaShf40mLtwayIsniOHhJmd+PXVVvHjRvlc2CY8lD75Ju4AdBzp34NWiLD
K9PkZLnkOgajk9S3zgZXwQdRsUV8cbMQbMMbugA/liPh1gm8hUIqQJ2A61EbunYV
3fPxc24ZKdMdeey9NacbwxsoT1k6ET4x34buCjsULSlxkW6EU9QiyD9lyIulfFbm
tPcjUE+M7wF7hIh6jBXIa1ur9kAChC3hiRz3Cyt9H3qYmSGZys/r4V6Bk0D+wmhJ
Tu/Q1TaXbaoEIZwVdRO39d83Zlazp2/z0ZEb9rU/C1rzjDcPOfsQ8bn60EB5N4Gc
ihwykXX193NiSP3CVOKPxZL70SPziExieCv5GOSeugwh2j2yyBpGjYVf6DZOUm7J
AMFHTOWJlynkHgc9gBdCUEzKXgJbeW6fdbofZ/ne0wIrEQQuWfnDW3h1cWE8vduz
sR1OrgSa1x14RdCNmHbx8FQXRz4fqEHLcznG/+OtRH9bJOHQersYApbuqVcDzeJU
4CATfD5m+buH6lbOJniQB7HiMH15SnVav5VFI3hP0YaS3V2r5kDmxRrX+OBFw0t3
cPkcLuBvax4Q/q5tlkDzh5LQk1nLQgKrai0puXM1FWFVbw5BRxdn/wDb+SFvLyuO
mtf2xVLT/K3UY6WcbtZmgpEq8nvcHBI8EDOqf1jmk5duj2JE8E1zQ6cfTuY4IYSE
iIoY76Fk268h3VAqAc6jlFF8fiSfujbWbHwI93AxmlKxbLR2j6MOnkuP7J5EOvMK
RKLOJ8bf7sz8uSQo71lfzaGZvPaIahFRtsPKRmN9ZZEgP2lgir08atxgxGuKhxPt
bgx2s5qWDKSKIxrNIR7f5QWbcGIty+M6Mn8pm/8rilmCnY4N5OSRgQyL+avOzmAb
iqFrn64zUxjDYPfRz4dfhIuH721/kTg1u78q8ZkAPxj5dq+yeylhvJ12/3fdWRMj
Y9f2sJqPbQWMTvZ6pkKXT22H7ktBS8ghahoqkrU/lObbDIGONY82Vzxp1a5RwDm6
ldMhuEBYGmi141za8midpQ+6I19n0HQAezYFH/FcnJzeCLEPCJjFVfxflWSVx8yW
7W/Az0UVKw4gUkE5RGEPJrtmctY1KcX6XTz/tjPsHdHGLOXIfuRZSO+aIMFVvYJP
i/0xLd0F2eHJ0sEfTyCYMUPOt/+0F4eUSJfnaHF+zIVEVm5n9YdOWYgRodGkzlFl
u3G30pGpe8LPXyCPhzFenPgeOe82WtKsIMlwucperzKW9xy3/lY/fXWkESP0c6al
Oew1nWJbNN6v8rnnkFBMAJ2hAQgBQgBR7nkR+T6u2PYYRgmELASG3GIHc5H6NW9X
DAHanBzQacF4C9LkdIfG1TO04Rw0k15OuFwEUjRP7xk=
`protect end_protected