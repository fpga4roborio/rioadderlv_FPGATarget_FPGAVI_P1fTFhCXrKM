`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
ddtXksX2+yylW5zu6QL2Lhnb2d1sD00763mmSITNX595NcHTEkwn0zB1Dry37fOW
FufOhVzEJp80NC5qZ/+F0Vk7Ik02dIR0elf3clrjeJRK85K4e3Hoo4xn7YbFUIms
l/8VZSb14+JVGURjfswrIyCUotIzlzVYZ6gzoZwDXIi5gQIBf/gI+KxNXPaKV+PQ
Ufys/12rjO6aI/pPlqSm0hCvftmBcnezN2hk1UeXgOIuKZnogjOsf0iJVX2aOOWE
6pD/psybjbnsNB6kH5uFTA5frkzIzkzl5d9+YDm9OyC+k84E83I/7/j+rk4L2dah
QJOvksSIzN867/4Qt8qYTQ==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="MvBXkzurAa5VTw+1JJ70nePUfoQXBvZOku/SMmg4TwQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
oRtzZL4VJ4iwysPsC8SXYCzXS8Fw2gtZTOskLcDV+1B9Nzn1zTyNtlo6lNICRmmK
ZRVu2BmCc2G+fmzynYlNTnSa7C0Cuel6FYpxCBlOuk3OF2tzAmLAuDyOH3Z1Yjzk
a0aHuoCdIRKv7BrZCdALt03JeUmXKPdOmIlkVGFl8yw=
`protect rights_digest_method = "sha256"
`protect end_toolblock="Jn9CQpRhJt4rnzZPRk+dOpzAubz7omckX1MrFd4p81o="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 3712 )
`protect data_block
gD6l00tciPUa6pDNTk/+t0OO0nC/UTtBwLB41d4inuAUA3i/ALrNyoJVcBnAmEQW
ptbcNp5fxEUJjnOxnedyZEuEBxWRieZFQnkRdF269oNSlzD2ys4W5hh5CCMd9G4i
s9MsFQakgYlQITYXrJInTztCt3ZOYDMTn6TEWtGuy5POF2DOqkzN5pSZj8AGHYSG
81Qc48HANgApmuzQ5NbLAMX404Oe2l21ENKJQh889qIM7iMEuWVJHvK+VzjxtiLF
wftQilIHWV/bnOe5PzYUOeWyaAmtXC6mvHItgSU8zaDY1Ywti8eKJoktT5f/vsnR
rCgCoEOL8sINpzK2H9Bb6Y9vVZ8zKBiCnIhpdMxNQccnxKzZMwLerxMvMuyGGGB0
oJ/O+WXeZwMbk4aBZsMu1sJMS4TKpyNKmH12sW9/HJ4PyzS4Y6G7BAbBsbGMtJJm
LkL44DF+Vayz0BbqZ/7yUySrPkCBNjiaTYAk13UZaZe9wHtyjg49eGD+ZsxSyBMj
NPgCnkKYPf5T0dPH2HY2CTJm+HHUe0s0uoCpWoJMTPxGrlDb1sk/Nnl/AUVycDxS
ow6EGoTtLpQwe/NJhdVHoeDlrz0NfT+YzU06WLJsKfJVVv3q2qBLUrv3dLv1vAeA
uVCeeVxQvg0Qd5AA5fJXCh+m3p317lSJ9YB5B4WJwLfC9DL99G/NmctABKXLXMFe
TxHvcNBrkLw4IqjBC4xs3ndbtum9Rb1Jyef3xaJ4daSNTS1IFw3SpBic5vgZh3Mm
n36yurinzFLY1Bg5DjctCNS1RNjhJaTF6BCuQx60m1YBHG3tUKhWyEbKNyAD64Ju
i5OCCNaeOl1ETpVZ6h+wjPJzirZ/rtaDtU4/GpOV6Iu4iRskTdLHXMCYkFXCQIb+
FN/RFfTHPJTzk5luZ1G7nEd4HaU+LK8mTY3mDHN3j3/lmKk9uE1bn4KqKxc2y4Ah
AQwwZYh7sKfp7ijfSsoJEBlzUh9wakcj5GZtKpgZl+mpDLA1M3MT37zJTLTsNgX2
kZ+n9tlNGBdoLYF6JG9eVwCISBemke6re3tIo7hMHLf8O7nG4LOK/iMHi6uq/V0k
XJV/t/WYsmRfn6n9BpGa3JNfZ6wH9fr9YWHkJByUMgjIZ7a++q9PNSg6GPOKkERl
cISs2IK4ZmQbmAo26m3QeDy4ObH6IidEL0W23dnu+xNPgS14P+DY9svBMgWE4dSI
LYCpv7BhTNfQWW2AV3olOFuTLgQDKdv7vxPIxbfCC7UywdOvEbXw3jrws790qolN
GPwp7BXkWd4Nx0TD9Rwt9V+88Aekeb1i7M6MaGxtWLzKyH+5ucmbtVjcu/xG1pmj
IhJrtof54M1o0UtcE5Gre7mmjFFqf5TB5I9Q2mSgXzdnzZdBYq7v7QxxKMdoh36P
/59BuDfbrpOTMZOL9AvtHI46FDpEIPKGhfjWM+ayIHrk7naoKZ202iwYonxl7NCh
SI95J9aPCqk9qJF/K2LEd7yTyUpGBEwZ/KnE+q1WllzM2nL5ZdByMJoNChMRpuQu
mRyNwZmGqasLVZO9pbPGGJHi87qAbodEimYo2tNsS3fIyNXHg/OvoeIgvjNTlNxr
VXy8IHrXNGDndOjhDGv2aTxgKICnUf2bZbhs7M9WUaPb1EOMQTyoIdIjx/0k0W0B
om0V09Lf/fvTv1USaWPChccDCxALAPcLy4qCZ0t2xPLlTE6JVAj7P6OHTVFtsaL3
bBlRp4/PunKE5E9/Po4N7Pp6KIDMtT7p42326a/tDn67ia7Wvhm5xyeyyZGOFfsO
OEvOyi7g0k7AayMeRHruhWpNUrihnuNO7fnhnRlE2HV8ULUDPEURwXXS/+mZfuJt
s859+r2Cr5fdSIWBtj/RjZDZaH2Wwjcj+8tw0nVg1Pjfsy2WAqXCSRmXneAjOEsA
2GGLaGfw9aowOTVAYCDGAtuKLbrbS6HrQB7JmMVdupnIkkSsLTF/N5a/knHi0bvs
eZUkuVMsl++hcbBMWL8zRn3Ynpty521Dp/ef/TigKknfQmS8fuQYdR7ebWKD6SlF
oO1XyOu0YtPiNL/VI6Sx4ZkiG9Ry4fHYSFzhHOdiGXrfMetIIu6Os1rvVgLYWsRv
XP6fEJfOsDyX1UdiPnLHxDEKeUZeg/sXM+Zr7iJN1iMfEa3HdgWYd6z/nnneZbZW
CLuWPALvOkAdN/ALwhv+UsEK3EZNZvK+MRbgCRC+lnsD4GwFHp+lFFSSyonidR1O
rbTDTqMtTof5QH3HaqhFh8nwqrDNlNEehUkOLnqmEVS982OVm8NyzA3HWz6z44Q2
193QubIeQGwUdAgNf4ofYT+zO03hSfbm7Ke6QsL78vgsEgG9Cc+kmAe3N5Gzqx3X
nf9W4v7qFcSjj0/46F7AobzAeh6QOrPAnTk4xxRHJR5R9SwY9RxEvsB7QIA9kDJC
kwFKYGw9CDbxYLxBRyOPvxoitRs1zUG449gzrGGfgfHLMvy0jL8X83BgSWsfJly0
3lo0mBnUhPVFrx958gcIGdBDdkY+VSWyvB78calxqJGgMSldEjmcN3KupUyDRTqo
ZcLKthELrbKxIAd1UGVkIAuT2HCmfi68z29mu7WczwN693QlVCne6tH40YLRMlvM
zGSIltfNb13GvZQBqACoxPtl2WrR1XmayWqQI2Qii4W1GG9Hy8FNQMrtNzS2Utuw
37yJl7a0UfD+onPy2WSAeOMqwVE6XjfoziqqPRjf1git+yUAtTMbrKei90m2Axr8
bGUZWiZcVUXdZOje9BF6yB/FcQWHshJYlPOL2Z66kJETUwcpZVGVYDoKrJwQAAk6
i6OsZ5iKJ1uMWmyz1Xb0Kq5BRMrJJs6xk2PxbcVm2uQaegF7K9a6rEeDXEyvX2HX
nwcTssyiTzMslxKGVXLr5ay0glKjCHMF2EMc8jhHiDyJqyvdnMPPQUEJDeOjae/2
43zp6AxTduLLMivuHzv2Q+TL+AOQoQsLxd41C3C09a2QTkdfRoCStI7Ae1Pze9s2
iLEChdE0pwGwM8qe7pCdLsaxr7Wlizi987DNdNMGuG2ZZdvRS6yFOEAlr1OOpw+v
OYALX/E6TUn7UjN4Ham8VeezUDi7WLumEGZM2O2M40sGEE/FZt2mc/26CXJOZBFu
Zsalijz+ZdHLlUV5FgX9XjNM/O6t6/VmVF2kOTdOZEAuVk4LznX5FyyCOpGQYLuo
o+v/rmmDxRk2ioH40R+AfNkjw/JXIL0e+lwqlRNRbJEIgTZDPFGG3BjQss3jbkOW
niUlM67WWTfJ/pqfW02Lc41DgBcGtI4wJksSt9u1SXYlge8ftlXZ62KwYbU+AgX2
ZdRUMpuOLosxKsxsb9tre4ty7u4HgSwmOiGR1RxyXgF2DyF7bFjo4JQBWnkARYlI
nPFYW6o1s9FECQM8lNRcI0gS/h50INKIMNUw5sl47WInsdhBqe/CbdIWnbLsD+U/
4LsVX0/u2EZLNKgp3MB3H8umMiNUn8Cx6oYmutoLfHZyjQcn7oXDnmcP4H3kDVbZ
S1lcdVso15xAbCQ4ltxdw6V0tytoXVpac2tUeqemocDwq41JLOJBLec/ht1WBfnU
DVB7h7xbXWIRgt8MOgJrPoYxtLmm80gRSuwGjkvjgnPmxg1fCChXqW/wZKJIubgi
jMtNjm/vjoPxxwXKzun+WseZ0bXRnRcDFjPh0+yXGYLTbLU+dOsZlzv80WnQ+um0
TkZcfFUVgOoSFlnZxhgSNs+5M/5rWwTLOhpqudN2WaMrKaDh+yRi+8gAA30uu8hO
djawqFR35fnb71E4MkAF/AJUJlI8rBNNb3SvtnFLztA3iP6TnLsiWBQ9L5kV6Khn
29GYXn3d1ohwvT5o48nduMuW6dWmK/8IKxjaPzCdN36YZ0Sg31f7yBHZOmn/pmmB
7STdNBJdsSjTWQZwI04Yc9xRGCd/1cXh8faG+NGQONvPid3LhCl/Yg5CefNT1pjt
JOO62NOjUWnKvWMYabf5nwZUU+7BnxbpY7W1itD+jYFwHqAIJZ/4l2D1RJ9wvtpk
6hbqta9fcRRK53wksUFgWgw17mvuxuGVXb1yIGsfs4jQ53eTPKPsgvRCMYHplUzm
1QP9aZgJxA7zS3FuMFJr7W3SPFaeGFCF8O0CiPbsndkI0990XwkbiPN8yZUVg2dM
kH+EAwYiKcUV3OugY0E2PZoFNpufK0fLHolicUftpZQ4u37dO7ydDhiNfhUFZfqQ
QTEaQmybMVj5wmyovyHzdqEt8ZMeHS6MMgCy8OmU22MDh4LPFWMJrmppd7jlUT2K
k6ls4kI4mG6aFrol9MSa3jndgmiD+0qcHjplkGnXLZYk7z10cuO9v8KDvzzk4flX
PXV9C54mKGLRVG/Sf0p1UrhQ3T4yj9ctns+yNkrU5XJ9xTJ/AJY3YOvoSzH7fkAe
ofVGcFMAbOXUIdYnPzYrGB6d8OYfzibPxNkNZoB2KbRQkrX/Wl2XTwz8mXW+THGM
rT/KbEtdlZXNJe4ZWz6a1b9iuGihrEmQLjPCw9ihihUfX0KeNb+WyelXqLleMPkQ
dv2XsgeixmIdI799Gpddlon2UHxnNFGMgVB9RPgn6aeEe8B94/p9hQttqcL5R2f+
R/TqLdZy1bTyLqrolYaXakaZPUEr0BcQ6/DTErXtqj942EbRFA5PDKVI5jma+vWL
oVJFMkaI+xY/2Pf4HEUqh/KISqAOtP89/NHqPLrNpQQTRV4QNmdRRimtegJqHANi
vXxvYGwWptekJBj+MWkHUnLHotNDd9d36NDdHQ4n9hV2925gc3w7yUpgt8QCj4Co
qL7zRNgL+lBClZJLmABDH1JqLtlKCo+aDzs4UVmfa3z2AbVeuTObjhKs7wbG3l50
3wtHrUN+HdC4UlAbNEVBpgVa+l5QeXM72Y6vA3pdkKSL8jkcOtkPPvnKFhHBGTkf
FcSu4jqUyb+SI0GkSJ0s1w==
`protect end_protected