`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
ddtXksX2+yylW5zu6QL2Lhnb2d1sD00763mmSITNX595NcHTEkwn0zB1Dry37fOW
FufOhVzEJp80NC5qZ/+F0Vk7Ik02dIR0elf3clrjeJRK85K4e3Hoo4xn7YbFUIms
l/8VZSb14+JVGURjfswrIyCUotIzlzVYZ6gzoZwDXIi5gQIBf/gI+KxNXPaKV+PQ
Ufys/12rjO6aI/pPlqSm0hCvftmBcnezN2hk1UeXgOIuKZnogjOsf0iJVX2aOOWE
6pD/psybjbnsNB6kH5uFTA5frkzIzkzl5d9+YDm9OyC+k84E83I/7/j+rk4L2dah
QJOvksSIzN867/4Qt8qYTQ==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="MvBXkzurAa5VTw+1JJ70nePUfoQXBvZOku/SMmg4TwQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
oRtzZL4VJ4iwysPsC8SXYCzXS8Fw2gtZTOskLcDV+1B9Nzn1zTyNtlo6lNICRmmK
ZRVu2BmCc2G+fmzynYlNTnSa7C0Cuel6FYpxCBlOuk3OF2tzAmLAuDyOH3Z1Yjzk
a0aHuoCdIRKv7BrZCdALt03JeUmXKPdOmIlkVGFl8yw=
`protect rights_digest_method = "sha256"
`protect end_toolblock="Jn9CQpRhJt4rnzZPRk+dOpzAubz7omckX1MrFd4p81o="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 12432 )
`protect data_block
gD6l00tciPUa6pDNTk/+t0OO0nC/UTtBwLB41d4inuAUA3i/ALrNyoJVcBnAmEQW
ptbcNp5fxEUJjnOxnedyZEuEBxWRieZFQnkRdF269oPlOeZuJcPalp1uITIl2nMO
J84gq2U0QyfHyP+10pDbCmP+MiwycgYidEj0wEHjy3GV7hXpcQ8f5oEbyRw7RqVN
wnfkJ30+AVwY9BxnQNGX0yKidj6rGpCnT0rcGGozgOF3Z91SIabIfvGnRedaGDpC
zPOjMHmmiEye4uZegrW7oa7K8fPDGZX0dwauWLXXL3fXtF5UMvm6XLhmzgN5bFOO
9H2fZnhwkaB9JIVD5Oh+znyvvkuP+fxITLXQOjdfLBb4q6dFxBygvkOhTo0pk53O
HAtuL+Xx3VHNNB3ug3jrPpFGdGvKQmpXm1YEgSh9ygx85xtEMxz0UliXsDrXWpC5
6xz1fSLBWBsnknAg47dr73xv0S0Ppo+l2ka6LWor0xwbBh0siy1DTXF3nblxu8KT
Sr27Ej8M/aDh7/pWfYrCubYSj4ijnrVAhahoraUl/RHyhLPmMkzp4d+Va0SUhP8+
U5OsgQq1M3e0FaITnJjRU2xDCH49cyrgA4y4wK/t/Sv+EpR6SpDJhIyjEB1aw1MV
MODyRskZu5dB0EzC7szNuS2zB7HlBry2BDA/wOgNfKIxmeywbjOzgIUT7hDaWMOT
asllEcq5ZzBwLUIxERaaeROsbNfBhOjexyXf3miS2sLeG1m5P5I1LOR8yeNZKgKK
UY5mKoY01bAQjMSymbyecKDEm1300sn8cwxYSXmQMFisyO9oobAkb6pWgz0Qe3wx
tazdXn2URBTzjCStLI8CNXEsJu0oHB1f/iF4nHZIeK6xWg4rN85agOov/qYCHo2K
0Jbx9YWFjCZzHl1yr4mwSo+v8EGekkzznkpD1pgpgBEcPVGn+5Bzzbhw2CYdnpmr
mSxKQeH5f0C51vni0KUmThApv+JTe1vOMSksTagi9r0Z/R8s3+F0dl2o11cuxQr5
jbGsLjJto8fXTW+h3uUD8bzx815c6aGYJgYqyijanL5beqbR12WkWSZN6ZquQvAV
KSLmIH/ZXLF3aaQVb1SCva1Jv3SJVZht1hqjeD02yrp6Nwvvi9QByHiFD0SKSWS0
1iTi8j/ZoeU/mcMuiKPv4LJB3ozuyHZcIyGrdTjr8aGs0jvddHtihanjJLwt0Nlt
CnKysFKxm88ia+bzLFYvzghGhdBkmYU7tn9ZaywkkCqpEFyc8yTYZCwrP3zX5CX2
XDldczAseL+5nNZ7Jfq3gDnJdW7p7ksf4txc7W5x1xXmhUtkIOOozEcVdpsXd+5j
u1trVHryShK+mtvvQfy1yoQWo1oEQKBWLD4UCAtYva2VA1cCvOToMWzP/2ZGwB9J
PY8d8GQj4DEm5l8uls8CQ8Od+zUb6QRaJMIh+xoDGVgh8Rp0XXqKuz4N2y7X6lqH
+LhdLw0bXc7y5zOk2ChcawrHeI/BJyVuDIchS7p8BAA8ItWFVt+k8U/a/Rnz1GOq
ci/5kZR9soUnxDqVchmy2shMBmalHuBpmumxdF8ZiG4fvvxAsBV9F+2y9Q3XZGVA
Yem+qjrfGX2x2vsxfDVEOjgm0CDcInunNl4LtoZPxU5+8jV3hsncNAQsJaG1MHk7
moKwGeefU6XraWYqAdAHNu/odADxGh0tN2J4ypEqKg+fJSSjgMK9HghSQ/s5tiOX
YzrwVNN4nFWN1dSHVAU3w9fLXF/66sijo1PEIbf+38pW7rjE0nhg2H4B5zjqYBZJ
lElAkr6tqMaucXijkc3c/1CSL7xQ5ThvRMugYaZXF1rsSJ9Ru9n605tQBhJqhYju
GN/6WEcEdlnrra+LK0G3V4cG1+WDZDcGR4pbY9QvjVFHecdFsaJDc86zbg42DhY9
ViVELUVzTVdKAgxZofUckVQxaDA+UlfWcm3g/InzdlP99vw1kTtwsMg9qC5d3QPs
1J7s1zTvL6U3XGHZjn5ctQLVIWWFDzyzE4wdqZmQhtNifAgcc3+3uniDFE+V9yOG
V33uTCB9xLvGtXEIBAF+hfNU/RvFjgYIwjjRAsrR7r8O0tOFEfotyGT92k1ycmN/
eP3oxNq67MmY06VDTV6qMdewy6RvZfKnAtiY7ehHseRG3/fMadklwpsjGd7xjmL2
fsDOvB9TlIGT5+Vmn9vABJ1oGKLLaCLsPOJC8gAyaIergh0boI6D2cmil/tDm6Is
JkZvV8WG7yBTcguzzOJLDyE9guVKEu9UotEqGqEaqpBAPzDypWhhPNHO55qCQN7e
UiJn56yBldozJcHsB9Nx/0g7bG9V+tHh6UQk8BcvVwctXJ58g4BmK/d2u3sQRVhq
aMBFAXz5nUThvH169L6J7ghFte0AjVXT8IesC9lxASNBE8Sv28YUo8GIDbDs8quA
ifAnogEhC2CU+zVEo6SHA3CgxO3UA/os8UVKVTvk9VyUGjf35MNuKwXzYW14MJCR
MkHvW+KcmXdxNCtSczUOb0y474y/m69zOI8JIc9HAaNe02mPl73d+IOIqUxZIBeP
bl/nAqjr7p0kDa/48jt4QFxd0exaBXxl+4VSFWOGMsjBvRs5uoDKUt6P39NN3jIW
RUf4+BCLuLMONnb2g9+lGhcyUOL3aAOqkqnjT9nypnbSHtsBc4oyJz/eNEzhYpYm
4cDr7fLDVQz9DmUy8wJXbqQTVfv4lR+jzXYaVudxWIr95GHJ/mC7cih11fJnNlVh
17phsOnKr1uG664yn6iMvZTz1eo1/yKw92y+w4jFJo0h+m3rYcrARm5/dfH5YXmG
OPzcX3ulOyCiRilw34L/1bcQ7wmIRscY9iQkf9FaP9/sjpzt+I9XmJBrf4HdVOQ0
9OXnzzcKJF7cdy6+FFjc76r8XSAStUZrdNevl4mLyjwmL/NOtuFwhmOks0C0QquP
WpvpqvY3gPyMrEHVXEsrF1at2+4i5r498iF0jJEK+UDP/Ky+AIUzntL7hrHCwbjJ
BYN10DD7a/gonQX0RN30pP6Bu2iZQ8wSZieag8SQH60Qm5cUqOIwtEZUHQrcTkqb
gnf3BNRuWbvltcOQgSWB2cCScAx9PSKepfbKa3Os/krnuPHTSbLBMb/60P0/WWi2
n60Rob6tdXAv8m1hOAIbDs1eBj9U1o6tFj2yH8j46I/Q/cZDG/k15VLJAtNYCPk2
Ubr6TTvKUjF93Oo16CE5vf8L2aA6wX5tc55OyFimlTvKYNIDluity3pRtpFnVBJb
Sl09rbM9AVhQQhFdpnW79QD4jtq/dVlNaExR3v2dD9f6WA7UeCZzfxL4pKPZMgui
ijtUXSUmOYdESmoyBnNHePuh6ycArZ8LEozSvurhkKFxNDOXRRDQSUrJz1rxSz7g
+itZ5AP5iOq6ZVLQb/EF6Cny/CfNhYu9CNsodIClPuImIPYaA8Kx3oCuumxiJZVN
mcYxmho7JJ1fwdASUBWphxMArR1pbMlEzS4iX2C6PXXjGGfgdwwIbZnHctp2q1yn
cVHTaNdD3Wm+N/fQ88sidVvTWdxsuOUUwongE8eMwxFGhxlOx9btsfMutRB8xxXD
AKKYS/cYbe4n/5iX8BQYOVIFSdl/fzDdjGUsDD7Opre3XSeKGq1dHQuAhYKQOmvd
dYLjvd+BdjApPcKe/pI3HZb1YZ5SkfHS74/iBwpZHU5k0u1QpxsReFTLy9UcKkM/
kZKL/mu2e8CWG3MOuCaMsLrraeXDtQQgqNriqi1zJNcoIJL1/atERp95P/+MtYlD
1UOkQitJoAzi9kjn9SrRZO/NnXLnqAAeP2FZB5LfvVwfC71P68bZmbPu9O4fPkNO
xtttOXya/oYCuyBEk3diuj/q4SV+c863+2BlbVkJgLoelcgPjL0r0b0E6nTgXiyN
+WDBjNXAw90L2nGDkjJoGg0oF7WKbOCAGfCzqRfRMEBk78zsUpnBxA1l1dgp8rdA
dvCCYND+tNZ8fSmuCJc34lAg1871Cjmcbbz6zCIamqDksxP65Vsu4iyKgvv+j72B
dYfKTLnmErmeqsluX+Us8WoQ6/RtZih8Sxf5Lz9k1sbt8ShvAfHOeB+9twZ54oFT
03DLWiCM9xZUwHhmSgv4YOu8AFbKVQGP5og7z1FL+tGlhYLOA5N7FTKEH8geAUc8
XHNd7VX6S0Hw959v6IEZiKFSlUhxC6WsDiJePFluTvvg9S8c1o33z2qQxnORjALU
QAUdxuemgDiATF8v1R6RUCh84M27SCm6cyxr8AVKp8/E/V7IlIa1vs3yi0AAMG3k
DVi9Hrq4CTLxLN3F9mn/VDo40JJhYcz0rOZRNlgWxzkgkbdZVGctFJCDCsNR+NVH
ZV2NGNgSQXmhnRlLTUw8MQ0+HVYl1ttOmKiwRZseOlONyDQN09bEQghI8oxXbY9H
n38vS9kzHI170RqJQoxAx8HGvoiB6jlNGclfy21uH4O1/nhWO5ZQhv8JxPCsPbyd
sjbFmnU8ysW2+0mhhi+WKCwVd9K+zzlQ3rQnCI5oSwT6sp5Y6EhN+YJpW7buy0/J
vNtEvOA9JeSehODWaw7zprJMEq4gTFQcQS+sf3/e76buEjtyZcNI7IMyVXFwZQ8x
pc/ldB1LnFHnvEAUjV2dqbczuAIZy5wd2taUll4g3+R9ibw3J06AyApVbIS+0zqg
Sk+AqMZtCIptQQhvl2lPq/FTLWYGV12Vh9OBfak3O6gHnrO02jclf+5iOEp0haeA
L4vAMDvMWg2dRTfXxLKyQXqo2C5u9hvEb8GHMi0Uz7uTRHBCOjXeruJHamMkFI24
DkEndHy47x+BvCuNSf9UwhFSI3HDoYQ4Vty7NTmJvqBnqf16kQWDdYiKa/zrQ0Un
+8YwZaI3oX7R+ZezN1rJe9Friv2sHnQWF1C9h6QOsXLmq81HwJCvjJYbBqlByoRo
431pKkKz5CA3fa2OwichUIfp6MxuESiKzOKVAfogaCVZ/GesVZW5unJu4AZYzJbC
MXEymwd3lTBaBXgGXtTxeW4eF+rgNx1zkwxZQtVfOUOIbRDd59H3b8M9olJWL60X
tx8Ko/D7SaHeW0ySszsekrDcJMXGQwGd9frD8OCso3ZMvBVaPWriw5QLIPiWtC5/
ncXrXdHJXrRthrdBHUd0TnSABPA60RQvOppycsmteq4SqLWk0C/QqM66rbjjEX4I
QiJmSIJdp5sENZnWUHf2CkcvFLCwRSxTnN8WDLCC+1VvIjrbyJU+ryPT/MV3VQsZ
uLy1CkV2RRsSrbgi6SHRL5jCnOvU+RBM9p65TYAPsV6ejkj8q6ynG/Jq6TZlATyU
+0xxrkLtxQwZwt+lVt9u4EtHnfvpt5AZ77CoHk/ycFRAmuoEYIC342zLHNUyjJFk
X5cbpleX7O6upq+/ZXNzzmJT662HKBiam+whpOeVtEojTAaa4UEJ4NGwPrREfIhX
AhQy6/HZvwQX3Rfyf2vfXHlDED7x3/9TJwla4irILoV6aBUWuGf/59qbAoTrkx5s
9icLr2GB1OaQbkflq1yITIGkmQXgouIfy2nN+hVRswAUeWaqGAHzzKaxKFCBE1C/
tF+5HBtppC7YnOuIAey1UJq5bqEC6yJVqps66brmnmoG++eyySLoe99czQFSpxiM
TtBQCe2lvr/25m/n2wsbLUuppLrfxzh4Ns/nHi+d+UPB99D2eekevo08mhwxaqdV
j/Hq/ruAxOUI/SZeBMsQ2qqp4N4tsZAMQ/xWlNPmLSWEcv/DLZ+Jt1Z2ciCWMbsu
sIVy0f8gJaym6lCvoVtUK1LH2Qa/Zx50a+mOB39G4heGKuWtj8iub0g8gXX1yrRG
Tz1LqD8hAkm0mxNg+JJOy4mgDdhkhC8o+kZFYVmOIZARelG3vbSGRuPuDEeDd0yz
nWUJdUigUBYHSOEZ/9GGUCOGiTu+QET2XyhtHJRixZpCZeM8lc6WddwKlUZe/tFS
0NgHKn/nd3+EXxF6hN6ukCrr5af9Ev7B7RKdM1PCKCSxwMFbNKlQVVKu9sgD+e+l
3ucjYV+VrqGDg6vk+L1GK6swCwedo7HgNbwY5nq4fz02En7hD79x2SzLn7PXO20U
Qs14cDoX9scGO2QhdWKCvTqs0iNWCV9TJnuVsOL76fZ/R9KE9sdQJpdCp/OVej8I
6myMhBNiKvq+jmPv1eLtryk4dqoPBKn+a540bM80bQbV5/kumqEvk0XVv1FsaUa0
J/DkXtl9nkStOPyTGfLmmXRWX6PjkKbRWVG9536DR6aO5HaLNrk7MWIhJ+8CbL+5
mppfBYsmMPLz8O4dQhibH8JkTEc6kJ66ReUSHkTpeUiy2XajqwxgEX0MtVoMu8fi
rb3FQJozH1VHjlyY7B1UAyNdWKl4g7+cU+Fo6OJbv4jF/tShCIUGyU47y6g9zyjm
tuMBdMpni7VKvWDRf9z0FwIwOlqB3S85l2EOqCzEaO9B9KpsgDXTRiWrBihnm873
upP4+mpH78sFHa5PuosnCSr6wGyXf40mBXyFvLEP3GUB+0z1Cb/zlCiJswicbNEi
Br13IQOFJrqUxNcWj5/WAw92LcRy9RAtNJtHfQAKcA8LytqCXSVqEdWVOMtVVEp8
3dSQ2wvPadmtFqbJtWuRWei/EHZL3PJxVEfSm+88c8Rg/uGvazq3LEDX6+a/7TUJ
WBk4u2lJM4JtolSlZTDFtcyyZJCVGbOAKo50qq3eiVrIkwSs3pxZaDeSRN1+7bQm
c5TtPbdvT17pmyjpZ1YBBY6zpNA2TIeI0/nN7qZOKcquqaqBc/xIjVCoJAZ83ABN
PKZ3foj59A7K3wGYTTepfahPGVmpwe9BrHTLSfYBRs6XU4v6TEQ8VoME/NnF+Ewl
yOkSsD6zig3jfzUN6QvAbETpm9T77rBQ6eFAxJ5Dt6vFklZnxWzzJfM/tuiqe714
qMIqygTrbjrRW5vjMXl+iQH77z9YIE8VN4yqRi+TFHaxgN5gIdVF/21J9ZIU5Xj6
K+9BcNsDzS9zxWtqmJGge5IeAxlPAfO4LXMR8YfxyDgXr01DnoWBuW/vfXRvKYwx
vkfOJNAWIbmezu9ri8ozwkSsWB8rpw50rY/zPxRVr421Mbj/tIaKSqxpwltUfQcv
k18sS+vdaQk712Jhh2Wicw0SFXXAduSCI6fZsrF+iyz7CYfjUv3u3VWx8IEzMrgW
yjcVvan5Ywtm4q3Q0IzXP0l/px0X0nJAVYqkHnWhtRcFsNFgsZMtVMayq1dcFv/i
CBkyyGfp0W1LATf5hBLuZXsMBP3UXSfjWLidtkQXILrgSy+ytRDQoa5avaZiwT5W
dDGSA5HAAbWR4gbTHbF5SiytlTM7R4C2W1+ZZ5JXVARpUW2AhjCUCPLUV8G/EqmJ
PtdbMvlBArMpNJSSXj2vU3UgSmaUaVsFsVJBBPksUKkjQNj8PWC3lPoog7Fj6pAC
crp+nd+maHYroR9g6umtC5pVbTA+o1F1CvYjKGP/qr8y5PT5YEHp2UzZ28S1GJ/a
4qAu+YSDGWhDQ9XFg3tlDi2ZaANP6Us6442aqJ9GKrM5C0xj5CZZmajdxBOGS+yc
uSBsecSw3s9r5ZbzLlTRB+k5jFzrmChR0lZfpqfuLxw4h1FHxscaISsL0/uDfVGS
LbVxZbAnwtVOkgSSauW4uJM79wIl9YG9ET1oOE/HDNoVUBcXHE7WT97WiGtMOt04
PaThAzv6Y0sw8J7P9Z4iw5OHlT4ly+QtPAPVVgf8yUDMd9Sq6zA/GlrEzYK8ZQ/b
xYabmzEROfc7Tsfg2rgh827HtOLNzdwgLVC6UIaFuQXQCowBYCsYscE62Fc42GDQ
8c7zPguoHSPRAAoY6x0jaM5Rp8scF+XuEbXMxWv25x0G6fv9HjCgJAQKMhamfHnt
66SNftePYQQ1n3ddJX2mxemoDl/0ulsLutbpetfI+qfrJvBy/IheY4o+RG0+IPBM
W1pjRzBJCoaGXw5c15CAlS3r09I8BQmKXO+81Mqd7oo8BDYeqUo/yYpnhh36Bx9/
Eb2wtLFMHCkrDTlhlPPzj7wEqpXqlfxf7yjOgQS1AKydsthsfpee19b7F6ngnG39
XSdBCJBhsRaGbskBQ4PyN8ta161nilpz6DfdglMOYVbz7jKkK+LHmyugDXv55Xg2
jNSivdbzEEogpdOp3LEl3ti3XR88bAldh3r/Iq9Rke3br/ph97zt0DgL8eSxZ0Yq
MnQDvWjYG1+Hf0J7Iw8M/yqwkZk96OYykL6+L2Hl8UX+HmoC6d26Rk1NtpMJQRbc
MDWYWGbleHGoORDeKEgIFZEIgbjkgY+JYFGCKWfHrsLoGIW/Unt3c9iaZPe60VDD
L7Ol4X9yIyRXx9WyPX271nQI5GHN5n+6bBMSsevbjWOUG6Ny97/jaDbw0TzO+XE/
EDGkKoULm7+AEaVwPPMxkmymCYMS/hRVgeh3uNEHAlxKgYYQzK/di3N1lxG9R+Nq
lsk4Sd/KtupckO1J79rKNHfGKPSKml51ZdmT7wzY1FWSWQmFN2pLz4WJZY1M7H43
lTNHA69BMSTJL0hSVB5C/iL1D09uMo/+Q9ifFTMhntVzWtPO+ZEjD6vG6RebFgPN
YSFqZZ+VM4QZ/hACw3DFZb9nLf27onbZ9VN2gLKgW7yJ1ZAGvOLi29woJXcCT/Lu
UMuTOGD2yp/SCRfU9tRIucOmfe3uM4+kO4vzXpcoWXD8rJvn/HB59aWAdQH1XR8N
zkfhcOHwrYkTX0BGNRIQbItPwpUF0v4M5o53BDm61qwYul0xxKfL3UyTd00lEiVQ
P+21iv9MyGIkC3MbsH1csTeOZh4KbL0nFhapLTCthnPZoxxl0QMn5cXlmOgLf5DN
HecDd3CCu+Hl/Qz/c7xSJg+jEMf206Gg2XvF3rZD/LveUqLmjSu40qhj6PnRIBtC
vfcqajaDg7WaxBDewFWoCWa57D+kwmR8j1HYUZL1qVWUXMbv+xDOuvbQbH9UYJdn
T7XfVcwf5JcaETbw88TiQvFh+GBlnIHWJdk6wLAE2kKRn+tGEgNdyyDAF/4A4pHe
3/Kh502TyBGIJ5ESaaSmMMC01+n9G/ZrR48ZYio/+d+DP4Qp0EZ41kk7ZjvsvrE9
ZzAIckO6cObYeYst3sAv4vZJVtsVG2czKRgzu5A5CAjZjtXYUn6ebEvh58xm/4Mn
XznIAdYaVQCrs2C67gNTn7GpnM7H9YyYlOK5sAa/rtpY3bBNMlzIXIgoIMDngz/p
EbKAvCWQ+OnekNMl0GOFHkc1bBXgDE82grRo+PfV3qyJQZMd7YhLA48pjRu0X8Nh
/Yhbjc/vIKeVwJ084WVw4Meiv8XMuVjL2OBPIX0+h2FOj2exuMcsbvpFJdHHqx9a
cgycX7GfvjGdKGjjPSnOb61Ulew6ZMjAJUCfOytNB7nORizKzi9GRB91vDKkB0zo
hNlFOUl8m+7o4qlv2HyatBW7fuCt2j3gAOb8TLjRSsOl+1+wLLum/ycQD83INTbf
SBYxNs0USdKjmLCrQRfAN0OsLOMaaE3Buqs5YMxlTLOdF5vPMp/vP2MYBRwVH3o5
ggXlSbTsSSE6caVfZyJbeDC1T3yBV9+sDo+zZgtBN1EjKmDfSlhdLw1u7Y/4Yo9l
5vtCeaPlafGbFDIX7jOITJ/b+x/moBGwb+lb7s5Kv8HZC/1p2zTxcL0MrsMZcFtv
LQfFoJ60aICW2yflOc9kAsF8xvHs1SSp7kJ+ctyuw1TUoFydjgbXRpjPjXFeM1xZ
q4NM0TK4aRWKEko1eATVq3LPa0anRzEEBz2H5j5XH0reA6FKNG1yWtMEmGnAegJy
Lf1YALe8og7Is/MGgeS3up8RyClJou06gUWwlxE1JZu/volYO65Cws9K9ZhLvhx5
rdd097lY+qEz3t9BF/0yqJ7NaawrJuVT+2OixU3ytrS9uHvmR0U9QdkBiSyLVOm3
0N1JRxGc02eKHyJ9UNDedZRU74BV1aN+A/7kuY3EYVhaP5tZkMOT6aAZH4tQjwLc
jTDxqbp1iP5ZBpH4pxJdu2NU2Gs6tUhlr7/eD4+RLCXHnduzo87/cUhs2jjJgpnU
0VWh0MIY6gDx2eDpQ4JWPUKEuHQEGsHsM8JQF2dcqPDRwyzuRugCyvuC0zNry3pe
E/6hknoqDE78iYJ1IZ5V3LDWqvKec4DyERbzmD8CUDJfNFNqBAHsLEaIXulw6Qvn
cNlQUEolSZ1/qIQJTAipfdfi5HgaoQQzXnYj4DVrLeQSpgnpIc/EmWsGfm3mEMcP
ImctSrgdpLK40+ieYKpNuxgICsVPb8Y5zHuXSNMwe6JQOK8oJiIP8xHcZ/bM9+VT
QwANqVq3vvymppMSlYHe73W7rchMvkLymyfuWhLftU7LWXVWdlBa4AjHXAzvRZR8
VCF1IgUFoGgjvuNoRzNuqVOe4Hn0zkbeU+p20z4GwqJATCLkAGeONmWqiBlPeOJR
zanrC6RpquO3vMOl9pOfONoqHj2EA4Fpw5tZ0scuZcAteh+bwfPDu+kh8+hnK0dG
YBm8goq2EUuRTAXUD47iIx9beORGUrlqwgAYYeEa73f4auBb6yduGWNM4zjKo+HN
1o7ejcQDck8R17GLBZJ/ePmCxR7OKUiMz+gg/p3XK66leauITvfqlmncHAee35s0
rSpNNVMeMSNCNEnfXme0As0py6vImitniFBLsZH6BeFm9oUIaS2ijenIhJU+EfYc
h+ukmZFJMEmjDQqq6yr+WeB/3DFbqCA//52+I8TZVy8+F56EFZzdEaAbEQpYqWc4
xDnZYUjbuOFgT1tKEyS1hrQbQHq710t8f3IuHKsE3m7Mb+10oYHLKPPXBkK81+Io
fsVjO5WlkfysdTS35YyO/sNKplad+Hzcq3DDKj+f4Mx3OeQzBbaTPsBrvmfXGKPl
A7eO0Vvk5Zz68QzKu47wtFSL0SSPdPASmP47ZPSLcqZa7vqJzSitgS3rNnDU1otJ
uZiwQpxliNILNBjS0HM10nkCixPhOqOHKuN4zpV63K/56oT8kIH/SMfpwPigK0cU
WtuR/fMYtKQsz07CnjgCTdbj/EW2z5IJfpZbzG0cL4vwulzbdVVAhHLM7Il0UKpa
Pp7BD/9Dh+OEJJhQKX/ej1f5LzwMsfU8DKzyZp93Fr98peqhCLTkmOoClgMNNZlf
JLEGDWmmspL1rZYBag+QIZotKbVMo026+mG7CwZfAfne0bBYGpfQKdo0P7nUVkAK
lXGSzYvuHHRalwh2kWU2D03B/1Q9mKgaH0tXQTmN6YqnN59Qhw05r9vK7Tt7y+Mp
EpxP9m0PwxxM9plGDj2ZLUaGrsZ/0be02hpL5xKk1g8xnDA7/VCewqKjkBgAFcgw
WE/ZStFVdoBbqNV8YwY0Vxq/HpJKisBHCvtlvdOg0ZfZLy4R/lXt5xiEIqvi0hPy
03i5Nmw+ggLsmBvBPTiJhbbIUsbjzqB4E48Id9QJt8P+f7k2TVGiw+4wJgCxJ4jc
URygCN8e1o2lKvVOjsC6X88Y3mLrHjQKnBgyZG/mSSaOHY9pamq+53M0kLjY+Pcp
U0FgcVm2kcUJr8fG+Phh+yN7i5vqjaIbT2I6eQAgDVxepCDm9hD39zV0u6scs2fw
e8P1ciLMKD3n5Ksw2WFqHYR3L2/aBsWTLfkmnLiuwlyHsAQOvad1gWJIvY0AlWep
1gwBLBubpKGHJ54WHswPP1ZmXtKvk9PRbQF3pu33eg54XIOcWUQBxQSEiiAKwvoY
4ipE5Yped2aWl9peMJ1UvdnYeX1gReovJOWmFomzzVB5RzOD4xk2NN+OruKa5aaW
llCRKPfwOZrzzUFfuW7d7R8sBuy/9enlCsxeipxNmo+r4ukb9qZyaV+s19SKrKUF
A7u4a+gHX3+GcUBaWQaCTjWlCeeglXOsRWpkMEeF9WOnP3M+Eljd/sN6c36lUeru
qreNIVSkD8PH+A0PwL7txCz1h8ImnQrN6hLZCwOWI4pD8BzuueFSoUZRzJxsE+4S
oQ0+i2jNDR78nH5gUyX91ZuFcCi+UNdlkcHtxkumv4TiluMCB+XlaAuhiy5FQUjl
hTiNQ4b/Ym18zKbihONto9WwVVsPFuJhXY97MSOPInrz8MAlV2O/BdpZRIyyPOVv
l2/9+dxNuTAdllm77ykgLvXMYa18Qp+LgmrAvrVqtEeNs+C1epp1sXBqNj02VbQl
9IQXqOo0dv0ZUIn5UQiTqgrhuO/6U+nzK9tCczgzm+muI9LYnq7R6BgcsrYGjWIq
zezHPpnUwx5xHezeQ6CkmMuSHO41VnvABQIyZzmQeZ9eOzkXRUWN6FvJtq/dgf/N
EXeob7bynOkHoHXfAadxCaTK5MAM+9PfCymrH2m1gk/6P6qbmdC2s52HHhoiPrzQ
PbHdCWNEpgb2eeaOzKS2k+Cf4opUAboNMbRBGaS3Sd9onGcxTgllZ1tm3dA1NwDA
qXoBNAaiRTXbJX46LdubabOJpbzEPSFNLwcT/vXpwqJ1G9f9/roMzbBiZin8gnY0
7xGj7fliLFws8yKkXGy93e6RyZIcjVjirw9/HuGnupu85bMJc4bxYM2zjJxSxh0X
owfKAEg3JAuJAmjo/Ovzo+kHV5bc6RXQOLFlpiVA8oBGWMwQnYCXaoEjpGstBC1y
Ehlo2JetRmWW50cqFDdnbAs80gGEzsvCsfNAzJdRFaNzY5Wx3EUPs1+S+yp04ANS
wBnB0KQD05XsclpzzSziwOO4aqOlhQ3WQMc3uStOUo5va0ve+6hYKyGMerareSR4
WcZSxFbPRJR7pDeUD9xb2BjF/A054YbpTnU5EL4S+sXIIU5K2m9Gzaq4ZuZZvEzm
nkew2NaBQI11CqUts9ywj9wqQsKXw7A275IS7V4WP8yzZwGzBjOmdpf9oyUFaVpy
KY22Y+TByKkMfPcXO1JggJx9gNJSWiFpdEfuYmL9RhPkrVI59iNNkiKqNgpXHfEF
3BZShYsqz7s+LVV4Jx1GM/kOfSbKHlWUIv8PURQHHK1ZepVPRvgrXGI45UwssPo1
iZetURBeHju5c4/ofF68jaPAGd7ySAOi5MhqiBmC+EbzqFOx7eF1s8mQCH57ugtc
R2QPEBURWR8fIf0F96bQzqcDqwSnZiF/LuYpuD32lrUpzYMR9J607n+cBl8UoedL
L+ZX0Jtvon9U4lGp64jFk1Od4WZNOvsdKv+6KPrKkq2u+HUQp5hy7ceomdxYqd5G
uepuBBWyaJUWqqVO6W2OeB2xr+bQmIiDe7AENdJhkCkTPZjaTNEgROH2qsxGMKZH
RZxd5aHdW7F20UX4N7MKuKvlvUXv1pR7RdtvuwBybUgN02w37pkFX+OyGMDJectZ
YL3eqFha8OzmHDZjyc43IzpHpqXZTSyCu5h64SbH1C1QkLq3QR3RIJd9UNPzG52k
T6z7mU0zhywLnuL5DEAK4Mz+RN9r+qDe39azmhiG8nogAKEEXfl3D8x9MgQFdPNt
UH+RO9a19YuR/Y7diC/1Xcmu1NQw83VXwXN+ZXrWjLaqGZyWs4beNBFMyLUgKKaX
newCaxeFJjBbptXbw3Qj6D7LIh9/QNZa3UueBv3aD6BPEQsOgFE0qEzw2aHRhsi/
cLXQZlips2nZP5Cjlb1uknXSBd7Oc7dz2ZMquLBCe+NsUq4iWyljJwaQROfBJmU/
J57x8L8EzSpcG9tH57iMJv+hMN30Y6BouJOHQoTy5AzpBZGerAYjgCfKAfQKwv40
Szs5Voop9JgMVTAs+b51nRtdOInL7gzNlpRzDQsL2HB+Or8WU2b4AIdh0k9KMCSi
KUCMXTncR7/viXqLrv6dbBvBLaDcxYNikatT1PNiJj9JPLLpfKnvZdiJD7aWLCVV
K9Bqz1QKola5QHqzHLda+L7lMcrTpUehtMFpBOQvzO89UPHqbe0uAUvpo3Xhsndc
H+P5wJp5e+yGmg6wJ09dsb9RpsrkP0+IkXId4KvWhYVBlH6/6AiYZhxmosffkNKi
mVYGcJN6NPBY1pnC7K61lj3aUdVXiYXxudppz4SUdRXyHtCD+MQilblWyerAjOsL
P8wSXVu5D2+RSAF2dhJWeTtqhphNl6ak4RZPel3rsDB0hDJtsNxe3EKMmxddRvad
QAKWGDT8Bi9g1NWKUxq5fZcOLcChj3Uli3V7O3R2D+naSNk6rKKapfHivSwZw1g/
MvUekOBIobs327ZDNnu3Ydp3u5/Lye3oq5dryIfEqSvjx2AAGfcRqXuFFQDSiu8H
Uft7ccjdocv1wp5bFqG1DDfm8vAke9Lldxrx8aQRBA9eOmRPAO89yAnyAB99s6lN
fckopUwH4O/XBxYNzFvs4ngY5+hF30nNxZ72akWi2O+9z9Ay/VI9uK/36wq8SQDK
6uREojPIXrcq136ARj3W3C0RBJsrD2j/wGxcJHrhYJOpAk4CkuE4MyZJfWtl6OmR
E0U1BwBaN4g4EzR42zXdzzFbXPi/LX1qRo8cmrCHJCzqjAtK6XyGsBg6++VIZdki
hcGhXsEWBCCSGdf2baGGTwaxzwxALsKvlKp0lN7QWHhc86plrI+DXrJXz1EVJm41
OcFGsdQF++/L7xUmrxSb3KFARLugkm9JGv7YCIgRL7FBKh2kNS93kNcBwLkcZu06
1nCfdQg1MxdlofBknCA4unD5X9HQRcS+zGiKEDsgq3cGffFQv8XLP8B8jJY3r9JT
KEk5wwrrUVY5Fd5+IuGympdNLxd22R/yaBznSFwHuVqkH4eqn/UeLXMCxULg0ZcK
VDcYjIT81AAhBkdHzI1g8SBQCiQs6nIWtt1R/OR5NuDi8WI3vjbWtuSXrRPk9kIK
m1UZolPNUrnH5ITcD5PdvrrGid/9qVMDLtDeaj9q4x5zBHV5UiQiicB9LDuwH2Bw
Etilwf1xr6O3yoRItCrsrxs+LnCLJJqrukhPnNPqQpgjJGhwrpAUmAHd49wbRrD2
8b/ngiqQveO4nTczfrMOoSqHM08mNQbejhRb3GvVe4lhOpR3BTSc0nv8e+fP4huf
uvHpEDaFdiYZNr6RaEp568hodIYaHVIlk6r6oh96C6xb2fao9WSXQp2uo5RsCl1v
AaaMqhpigqiwvKlI0hKajH9Zed47VtG8NDhEFYKNCeT3XIacxDRSXmHHmyb4rIYZ
ujYn0IDjgudKDxhpcV+i3nWCHapGuYxEPzSVC5prJuRmM+KBX3D+1vMIkdj4ASpN
oX7Yd02nnm1n7Vjxm471WA9Y9cYiZAdSs/dyKjO5Ab1chL6kXPozoAcpfCupMLD3
ferR/2494r1Ao5+zDsxwnRfOzf9DxPt66Uk5hcIDJeQjrTquEYIDjhzXWmAvP6jC
6VkriPOg6/AJzUnnp0KSwg1ydPKhYuj6uAfMYtkWEfoLzgrUnwZT0xuZxJMaNalz
ExNx9ghWd9ODLaZf2faHcxbnuttOQSHuUr/BZVTjfDw1tsyRbLK4SIR3M5pTlP4x
nrGlWP8JYf/GriAErxS8tp2QxBRDxWm4a8npmlNvgatbrQ/0vZ5VNs/te1jHB0po
DjcG6IR7mdd7ZU9St6S/mudZSC6T1yTc0QHOa3LEpCSHU6Vmk8UBwbqHsfugj8oo
giD6Kvpa4LJaKx67WnnpvGKFZMkaRGriooJbMvg8e9vnHlc58Uyw/spG3dpa4v/N
jUgL9qYFzkWXV4eTeWrypOV98FW82o5KkcMi7nmOCHwnoPVkRdV3053soa/Ywg4U
OrXUEuN3vic/SRx9vhcr1AFy9n9r/VwMiNtUcyT0Bdo/PrGe/v0c7t5wCT2Za2ys
8lvVz75y6GYJ8Zq7zOlx+D+vFmb3nL+sCUFNxaw9gmey8O2UDov4AtbePgf3Hd/j
b0oL+WCYXJHqZEdzosoaV98Nwh93ZWYM/2FOr11curX3/ziQe/pDW4UQ5jb6Rgae
uzCjh+efdQO0L8EfqDl7s1XHrtK+kLx3SNybKQhwoBgEYFXd1tivpvb4hT8e02Ug
X+Tiywpr2Vrl42tQ9wA7PUaX+Nc+kRazxF5BRzdEyKrcukAoHHS1VwuEv8hPulGa
5rQ6OdxchUGAxZUfR9yH9ua1zdba7bXp9xMThGLvhXW5tc5UHJHiIpkA9xSmsM7R
tRslYc3pN996Lk6ftSibnhKZpL/Ey3H7ZQjEDrW2EB+swlVVlHumI9CZNQKpEWz5
/ujI0PbN6jDI/yXMxamgoEv72dub7uhjSB2Qp/VGz66/jU/q/4JKWxLa9PBYYfLn
yPsS0xR9408XjmXIlQtHTXS/lBJiXNETfYwP/8C8P2AcHfuQ0PgTecHV3YAfN55I
JVTEAdr42CAy21n/qK89qVPetbO0NK3hVAbMjpzsWcXT3E5Xd7Kse+1LYNAuy/ZV
q073c9tLp9c9qArj9TdVrTGm1gU96yKpt70yedjajkZ1Gm+awL+/No3xmUpoPdwY
nRo7FyMcAP9g81fx5aURLxlazP+msHsPBuTUgLVh6+YmobNIvSCr273oboQ5lR3r
/6oVQfVnVlGLdhmQHc/rm6DVXWzG8XO3+F5lvPGucx/EsGcdf/GL17u7xzP/oy4B
JjlqtAdwDPOXDtsLV38vB2OCE9yrRXpvsOWkOVJs9lam+v2WlJE5pOQHvZH0nDHZ
`protect end_protected