`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
ddtXksX2+yylW5zu6QL2Lhnb2d1sD00763mmSITNX595NcHTEkwn0zB1Dry37fOW
FufOhVzEJp80NC5qZ/+F0Vk7Ik02dIR0elf3clrjeJRK85K4e3Hoo4xn7YbFUIms
l/8VZSb14+JVGURjfswrIyCUotIzlzVYZ6gzoZwDXIi5gQIBf/gI+KxNXPaKV+PQ
Ufys/12rjO6aI/pPlqSm0hCvftmBcnezN2hk1UeXgOIuKZnogjOsf0iJVX2aOOWE
6pD/psybjbnsNB6kH5uFTA5frkzIzkzl5d9+YDm9OyC+k84E83I/7/j+rk4L2dah
QJOvksSIzN867/4Qt8qYTQ==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="MvBXkzurAa5VTw+1JJ70nePUfoQXBvZOku/SMmg4TwQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
oRtzZL4VJ4iwysPsC8SXYCzXS8Fw2gtZTOskLcDV+1B9Nzn1zTyNtlo6lNICRmmK
ZRVu2BmCc2G+fmzynYlNTnSa7C0Cuel6FYpxCBlOuk3OF2tzAmLAuDyOH3Z1Yjzk
a0aHuoCdIRKv7BrZCdALt03JeUmXKPdOmIlkVGFl8yw=
`protect rights_digest_method = "sha256"
`protect end_toolblock="Jn9CQpRhJt4rnzZPRk+dOpzAubz7omckX1MrFd4p81o="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 21488 )
`protect data_block
gD6l00tciPUa6pDNTk/+t0OO0nC/UTtBwLB41d4inuAUA3i/ALrNyoJVcBnAmEQW
ptbcNp5fxEUJjnOxnedyZEuEBxWRieZFQnkRdF269oMattoASwe7rdT7/z0s530p
crDOKrnij5bic1G6A9r3P3EBhs7Ojf7Pme5l51mcQbbxeXKOtHX22+3kVP2U32+Y
YPcjNc2CEE5pemfmN5uXMy++bfWy/ZGKVP6P1PoJpa8JaixrdT/v/5IxmCvQ4pM9
J3C6lB9JwawpyC1mvNYknukbHvQuOHr3MfhhADQP9+hz+aJEN/3fhgxpj2gsrelM
vJ/NmfsLosEXMOneqkA4Ea/xmU41mUCnRmMDWEIxFHeE8n5KnLagheJLOaz8/5pD
fLngpim0G0aJwus8cERkPloGsfJLv3rPeWQsEYNkXXn9aZMiz4688aPoZoPBjN8w
c8m+AtJcBnp//vwio1oLCxuMqUEoD0465qYs65eyzlGXZMZZ0E4o2FuNFDhDvfkb
gBqyww/6OxBgdM2OyscpmzoZgB7vaoNHABZYjFBW9zyhaH/WP7uig6Xr6epm2Zzo
tF+fg+BGuTmp9xc+YENzz/f9ELpyNsAB5r5HOfHv7CdPMUZbgQWylF1uXUoUHuGG
AJOu3gRXt6Bs8i47sW9H1pFk3s2mmmR3nA21olUqWgKarSNsQeaEO6jLDTItmf9W
gkLhwEIDg/4SMJOais7VHA94uJY1EkTbOfd4tNrcqmbqsWPAdKfwQv4ZssYD8rdF
4d/lo7BLwQQCcF6xMhuFx4xqnw2tntb2ahmcSgUNdjMeatHDh9Kpb4CiYyVz4ANh
6JQ35liCGgWQvbk8ltHI0kF/P3Mo+uWPZ/qrgD9EY+B5HkKzJShNTXo5a7rL1045
FdRvkgOMX/V6/Z4zwNBxcMQxFui4wYmknz53gg5Jml7KHOriij5KlEeUm7fnKUfe
q4P6XCHPaqZ1krrld6EtdHVvxnTHdcrz5vivgdNsMzMmaNTdoUhVx9IRWe8dUezb
vYU4sCOoeL3KvKzKJrKm8U53eBLlug3qujAO6S/sxBgftsG8GofXNXwGozubmSeS
iR+fKtblJc9IXFBQe4kyWDwqMDOxbBnpNsb9IjSvcL5kErdkR8opcK8Ien22ERhE
HmvkAhWWZ4IKfOvWTOuqpD9OWT7O14iMfodDNVKoti90GIF1NlWYsR7URDRzq5wd
Droq3oPVSkAzgxojBHTflrcbnzo+knZWCoYrrOHVlhl8YGqKwpnrWIH+Qgbx5qtu
RZjqkIL6R1OBjQSq/mG/qL7xb48hIyIhdQPAuHJdVF+qCN27u594XHp8StjA/WMc
rsTer+ZtgWKhrTAQ2St/7tOkV1OBJIgfnmoGi1As7MZO0UnN9wmWSSM7Xa/N/aep
jMghKbLBsLmEwfDtnloYVNAkaWL5lFy7bupRfMJX3S4i6KEp+Cq89OWKqvgZnjwn
u2htn70nCQ52Kt9IwxdTv1VkzpxPkWfFHNVAoe+t08plMuFhq9E+FO4Fv+BAu3Aj
I86AulcXZpX+NYqAbzevGcWT7aiup6WkTTQZhGShKy4vZXmIh8zQ8acbiTQYjtaD
jSpf8+ZIm0m6mWmrz3jybHIXT1x66LyxJX9/lrlt5gzxqk6F4UICCRhw3bE282E3
2meQkc3Ebvtfj+pd/X24PS3kfSFLBPYlIY5i3rG06ZpqkD/cZ8Os+Q7cRkk4hlfC
ze2HIyKfvGhj96qjAPDhU3xFAf5dBgji+YWkl4q+/HGP6RncbDDdWffjQtt+jMHE
B0lD7Y+s/SC3lRZhiPqHleJySH/XMKJzjbzi9FClENv58KJgGh7oRqIFutjNSq7I
JVdlK3sbZsEpDsBphjN+Gv+ikZ/ZXAX3KMafn8q/EUuR34G4p5Z6QU6GXPzzba7T
c1ZazdgAx3Qdjl3YOnQ9BzD9KlgqliyAqJcBY05lDAoDRgYDu852YLAZg6VrkiYB
H9xItrwnuuCVa6FKgL9OdY+aiWf01KGd3SxKgGZGNnereOiKWlAVi4mszMiVYreZ
j+43eoBRzLIGRq9FdLjy9yZZvm5dJH3VFys9DOXd1zhFvUB8ivHznEzZlOGuU+ql
hgz7y7t+WMgTlhMySAGo/yfNMvgMXVSLpSrtZxHpPICw7JBXuv22TNpFA5tj61ME
GmofbQs5VtN8oZzlodfIhavpjyCdqvJo+YQ4oSpreZVnQ3nyhBA2Ln92pyI8mcmd
XYsewUzUHjOCoy0r49AKgAJptAQwkSALpkyC7/LSs7bHPwzexHgbfY0B6Zb959qE
tomIFwdXTziSuVraSmnFGooAK2NG7OBDMLqhpc1zpcx9jsxWa+ivnEKoIzbsxU8O
FeECrwg5wpBji4nj3Q/X0mNy4t0TulrAB+gByYhqV8SAV1kemOGRn7xD7BojQ8eD
nOd6dqiAw+ABOgyY6kBTpEgIRbezs/GSmy/qlwJzAImVLz8vPAFbsMDShrGKznbH
/eEC6GTpyAhkvReAy11z+J8VCO8wzSID9puOzKE9YoZwRRzvbA9uhLVuOJpQ5wVC
P/2ZJnNgLPFoNaoOQVxUSoaAvij2C5LXuHpmI5ZB58e2I4fu2xSIKZBBjv1omGBB
bKCcxGmWJJCT96cHM3TtI+l9b8UH0xrIZ0DKjJyXX0eBznbcxPeDMuEg71uF/H3I
VSTnhVytPvXiEMh4ZXpHJo9Y/QK5iqYDbhwMSI1yh13kdBTcnPByaty2tRakWALu
X0wqkTb8YuQWWObj3Tb4ODJPoKJyeKk1Xzw0ptZsjyBQDgfqHqndEIVXya1GoSjK
3OMM96OASGUvSzNTDH1XDIja6D2XjIREiSl03dozosTX7HBV3WRk5HR0yvjPlrkj
zcmYgCWEs4u2BXLlrack0kYHhQe9BKttQqSHN9kbc9gYX7EAzMTg/5t5CBGaV9Gi
R+kSjzdXKX4vdJsJ9ZHxhzeaqwgMTi58TDvjHpZQNw5MvI57gsV9XEH5PwRTUuFH
pEOZ+IqAY24BEgLWAIb2WHmeeMph2rE4uRW9fheno81uHQHmUkfiI4wIyHB/2Odf
3I22/+aG3zk7vSPJvhylJktqLZ2CQyMfxYzG5VBJIDWpPDhWKp1A0RQglSQlwmIq
ooQPD6nHisLYRwvX0g1pR+DaggLOuvwS/lrmJmYRBkBqAbnKJQUAMrJvUW7AeWMv
W+cEPfZORvBnqYxf0/ZD9cdEmw7bLTuyYBjBejrJG5HBFhMHeKkDqouoNl2p22KJ
HEwOUg2LGno8TcLhQar6bXjrzPyfuiVynqhXmWzTWd/GQ+Hzenl7Da5O9XQZoIRa
n2jP8xw3+KNAVChjNLCn9Vf4tJ6cfXUq8l1WwtDwMa/3r5zjwFGEyf3LB7U1vwmV
xJSKbR65hY0SzmjFQNTS/JCZlnzXwwVVB6/lHgvqEWvxKIb+celLDE0UNjSEA/x2
Kb0gecgLVf0hUeG/DINfIpsuHd7LjoHja9f39or4Nhzryv7lUBbBms50LYTxJiUl
HMlIle2v8RUawnyqIWJRZ1afYYvEfY4bZP6UvJORpffr1QHH+DKSCXqVuXZoZlZ2
9B7xFfEpdYn7UwIIyTBBEwgTPnVSahcwnpSslHtQ6/IE1K27ms+YTPP8lVrqfyB7
NFzhtvhM7h6AjodKU0+7ZVD5uhXFhfZ3nCLF5g322U3gvkWOTSMe0P5LTtdcNKAB
ghZdrHESLWoV57WpxP2eOR3sQWxr9CS6YbGgrJmvqt9jNru91IesgIpRIlwDTbff
P/0SNUkI6OFWjoP1/LZ+q56o21N2r7IGer4rZaU2+hP6meGAlPYeHbM6/sJUnnuN
ZWYrWrAhlUd7MIARFvWsptbjDIiayHqFu7lK7ZfLdTnEGv5ZpEMZYmwyp3wcY8Gk
YlPWwQy0sjgAxRtCeAnparrS+v/LkqLjXYmX5aFJuy3NUkTqFM7ZYRmNOhbi5/pK
l8Yj231LAKVLY9D0+pLLB0L4iYHGsN1I/CqDy1nP0xBrzse++gR2z/A8BPzRJmfn
SHahAw+twO83rMUFGTBRNHZiKTTBzGpYsi4PqqYMmgG3Kqf2FqtohPVfTNc+yhyR
CcpyJUVUGtZu7HXE3WGafOvh3+PnhJxIZBBY/rvkdLlqQUWORmObbiLAU317qCLW
NnLp9Q+ncJarzGpuBR8uIpgI2KQflIKVnKFI4jOF9C+oOeWJ49cHUJt/Uv8+2uKF
oIzEIQlY3eM+zS6jnImsBMk5AeMSjZPVEp7DhXKs/iyXyHYars4bfucreQB5AjBt
1W99PW04F3Oi31z1mLs4YLCl6uyx5SUt2QDZTICE5nIGOCq6M12h9uv/1wnY7LWx
TTDDNVsprUpSvpMdnO/0uMdiFEJxFWoeWuTU14FIgYGCAtXwKd4c8bsbLeBgTjJM
Jcwlz2NetjNJGVXhXuaweQDHNmGOHQtX9k0qxPs6b9l8HGz4CnK+yih4hi44snUT
dV8tjffUj0dL/ZfQnybyt/o/hURqNd7KK45qsakyWf/Pwy8yfqboKdnFhSGY1xAc
2ZT0R5+zcgf+u+ffXbVGARI7DqMJh2Ux142NCnZxxiJtHjI3W3g2TngvGoFnHxGV
O+b66+X32d6Sbc1bcSvoelTCC4xvCBWzx7CeK7wU5XeqyDMX45P68Uq+s7/Ou4dC
obEqYwZfLQ+Mc1eBMSOc1DvEWyH91JVsd8R7d5WqxtzcSCh4QPZ5jSo38PdQKtM/
+y+MJ0CFBlKtYdy/SrqcCyhQ09/cdypqJgYuZ1JVfQ4YUo/cA8Y8REeLyCX/Xgeu
h8I12yjawKEi75o3fYREPiSf1KxGoy8vVhw9Zcx5AmEM/s7uTJmBwNnmaS/tGalw
g1RSLolOTfAVzsgwuxkzKVC6EP2x/xVFWb+KsnsOkfABt4fVRiC5HHcQHGSBtCXs
eDC1G/FOggVOQ5+mZMJuqiGLTvHjyMz8otdCsC5GMsorB6o6KddHDGa6HBl7prRL
A3T4OKo8O0kWKQE+CY8VJwQMFRaASVRfagzAYcL3qiR4jXvlCSOhDu1cSXChC8xV
STlfX1EC2+4fOcG7WwuAtY9aU65QJrCYlh51ClTR5/RxcAUHJChZlmKcuKHX+pr0
04ribSGQBBDNHjEHcvLl7HElQYPhUkWMUEkZq2T4oZoFjhP6DKkL0dshf3rEQ+wZ
i8z7Bz6MBuwHr3PkA3pDY7hmWGDLiZD9CUEc8H5g4qJClZRPS77eLY+j4YOTPhYV
18tpiVXcIV9VVZ/ftvVirQnF72UEaCVRZu4a+ilQIBlbvKyL2dIROfbrsa13fnbD
SrSIm98oz1BdZg0c8hLVbtLluUS68iWXJ/Qfy+lISsVHoPzOApauwY6Pa21E9lGw
AWfOdI1/fxZmza9CTKWDzm0IZs6IlBl1wkry93kjvVKl6pOJXj+YzQ1v/s85k3Qb
SvOG9E1oMFhI2YrsQytB49HY5/U90bprxhslq9M+TRJhftxJzbExw3xVNQjjK8Hf
Dl/QbB2CS3IZ2Ei5HK7btteUccDPF0dlQD91yLT+tTSwM5J+EK8y5r6vzoMtEn/d
VOHTKCnFCfeoJG0oXK11MjuaeCZ7a8AmfgZJVd3UMtQFy5OTDDSulkUZzAzCwEwq
EGTOw0mlL/LHtD8GVx0TlhqfTmVHgAK/0FAtEvjhMXQfdDBveYPnnIM1aelmjrwm
9vXoog6n2Q87lGi+MIrFjuOZWayZjvN2PqmlwCUKZ4k6ck6uDzuNUEXAL3DgpYOa
mYCSq8bql8u16uMWiTJ0sTpcHssYSk1SnpGst3D6gY4QUCeVis40FZHv5hmYhDW8
kMiGLr6d6LuqvnzEheNkgj4I+DxxIP/1HcUZxpmzcTtW6fUjHXbnTLpqBdSjA+UU
hlwDW5tfvPp4giYbckV2xOfl806hgjDHkLBOo6e5i0ir6tdEUY80RM+kzv9EIk0L
MMEnN59cLFYp5QvW+Dm1RSz0fFpedKJlWNnPCow1AZEG3vkN4evQvlqclJVX6SW3
YZSVrxEznibrL8O/qeq/sscDBqKMg75LRsh00e1/f/bs7PeULM0XHSdC7Fr09mh0
Cnrws76a9rsuxFhI70aYovyl7SQMgdq9c2d6GsBsCBYrhxZHtS7eH96fUaMQ3l59
KJlq5YFDXOoegecCIHjo1cpA7WJUc96cnpa2OjUsW6UKU8ucW7t9Li427HoP6bXF
C1DbFLFmSS/0MbtCtXQFv8dPDrGqPxA1VCl++JPNOxzd+k0dylIT8tgiZ/Y8Dnnc
S+N5qgAN49aG+uTNIANB82+Tniohh28UUEr9a/d+joRntyCp1J4bsOjmiNc8QeIA
4ZoUg66QskCys1YHHxDA6r84BBs6dlMkVHqDb3AzGX1sopvRuFUuScDG5CiGJuVU
guBuiBRomyDUzw1sWpVv+SP2VSaj3fvCLvxJk78dqfzC/4QlzRybkeeDEyVRHjSu
QwXHr5ep2/fB4twY/DrZ0ZB29WPQ4VU1/ZfrqZugnHSfQSHxOGWl0sZ1iIzZnnmj
GL4wPa3hIclEWJ2UzX+8LS4y4Fs/x3Q0MMUjhJGP+wuJbQfXuS+40y+jBqi98zKj
AKudqLJsv/ihwRL9YUfGp6h7iF9FtNLFCTYEisC0hcDZpWkcCHSLxxU/CulQrQCE
JMboJKwyIvAop2mADNqdfdO7Zcwh7kt2UQgiBNwscH7y7FCUAEaiy65fD03zVuVZ
t/VP0NTjg/j3D8g2BzB+WhyGTuT+ZW+8HbHqqwYsCeDe7zAJlosXdOsMkNK9wQxi
LlVuDyvKPs35KljtBXntAmLy0SRDGfQ4ntrQP8ZDmIIVWEqPKRcEYLXObmcuB9XJ
vA89lWPJBigojFcSGwyACvqcdVB1JlbMKzNIhVu9KG6h48NGT6GxV22wj7poqV2O
/jtSvok1kWdpy72xWJhSqgbk/o123MRXaaIt0oGqqIWzFxOsk/UR/8WhoV3fc6cm
tT5IeFZHKMotJcBNGwRHDx7caTgsLzwnxzkfKhNn+JYO/fidtFMBDX1Yuv8Gzy30
YkLtKZyuQu5Ywqr9foKe3vuVWHK6rOUCi3K/takW90I6sDgpQwSG49O/DlWElTs1
Sz8STpApV1jJDrG1DX+iOMQjjaU2NSj+Jhzn/A0CDUT/eJhMfHRlyRyiAkYvIGFt
J9F5EeNjjuLB39yJ4ZNryjT1uZPN4gbt+xcur4I9vLhovZc+nYLUkm51UWdmAjV5
4P47ydsjEajYFi/2Pazk0OIpGEBdRGy/cAuX7VxFtPvi7NnWIz8EMHbd75O/Hbk0
TyrkUa8nV8vZq7E0kDSpKBT5o7coZNVa+QRMNp1j3CBDBgCEPsCj2F79cfggOdNm
UN1yIBgiBZ4ZGgYcetOjdfose+ka/bMn7OA37bMdTB5LrxxYAlVFVcepPvo+Z9Tz
hLqpPSm06lfDj+5YgMTzWoRa0hZSygPZlxWZP1+p8Xpqznq4gV+y2KrZsN6Z9fWZ
MReZS/e8TkHOAgaCOGbtWKQ83CIej3TxYNnEwIoIa1AePZl7u1RnUe/hb1UP0MsM
NvDHFzSNS0lBqZ07qoTUxMmjPxUMCqziO05MvRRugBX1s37I+1IbKmiPPXUTCgtS
HQpts07ACf/PWSSzSxE+SiGKCTSWdgiV1f6AcPNmBx6ZOFzKboh1yzFI2/WqnVDW
i8z7aS5NpePYxNhUs6Z+hR6QYFN/B+CSCFPhDF26ygxISwAoKEgnVdLJ7Nliwxa3
s2RgMlTpYrOSxvinXv0O2uK9BRK51Kw0L5QFn50CTcoOxknYyUlZ6pA3ut4PVtdt
xV7gB+U/teA2w0AGWjUWDuYQk7zl4C+KyvHN/aa6jhyNT257F7ZMjdWb2JQa62dM
uDOdMlXMoiXvE+FAVBCUYJMrG/5mzvNBHwEertIdKbQgPaiQfNnumOtz7R3/lGkv
8T9yc2I9aDOxdmn1/mkslpJQEYIsAs7hzS1Sr+FjwBDgb1edZGn/sfwiPZxW3bi0
izonxOUAcMZNZOGqnbcrX9prHQB6XiZvsI/fC0Er5dKQPA9TjrG4c3EW8wSgLfDk
prL+W0u0y0EN1aq1MzbcDRwACGOWLsppW+009S6GBAdRLunuavjLkxf8nN2uVbv3
UFPU27Y1k6dnLWVDLP+VcwOgWH+277tNpwbHpKISsguPcxVSmz8DcgboNP++1lAb
NLm7zSOQed9Bl9qlgJrA0KDuKd2zCz8AtqYXgkPS5dslebZ3PsftLliXbNJE9GOJ
mlYxeayEZISPuWQrheWFril3rhYqKEGiBWL0a43yl/zENzw51rv1GhQc5MstTbZP
OryUTWqtf1oLiGkx4D8of+QjSPklh/jzQILKm6EbeHDZSwOsTO0/dUpYpWrMukxi
tmMP8lBC1KAwyooW3b503IdiJuHd1iCE3FeQZpfAOaPA0TOJT63fe9RZA2/KiArz
R5Yo9B2dR8cOcVg4hiqkxEImP16HQwCzV2trircSk8MEuFZ5AO1wherreQBl2QGr
IIXSH4TTlbaK0o98IfqwTmn12ml+g/x8AKtMnQpS011pBJPZNbo8kVsKaOltpCXs
comIVOJDMeN/1rJ0l3x8nLhr4REnDDP6iUGSwQZLtZUAxy/7m99KbxeaoSNKbqw2
3k7Evnd0eAM2zv6bRSRddqXl5fcfPaRbrlKVLxe9sjm0QAZgpbjsjf/9HrWwY+hO
T+mZQHyzt5FqN9GLh0uK3VTv9q1zdS89khpny1FVNyHVK6/gfWG4Lne154MjGD1Y
pblLrhMxGWCclAlyerxWte2TO4RqlVf1QbS5wrhGy3lYf5bP8piLpkme9NPt83CZ
moKs67/r+kNxlVGUwT4/Lam7TKeftHpu5pop58lZWCnXQ5WPxpQaq6+mh0hMhgj2
MO7O2UT3IevW0UjmNcgl/0gdqIuTlC0XgaOX6j8Ip2dxyHWf1B7uOA1/Uf6TyjRa
YJ5Lj+zTB8AlKbdHgvui/XXzZbl1UdWqkotK9+Wmx4hucE3vhmoe17lU3EvIUbe0
JaCoxWOGh1isQ+HkMVGEEroymX/5PyUrMNO5lIrQC5OEIPyDU8VZ0pb2YGuhXXj4
9/aRv704wAsu4CmNwnG+ZR12VhWT4K81i0dDnfmb05Uj8iTWEMJm4ToHledP4tPl
A9MsiC8Dx7Xbgh4mYX6LkAz/TwUc8MQQ88a9Z2XgcIf2WF3G7pLfbaQEl3evRk4D
jPdnIOBQPT5qcd27IJmARpVne2dW4YSCJrdSkKY7rilAqTLxwwTLEC8OoanRfZ+p
/B4bSr222O9jQgo4bRRn5Hr2SB6zoqrCop9uBpKCuafMnocLAcClzclX6AzzESVS
MpMUufsDUujK3hqATfokenpRkAfdoKaVpyOxIXBU0VMAMix6jCJK3QUMolimi+F+
x/F8ZUnOYhUTk2qpSOMZVRP/qqfpj9xpgTJHqhQJvQM4KqXZPqrljwjaW+LDhmWN
hKyAbTmnVnKSmE8hNlwCabBd3baYJJKbXQiUGoN57yBTzZ/gP1Emp/+7nkZCdEC0
Sokgbn3B0k1ODoiABGGA6skYLbjbCyEH33UG/CGyoDvpmyX6E8NZUUrE/1JnUNx0
HYeDtA+XstM+NEx+UZmPY7NgUrPrEFWvYukI8T+l5vQXr0d6/tIzMjiXzPiR5/dB
xugZBgtFbnArIHDglVPGUwLrFmSci31B2gQ/OsSb+YuF9t/9MCAfCvDhUWaYsTOV
mj5oQTpnxA/OIF7WnRnX8WrGJOi2b4YKHpF3u/pZu+tYi/MSnfEr2XAHxieMk92e
e1eCKjD0FdPofnSLUGXCwsEoDMP1OsPH6/0vW0TUKwhpRxw9zCvhGGRq5Uq/eh6E
394gniShU62OvjTbBCJC68wBuaSmRQjmeJhmdxQd1ip4MRLV8MyKJmCjCuEeaA/g
+M9FvMM5CuabEkrHqIQYS09Ff0+VoF0f7wy1ubP1Crz5+CqJ6Eo2nnmyb05Xe237
VVWAMviyNHh3Fn7nY7vJ2Xw01WoZq3x9EeZz4nqD69VKtTkB/uc3/bCv/3vJC1R3
f70gfsNQnPdhy4mWtGpF+7g4edg3nlbuSxG5NXXXzvXPZqIRibQYlPTCTIbKC9O3
fwTFpgDOdpTN6NWUHUGSVZL41x783rQX/6Gb6dJG9fzroQKy7A5fzGQJzx40aeXo
Cm3a5L1eI8lqlk7St76kk0VTNfKSliMnkqP4hN25TLk3AwqbavSDxywJQ8NoUCR2
pu7UJL1dGZkJNoiNWb5tdmLI7Ldx2uAOesrecStkxiwyyPLKLTPtMS1rZ5z1hVz1
OmGKhB6pvmwvgIesvhXQPx/IAcANknr3BQo7ElozWZf8358Hta2hthBmNQYryJ+F
T+6owAHI814qqirzdGd0lcXMpT7S7r22TgGK56y7xTHH+mifSpbuixAp603iQ5J5
lWmkEKVj+huCLZ/4jicNWZEMekQy9p4/mGhvVQmVr1DBS4FuURGOATLezTrkeOw4
crZi7Z8yn1tBba1S17mZ7d5VdL8WKgfy74IDKiMCKZPJfVNpHRerZVIImwfkZwcP
/GNsjei3L0vhBMOct/OeSBRHViqkS04kwM29V7cmuRCMtFnt8/V/ykvGTSnpd0Xr
e2iP2LkV3nxQdJWJHgD+YXNOXDHjE7aP94TpRuL2j0favWGltwMSupoPkIB817It
MyXVNYBHgjfZykTxTp706wAbtk2h6yh5AfZG/68YA6MuNFJUY6lNLMcGu19Ad9ns
f3ulS+2UlF+t+mmMQNMwRY0he1Lmslxw3A/vIOvHLdncLSOW3Qh+h/gVXAb35lH9
0VXUaRpLw+z9YiaBRg0jh0INAyq7lbiiNZMQWwwcx/Y7kVT8aUJJn+lwR7WVDSj9
fmIpugbaMSvgi3T5o+jTVI+mhsp9n8Ig3xaqNCt8Y8jcVw3HhmA5XGzt+Wowo348
3AZJHyGJxD+NO4NJeZJk31doqIOc+MeKJsEF2WZX9HZiseggtT0NFG4+NI1GOAHG
78cpDkbpRwP7jxawuN/jTbdFFRdKGTSyqcG7HKDS9+6lY2wrR3LNvVrF0Tkjn5MO
tsyDr0upx+lKwEl+hJ4T0sOFudXUwD1e/TxUvkRG09fIFd3LiLYaCT1FNjbEnGD2
usJm5ver/GjVrgAma2RKs+pDZEmSWIvAnWwCLZYLos+ASMGOv4H7b7aoe2UFlOCF
E6UzrTYpvVEoQfvoz1mYYeGl/GSano22IhF2noIV0XXKLuX3wC7/elLZ+1k9gSDs
6qyZCmOPDAb+tAZURcfm/4+4SMD+foGs5MqQxxfbZrLGgzxB5Th0Ozj3fTZcySpE
f5ycxUZB4jEEXwUJirM1fPDrWSWr9e7YBePOEY+0L0IFdiK9Aa5qkr2jCjcf07Jf
WxfQMONDSJvd3ytZjTTzYEn33eXcEMmE8ghNi73ZYpHIVnfso7739idhd/6vKGag
jPbWAEwBPmmsd+K3lPTTRjLSqGicSQLPV3LCRMYpS+93NH2xvywYy3LhNK4L8T0Q
xgzlmo/B32R/AsKfM01lyjVpP9XRPob1RtBhK3idQsmwxGLztTMpOKXZo7ByQ1Rd
JGSL92+/Z+OjbupFGa7TddZpTvlJATaesmpvyQfxzYl7JCdM4kVAmjpWdIAi1C5W
a4QFH07Wjzs0xeiHoRsT8DUWXOk1EUG/BeaeS0DDo+Q0LqxSu71OAfn3/8u3aFrU
xD28koCq65LU1/wTb5eLNDoibqOsw6jAZl5q+uj7y1vIGvCj6k3F6PLp6HfGvKQD
uHw/x9DXNyWaiNbJaMP/gUxx4OVXJxs3+xXIHUaK+lG/iVw2QQjMpc31zwCO+bpE
gefsqZ37iKNcq6ZYN4orMqqnDvM0Gt+PPT1qdpRL4BG1usvtde+esD4NPmVMajMn
Kk+YZYxgh1+xsX/l/N+ibPhoUUokqtI3VuoCk7WHz8ZwgHAPrfKRvF410XXsyb5q
Lq4ps7HZWAiAseG0XrPFt/U8lFevq7TjgHmhYedM/k5lfrXUnPcI7z65cOdc7nmZ
vzScMi/xW3iBrofejBpH/a58C4ODVW82ATXl2G5vZCD0g0IPVJc6V1zKIAIQNfuO
Ra2+RSL3xb5mygf+bDBY8dLBH3hadxC9kBsxC6nalBS+hEVBZryjxhTE6TCZaKV8
KlB6Pq9zaSu6R+IbmXwkxkPBS1LAaYttxWO1urb7YjpREytvfqDfFI/U2qKDP4/W
F5G2pNyUY8I1wR18bCmPNOPypLiNUlQnT55sVbZnqCeybHRdlOtHPG/AibPNxtkN
s8JZn229Pj3RJst9nIkEeXq7XaX8quWPJNB4BpuqjDAwrag0OPi/bQYU/49Pewgs
3I42jvG9IccFa7dDfr15AkLQHxqSPDrQqj89hFkIR7fvBfimWer14cm9gRsBykkp
0aVc6Lmp7MH76baYWNV/9VlzLVPiGJlWnczszlLDqlwGLbbh27BtybsXaQvs0+I0
y3tlNM3y4MwcfYS7dKBfdCMaY1R9mY4O8HrtBnxRn7Zckg3+EVG5z+aFPQ/yAVoD
wkw7rmjbzyKkGFcIIUy7zpVqEfz4PlqcYnIvl4YvQTzYDKzITJm/vfluhq0sXkR7
RIvB3+ovAaAA5LIeHmKN6d6DbyGB/BMqwdghlidzpAetrbBxs9IhzVKHelrmqjyF
0IMPGH762pYpDWk05OwclG126Q2dJqhyNnQOOL+8yNLDJKNJRTHUBYPFhJGUyBE9
s9NbfC90Z0s4M7HP5mnkmAW/bWVHs3Rve6Eu2W960HdSit7k49lXX26TxMn1T3Mc
S4Fazj1IwxU3DWq/D0yKKsuSLfaqGGZszGo98VTFWhS0/ogZweityCLc0rqEVh3N
FRZntfVZhPhJOM33O5S4CyGrD2Q4FlWt6SjE629oY9aI+Xn8KnZxYA82I9rpw45f
nKKR7C2WpJ8Z+AmIcXNWedrCzxih9JgMtOVQAi87TP16F91KbRNKaG9JQCdKqRQH
G8FB5G6GWzYIYadGr4m1j4MCiykqfSwO6Hg/U403/o4LkRutPYmdqr4rSRGqCAiM
z0hQdXHhEJuPBENHLAKp8ToD1xaYKjEcGGl9UdVbdwJ2Xyw6cUDedc45q9F/46vp
jz7pvt2Q2+cOUojL6z+u0rD7gDRuJ4SOxx+LOsryzTTEgDLVLgcP6VlXinrtHqEe
XyD8An06ikKkpQStgt8GDUelnqz6JnHkfVf8gic52GAdQNpTmp9ZNAMaQKvPil5A
93AIO/Tcgs6++aaMNXcB757xuaXXNYbOE/fEI8e94l888osM7sFMcrOJdQat9kb/
5s22t5wbaX4viSIShhRqKZ8PF/LKK3QJ2aKnLvYY7eLnhgl9BTv0zZv13SExYC5u
pA3zptC8i5qcbQkNxKtVpOjpBt8U11q52dxBvglFTe8LrLl5jmgbQ5O70CNnShua
OJkpeE5In5VfXjdFMluITmnNmbbu91kdu/LSAs8i02ctFFg/wGAls1aupfgwTu3t
ismc4XPkYQ/aQ2RQE/6Tlid9nhISBkBzu8IVsWQZRqFHw+TPLoqkI6X36QuBHswR
ret2LuRP+uprmrWfT/4XHp1hODqnCMmvLwy4ilQ+rqCnQtOaaGgBG/dCE14v6IpW
uLncT0zazcejX/tZbTn+phj/iDkBtaTwFz42ZH3nAhYBB2doo0lY2xx8obLz+8hX
gtwCpWqHkTgWgrs0AGMyTk4DMLSaBzrtFrNfPzFF+kljDYvVphkob3NBbi6ePnaA
vkcUqhvSFZVKFEajJr3nFFOekyPexbcwXAeSiacElF6BhxA9sQBvC3Re3nx0Q0qK
zW/8qOh0UHNx0Kmn7XfunrvOtfgZxAuDfTFVkcs1+K2ajyj9IoymeHKAiEEjxQBR
L8PMgcfInzJNIwCE7//W+Fi8UEs+V9mpOq+aKyF+pY5KeQWSXurfsC0GMZpVuUC9
wUrQoP6top9ck+a/MJLVFE7oqgD/zvgx97s/OPUpeEj6+S7rMoJbYLZaTH2WwSLF
KenwbBEj4IPHmRHbKLZL78rfgpzfFecpargjWoU/ghG+uUEZUSePHhAVR+3wH1+5
BObiZWpqQ1meVuZ6noyTuFTEvV2oJBleoD6kv7mzyt/uZwIdy8YmPpI+0vvNCoNt
t7lJ7ahmIfJaaJT8gtySxYnFMR45GjLM55RpOuhTcwxOECZifGMo54x2HSR7i1MJ
Oqy6vwbpBfpzO9VBDkRQUtaYg3T5/Vvj8RNvMbMGsqutR1YnGqRIzD5uObOCqnKx
sY7Du2YVu6Oj5t4fl5V0AqNHJZQ+lZLUWDAfWwRwtmekkVMiiMgH+1vh1qCKIC1f
yJcdOVOoX4FTnwPRektGb8G0kAqw0BBgb7u+5LYbbtv7L8tamcSdKy+eaV4brh8i
MVHeyknGDjqYGsW+ULlKgmELiI9ONsl3LflO7ZP249x159J98omKKnm+fi4Xh3UR
aIaOpEYtQobVBLrFo2CD7oKDtCqvo7KYAzOMsHXwExe3Ko0Zpn/Dbq9HP3X6xaRr
JJ1KzRxb724fGUsRZOqJVcWIVfWMRxH9pAlp/oyFE4K+jOuTn3ify/P9dYGjMTJ9
1/hU813G1v/3S78H1MQtHzidN443y3T8+W7wx2q7IoS+Pl3Mr4wBpe/RJH8exFPB
HN6V76S4+KdMi5CE/qNIHRC/6eNsv/knOCZUPInwSlk0g+9A2MjKOW9zelfGoU/9
A9gEUlId1KuhzMOJ1HbB4LpB2P2IJeT52xLnf+vj949fcWB/kyAjBwz8jsZC3zEB
4OPkd2ARysJNnl5kBvI+WsAPxLQqE7fDDa4mwakD5WlT467ShDuSyz7J5/2jxBVt
beGTLqcI8kVDsHm4EgC1jrCat1qqQyQ+WWVI2h9/OqSOgum1QMfZqFVPlV2jXDkb
oLvqW1PIl/kLN8gwxxul37+V/Q1hhBL3zOdwvirQU5Un424zYubV1zrX50IMa9yC
dNNGBxHoOUbBVsHBp+BuRhRkH2yS0tjjkvjiYVxUBSvG5gkBgsKuO8kg6IWWBoh0
L2q016SY8qyP7SawoG0biY1QuL3aYMHe9kNdwypUIZmWbNWPEvtcQGi+5HHRcWNF
7118DPm9FWjZKllxe0z74NWktXhDa4WQJWdvbMyI5f5NhE7vNOWxAxxGm91uwI3W
BRE0cDYlPeS/1mWume+N9w8oRSCIrNY8J1ROPH38Dk18J9qjiX32/882WWpu7ZmQ
+hhNHZqEkEV7kDbeJEXUYYJz/tcqiDbK4+Ap4AlAiGfuQNIbjKHXqnl891eKi/vf
B+Pk8VP5ZaoNP+yMAVzEACPfS8p9WtYDJflTv4kaB5T0yQzxLaxmNIA5JF9Z2qfY
IPjmQQRE5xnSC1x9sJLf78QPN+H5om90z72odWX6a55yF7KvQWnxuJ0QBWvTLZ0m
VDeY2ChPc11zXzKVPJuYRKbmrtyWD6BRce3OSQ59R7BQrj/rYLWIarKDe8ecYzn+
h8vdwJI1ajdnailKXw56RKjDrLSHVpnewO1w3WcToO2DhOWHPTK2Oy7L7NLiQ80V
Pp9hN1az4RXlZXGl8zu7DUnL3N9k8J7g+jRARgrAn4LnTVAAKX9+6fEidQGE6A7y
ctYv9seu9JE29oF0NpXY+u+8RZIiL9JTmlr0Im4T8Uc4hGxmr/Z1FSiyvebctrbM
FTZp8TcepLVUxGsZl/DUR8Q8rgyzpms1+qVbhxY5odlMTdTwQxGqi0SCYn5wnGAw
FQSAQ/R+yaFWVR/YgU1RIyPoElJH9h/NGibjPlAxms5w36LYSPndC23hzcEicK3x
zIBiZqN+zaYztXoZwUD1zvkYVAEF0rG+EVfJ93fdh4lULw9HWlAc0fIOFgRqXL/A
ti3crO8OmxfWuXMe4nm/EJDPRrLjyfn0uPvk8TINN5r4oalL+C90nv6uibmUVNZX
P0yqusUM537qsqi2QxUEuPrYgTdmean9hwvRj82UdG2ZPXcZI8csHud5IewxT+j9
ZLR7VwLHHW7QiY2x4uxSMn6ysj34BnTaeEjoS6lyydJCQUq66w2xXAZrxPeWMWzT
Lu+09xZ6W0KeSbGZtokEand1rg6TUxg13uo/WxZ+gFK9h3avp2DGVVASaqgIIvVj
CP5hXWcVg76oiJUc/ptV3n2geaC1hYN+F/E8XKI/HoAO+YWWoMeNovOL1OXdZovH
xci1sT2ZesLQUXx6UPFlQh92G/PtAUqQUp6sKgYmuxQdvz5ixMboTY4rwMCkN2C/
xZuGXe9CLy0Ixfhk43N1DZab8RsfNzhKg7e+8Rd3mKX6tBmy8T7cjB7XMgszMrJV
KJAcHOpUxMKnvbXWrXLSybIKApbhnln1abSXOyB5l4+ryZ++Eu1OyH78yatHU2wA
EsCuJxFPk3W+VlFLIGdDhiiDhCiIpHElQoE4LByElpBOQ3IhZ43ijTxS1upMuoff
HqrCYRpLWEbiADUzHQ13Zcl7D129hIQxaKm7H5lb0dOC389FWyB6Ll9nrGxmTi23
CVCeKaEawsPjaYxVTPcBj2CLYgzok7YKUEm4fapNRXhsYtHYwmAaDt+aW5t3c1KQ
Bo+Ega2lrGY3YVN8X1Mqrja2/9hIopfdAh2OxQvwNuqGtYXoaZRb2lv9drdTTc3C
Ua8qlCVnXqaGE0WQEM+0v598TqSgpIRXhH5Awz94bJneWx7zFcPBgnFxVqiwbkqF
ruwsHMeHcrcw/GXfV01ekvPv+V9/mNYsLKP99bToqnLO6MtsBK8NtQbtx3PchQxU
MKnLPyq/kntFlIyX4RFbH8+vSO+u/eo4qyFN0r1rFYPr2GieCw5LYDyE8o81NXqU
frZiGlerGdobkS8RdjWTz8WfVR4cvqSAPxhkVMosAzkI8VpOHd00/QdbSs0Ddx+G
CBc2cIy1vsjLB9LNYSB0DLshLIqbOg5HYmWpCGfNXOzrq2a3Qjs0sbmFFf+9kULl
4fRDN54S2Q/d3jdqDD4odu2LrcSDr8kopzknyKLwDMtowtzgcVu3WlHA4Qbh6nqq
v9UjP1g2IP7puV9iKVqfAUwnmjaS4VyMRiXUrlfSw4eopX1h9OWggQN0bt/6xf6F
kWZcWovkN477ljGeGEs+1g0egkQyQVV0ziJBoiiSci4GEOH/w64pIbWQ67NE2r8K
mwsBbIUgvHCP2yJlv7yJoYgzQiZi/H0jOOW8esLc/+iLe1En6ijdmZN4gsap+Kn7
IqtWqrWI64u9P8xDFBHjcTlKY+RtByyIQyy3QjdRflUTbLtZt09PRQvDSQd8oQXd
nbyU2UCtF5MCKIhGntamf8fTLJxw0athjNnZ8EOhkJd/pyyuRmXQzho7ExWIyvq+
IXShFwHg2DNrWF93HPy8oLbGxgfKpe0jjK8WPHjPp7TlfiBoE2X8OVhFkNX/uUzU
ZSZOfUgmIg1aBRPUYbgZEcFsfOjWj96jzM28/pNlEDT+FughGtYJN7VPzOJMmeHd
i7UZd/vm80SpWW6pdDLs/NK9Ws71VQ/wceC3zZbnjfx2DiWUmaxq5nbsQfuBSi3Z
7Q4ZVEuTHcuwrkjgjMKV//g20317jT/ATMZ7AfVi6Q1b4fvDZrq6ad5zwFCfT8Na
JLsJ2bM1ZnxfJCH9VRyRmNVOjDiuO7qUoGtPkvZO+ZeR72MvEpHuWp+gPOeWMIaa
prmZE+FH2Gm5ghyl+jyNQ6gp3g2DyI1DNv3tpJWn6M5dMUQKVqKl5qqROOlRAdNM
UhZ+rbcqhH0u2Tr7d/un5QYdTk0deVBYwfK3ot+qtjGxn8dTwB51nJeH1RCz0AyV
bD2KWIgUrxhd4JNb/j0wHF+oQR6xJjc/wUZyAQn/4ztHttpYKqCGSZALZzYLJMKr
SYdNaLIwagysfGygwrFDoOSCwwLVbaDVc1k1r4suzDRmbrT8Vdygp9sr2oVHOTTf
1aF4KBOMP90e1A1U1GRo28M0bWl017tk/BGfp2clBbBUUb7RzXYNFS6E8y5FiIH/
mIV+bXeV8bvtgQXqW3M4AS+LYdRm2QpazV1OXbupFUgPhQJvaPScHzQ45nVIUMJ/
MTW/lk3DcCPOCIAYfg3RGXochO+hC5JD3uY/Tf1PRObpgkqMRcARbccxvB9G5J+M
pIMGCkLfhXHegnl8gFkQt7WINK6Qe2p4Po86+PFzprUqrI6n7JA59yUdbhCa7bJW
dm2Orp22a574VMJPZxfX3wsFgFo650imRk+yhNR+nLhG38i3a+mG2vGRDD8/NIET
FBfC7Rwlaju4ok/VXDwLUxsMscdQRH7WFId+1su146qbH4vylGq6RMWavfIIsjJ0
xWJhh+jTIxP+dyka4zsR9tUhIwBwmbU0vbuZbSpkgQ9xofuYGjvIdsH20yQ4gb7c
kuSfIwEOkiQVLz59CaSKTLjvdQg3R3I3JQEhkiaHK/VuPyWtvMjd7LFPPhkqTT2X
0COJRUS3iWMrSiSUWWc0XDMp8wpNI880vBitD8ItMXdbqiW4vH/qd/yj71fnhDOt
jgMAJEefKyEri75jFRK8EG5Al53gaNCUbbYEFsh+7axivdqocNl+pUXHBTfgjBUQ
nC6sp98WGQ9GMOXfSW04AzhSooCfho1vKm9VVzeDucvw9nkDG+bKYc9aR8Aphbrv
85bKqFaUgYYvWmufGZaXiWZbSSRDLKN2q/GDWN9lJ/f83dfTJJco0Zx9EBPx88aJ
okSUUtyKU4SyE1Use+zjDiw1Ytbjv4NUM7XqTSp8GflFjDuwyO2faYkeVKD7j6Jh
pzgqrMqM16B6rMe4yM42N0J6V+ZRe5vVwzpVdjGpS02d03BXNfkkxaf4xP0HkHtz
tCMUDfwXdsLMqODFkrtWpa7614LbXB6jRstg1J7k+UGGyRO/+LWRmxUA/xYXdjkS
hpCOP7Tmk3d2gp+zV0aNOQJfvD5neeBTz0us4c0+N8tsnOkwyuTL+cSE7VKMjDsI
g3GwE++hKXaij/OwH76EGzxzCZ7h/mYfLEalGBEtV5tLA17sBIg/bzYYnIQPGHHz
Werm9w35/ITdFgR4NBPyV+vUmpnZvT8S0VIbV5RPPLT7p0tz9aDLtMA39VzaMwZy
i29Aw/b9Zsidd83PtX7LY5WDRLiF21+Cooh1J37TAndjCYZZ2fFUf9EjL3lMhGFM
2Y7gWxSdNRc4KmSJgjtw9rKDEdTr4k2qxtHi0VJQ+kOIoTSIvAsjLoi5lM20k0Jj
oMh1ViuvfEQPywWn43X3T6qOjT64fkpQUTgFMYnpRWYs6FS1EBTp6MGOalTg5Cao
j+DsyJIrkzCBQIElSREwbhRptgGL9ZMULWYpbIgbnLOApMEdxYzFY3bkGljmCuHh
eO7O7c/hTd4FvJuqOMGeVHOaC7qLCSfqe4NvFtyjb+IjPIeeDuy7UhQOAhI4YK/I
2FA0NGKw9jrwfmNUj4txvLbDZcii8+Kk/RbiQvylmjW9UdYoh1feLay0jADSF2ei
ZwSk0HbsWbQVt/ZTQ9MQBIfxCLqDA/FT2xRLVMXJ/4Yk+SQRu4kJUXA0aTc9yWlA
kOutC4ofB7kk+2ktZYjcG4WprxKeC/fDoGXlYncDTHb61qaKW95Z7Roxh6rDT8+Z
nkjyTdLf7WZ/ChWsjc9WIQutdC33/G2q68JI51PbRSH3bT5kmakGyOJguGg4tMxR
Yt7FHVC9Otr3XSWqV5BO2rV+RHU3qVifGxJyynzWy0oQc1W9349kZpkjMM+uuhpt
uxJ8RV9OZFYQjhF0geyh6d9DXXQmZ6kdUdCCRlJb0we0+w4970D41QDtkIHWgcAZ
CsVpuIHSSwY0dJAEO6Ij+qOJUBhV/uDmMyaDKIQQkSr8TToJxdLGgMK5U/mVK3Yw
bzVLZF9W01ifHBRy7s6UMdomL/SnwpWDV9DDyru/djfV327I1zvGksxXkxF6srQu
F2PstoYeXaQLtaRfnkop332VCvrgTi5zQTXMck99PRSlM89DC/lkxjyUO+vUJ73r
lEfaoK3UxC+nwKgepTGb4xsye9NuftEwfcgrJ9HteItxlGvp6jOBKgGVgV2e5rE4
BQB755eMQZ6M7lX/fBFLpaHQvkhOOZdP25uAU1V1YcoedzBU+kosP8iBzjQesOcO
EwEa+m8fKclewDfYRSDZDPm088lFduMehaqz/goJSMv2N9sm+pn+A5/1FD0thDeL
jRcRhwo+p8jL2Eec4FkdTQl0qJ5y8b5Kh+Yoh2e6P3aPfOC5DsejMOt3+4MTaIvQ
txAiKtJREHcx9i8tZcsCBFlRvfoKn1XZH/6sDwihFJBVI0P1thFZpRmd8Viby4gQ
GQ7OiMwprIRBMANtufcyc+wUL4EwfbQQmZISYS2JWfbvdyZ/u+sY7Ln903wJk03i
pyaDIO2weX1AYe94OLVaXzbnxs7fTdigi077NVLwAacH+iiBqXm424eufBObzMKn
LCSghihAkXu1ARhFZV3UiSehF4+HXCR2AhEsmCaSbgbZEO0RjYro9bSopwV4nIDa
NEle1chTmQRxkHFYIUmrSfwkwzvkWG/1utRuIKw83V5K5aSecxwDDiDpyTTgrbD0
gP6EXp/U3y23IZ1AC29QnTKgxNX1qjLzyDIURGWmSbOg7W3NClrWXfTKwnh2qx1n
dJalqOpR0vPSoRciEUna1qiJYimrn4IgAVQWc0vxm4k4MRpTTCWYNItDeuxFukhW
GYWjdSmyKMLbMxdcQJcEdzTrR+jNxrqsx8y0X2y7+6GH7hboayoPeBt4FJCXMEle
yjSudxfDX+/WmNVnBTNyMm4asFnzoWgZJeXQ+WXMkeAKR6CNiAAWOk//4LzfKzs9
rHuPoCijlQWNuQpnwszgRpmlSPwlom+y4hSaXbF/4oDIrxDZ+wrh1cwq1HOsJKKv
rKLPsjFVBHoumQZFOOdkWngJfp2MNsa1fJ1+B+1M+eKw6SOkHORKjuMfyF3DUDN3
K3a5PHPHa+bkyG/eY+Cjgdq2PT64mZXO0kjy6A6fKyXJbrIxa1iSFqiqZMVNNqD7
mKNvvzbgT/lBoRLgMiacqjtBIS/cx1r7Nl9FTo9GJREmpM9P0hPwSVY7Rvt6J8jL
vEwM5FOfiBIbMUJHgpAx6Y5RxiuXaNjk1FlZ5Yan8662ehAt5RdGnuNGwvR15QuS
Uzm5LIxRDjYQAVlbtBbexyqMhIq7haStaOz1uQQ8LqIfsIxevGhmwhl/ddfM6AgD
hVgDYfBAY9MkXGkqnFq4KVPOOjjFlMQcoLvTsUnDMvCeis50RsAs6ePOWFOB+aed
jwoJhdT1SGCLK7kz8WFVfhQiWNFE0UmokRxalZbIcSUqOZ1CzUI2Z+taH9TAkFiY
aJ7hncxkgGqnWNHSSZ0wa+RnLFaYWYyPceupLtjs3m47G4s2b5SW31iwhsmmTY7b
BZ2MCT+nkSpCRro6JCoqKG7IeLq4ZGjjR/UUli/O5WDALBTy4vI93+zE8Tr5d5YV
uwk2e7ye6sHXKnv4eafmYukYumfqfi/eZjiQCTRNxdS0HjYOMpcsx+dVQRJxJHwU
Fp8IGJ3jda2jicMqNJ2QYhxARif4rpXvjwCQD9KtVMnpDcZqMNizOxPcfAmv6VRk
ms4pYazrIEa441/FXNVONzrLL3GgXhh+7bs/xTgJ/dwuec1VV3x7z/c1gmYZdgXZ
HdfPIMX816VjTrUTiUAmQo3oRO8B7w7Npedkbwgsa7JvtgGS2iqoiK5DG2Dq75hy
k44EPd6TPhiB6GL1gDjiwt29hqlzqj9M1Q5aNlPezKJtzouTkEjuD0IHlvh5gNvG
6oA4ZEUD9vBZYQrTbtvVvDWTTX3v/I/nOIS5tqEtEUvsZCnB9qK8kCzvetvHydW8
GIpCI6SylZirPoJhS0f3GbXpmkCcSzmjsAow3yypjd3a+lyQ0lzmmkRrmYuIp+yY
SGViRilvv9N9z4mVnGRzlImkpnkazaxK58DV/xqZCbOja/Uy/R/6O3O45xCwNyC2
kL+ZIakg5XdNnjImsyRrM4zoQ3MDQq6PMZT9R3ZaDoMdz1aEuiAQZiHy6giwzOdY
m4GwRGYzZxKDmjdsMyl3UEobSqMpTzFpRrAvcUgIOWpxaymgR/4qU0EbBNV6bW7S
QRImQIRuVSuAED0Q7ehWwiEtVLp7RzxFm/NXsuxXfluPHKyDG2Af2OGJBfEEIKIW
pOs/ecoaegE6L+n4jd57rRPHUYj24gsIS3svljcvcX74lvxdXvXetCf1iqxsL6tb
Of9iigC37DUJ3NCPhpWKOWGHAD+JAm3UxK4tGSTVBfoND7dv7KfG/AD8xPohYPQw
n56DTTi77528CGqccBOrZ3fcKsirFMSluyoBoGD6DxS/6+hrQEJ1fz9bjb6jSBqj
wSgyTkXYHYyGSymggUQmBmiPTw0IbjlAOCKYV23U8i1j4VaEtivLHuNWfmTAGqEp
otzM5n1pDTmIk+ctBkchnLLyKk7LNVEwLciKeXNcchLBIcFxGxGPwl21QXvi7M9w
6sE1ckW3Dc38XhkQF3oMkAQ2Fa2ucziGLTvoVhSOV0SNJBzuDXMlSVUUuA9cJ/kH
m1iCtpCPi3J79+mMmWmQQUrfP9GGnIqtI27eOeg/YNH8eP+Wo3hzy0OToz4FpSD5
YLQbV9+2y/u7uuex0WbcDMYXQUiZ6BsSK0nNS1YP7ri5SpXh9hthEVpukw+Rflez
VsbQLIZcK81HumD71iqUxKSamzZLgiAXasfdn81pfcv0v/rvGiuPPsUzv99dgqrx
GMmxTrfDnfOsuyifCwgEhmvbUBvZ1jL9rumpzjDNCwxaQKh2XJjiVG77ar19+V/F
8JBsYk/8k6spnxMyVhrFKSlyG8FnG/LO7rM9CFZWPO0GXmZxVEYr3IOGScCWiSvm
dMoBNQ3WoGQwqBgsARqYvfuPVg3liMfTBr6a0uCMpqo+bErM4u1RsPlAZm+VXLmq
Aq8UpW/lpVg78wmJqVADxhc01bgrO/OTBR1V3xJTQF9WpV7KGTXVDkP2j/eGaHiu
j4cuGZRrIl782UNBhdkJ0sr/O11geJ1I59a64gmSZuUMI42xsCRsvyIvdrpC0d4l
nsjdPce87KO4LIzXjcIr6ykEE+m4Dld4SwI87tbrk/rov7Tpkqqv3TuVNdGA8shT
I9V4HKJnSJEpzy7vLwOJlU5toduGlWLllqbVJBop3OYrGInLMmpWu+srGpTMxoYe
Puei7hINPo2QGw9RvaYeHD40kPy7YHeETobBsgtGqiQw0lUh9WYsOJSd+OAStFfx
q93NIiHHPMmyhVC7tuM74eOGlHnK9mqEoXu9mwo449xV1GFrL0G3cl+HkPCDw8Xd
eFvQjmhdK8aztWhVi2V7Dwo0/9reo3oYLvWIb2I/nWss9fe4j5t+xOcnw25/wWAT
OY+2LwQgaW4SWd6wUtTubUU840OZmXVY28eEj965alY3ix6/IosjzrtQZ4I/r4MH
EmBkBDeGKQIhaDXYE+Xi6H1BKiwApGm5O96UF91EY17ZYGywfizBiW9BDYmhk4BO
EqOyB/QUrMfzOhV1snmPfSDvgFC/+UKFd2skoWf1Wp0VOJAaFU/dRNUuF2Diw0NA
UNgo7D/Y54OcQvnclUF9YsXDWPqnn4pfzVFD7/QPjHGzZMD9ZB+RjDQQgKo8bnfS
uPmFwC4ykypsboUtwakSrXa8R5AWQVHl8raZ1CjdoseSiFzWp4hXubcm7uvzwcVV
biMg9skZAzDVKnMjSfyrAW/U4+I8fOC9Rvw/L/jcNWBAZff+cRcmHj8gvJHXsGSP
9EBXamfm8JS89Uy6iTlU6RJNnPxIwHSdp1U69ufRLCbZ1wA2pECvTD7njebVKGMc
/8jxMogoBs8loBabzLPIQbikd53YUdh7yL0n0WVTufjznN0Dsz9xTaCS0tFRD34s
E4yIrWLOWl8oNAqAGPoyA7JiabhIq9qpS8eJ1yRvOK7WQx0zpuYFwvrO7foIiXnk
o999tXKKed64TXSwwMrt1E0K7Upbz2tc+MzLP9zE0y3wv/mqpGiUuYvDo/dVyvVA
DxkJ2SJVXUfILb0c/xbZVY1qmJuZaLhPq4jXHig3OVJHaLru3UoEWYfmasluNmw/
jTdrPuOGC4J5nq6PWPgr7CfDizxmkxRxRZ+FxGciCFjOgq754C169CH6TIr85/TJ
Agubrhl2w/MvVQ0hxDUdAOdRAqLnSamgnd+iEySNJU/lF99RCYicOPSVpDNea8Q7
cZecJupfnZXAa/kdiBqXU7lnRSzzAxcxeovmR1VfatibkBOQRQxdfKuhf4gHJpPr
4oOfdQN3sy9/ePpg9U7/rhzRcU24rOsog5ZncVXr0PUe0mqpXDav2jPy/ApGWxXN
lgasNXRiP0XpgE8yB4ffxZPUtPGverC3sT8lXDl1eZFC+FBJQOQy/Qiq9OZXtkFO
kdBjw0JuFYI5CwrTqfeKd7DzGaJ2r/dg97nn9j8BvXNRsdbb/w3xEEuB56A5Og8V
9qRLA+Xl1nslJRLLfVyc3nG9ARE0f+6zWeZ0EN1otoVfHPub+6eXf3+LUwndWd44
ukHK+HDzOLcqCgKIPuN8UpR7nnTUCkNimUmXxdYL/X/j+nI+CoOZvD0WiDl31Lyt
3+hTbLFhtWzu2ozkTi8I5ivcroXsnZDHFwHqzaWvlPe9zDPyEWisS2FbES8pMZNf
h5vPtCi3jkCfEmw7NEHvTMHUrCZUNOqyklEcO6YXO+eW0+eklAJp7dJGY2tjASjY
EXC+/zXVJhy9SbFBuP3kbGKMpp1SK75XgxoKGH4I07iY4+jcyD4KOmCtwSPf9u7Q
JWop1NSW4wAXXzWQS7+W5iW3TA6iLM2bkVxV5agwybqnTjM6+CL/qKGK77LlLjbs
wKMr9L5hLslqHwTJa2n6zAYcy3q8CWfytbQS764O0mpvINzVxDahVAzP80F210uI
A9rKsQHGqYWofrKjeVFwSgkkGFePSjYqaSszJjzTy41QIF7+3/asGEIjMkxtW6d5
Ksh0+VZmp83w4Zth5Nqj2a06a7oTn+5PLEzIuxtBTwvSY2Crwny8IIROAVOED2yz
rRljAgRVhtH/qrKIXJoKYalYQHwJ+DswbAtHSkxgDDpRA5GqFfUUM9k0pessFpMY
39mlbpIrpBf2PtbHJ/9QC0kCApsuwnm4iSzRW8qEor1Ge7IyeP0qOC6a9M+4c01D
cK4xUDaGeXlFd5f923grkK1Fg5DOj3q78LZSX4d7tJ/ws56gP9tcrnkKjttvZXVb
5w9OJRBDEUNsSj1B/hLijLybeSEQ9IgAiDEECTrEg0d9i+RxKEwbwNb/uHy9aHtM
CHcILP2uRzFGTkcsa+75Wg5PsbpGqBIzZykfB48/yb+LAWBzQwDPO6Q/PUEgHhwl
IBRlfhntgFztXryhd70eQJHzRxBP8uzz9Ze/rHd6CNwSvFJ0SaeMpE4fUUon0LWr
JxYueHraDh0uobJW527zhAWojjos6vG3GEg7u7Lf/zzNJCcm4h95Vdbn6kzZZZeG
YMGJ0Hr2sDrxWF8VWCe1Atij4TOHwtnShoADxnfSM4W2XphwnUQgOZd5c26VezaA
myC7YBcjXxHb3J0rEqrxBmA+/0HDFReMOxEiESL1L7m2FB9KtvDb+Hec+PwPCcPf
SWig31uQEFAYSW6kfdmggGwur0T1A/eRJbK+8nBik9i23h8DM8IiJ+OI/HWlT65z
N1NQ9IMfBCFhC2r8t0cmWEs2FtJ6zL4RDZDcg1alqMQnZi+adRtzd19/GA+6Hh0l
yz6Xb6QHPbiwJ3JFlxIFVT54gC2fJx2vd0srtq5gcr3dzVjsFeDpFXGaZ7jj1ym2
dVCLDUw9X+E6Ms/TV1vzmeEElcF0WmrIZ6RrXidNDC8kHpQM6yVaM+2EXBagw63z
PnuppkiSwuDmyxMoypmLI4k/cllxo+ekgFLBZjEntv3z6Y+EaWvY2S2d5R3XmCZ5
oh0aZU927QKZqpVkyccrotELbyZzoIHjEFAcgYsDriiIb6SI4ex6Umlpi4mxAsZj
XDmoascgEIBN1IvXWhrCrNAPdyesaqSHslQg36kLcC5U3TKYp9IulocpfQ6XDJNt
N/AUfS9aGj3tuVjbU/qfLKBwMyKl0UxX30B94v0GZ2kxPuQKHWrxp+S8Ydl+tjxl
ODtTW2QLZir7nmlL2u2u3LwEWvJWZCnh5IFEqsYWRdfqBJ3Jtd4jdZ+m7z2R2MPq
7zIjLlaXgA7SdGhSJs2tj9iNL2Eb3PzWnYA8Pr8Sn/skxM6P2Om9wRfQ0tCXXQZK
QQ3iuIj3JscGnfsQWZu8oyxEwKsZ7f0d3vAIVLD7tc4IiDeGr7j+JPkBlvFsSW91
IOYERk6nW/EKsDP6xSSVKZ220V7+xT6TKq3TC7xGdZmAbzPza6IEFkjl0bJ0pNia
MPq9C2eayDI4nwTNdLgVy3Z0hd6Ql4b1nJBnMxsxpUf8AtcISAkPndGwrqVQnv0d
bwaIHoDm7Cj/c+rHGpgthK+pq7AcQ6y7rlssLCsW+76Cv9c9riT+jLqXPIPYx8AD
XCQP9yPeE/P76ZhDW837CjbwAsqaaAmnb4Pu1VG69YJ8yn69q/O7V3BbDATlJn0I
M8YxETGznZOz3SCU+7AhvGkuYlzyyA0kPb+TfAh7kdnELd+67ph/lYRLI+1WJC8t
1fei5p/Cx1yuMkMYzep8Z2z0dxcmXvAImO2cbvZjZ+mEhw7lLtauNlk2BOdmVSzl
66KTH/iCMM+jPoe4cqEApuVOAOiPKr6kwnLHFg61FZ91Rze84DVTpsb9rg/VKaCt
QHA4EXbD7cNeUOmVKR0GjO2XQTyjDa1eNpZNAYwUUtMozDVGOVQo0YimV/a4o7Yz
GwRx9CaPvktqAepkg3ePmSr6HQOHbA5IFdgzl24uepfKgnvoRE24rPhhMLPtvQH1
J8zZmegN1Q1/4L5oWlL5mO7FpowKNFaUA7kJgcpp7sWPBtQqxXZORU+nb6OABEL9
C/7LY1QTNVSSQSG6AOOK3tWoWOiPtD8bcUIYWeVQZNJLJW9Tw6NY+WpHyMvbWrFx
McVsVFmdjzlwiXp1+lP0Wm5p4DRwvlTA0hfPBil6ox+pa7s7f0tkSk3N2+5EGzct
uiGzjbb/DB2uWHwWdWvq9Eaj5HEUlVXeDuAIh5iQqGFly8OkOcNeEvK+4QmUYjp8
8oLy+0PHolxA9D5rkhMczrJ1xDbBFj9CTyphHAxdsid3eMQ9SX7xRfMB25/d1KnR
NKGOchgPcUGG2fR/gW48OI1F3kFV9smoV7kAfwSuxhn5a13oM02n7TdWfgMNTAKF
BU6hBbudO2u+9jGQDuhTXQG9jvPASWbPVN+/UkQxyfCArwgQzX+nYIFHmJthFZWp
kBo6m24en0UdDf15uI/YZ6ZlKLhLumvngM/DWJDIz41Om16WeHgOL136j3Q6B+K8
bGFgv3mXBsW9UoZMnigQyRjS6rKS5G91fzSt0336jxYja+7adhNeU2Q5wPpG4ZBk
8aVgp4xvGmUwsmpTfUln88j/TUOHqSnjRtkdpyfGkK0X1/PQr2FvI4BDsBuwbiLG
t6nZBvtHVX/VmySb8XSm/+eTUnpat7aZBzXMvz/1SZgHY5GsdbfF+5f6K6x0B6AC
Jqt1pjLC7BUd9umIP6PEZC62u5xffdi2NKQq7pFXhTmWVrmzr88Vmcl/a2BmmEJw
Mc75KYIRDRzPe/tOePbSDuHnXETYe78rvD1ouyq49NwPc9f8A0ILfC911dZVctzE
W9X7KKJR32KeT9hDZy3SvjxCpmtrvf6W+edQ82Lj1RVllwu25T6XaNWNpO5UZied
RWzCY5FbdBlraAw4AimVtGaRYb8cLJTcg/T2B0ewoPUOKBVBFLlxyOiR6pXSjCY1
4GKMkw608uPyL3gJQA3Xcxl3KCv+a7nDU9Zded719D55Okf2Q4CAt+bSqTr0CBuG
IjB7Sd8kd1wK3urmtirl9kagD2yrMXPyNr55a6jnoMjTI27HYGKzaFMOsqt/AuRt
H/CclyuHtXD5Tmm9MnUp7GZYe6lUDB/KCgHRX8Mfy5NAPief0SwZyRR7Tdpop9cy
9XNpJc7hyECFyZFRGvfT1Po2kF4e6dKwce4JXGaffkbZeC2yhH8IhdJ8KBxeKAhG
9pdzenLUg/xlF9bSsfeuSooeOeQyLgRulozNHdHqdw1eMFoXlks+0dY3hgdpl2bF
h8LRgRbBtw9l+S+5kmHm5i01jSqHMk4zm3dbZ0BnOmXzpfxCA84ucwf1rOfHn2C9
g04EhiCLHDzJ41dMRIX8cIBDZxV5Nd/5Bcwb4Z4AadHPIexrmQODAAdNRd+Ay1PX
4F0i0oN2iqvlZqwcQZyrB6UhAFJs9S9AyUrTk8C98ShfgiAd5zuZmf49hOO3tqIa
1p/Uu/p54qKInNOociSyLH3O4A208M0x1KzOdlIjy5nMzfwhzI/+vqooqOUzMz39
fNFTRlzWSfpeC80xdR7dztRelUr7GREiX8XI7WVHsx37+ivoz799KOISwGNUWJmh
1qlhAE7Xqbr3pTXDvcVKHvcU6RwNGJKWaNT9Dnj4zt6anbS38baqMln2rNAG0Z5j
vqMAszneHkQ17BzcXOgJ8OXQDtRzkeSP5/EmuDwSIzx22fGQ+39gI3D77wXw6uDc
BEJDNWmrq1KeSdjmkLEByoNYCUwtJcx2jw9eIkOudHs=
`protect end_protected