`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
ddtXksX2+yylW5zu6QL2Lhnb2d1sD00763mmSITNX595NcHTEkwn0zB1Dry37fOW
FufOhVzEJp80NC5qZ/+F0Vk7Ik02dIR0elf3clrjeJRK85K4e3Hoo4xn7YbFUIms
l/8VZSb14+JVGURjfswrIyCUotIzlzVYZ6gzoZwDXIi5gQIBf/gI+KxNXPaKV+PQ
Ufys/12rjO6aI/pPlqSm0hCvftmBcnezN2hk1UeXgOIuKZnogjOsf0iJVX2aOOWE
6pD/psybjbnsNB6kH5uFTA5frkzIzkzl5d9+YDm9OyC+k84E83I/7/j+rk4L2dah
QJOvksSIzN867/4Qt8qYTQ==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="MvBXkzurAa5VTw+1JJ70nePUfoQXBvZOku/SMmg4TwQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
oRtzZL4VJ4iwysPsC8SXYCzXS8Fw2gtZTOskLcDV+1B9Nzn1zTyNtlo6lNICRmmK
ZRVu2BmCc2G+fmzynYlNTnSa7C0Cuel6FYpxCBlOuk3OF2tzAmLAuDyOH3Z1Yjzk
a0aHuoCdIRKv7BrZCdALt03JeUmXKPdOmIlkVGFl8yw=
`protect rights_digest_method = "sha256"
`protect end_toolblock="Jn9CQpRhJt4rnzZPRk+dOpzAubz7omckX1MrFd4p81o="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 10128 )
`protect data_block
gD6l00tciPUa6pDNTk/+t0OO0nC/UTtBwLB41d4inuAUA3i/ALrNyoJVcBnAmEQW
ptbcNp5fxEUJjnOxnedyZEuEBxWRieZFQnkRdF269oMWYtveDYtwKRcQUYnZrNC4
vBqptfsHrtjSmmSfDQQshdupCcJzyBrK/SKny7qJ9zBX0pF4RlgLIOsp5Nq6fRr6
mmyWtIuFHC9okX6eHxRP8tg7WjCMSqh/wMDtpqF4VBjWQzraDSlQ8NPOlZnKi4gQ
wITs4qbR4yzKKa/roRwyoyo03cYfzDYkuHF1M26ME8JUG3Omss5mzrOrC0y3xc3G
lacg096tI48SNa9GevBPP0vWjRTFf77VhzIiZjMxzBV8fGC4/vzYhmfoZcLSYxMJ
FJaR4DRPV7TXbvpkBbLO2L3r2LJkJeD373ICG5Ed6Oh3L7ezRWD68cfJcFtyRyWL
S+hHaXdvQ5FVggUn6wEglOG+94iKP025EkBkpOWjd4+v5FECgpKFWpQuSVdLYaVs
VX5VUv3+YXrWML+TR4qplJmstUJD62QLdgzMUZFa6EdF6rGZLRCsfQAJh5qj9P0n
70XQHl/oRvpVGw3ogBFcSCBFc3KbMnWOIl4TdE/iZtUfeUXO0FBcNLjdPddaVL+D
17JdD2xSr6CanJHxdpnGcLgSycZTbgYD21DebRl9fFcHjoOUNLI43UUpj2zLfVSu
FA/jrmM9HlQWWHzexThTvGvuFWxLykrLzYKTFPyTfmKfl+hokCXZ639xvOIe8seD
Y2DSevN6L8WWuX+iP8+saLaMwNdMr9vOZ7Ne6f7POk2+SwzxeS4s92YdBbIwL6Q8
UDxsB1smcS+XDKbMoH1Op9id1IchcR4Gq0Nvhg7rDrTGxaSYlrWaCiJ3w9mxKhU3
sXtfVotxkhHrYBO6nCRUfrX/Ih3jl0uX7/u2PmxIl9sNuZoTmDHwkv6FTh4ZaHbI
eeZPqwyEYdnjqfIw8bDKRT4vT9jv3jZnnDrpDsq7Z0IFQ+JZDryriXmkGo2XSBJv
trHYJYjzzpxMi3Nibuv9C05wDnfXkn3PYWuLhnCNa4ESWLKg7rlzGaZAj2ebn9xE
UG81Mmf1sSl+PUWYq7D+HFpSn4P27HjBz97Sk2fZPPOQv2Rx2i+Mt+UlMx5M8mef
eXSIa1HReLh1OD3WKWCmx3TlrGhjHay8ctRmV3KPeSF3hpgqPH4XU3Oda7JSpwuH
AsuTu0QlpLCBZwk3UcAH3IEZC/WdQ4XxE+lbijZ2N4d/K+lY90i3izU/rO8k/eR5
WH888CgiYJV0HbDaP0IdzQPIm9TKtP/iBHYZKOP5qNw0P570xf89edJa09nFCK+z
ci+txVPC9C2xAIGlfUlHzTGJt7nx5ByVPvExreg6F735dn/UyrTTgbAK+S701llh
wYCD7SzZRGP8CJlgfFbMj+0o+fKep5Kqhc5XtWFZt/UITBszLpFgVeu9oa2gdn7h
wEcZcFJH9HjG/8EGIG/YW8N6NR2fI5wUP765s/fx7ju8qQThibaTeel4pp/zfNEj
9jupTAueyw2FEfAQhqCT0Okzai5nxOp2MsChws7Tlr3zbuebHv3qV2kQ9Tc4PlFo
ZjvGgaaXYFlmLDtY7CAX+pCB74/CBgfwWbafdciBHmoLyeTC5kgd1MhhQz8V3Sc4
LCsQq72AebdzqyjXSYBQ4Ml5iQajX5XBdLopAlYn8r97E0n4SKkakeE4/YdowmHA
m/C5tdnqzcFciGTtDyJSb1Hl8NVEoZcuOfV4NTll1umMPzO9zE7ZWPYzbbCejC3o
aLvXrb7idIng5e5vY76bkOPw/38NNZuX4f9eygWoqg35uDshnwk1JeiZDbKvAU7g
3K4q7xMioXqPmQPZTlN5ofpxr5giq+ZWfBdhu+0xz36p1OuBhnv7FS7aMDLXEtMw
xPVGoZ2SWxqPNpYbfBr8HpCds/Bbec3KuvAHxlcIA9ICsA4EvuzLyADcA//ypRC/
Bke6Fry1b+FxyuXfR8BAy+2jfX9NfxnW3QUKE7XRLt0WhexGN47kMOA8sntka7Du
8SDnc1wpprE87eeZEKniI+E+cdkHT/0v7pnZIw7p1Tfem/cKvvRQUeLRMO6+XTre
mFf0rNnhV9XEyIm5jQ6JlVK6eIGyDQUmpAoiEgeQFmGs64h+bhwplYKMzllzJs1n
E6bXG3Zx66MEYxaJh/BSisrTVz8baz2CcyYyJPpYkjXuJRXNMzx9fsHcLGsO5+6s
uPRntHN6Yvf3RvV+/rOkdiEnved/Lr3mXzCW7Rr5SwpCR8ZjvTLFBXzfzRR5OQhh
zseolywJLiSw+6O0M/pdo72oOMF1PI9OjOAN46wphWH1xGWflWjgve3jqmkzRLH7
gikDM7CEW3XW4ir+npsDeK4PAfSIZ9onmuAcVTj04tO/HV5xVpI6oBXmu+NZzazF
+soQu61RssBNbaFhK+wfDNrkvfgI6po53rdIfPzScRferaXApq1xAUD5AWTu0J52
b7GBg2xOYa1BrlN7Io6yJ4zNQafu7bdGcPSQ7Ki4AdNXpp4Q9ZiTEpRLLYF+Pdac
KvZYsv2h2fObF74zmQGiWIFStbIfu13X0BfsEsPsIOKxsxQ+UWNKk/FtyNy9fT2y
8qCfd1gIuQMjkiKNPOxF5u/kbVyKGCy6CUeNed1cdd4/ylngvqOnU506pc21yjqB
xGTWFzE0bOGWU9GymdGPWVo621+yKj33xKRlAI0jZIiRzbDXgXGx+McPNSZF3UV6
QR7+2pucdWSQ8EzWq2SeZoU1ONIon6G9p5S7BrgDX/LtkWuy1X+EGQ2y83tAZbPc
RmyNOKOI07Vtf71gAM9w9g8QIt2XX+oRuk3lPHPQiCH/mT2eVmYGFbspt85raUjP
YGyjzrYqTZl8xdYilqf72nE9sLppXAfZSX2PUMKRLrTMD3gKISJ/PR+UC03DFiwH
+75p/e3ELE8BrLybN09umurRbpVNWd6apvuuwh62+KHzS4yvSaoQrrUA5xIA4E/a
um8eSOUBCdD1Oj6dyhTCPkfxxNTZw1YDqnuNzZ2mV/Bwr20I8YQoKSfRTwJviMHO
vv9vPKlrQAiHgTQTDaS/gEuDQ5UZET8jYW8E4T05YAxE+PSUjRfifRejvTZSX9HU
kYDtdd5S78eqLBnZbG79O6tfaZQZlUHi1cjW5HKNXxY8gMukTqDI/eC0ZwpYCYk4
9z91BTieMEcjI5/P1RtxtzcWUMDD8yHhJRZwFxs+t/xI3XEj7vDx7BscHmjtHyoh
YOFo0Sq+18D1yJpx8seZgpSq7gvPbpxIYKwmdb25pquCPvHyY330IVVvhsR4xt3H
+uHbmUHLlEMh5Tk/WJLk9pvj9bIYIj3kvFULo5SsdcjI9Ro5+y78rFQ1JNZuD6i2
JAb5OqOCRzJsYqRr3gWBtX3xYO+q8vDFQLD83oC4d4WujJL8BOcgBUfVxBOhKgjf
wYjwlpkhC5eUwv/Rekf2vc4CBzJJQNKRx036UnfSTiG6AjuSRSclbKV4l3aLpOdM
Udgvh85yYOx2RwYUqsa3Pmy0Z8cgPE0q8gu0b9s5LKeXS/jucGmM/ccHIkTfIN/a
lXANKJvQYZb04lOYK4UV8C+NEM4q99fhsLkO3ZAwI8iCZqGNdLCdrh+VvhJDocRn
UpOl5eD5//tUTA/f+sAunma8f12iyQri0kEhizSMzyIP/ni+fPat4T+K1Obkv5Z8
fVrz5HiVzRsTMva3wiHCegq9oPQ+tvNXvCQLqFWLXxog8Iw4ZPnIHMoeAdyH9GCg
FrZ41SahndSa9Q4y+ZXUypSEhDGEMfeHvv6rlW4j089u758whcQpg245dYKpUJf/
phyJxdPNobIPeY4YI67wNO0UGrSlJy/CtISxM6TpRk39/s1lwDfaX3ABxZwoMmv9
+v5PzWeH1X3OAMjFO0qdopM5DsdC55P4qWUZNMdIClQ2vk6Q/+s3WkK8KWvEGSXe
hc7lcpEy/Gsti1enafwbzL1qshZluX6nhtafvQ3fLiZe/vKAb2PDEe8uVBCvjRx5
eDmy4MbUolBjFkcJY4KkdXkch2XMohRpyUSYrXdV0i053YSQ2NIcQYwmMpmrxYCk
1EInxHREN7atXBcrwLE5IgPlK4gRgQVh1FO0F+N6M6H16hz8a1MlpuP75qESbbAl
uAA4juuOcEXeVhzPp2J13TSwMu63kQ1C6qSw5pzPB4Hgw6bjRbrHjjLM8voqqkxH
upAHT889E0361EmZJcrG+oyS6ALBNSZquMUSURKCBb0nb4RV1BRA8hFfRfC4kQ5F
/x2apiyAoXwrrLiW4uk6F5AGQz4WJZV+bjMeXiU3PEibWjZTNw0dt3TPdlxQbPVe
GI7Be35IChQCnIz9rCxTs8P/FuQXWcvnYQjfyBCy/eHWrlarLMOJelaPR2If1a1u
O3FdJ76bvc4i3X/DUsNnWxz1foc+B9q6e/kupIzFSsWcO5ZG0PRnL+CGaM0K/WAQ
yK48SNxRMTqCl2hKwQMM3DzwpWywjUITDRZ2A5Eh2sAIiA0taz3wJs+zGC1sOFDF
hqNk1X71zsSCoze8JVzmmYAxgnJN4goCVd3jtH278B/77noa8F4Sf9IBeu8k5YNR
m2Ar/JzD4M6Xk3WgluDYJqW1hx9NmYq6yiLN8LZY3ZgF0gk9JnXa3/iUZPjaYLhi
khdjEuJKo2iGHdLFM5FOLVueh+PMnZTNYyc847TXbnDN3qBA3IfvVhj3ZJQCoEc9
yzn+Zl2ou3j2Zbfon/cxp5MKAigYgfN+XaLNgkt4fxgR0TqSVQiyJKNtv5wIC+sj
ohORy4UUIot0xGrK4wnIoHS1QaF67Vx4gYYmSqjmqQBzWPZ20Q5Po7pNrZLru9vH
zBxG8hzXCKmHDBFvdwVROAttRsvBXyeAZx4PR/sN2B8wTkN8vzUqFgOaTfnM7APb
/44FPtuGiSsH2yDK6Om//2liKXJlToXQTGXoWOgsuUsZqbdFFoWo60OY6J54FBCj
1DwmNmfzBOTaKz8AWyce2R9yHhvzNkBeBMvAhnRwEDrYVcNNJBJV8BtRTAyNRtCq
5lx6RN/yel61p/H1svlghsLPr9oNVMwZX0Lf8VYB6mGiimyG6YgafXRyDVGVzrA3
S2Q7EUVq7hZT2yj27Spr/TmNV5bNDx0g/FuKG/GVH0YFZaDlNxxR6a6OvL/Z0wxh
qxgtqCuFWw/nCQXsd7CboS3bn7IC7WUbkZJUgclkQ/eq9ubxfrRQw11ocaiydaEs
4Jx2dsnRrRJtZ48FGAGHYVqnl5dkNfZjItfkA3qjKEq8QzAl++rEsk7+0Q4V8lgy
rsSTJu2sX+PY677bvPdNV5zOmJMNYyq0XvdM95Y2oKzdxl32f8o0xicLwF3ZPcBA
5gld9k+Bnrav4pkHMj+5K076nsuYg77KrruPjBk7hDpi0IetMLE4QLKck+lsKThw
4om7XQ48+ZmcV2RvKIg5fFJsvyjhqk/AXyCseNoP83Fgx6sEbhPjQmJnGreAeb3n
oyexX0Qzdp2zalcRA7e9CrOwXFcwHG0CLD9aihrT8pC3iAco2hZyLuE7IytuDRGu
g0UdGyC17AHFHbKpndqo2aiFn6zRZl0mlN2Kuyz7Y/uHwg0pehG9JRgdbxQ7vlzR
eohIuGIG8ZJbehuQKk4uxGonP8/6+sgv6S1nOzSDKrvu/0HsDzgEsguIoLqxyU4E
WN/hgrk6G5aulLQ55xKMCnWr3PbXoqdyxrp1REwIUkTGcK69S8dUKtGpFU7YZqBW
BaC2XLevDACi+FoIEEdg8qFHF/KbNHF3RMZrQud9aMkTmqGa8VZrcm+WIYrr7TwI
9ip+UBYyjRZ9qX1iBOgxxSRSlAJXLp6Spr76/JjsMroGpq98lOUPHp+6kTiheXb3
UFKcHOEq+daqVG7/LRqExNyfGRmFmoQ6kceErUf70J70DqwU3KbW1g/FZFQEvXs8
4EZ1FbmX6g7LyIOujJJ6X2f50N6m0WaJxpUXMsaqqkQm+331mq90qYuXmgdwAf5Q
rpM7xd6tdCnVc5NKW4ugQs4qVUbQVPZAFuT7lROHCua8RwvmAtz6FlY7ECIN8Fdj
t2qAH1By8C4mzP1gkLSmJ4CvX3r1hrQXEPaJUeCqvW1IxG2Fx14xQXE1YdA7YLee
DQCbcB9zmz6ZD0GUU9JEZBLTfOIFYOhxPHDBYtVit5Me+32QqUWrk8EpIaqYy3Uu
Dpm37hzJ01nUptNhidxZgGAe/k9TZmOXCthcMB9mfp3Glajv5Xud8BqB3YCOFGFs
xSmmUiVBlHJqxZARcDqiS/j8ekV0a3pFI+n+0y0mMtMhmMi6wfzWTtgspek8aRdF
JESo3GpG6PE2VP9pYqZ/chcDg2HcdRcNyb2lLXImPXDf6PPY3W5jB4pznFTNBp6L
sYVr75mEMSeR/RJOxQJw/g3GO/+4YkHcYYd42J2RjKi9i5kKuf1qZw8JeNpqno+G
bUQX80FbllB1ZvyJQGXYe1/SGh03yAzHpJ9o2vfQ+G1Sw2KTZWxxsmfP/3t4ZJ+q
JtLAEXABGejZg4d2iX4r++YrBYhXPX8x0uYXissZfH26z+7Zb3fzJ4RwoiN6s8b5
DOFjKgYoJkzPq59Zdp7eUAW+QoPl3OctgZkkwg9Ct5iUB8mIytUxdxTThB+bhRhu
Vlw4Kl44EsC5ZGcKmWvsOMxqyJ6EUQWaqlXeW9txndIUgMfVOd3pOYc67Oy7ukxG
lfm/eqfiOMWgzWTaKzFf+rPp8Q+QhTeyHAZh4A/kx2qobhfIXkK7kUl2gncVFkkM
2iSg247r2SmHlWu034aqgTz55kdqSHbEfzCva7fWNOE89Ua1sewTE52HRHbz1uOv
MRjPpVO/N6Jbb/+ggPIud4tjz5ecQ6klGwm1+O+9kxfgGWH4JsYWx06XCReau+6p
aMoVx8FO7A0XNgudRWwhxMW2bmdZ3VsngGvDuX4uXK/d8q1mZM9LvN5KaK2LrNyV
CpNh+d4WVDiox925r7swu9M5BamjTcHnSSPrmt7vtBwSFzPpTB5aXNHb1XjYJ5nc
VJs4qYI1ieUTwn+iOZ785A+MxvlAhWbc9qea1jQZWsgWd0usHFI78IffFZrdgieX
gP130Z7A2DO5U7LbCXXxjBv4xAoJvIIeSITqi3aeDF7eAA2MohprIX8TBFSxR88S
nUxEdoiAwKELch52LpKcshOaNh+W1hU/y8/Da+LLBu6RhT6k62z11A5o21S5yCIo
cSTvmqUA+JZslNBTVXU1oLbYFmCAlIy4uHDrimQRVehaEjvuZs7pC7WqLSl2f0eL
90C1lVVb11EsRjJ8j/Mn60tJbNZGXk03ecYidmJl8HYJYGdr6RSJT3RXhRWJwH0v
0lURBzSVO3PzRoRmF1Eun0LY75nubjIiRj+sKZaMvPhU/iWgkjRtdTCRcsbABML1
WksX2e773KR2WAM/qQMWOyd3YeR8xHBhegCTh2a64xEoLk83RcuBoMMKQhCB5gIg
CemYwaDdmMuMa5I6lrTAONwOprK9A698VqVwT065HJ7cHkF999ZO57ff2PVSMqqp
cM5j9UZ7C+IpHYDH4VBBxMKC8lojOw+HV0HYfVxPwSlZZvODz6FHAQJVrdgNHw4v
pPCKxApLGrR8yHWZPZHpQSCaxB8XeTfPF+c3VLUXWVQN3kS3nvo4sYxDsI1aa9iV
GaD7uV38gZo9i0Kyw1eVsAUHfEYPw+888lNgtvtxXluaErW9gyOU19JEreSD4+77
g+4NejewX1KOf4aDJCH+13ZaO9fwPhBwTGugq4OAeHEbkD07gRPC1WTA0EvcCbGA
K5Lf44tAEgJdff2VYP5Yn0QV2NLjm31fryvUuIPvqd8ZKlbx3LDM1vBGzOfGA6N1
obpg3k9VjCUQcKxTPqKFqsGg7QzNnQ20yKX1WgcodHhugJePMxNfPybrgIJg1LLd
aHn9W4ES7WkObEynGiPfOj0DPzR0ee6+LxbeAyOEKjO0CKL2danoGkHJm11JCOzI
GueIGW2W6lvGznXLF6OX0Cgd56UNcMf9dmf++l7LGitjZ9YHbdhzDtg9PLEOSNEr
aMJ7JnCJ+rhXrfHBoOEs+/beRSC4SJMZL40oKVbVheElWr4/xEDgQ+5bcIQQMeXH
O94/RxdYL88LQOmr+2L6fJUslQPouI+iY9DPVIiWetCECKeGbeFm1AZr9oyAvrGv
/92xwDLElLFo+bdJjxSY4EuhoFF7l+ngbQpxc2HV1qCbAabSwRVyd2MLf9HEhkZk
IcSSLTKZxwV2ZlgkDM3kpLm4OqRYJd9uKiQygvbdFdA7lUB+j+rKC2ogVM8+fYcZ
CF5mrSdkyj3oOjgOmOEK4azoA6/nbd2tqZPCr8msETSPLrGxfUZdVbb+Jv8M/Wfb
KHZp2hE4J3L1sM5vZzG2qzusWp/ysw1Yje6Isrfabzcz8HwZ9SeqJGcltN7d6iMe
4Q6fxp/gmiZBpTlj/wQ7EA0VweOG1IX5hb5tc5UavvlWvYcDprMS/EynwxPq2cyY
UOXxRyRbP6yaOvj4gV9undxLLkAY570Pc4qtM5cS92eown4cOf2I+sZoUWCx8X9O
UFu3D7cg+ZiDBW4bc6ua9POrtOLG2pwvmtwH+dELtLAY5+1MNnv48uY5UgGh1nQg
9xhvf7PGov+l9GfjpKLUGAmm1hV+YjbtET1SulHq4DRzZBTP/J5+Hh7AJMKAqmRN
658EstW7NLINi902gqZvE9I4ADLTU49bbStc9ZCr5o7IeSRnU0yR0aLdIBnuOrc6
XrCMcFWYF/DW5MenwQrfAcsjGcqoQ87R3sddmyn61weOcv7xfdtz6bTsPqf1tgLN
JusjuJwg2u8Wbn9b9bFHCFHIopbkCb9SyLf8gD5ix3XCSRRJqaHq3YZzoU173HhI
Nte+e4qg+r+Yr8r6X5prVEaqMtyKY93EXRYQvIjWywe//CFXA1uN95GFTeaosnbb
bwh52ED4N8ExdYmMLZxBPuqlbvLa4KAyp5Y4xrIzrBsclHIDLYPOY9pFOT16In+5
Rw+srRpcvSIey5fU24hBbsLyXSdNTH9TOsCxq/4OIKG3dnCNInCUEEhAIWztw9Xq
rBn1Mx3MHJZchq6WqpehtuVuM4slUHNTTbHrhF1EqCdYoGt60u8LIYXzXSkzRVUv
7kIXT+NLvAQWAP/JD+xHQJ/dtevvqYFxTqqMHCSDvEClOMYp/a4nbqzX1IOoN2HB
dPQFM46GwzJ3NcemkgJZIiEaJ5VzWfFVWSxgFIsuKwO3F0FZeZ97HiUPReotuGWg
6UqxN0FCeGeAUrw9z+8bip/yU/fNEyYd9Dl6RyQllFCXB773gobhYkDiJu/Fglpm
IqRUTmetzGhDbWgwBA8VECuygPmQeiikZh8V2+OdavLRSRVHbLyDJgCSH+pP3wVd
EzRts1IdL5ji0nkIC2PnRWw+zgmGjLLt15Nfw5gsNni1KDclV91atya39tnlrLqs
JzGpz0pRt/c8ks7Lclj5xNdGCYPb8uhDnMcJ5KdXrVH6Nb3itst8pZrSDQn/bWO8
dzpruzXHJmmBy4Stj73U7xolDamCUqPTiqw3iVZXToiNMfK2GjUQ4d4YYGBmOtCy
ZzPvJOeGph+GVwxg554wX367L6+XBjK92ft6ppFALtlcUmt4b4VR0jCNp89IH61x
RoSnc5FJY5VGhC5TkaDk2mguJD+DaeKYguGALWiCT8m6EBKenMJGE/RKEoRIOexV
CkXBvkoi5vI2jXdaVcjCNiFnMMd6BmKE9cYZ/9yPYxyIw5/eyMFrdzMwNPwnBPGm
kdyoYoRDU58bEwCoPoHfdls2V7NmmP9taUCY5tzSmJzxUGKkl7MBX5aUTxcRxebw
tIxoNZFFMqzL9gMx7BPSb7MEF5UK8XCypRF3aFh4sfLvtsGYbjjv+ltkaj2eom0s
rZthIzaR5nToE2DG9zT5ZdQArQPRSuvvFACdvrrIJ8dyo35EdxwQeWzOIV2XheSb
PyEdwA7T49iNEClYfeLOW+tld7DcHduoBN9O30xnxxVHPzzn1mPOyby93xBDc+d2
TOeYV8lxq/zZUuVvwnfigjNGhhxZlAXvtFTI7grwDVUU31kFXCmgw3rGhqvqLk2x
bAoLcSfUCX79vjoP5GQ1TAA/8w9vg6JhaybQo3QNBbQntekj23mA7nATNhV4Q6PJ
8u+5whRZhR+azgP+0agvahb5Q3v9rdhSjZasEmJy2zBV3cd/lP8glrmMOtwGo3ip
sSKcAOQW0nhs/1GR6lcw9LcVJ0YH6LbdC2eWFBrB5uWJrmvrK2l/kaFoJ5S8Wd9g
f7wLbniByZZkgocFLyTUPUTfeBx/WZ1tEaUjdPkuloCfflCQHaaQVF/p9qrUEvSr
+yl7KsYkJ9MSYBVe0FFaEI6O2CYAYUE2tbRNuWdQgiZLfJFBKafiR6ijjPqNfyCH
vKlhvxDg7csMWXiU6SpAuA6CdijBwsMhpKJy/iTcI+QgbwGpXcALnGejcM9G03m1
lgmx30P39LN1LDfTRZjWMY5k21vEKsu/YmNWCyiR9QSiJPV/Db20gNy8YxZjwkZA
VcihDJugLpWdyQcrg5ddIK4GfVCtmF5P9EMY/J3sja3pI+mV11o+ZgCNUdTa4txM
BovNm7WDc24lZ1UvhttlNTP7x5o6+vLgTVPSgIAqNeyCDtcim1ufvxcAoIrmVFua
zpySWHS20ogXhM37YlAJfB0AWSEedlIPEtyJTmWy910fd/PGIJtZTBzsbdXdKeQt
BIdMsCKDym63PFdisoPIcidv1epoMz3SVbyqbRnW1DbRNS1PMuHdi9Y0gFgHZ4+U
ZZV4OCb4SRmPQ5NmE8DmWaE6oxgShzEStUdA+McncKhl8jKJJWYJorQxPl51wS6M
r637GpTUiZiaIWIrE0XbJyP+1dVaQJd8mHsYgZDFDfEy0nu2Yndvh0ORr1Rj1Rlo
YhwJ8LwAvoVB9gZDaDVdKfz624JkizUJhB8n5LEreWGMcLlUQPikPbtJDnUzqJ7a
4DP+X1htiQ+rVriK4g4m0t9CYiP9tGhJ2GZJ3VVOu+xWg2oKfhz9uDgBCY+EhjBE
VGR7TXZvtYitJe1B2uKndcDPbK56dmWdwaal4I/13s5wTI9nNDUyTpoWd/wZRRqJ
R6nDY4snZ7C27wcxedSpMNecxM4jCUuQDGdJ4PzaeNsy9RRKcCSxl8JrHETvdhnI
EWrUjJsG1b/jbL1gDHdi7SzFbk1R1bztKDr2Kuvr6bAgqnCQILtdoJp1gePJmFlI
sVwopNokNX70JY3dWX2kBlXHwJnGoNDO2KX1jX32rC2A61gLmJkREz78yBvaq6JR
RODeZgeTpJSvbLwOjC0rE0nwmWPwmNMTPTQewyFvAPwzffuNY4wWJiYoQLwC5vOw
2MG4+SALFN+j6i3Zq4Lm7Nkg2Lh4gj6ORgFZpxSVxRSqMn/ewQooHiUPoA9fphuE
wAs+oODaUh/DRRSadDa6g1QzrDGcd0gFlVfkLlqcXz++tv2wZjQpm4bGswfo1j9x
2cNFVA+Zc5Ug2liYaTmM9oaLI/yGxoIJZcX+QxKN3OeFCu17BciwK1EVk+UmJhJk
kp0JvVBlq/OUfBPwwtkBbmAXUhSBLrL52wau+39eEYlBgueaD2CqAOyRkAhEZlXI
PLLRoODyXHFPG8v/7xBwAePXe2Natcgs2oLiZRMExXnanzfW/9x557/TNPxVpFue
Qo8KAQJv//jS7NZ8+TJqJwX3SCkth/8TpuQO6BWiz9T7/OZfLi8mux1A2uzUq6d3
8H9ueyR7M9kOY44IqTGor/lvIv6psrg5l52wt+vmRIwEyDZtjurJnq4cqwiEvh6/
Jq4yZZhAvc/8E8vS0qMcaaJsZ4rbIDZK+yvHqYihLAqh1NLAxnZsAhctkUP2afXd
/48Rln1f0AlvGl65YxtZTSag3TpePiTuwlhEuvI+NIrah0WdGQc2XN8vsBUrG2h1
mE3Jw0nlaHudQN3ETWeKOCjLMkYcTjnubkw8wtVo3zXNJAwln/3LnUWjKgLOHXO+
LWMLHthyNs94h+w3sGmJH3Lqh/wGI9sxxQlgGd1KwtADXL4wENy2+Ikt5upJdTxN
2GrqjliKf9qBkJGhvwt4AhiKe6yyMseI8Tl3J9sI4NbDPAQb8A+wLSPbq3Sm9XBR
jE1rzjgAiV3j9taNK3YL+Ay7ULAJ1g2MnsgAn7Z19GqXQLO8owHhOrPVHXGa2pCL
F9fxDtj02bVFivEZN7F7rguW9BInK2JnLrsLits8+bPi3I6iV154JXVT+0YJmWBA
RHkXAz+BL9jTSD4n6fVLfybTPOOZ/saNCTeESRhqeXTJaMTHuQTtN/prK9ueLuSQ
P+k4WzisanXETYD0wwPTlro7HLSILPUt3IdrOTYKic0YlURCBZBZoobOLpZfRKKk
UllJugnZN1afIdYQu5eiMCwudIz4/M97VnUruM83Hzg9vSHTc8m4DcYRmS04kLi2
F8L6C+VigyO7cHvPIHo8khhyJDY5z3QpOtVIqJVOZxfco7yvBZneecqdum0STvyK
9H8zUw+Sk/uzHxdSMLt7dtYPLmLZBNPxOHgyBF+ZuIHdGjTrzQtmLym9X9JcSZMV
S+2zhD7Sto24kmUuGYmIqQMzknJilwJjdEAVYM8Wst/I/8BqO2CV4J+LOZF6sANw
Oq3TgXK6MtCw42HHT7ocT2s5hUkdQ6bhqhTPLyJp80+Qwf6WJMmYcQSUAMdiOjsP
CN3IbGoEVoWHWySXJxc2av9YDoArXRSFJ+2+j9/qJKG8mhcTnmbbki6RpUX/YLab
MtqC8WwO+dwt8qR8/m7rcv1CeVQgCVZKT5wSvBs+9Ndb4DQIfUMBLvNimXcsOZNi
iEu4J7iZ0d5IrngoVw/Ma4c3WajW5TBwA+h+sMtr0iCIrtZXgj69XtdyQdqkKpIn
f83Hrk8+AHmOuZcxSJyEIfSa4yPwvy+b7kfI4O5Q/OFnURGEIZEahpKYPlrkXoAx
33YCEUrCCoiiXngfxcag/5JoACm9DyDAu8CgM6vfww81oajw4NlRszBd301HF1cm
n5vE906n7EkT5zr07Nm2u9J/SHHO0eP0owCfPBoVSLTn2QsLFEAY9Xoi+/Wl8hHA
xkA6FvGZ8vs9QfeQCc5a4/aEAgVpo9SLbFhVSIlHGVqBfXmL+YrtFfKd/mhWysS/
1d/VzDMRRNx96g0e9k4FdTsGcD271U2yuVf/Fyf3VjEdSQfu+oUcVWoUfrGguSbE
ezyWSEhUJA1KCALEJblh2bX9m1mIGdBl4dz6CBh4J5U4ZK5l+6Ed9HzNnfhNSc6t
a58H8319NdkUyXCggXLoMScEY9R272i+eNXYemitS0dlZjQNfTu6zco6ckCh6PcU
M+tqwE7gNrIKNY94l+jDokGBXKizv08LeOTJ31O26gkYbtwz5rsUrCxSr3yeXBO9
PdA9nYioVJQwtXSc4jRvMu0himb4FK6XzXjA7X6AbJfV9bDBRMRLHc1oI50rRpaB
`protect end_protected