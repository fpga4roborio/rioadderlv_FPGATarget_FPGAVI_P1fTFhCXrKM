`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
ddtXksX2+yylW5zu6QL2Lhnb2d1sD00763mmSITNX595NcHTEkwn0zB1Dry37fOW
FufOhVzEJp80NC5qZ/+F0Vk7Ik02dIR0elf3clrjeJRK85K4e3Hoo4xn7YbFUIms
l/8VZSb14+JVGURjfswrIyCUotIzlzVYZ6gzoZwDXIi5gQIBf/gI+KxNXPaKV+PQ
Ufys/12rjO6aI/pPlqSm0hCvftmBcnezN2hk1UeXgOIuKZnogjOsf0iJVX2aOOWE
6pD/psybjbnsNB6kH5uFTA5frkzIzkzl5d9+YDm9OyC+k84E83I/7/j+rk4L2dah
QJOvksSIzN867/4Qt8qYTQ==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="MvBXkzurAa5VTw+1JJ70nePUfoQXBvZOku/SMmg4TwQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
oRtzZL4VJ4iwysPsC8SXYCzXS8Fw2gtZTOskLcDV+1B9Nzn1zTyNtlo6lNICRmmK
ZRVu2BmCc2G+fmzynYlNTnSa7C0Cuel6FYpxCBlOuk3OF2tzAmLAuDyOH3Z1Yjzk
a0aHuoCdIRKv7BrZCdALt03JeUmXKPdOmIlkVGFl8yw=
`protect rights_digest_method = "sha256"
`protect end_toolblock="Jn9CQpRhJt4rnzZPRk+dOpzAubz7omckX1MrFd4p81o="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 5840 )
`protect data_block
gD6l00tciPUa6pDNTk/+t0OO0nC/UTtBwLB41d4inuAUA3i/ALrNyoJVcBnAmEQW
ptbcNp5fxEUJjnOxnedyZEuEBxWRieZFQnkRdF269oNs81iKZawHwi+FHyfjdxUc
viVqhoAJ9sXTb+Hm30Bz0x7UauWSpiWvXQYGdNFn6V1lcoxThrXThLu/0Gjg7JRg
HakXsgMCHgpBXqWfs2MsqXb5AwaMzwwzt2QdvLriD/5aMTZf/iWzcwGyAdfEE3yO
fEYCZX91fIRqo1SkRVou1TTQMD2bdtlVOdshKQbOQn/bIfbLUkKgb1gwvRPkBQIO
3gYVD+m/yWELninUOpm3H/FV8Frda5eKR1qzNL9k44+zH9z9TiHp76kaft1liktv
89vTI3+VyRPgbO4YQ94jAel/qBAHz0b+FqFwGbcwQXauwxLV/VgnTVGMsT3BVl+/
rtimI6dSHPTgt3szxFxA0yrbUpxJAkhiOOdmJynK84rzJg+hYD5K1jrQRiRf3tcQ
W+hgIS427FTIvPrWYG51yjkrnYy815jeom77pVHTNmoKJjuX+Vkvv/Pr1z015V/A
6cgkb571rxoqDxM8MYUtlFTLDUxluwI0Eo/4z1ZJb70X0NZmWdjh0t8AeB2BOEEQ
hs/7EeaBUUOHnQ3tVc+tfuR2zGb2pSowudr7jTzRQ8oXK3zXV81HC0H1vQLu9UIJ
I1VQsKfNv/nGTTGaDitIoAb2c6dMm2lvZYZYD+NlivVA0vhu4OkB87miocC8+lP+
xNRMzrY6Xy9CwjJuL6CRkZcortpIkIYdu/WTgZv9hpuumHzLgi5Orcoy5CIyg9bc
zH0K3UISPE8KdkVRhw//Dq4HdtJs6eHiRcN+Zf0XpNZ5qmPFAfDS5kYpIVKvJASp
sEBTuhOALFCfcwyxmnXmWu2HMy9a8oFO0tptPtHLyzKSpORZI4JLaipY27cHD4FY
mu60tbIllJC+vEp6RTU2LGHjfAidKJo4SX8nJjvt/W+84BOYE6zrVxCGaRnq0Bl7
6/FzjV64cdp+OEpSXdWA3Ek/SCuA3gUjR4+D/rFBqzOrUysOI6Wpr4XuLUpa8hTn
pwzm6KllEzrPXFs48QM3l6CwSpiCNqSpoqPwZ9z19gg0F94q2cpzeEA7BIXAvAS1
8qfozXByW8lPuKPEEAf3pCNVOVbZ3MHnyCQbN4UvHILXO8LrnX7EjG1ti3/zdw6F
tBr15uYygVjSzHoPZeczYkTTbv1jcnMTHdTf0qVCXpXDNu+saifaGHOZz/31cft3
DX72pHmLi4+he7ww8pwmWgaxo5rLdsd6XiNK29ZNItNprrJQHj2d7ZlNFYhzNt/7
8goA3t8NGstxKfMayXj9epcAAihG7SP7+P09L23CW2I1Tku1ted+t7v5bVa3KV4+
UzvWeTmGSQ0XeuvqF2NmXZvVad5K9ywRjltUhrViUUEhadL5W4N2z1RcVq4drf9r
f4EyQ0OWg7kkNX4Q4KXS0RJe9I6ZWD1ihi3Q5/ROkjpSaBkC2I+8epLT7MzBl4z6
ZIS8Q3yKE0jt806kWKylmyB63b44O3R1Oe7hwB4PwG+rzH+lQwU40S6ro/KdXi0a
Fyr9SKAmPmDf7b9Qj2nDdUrxY3WdjeSuMU96Ln0LvkCokw31Tj77Xw6dwX1p5sEt
Zcnc7JVLg14DCicImNcTUQ72NVCjkmJFoqc4fwL6wTWjGzo3E+55jKSlJVZDXRMJ
WWlm+fQM8n0peOMcqbyWwNxTKwUWVPS1Qlf5eSh6f+QF/tMW2zFK8Neiz1c4urp2
i/DNa+4069f3amjxYmMj2CdBX6EjSQIiLlgiSw57wU0nw1C/OJ86/MW5xNgCQUlN
Okwa6XIv5OGdoDGJBbWgRCzhoec2h/3A3OfV4OG5ajmrCRQvoRO0qklb0TF5uD7i
Hac0SdIaN4UGIPq9zFWxl+YILuDhgbIVtCuuQLvryN67jgO5w1HSRNohgEby/GJF
HKDJky+0CQJjVwPSDDYY2DrflGgbp+Z74NfD4DwKhGuzPWnoc5weiinLCN/UEodt
IWDrAy6PFIPRY8w1ldrpfnwyTMrtln4z+TZm34Hs8Hb11b5hO89AIzgc9N6ZHg0P
Dxnos4RufjSAvtbB/91+QJxc8fkKNaMezt8ThR+uDFmIe8gS4icTwO1tTz5mND/l
6w/Bib5pEAJrBWelnFtEE4fYVz+56nR7u/H/X0WAmnRb2XWKk+w2vpEDN1oLM8WN
afw8iIQ9ZXVEwIBsytxDZlUlA3ZNx3G+XbvOi/D00haO6rZEiAVRxhVFB8+dhwxF
Hyrg8L2McNYara6HJCCqEZYPY8hK67+VOpvWrS4wrWY3UzG/ViJJh2k2xvEhHpKN
BPszEnyqty/vOcFaaDYifMAevee5cbB6g0uoDZ8i/mFZyIcCQBQ60go3H4hocO5T
y/9pR1sZ4ozuEb/6p1YCFU1tPJpka8xVCHpy59VBDI+KZljZTeLk2uX0X+Z+9xxi
j93vNlXlzgRHmVgJxfWDdGEIQsWdLgB7BhOUnU/jBSAD0rZpJFNHBw2DJXGKSePC
iZLukGdJaRU5ZDaZHHivAIx3n0FiWGnQOhEzYjh56AmTieKunQaQ6fA4d+KbT+H6
VAkhLiRNFE0YPp9uuqA25CiMgen4AMSjGRtAxf4hlCHkv/961b/C8IBd8nMlq842
/x0ysOFxXVZ3I2Y7gImKOyz9PYLCZqvPeA7ex2+GA97tJ03qiT/ZC3rBGqktBcBf
afLkDQ1my2ES3t7nlG+qNWQIE5NCdPML4hgL7+y2zY02k2iwace8q+IcXlJw7d67
EM3DxPKZQt/ySYNlUr8Jx/+PZp8b5XHkgRBgz01VBv7QDazi6JYV22ZK3ChHSErf
MHIEYhnqf1CVc/OZXboRK8OCa3kEE3fem3M/hds+qkZaKwXoZm8QiOtkXbwRWM+w
6iIWuxPufzXhrMEr4kkx1/BJ3/cypMKwkKsLvWrYK/E914FJetvXFxkwix8Y2hWC
//P9GPUoKU7JhZLwxcbRjC7KfOAgp4CBH3v3BWp4ihhOjWdMK/o9H0Kbsml9T5Np
6Lba9s2Km5tu8R+rpgKfDXVyPqPWV+/PlHHfnk9C77XvAqHsch5kJ8v+3JWAexc3
Y+6ABwc8hUI6jNMXtEH1ShksvaFCmERASvb6bQ3z3SFukFkOHTACCMztA0pGepP9
1pfRp04kQuDc641nFYpe/5qVvnwnVZaNoR9Mb+tdhqGKNFy8jXk/5QFVWAYNzNyu
C665JLxEcjrUy9+4amPCjI3iYg0fq/G4Z+y+rY41DFKu33veF5HDeCp6b/stQIl6
twlGlOsr9hoLtdrvFBM79tcQPF8ptZOwxJiVDWxqTJ1xmRfWhF0NCrHgrwmC+4ia
2Cp2N5nbmc6PFicoydMn3Bw2+nUz/OwmCsmJR29em7SONJs8UQAGNtFHgLTXXej6
LsE/S0Kn65YTyOTzht9jjSFIbL6ma/zEXnxH06k7WgC8fmCfgQsgQPUkvhP8M5gQ
3qddjN0ph7weY+YIkyx9cwsLvGUZ2ryzzeZ9NB1hhBcI/j4VGEfB+CHyLrZa/me7
7nOL1maiGmsw4IQ6k3cN62EQgjpO7eBeNpVQlUv0i4AEm46Uvu5hfTUsClz++mws
Gp3lCY0UreAz9RC5psp6JsbVqje5e1U9xLGx+lVq6wnIf0HvHLykDqRjCURl4b82
JOLyzD1HWHPB2qz1RGgKTQwk3pBQyOeX//McurWIGZRtTDEk3PoOGyjLW7xtN3vY
GnPYaQBVYE+bQwfh2w1lYwhStAXOj3T4VP4P2pS2QTbOuwxjpHnFOCkznzdWSKqE
yCUGCuROwbBZKofAuPScFA9yhR4r5y7l55ggbXWlA/IXPYYIFHvH1oEQkM8jBfx5
G9+QCPco+2zsI9/q54+GTCZvVdGh+0PlEZVqL5umJkXdQ4tw7h8msE7bBeYpCG8L
5QiY1l1JfndaXFImb3XRV2Ec2vVT0E7bYxEyA6hD5xfcNH04MC0Akl5wm6iqK4b/
EMPNc2oIkdqWq0M+ZtvREHbmKVRcd2qWFY4Mhb4N2pa7q/+KueIWeTlcUaDkFhhC
gOV6hMkYgZPfbg1cQLeob0pSS8X40rGrhwi/77KE5usL0T62706zV6CEOAwYcMVu
fcEbIfvZiotPXgD0+JnMekxR5x0Lua9q1R5BF8JfF5oMWwuDXmsQQzyDpa3KhjtO
4gw9XTBVrVOZLD/dHMx7bzNDq9ZFLQtV/imx6t7DvifHUIUMV/Faxld9t3Bg0OpW
c8nWCiN4tvWuD6xm0iaiauQPCokIisnRZ2rEYtE3gT9L8xLVUUnrahZJT+amW2+h
LOBgseBAaw+OZyjFVKthbJUm1Y6sGF576S5iBSELA3EWMsYI40yoE9f5cgWDuuj6
ifk/mhQ8R/lzFuaduHtWDUPeMNtSOdQQ84fltuGIUeyOHxTEB/eZifejYai9yZvT
GQ3oyPdKcvCNLSs7hSQB5DnWzavPcqwcNhobfgtnT73aS20r/76ExkM4HOUszKGZ
7NtgBUN6/ymRNxBF7F7gM/1OwZNA2nyzSKXR5aS3RM0ktEzypLaRTQHn4U48Gpgq
2wnfKTkPuSpWvtzZH9tUK7oEyItgMNQGr+Hrt0RthmS7G4JrAPqjD+YBWe0jth1N
gABWLtiphKRg9H/OnpYb7P4hxRG8IQzu0uIWVr3cWsD8v7nH9D/LA6pOn+TXmpbc
67IeLtpMyNMsHihHwkFKkV4PsJC4NiTiByEwJ4y6RCBAyxYkq0IJnldFhymo+6ww
2JaysrOlNMiFMuPDrlKInSCbbp+v5hvgM4M/FBI1ZW2X5toa8O/vmYN4kD2vZjdS
MNPDQ63BFyNaLVSwDVZe0MRTa7pwm1AVnJrZwoxTvECtItK62QKnRXZRFT7B5DU/
bTghdKRwxi1fn26CcOPJYSXyDjTBEAuacJl31p9r565Jix9B8hEP4C+ByHQkNQ5e
8rQE0zGjBTQ3kR/hmX09QsrOvwW7Y5zy1nJPkDz7aRetO44OiD1kJacqEXPJxcTB
1aEbpLiXztkWxaSiKupuVJfDExJX2KHHIwB4lDNtenIoGcroD0mxo5GCI9ri2Spl
cVMWRCDjStVamAsTNdNVXicbgxFCD57Ws1dfrGtOnlzTHY4mA9ifVWukosKz3JKm
mCe4Y7YaTX4nzz9ImU8jmTar9bI/R/QfQmEjEDt0LjNpWHqtjrv5gY0jJfRZgrut
j+UodN1m7ipdZe0YN4miXrYlUxMiLvBJrDC9HG/GyXLAeXsoLyWCt+pjlW96GhtJ
f+W+t4WgPw9rxc5pzIOGTi3m0LAhck2SH+c7ryQn/w09Aj8iE8Z1703VUS4IcBVv
/Fj3gRuK/4z8UEhjHjBREQhv72oso5DTdev+xfqeP6lyGsQpqdchhQkdRwXOU8Tz
1QuM2fxW7f51WqVl1AoPYKhIuSBCbeDMMCLEqPYnrw7Hjlk1GlEP85fcGCmXkwLT
kwn8pXeqPRXZvAahgeRyUbX0vDi35eCQXh820cuvWTPBvNGO1nm3qM3QRzHQuYa+
i77CSznls9QWOsnDFx5pVh7SvSaJCdt0Ef2kXQ7RUGo/Fku1mjpUHJHxfWXNLs11
u21Cd2sWwWE41JxM7H8bE9u0OItrBKIVi1NNotKF/bkvhesI6legilnX73i3gkrK
hWPzkwlyP+IdlPoR0WW8bA9xLomePa2FMc7Tw4+oRiXBmXfU48TRXoQWTK6UL2sO
3wMIXGIuY3RWzukcdufDOZ/9fU3nCuT0uGAHsMsjV9e8AaMqQU9agZQFwcUT+PjF
MiJsu8TCbasccVgLWXUv6/HZFPm/9IJD75VspLqWc8KSFU4FSwnOB1ZgtRM/xPTU
Sfz9lEI+O3BuQKGMDklW2uD3ZXDXqyAM8aU+TPkluQsPjWOp2LbHHzfDvn38LtrT
8ml2yk7Fy0xm1f3WVEKHZuzcQe6+2XS73InwITkXdQORwwpWLZjCAVAc6ofwGs+d
xawUf6eoqkE2mO2UTMPq4XF4VMkgj6MS/wxA8afAGzAtXrK+Yjvz9XSZe2Pp9+SY
oxxwh6C1LpUB+yIxEREhayDFWaf+ybOnhRHroGrLgJbAzIk/W45j8hSh1IbqWKQ3
7TCpn8tGWhO9tUXjdJF7zNyNLml7HJD03/d8vDwj5mv3VOsKJTPL1SXkxinrWPSn
Dzh7elNKLwJDkFPFmYUghPxEHqhZWN3P4Aa3cda2VkU1znIql+z1DnNJ4Z6ytvgV
HsqFzym5hLNAmi9odWp1C0EDXaFY0yvNJgS7GGgqQLsUaVthLExWcZvMzK7jp5Ey
vrBSYpZ3yqfBdy+tAQsHLP5eR8D4j5TaPsbo+VYcODoULiech/xgEwrtZv3RojAT
L+axemqzaYZzHY0WJPMl9Mcc4++842pXVsctxw1hP9hLnkBEa7kMcW/QSCXE8vaL
fDR0slCIzDnsqkWy0s2Pq3iloOyQxjW9pode6oAiTd3XVJZu0q78G3MGDBA5cGOf
k7lK9D8TqwkHea2iXYxnyiyJejUWVF4h9OWor0PIuXeivxE1wJC0vt93mWElGZWs
dD0VB+6TbG3iEG1AreWEHC/Fh1xLTXdfCfv4rokC5/vW9XIuXqkUzKzsTHVIa8Vi
AknB3rnAYzP3oqjtboQmAGZKA68/DYcjJ/4du1UACaeCj/zAR2NXjH8275fAxSZf
Tn7mdLy6a4boAKrHAGLcO/NCROjnilvkpBnotXtBFNOHfB3qMieCSvUnX5Ybj3+s
OxmCGWpan1zfGbxomau395ggS1eMawBfbeDCP2MzBoKs/S7h8DWJe6XDDaa6H9m5
Xli+HYC/9mY89YAEA2VcyrVZOnUkvC8gGlIHdQciod/hk2kfUFmA6BfwxZJoXL24
gPp+VWkUwucK5xsGbVjSM9pqAjkXBdd6t0xeg72Fg5K1hk43BLvCdPrI48tGW4sF
Vi2kfuz8YgdhmNz+nCL66ftBTAVmUk335CG1rK4oYrRk/II4VY4wtWkYZDNf1EIL
e3dfSTsj5RkLPK6fYIHWlrPQ280qLhFblu4gwcEGYMbk28eQhTZqUMXHbxoyrNyU
EYmhv3Efu3wsY1Lgo/saFsibqLpstCmlJvUOK4VhzVdS0/r31QHy8OYRE+AcbnFx
F3L3AlNmDrPXrDfQd9yvE60r1fp1Z+1AMaoXIIY30zqxiAI14zVze3EtDovejSp7
Atjqeeg/yq72plwAXQgJwiB8U8KEk3qd6/4NUpqcVKcZnpp9uAx5hMzriuxOGdAE
JnOWda5t8NGXbxTbU4O0WkXlqbC4VZIeQQi7ymUULyDP0CRy7QY+5KRqeri3GIsh
wh4RfqDhXwp4hdsrloJogMqsYX9DiY0NvYHMFlfTY8EUmKAJ63S+XdrpsxO4SNOK
MrXGyn1o+ISB4cRYEfCqN/lUzx52jmOnemXxWBrHUM/IK0aTh3iJgVb6KTeHxkJJ
x6YVaKTHQHsHtv/PC4VuqbhcTgUrcSyOCtgL+zAKjTQp653wfOrRqylAxEjRV2Gl
EYmJJsmicxgL4nbhpo/MkPKBXc6rqMz+6JGtM+uUBgZurbvRW2GMDdr7Vpyrv5fa
58/+CIF9WjOfiQSAyHyd4B0Ob3WlrUWS6/+yaAv5HwsB1hSWaHqC6IaJ5W3JSm5G
vHbgNXq8ZNUMPF9PkRK0l85EP6VuPA1X29nYmEAhFX1UcTtoTsOVb4QQFbU242Ya
IP38awiCzqYetGyvkpk5cu8No6JWmvVD0TGn90ZEhKs=
`protect end_protected