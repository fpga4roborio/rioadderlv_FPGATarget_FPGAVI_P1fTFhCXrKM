`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
ddtXksX2+yylW5zu6QL2Lhnb2d1sD00763mmSITNX595NcHTEkwn0zB1Dry37fOW
FufOhVzEJp80NC5qZ/+F0Vk7Ik02dIR0elf3clrjeJRK85K4e3Hoo4xn7YbFUIms
l/8VZSb14+JVGURjfswrIyCUotIzlzVYZ6gzoZwDXIi5gQIBf/gI+KxNXPaKV+PQ
Ufys/12rjO6aI/pPlqSm0hCvftmBcnezN2hk1UeXgOIuKZnogjOsf0iJVX2aOOWE
6pD/psybjbnsNB6kH5uFTA5frkzIzkzl5d9+YDm9OyC+k84E83I/7/j+rk4L2dah
QJOvksSIzN867/4Qt8qYTQ==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="MvBXkzurAa5VTw+1JJ70nePUfoQXBvZOku/SMmg4TwQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
oRtzZL4VJ4iwysPsC8SXYCzXS8Fw2gtZTOskLcDV+1B9Nzn1zTyNtlo6lNICRmmK
ZRVu2BmCc2G+fmzynYlNTnSa7C0Cuel6FYpxCBlOuk3OF2tzAmLAuDyOH3Z1Yjzk
a0aHuoCdIRKv7BrZCdALt03JeUmXKPdOmIlkVGFl8yw=
`protect rights_digest_method = "sha256"
`protect end_toolblock="Jn9CQpRhJt4rnzZPRk+dOpzAubz7omckX1MrFd4p81o="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 4272 )
`protect data_block
gD6l00tciPUa6pDNTk/+t0OO0nC/UTtBwLB41d4inuAUA3i/ALrNyoJVcBnAmEQW
ptbcNp5fxEUJjnOxnedyZEuEBxWRieZFQnkRdF269oMr5q4ip8/t5AXpPc1RyIFS
DXHbMYaJ0nw9308U0t9T0Vzp+LsydUNzQybGM9RmqMLSEh/1g+F5u+03JtcMQjcD
CzyM2BiYtSMh3JnPsXCwidRM2gs5RxYH0Zn0/lLZuPvg9Ylpr9QHuIR0VN8FL9DS
vWk01euUjbs6LM8BSHUsLRsjAu4yL2jWxRfiGHHEOGbA0tWEHP5wbg3LgiM3huMC
G18tg6EjH8n4Ohai8xQT3DO9iv0n2LjoqEb6eQxBmD9yxkOqv7whBzQ/pvsyl7vR
Gx8wyGbWFVkhpf3yU2RKQu/qV9lG07k5Yx6x6JeZQVgfzuikrrwSvXxNNRioW0GR
6R8bxXBc5S3KsIgta45d50hYC5pfwySXfAiN4uMLJmHJ4zwv3Hz32nC+MJQVeHKV
Xkind6HA2fUfLKGS3faDlBbW8kofbnDRsHJ299if7Y1ovOHNZ9UCYtU8xdZWChwL
22coCWNrfTBJK07Wh2jqlN00Pt5NBdH2rBQpr3xPz1/HXPJVCO8oYVaiL6Cagvca
nLF/05EskiLTHRxTwze+WW0EAfzdPlbrbKi+EO1SeZjqD+KgSg+CDAZ6DlbqjbFC
3eP1PRmt/agNZ/uzhUwQiSFDIN3kBJnwjvb1wWL7m+S/etnUrMOQ1Gu/eWoNubv+
IlL+7WIxMbtBDuYlbna1eaewvuF7UV4jKIrqKmQOXyHpvModBCEUCy7cOIV+h6/1
8Vnh3es6OyRQSxfMkW08eqoQxp6Cu0lnlVHfS5Am1oACHlnIqvir8pWrRCkd3VNa
tiqYVT0QMiVrLMtkHqI4VHRJgfcLwfgZF7VzucKPNXqmWtDJWIX4bS9bpCW5RsEC
HMBfZG6AEtjQ2jse4lRHE4h+zPhhHXBa2+el6XrLppvdQUsAraXA2A4108K+XTxJ
JJOTAl7524QXH1k5oyFEM77kl5BXFI291WQtKEFiDLndfyy9mi84wxf66pKfT5LS
9j8U/8NaJBrhJ6XQGFcCzqcIMeZjklSIhHCeOGCca+4eblkjA7Vd/nQPL7VVTKDJ
uPmKkGcRkXBZHB0oagpXTH8IfRGwq92a2OkI/CceQCFhmrhFs8OxI6cAqfkRH2Hz
Vt42oy0Usf531lOBNKY3ffCu5tyNG/coGZiOuZbPKm7TY3jN1tG7A3qp1zndh5gv
GlZalPsytI9rAaXfxoEr8Gf+wALc6P0g2HVqzdhnTLIgH3VgON7ufHju89G6ejbp
tIcE8r/6MprLIEjm6jbqzIaxt5XvAAaaiumZ2Zjqu8Rhu/Ok5nMk8NJk+zvNXpdF
0kj+I2gZKW32vudvSLKwKUuYqIL0swH+UQ51y9ezxozC048te+gtfworyieI5elH
9NvsDA44gpZYtHngRIJ3ZFTVo+EnOYXgAwsQboCvwQQ8M7F7k791nkH+WxnnXBV1
jPR8myHuafhLQDUOv3bQJCaTM7fxJ6D/SK6mdMPo36FBHig3O2+DfLYFr8m0KOKT
rh7HPgbSSJOA2ysQum2tunM6YwovYxNS6GeMHcmBru6IKl5CamENv4pmz6ui1E1+
s2AZrIjemMh5RjXadLPNN/mapGZpCTInzPxIfC8s2bLjEuPVEPCh4AWGmIm/3iWk
nOjxZSiB1+yQZCNNfrwMB/FVv8g2g/fCtX4/AMsmt+YUSntvWeFhQPJvqPaGasVA
FFlVJE9NWTFMFVLSMe3X64/Bl7gWwepetXhPl2j594ipLeRaSQuqDe260RBrzk5q
RnIbTYxKGwabHrKqNyHQu2FwaqSULKAhS+fuXrofBNG9WvlIsgthlHIq6vx7Rbi7
Y5LwI1p0R994zUB/xA/O4VSwLNOUXnriGV3agy2x/NRDOaKEwl84DuYE/9rk4G8l
Z3LprTK0GIdPP5sdtWGs5JWU+wgVP3jq7rHs/ffkXDPHmU/qviEa/T7naLzV+8Xz
ExYAH0Ubbd+HuSi+l9/QjnsCTs1ShVoE2gNsAEwF924zC/Ob0VPGvyGSVjKB9k4l
o5CrVKvumGWjQRGWIym2EY6GDGR/DSwhTeZaJg7NZaBFlOoH8Yg1thyWzCv0KgSe
r39vlTy7r6sa/Oyj2g36nPvQbxA2+cnj626OgIS70yp3MgOE7UlEfODoRMXvEP8q
KhWLQrXbOV8XAaDmsj91JvbWtHanOlIZhBiTPEA9E51NL4hTWTBW2Nw/Hh2A4/4d
fZj+/zN9fASs75T77T+JZw4SDBR/zQhslB9kqJU37tWlgFK/B+RiNQxyjLemNkUa
JrnnAjBTdG1VZoYCV+AMjuqH9loJ/8E43LeLzdz1wPflbcyxCmGfK59WvVBzKRf/
MGQTf2+n9It/6ipyiVYv7lI/J8fyYMUZKB0xpi+6F7UDvg1K6WBJpmKPrslAeHnE
h6sj6HOzZPLACfMxKUuVJtE0fEA+2JraR+ARSwsemI0pxni/2SX/41/SXNt1rq9g
w/53a4PzXt4QcDBh1aPGsG1dCKexdnKFHrLOM8xLQhRSaVAwmyBUbkmqXcYUDtBM
pIZJ0613vi/z4j3ybark22CDglB1LKa78w26R+AO++/9Pu2J/uJw+bYFI8uDvOsJ
CZrrliPtReFX8OD3RsRUPzN12iuVKRjlST9vhuu/CGbQ9wyT+l1Xfw1/ob1+YGb+
sjACRDgsuqm2JkMW5QIpDnCvWPzUzwPZs1pamiZLicfF8f8w7tZXMgpYmc+ymodN
djsIy59DLbvRL8UtqFwepZeJIO6/y3UM+rwWerIRBzs9d/m+7OITwkMFZgqhUEjO
mwqSniVcZp+IIja89E/HjJoIP57jg/6pFuM0ap6qUP0GR3e25ZTUslcZZTtxpIYr
vKw9vWiZVpJmMIdUCk+w41903ar9Kua7enl10ZXWQzARXRKrFHx8QnqAW2BhSF4m
Og5OG3cKce+1ffnnDuzbWIvoOotdjUwdhrueHgkXVUJQJXN8igf6DSMpcurhDmmG
3NYrCB2EY1PwkvITIOY6s9GwumNBsEH3jHIe0aEppPvCCzscalVE7XeLMYzfjSOg
cDU22rOWhmp5NYqSCmruR/SVhFgny4vpiVdbc3Q7zka+3na5nfkbdiyz9Xzk0TT/
alxmXrxGJpl3oAF19PHqmuaq5oB+irhh3gYrCOAAxmVCqAtns+bnoDiHnVXPNop1
CXgER1rL3WzVUQ5Er5vRzHKEemXMteNHyQeGGvh61a80LkEaN2U0wpjwHn4+Sv3t
tgF09BNYM6yvsplKWZC+6iCOP0+pxevFDRHvfDV5mJ7Q9MWcOZzXApza1/SUAKCn
U8PN7Ji3fLqWwomtdxeDAvZX35KYobwX5Uy/qTqepM3A6EdsqddbMS/cVNjBkZDj
o88f77KpFPO6OVbqrgWJm5wMvkHlD14rs5AHfe9RIs08uzwlpL0A/FA/PbjD0K0l
/aCBtIZm6WKlvQ/FOvrReEsyaHpmGPp8NpP3RCkZQFE6ireJqWgLQfJuNIU/o4Yg
a7QfMBy7rV/tpjqCBOoIbdlAJ204SPyivmimJkvlyhVLT2bZpdJ3eZrt9XvmIKJ5
y3fojPUphCbGqhhMEqHZi/uX1SWnZ9dBSmdY5VxrjJm1t7scVxjrpmoQEsynhuL9
/vWAk+fUcuzteuzRhbOelr2cZhD8pvhJp7IdkB7ufmYwmy/JKejn+O3b8JPb+14u
6OAOvobL3UAkmBQHi7LzMyUrxu6moJ1z1zeDtSOXJhBowRZjNslwdDZYFgG0ilp4
GqcvAx/b5ou2epWSHMdjLA9oGkuPRhoTZ0X/XS9G03lioYMS01eCxdp7qeSNBiKg
ONSaiXwETD75puZepcW3VEcJ2y9gSgRC5wjAx3oX6Vp1ij8Opt0/Q+PGxR/1IcY5
Auuk3IAP7xD0SPEnrI3y+KaMNSNwTdjN2w1Ck1wSlDavp7mVHFACarOF6ydTAkMb
GocNNOnHPDL0CyUDYCnnT6OwlWNZEC1O744drQ1d3fGNXRk6PfZrqNLsE/FymHaB
pIHOHdYbgSeWQGnSIzoWeWeZaLFB+2wDxUCWWlMGe7JQ53Hc3lT94URf+eztyYx8
uUeLBes4xCeO2O6vcUWTwOXwzzonIAFlUw5rp/jfPWBrylWsKvMpv3By2jtPqX6P
qcrrUckeVp+SmFuOkgQX5/geUPkTn9cThU6pt8avbSdSRMuGW6ws6eTSPWLDRKu+
iM/fmiFWaoeI3pKj5eVcznJR4Lq1PiyOk9YD11jGbXuI5lv4jRyCRznazDIJMp8M
zDdgUfztDpGkyW1nFysTu4nWE8LkKcCgCAbuW2UQzmR/7IKP9xhG3fFS+7YNSXQO
I9tD+p0/UIRqtVKw5P42PC1qgHz/5orioADa1AVGzXJWkQ6YhIvbO74u5LcxOe2F
1mzkZQDsd61hxOdYw5zSX/kXngPDaySNEptr23okrmONlyDF7wvgrhrbedBQH2dB
AYRlBYcKk/tQpBE3tACAv6ANYknx4TA68r1gDBPrUafaXCAiI/R3LdZH7BeSMcjU
JSeI7JPkKphHYllQhKzfoJoL7sdg2roWs8J9L295SUW1ig5PO+yazvmatiWpLLeW
hBVbxO87xNpzjbzrrkMh1dNcjzUNbG/HJ4Sd6J1mckP4Syb6AeGLDS18eLxqofLf
g4HaEogreaxffkSy1UI6amnShwSloo6SlIqt2/jKYfYsq7snB9p78L2QkbkdaqtN
j34gBgSWP6gH/n6L0vmhc27Md7/EstMA0zWY7NpBVRR55XY1lmGaMfUUoHotY8uN
0PQNUpY9KzyXFoqRxnwYAromgo65wpUAfpheB8tgDkG1HN5i/AGeDX0nldgDIIPV
Ydysif37p9cF+haFrOPUnGojKAOV6i8+5hXWjSGivLNan7KN1uql3XqM5LAQ8Q6K
IkfTOkEoeQljg7JOzcStnQT7TzLyM3QRcVqfjwqneH2xsKC81wSRzsDn9Vm1VTW0
A+XV67sTYnLd1XdTuozgrxk9fnkoBZ3PFJyTwQpdSI3QonTr5R9cZEutEphwPjrE
MzN3mF4jalziLviBGsxSLwHwQb2A2A/Tty4sFatD+lIDXkWSv9gN8y1K98W/PVs2
h2fUeQ8SMA3PAounKViOGesu5HOE7JJb65QxUGG41lTcvv7OF6r3PYat6rZ3WtHB
IAeuKuG+KKGUblZsYch68/ooNKaqX1PjbuNL6iU/fp3y9ZN1v631NLVJuE5e2NDT
Xo6hJtdXWEJf/67MjFeeAl9X03JyW4HaMX6KABq1B+Zgd8K19NrBDtlp7pN+iVFU
Luk5yKmA+JRXwSYEO1QBeYxieGANudZXbOaXFFFqRasjUcdlvUQh3TxVRxp/d8mn
DjSoIuHZnihZ1E5gmTKjNA7ZijGX3lzu7B8vYQLsPGgnubnXbuLlCdCp24338Ihx
jcAXU1t+wg6BKzzZusqJJwcowAKYZpb76fFRwxNsuh/wPxzdg/QS+U14mHJaNjIS
XKnTVdAsLNAm+Z6YvbFUT398rt0zcTeGsWthjCAsAj1Zya0vTpoxzzAaKXZK+Exe
QQT5HK+ZPut+4A0LXAuAnF2lt24XrIynuHszUSss6DLUdND1xCO64H7Zn6D9av+/
`protect end_protected