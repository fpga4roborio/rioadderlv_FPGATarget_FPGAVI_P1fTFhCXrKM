`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
ddtXksX2+yylW5zu6QL2Lhnb2d1sD00763mmSITNX595NcHTEkwn0zB1Dry37fOW
FufOhVzEJp80NC5qZ/+F0Vk7Ik02dIR0elf3clrjeJRK85K4e3Hoo4xn7YbFUIms
l/8VZSb14+JVGURjfswrIyCUotIzlzVYZ6gzoZwDXIi5gQIBf/gI+KxNXPaKV+PQ
Ufys/12rjO6aI/pPlqSm0hCvftmBcnezN2hk1UeXgOIuKZnogjOsf0iJVX2aOOWE
6pD/psybjbnsNB6kH5uFTA5frkzIzkzl5d9+YDm9OyC+k84E83I/7/j+rk4L2dah
QJOvksSIzN867/4Qt8qYTQ==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="MvBXkzurAa5VTw+1JJ70nePUfoQXBvZOku/SMmg4TwQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
oRtzZL4VJ4iwysPsC8SXYCzXS8Fw2gtZTOskLcDV+1B9Nzn1zTyNtlo6lNICRmmK
ZRVu2BmCc2G+fmzynYlNTnSa7C0Cuel6FYpxCBlOuk3OF2tzAmLAuDyOH3Z1Yjzk
a0aHuoCdIRKv7BrZCdALt03JeUmXKPdOmIlkVGFl8yw=
`protect rights_digest_method = "sha256"
`protect end_toolblock="Jn9CQpRhJt4rnzZPRk+dOpzAubz7omckX1MrFd4p81o="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 52544 )
`protect data_block
gD6l00tciPUa6pDNTk/+t1gcgy1iCdpjTkA/bOvU9JA+cpFEv5u/7dp25hHk7lLT
6tYtR8HgwcLXTcx68BnPlzdPHkVIv0lwXo6yhFVkYlDWBcqD9ubowgKij0UjlXmV
p4anbpVt/gKvAYRDYe8Q5F2CQ8AIsxOuOcJ2vhCPchS4QF3n7+oG0MKU5ZyzxTu6
JChvV/PInGqVYXshPMmGODJz/gvrQcP3GPxJYmgUbGfi76YOeJ1g95tjbcItZngs
oCmeHkqAEZe6WtZmTsWwy+nm+4G8AVih8EYfyWS0aTejTM4ZYxPj38KAS2aQGPLj
n8a2DUyBUcKDKqOhZbPxKklZJ41JL+dMl2Jn71qyTQGImDPX4Shktz8MLB8ge4st
8nJ1j/JGcTmpKWvZZADhZAbMtiHjRJsne8Wafp//i+Ooe3CSBBMi8qK27wJVbxfJ
pFoxHh7haZmckaQ+40S8anb5qHX40NJlV1SX701airCSdD3t1PAoLUiXbarVCiqp
NR84mrEM+F6OmzpuTQ4rOlbuCSB16HS3JtjQdjNsGBVyf/LF321svTs9ob3rn6gn
VKV9QeLyaVhR1idbTVP+N6aekvl9RbhfRzujFZRnn0EL0kiE4sSKok4grpLJ9BBH
cVrLJiu92WYvwArQ6em9JRNkNPrl+EuCPry+zKUt7X6/gdCSZoWSCdVAyCd64Rvr
q+KqzRwLT6de53IGN0UDx2fQaocsgkuLTUTqUM9S5VnEbCsMVocAb63FoHxL5/Ov
gzqCDuLprQPVMc2P8vkzEfL1SwMgILdGv6JmH0Dztnr8z2/HmjmmsHFVXeALR/ru
DvWih+HhcA7cqACeLTYKctdJRNvcA/CxmGhNtyGw9CDkcuKpp2Ux7xf2buW1VDmQ
sQVyr2wpMwLVnjaMisVdfNZrm3BaBhgkut7nShFACWSmg29j0yf0LJB6MN2SZs2+
Z6JIeXDsZuvK3W0GcUZIGmMr/BdwSl2WezdHRQBY9Wp/K0DcYi/sn9Z/jc91p8q1
PRAaxnvW7B9e8gxzsElJhKeL2ObXa6Hg1JmGYDDUzzdqVtDnqsNop6qKhy9vqSWo
P0h9IedQEnic8n+eGNOiDGDSXi+M2S6SgRFnZhUN+4r/EvSZn2J/8diCk/dAaGy0
jCvYDMtzzjEgrnKv2QwinhZ8fE0NXES1rYbBdzrY4FWCjWVTPEZd/rIPNSw/C1UZ
DAy0vQflJ1GdSJKGd+2C4gW7vFc6CElhAR93aE4MKtnZPnAfQ3U6op8aAO3Cns7M
Cs+IHNf+QE7Qopy3fu6glcJFEiTQzYqkoBCZTao1pq639bHITOfHQzy4Jd16JT+b
bMtYT9ubuO6x1Q8Lrhg0HMyz27fB7HJQ9LxvY+hjlwDBkrsM8dfi/uwOa6bxt4gy
IgyZqTgzMGGMbvmPMKZU7yLacLdwXAtfNsCVMW7+5B1mDqrcQd7zuzYeGGtMOm+K
40e8R51pNps7wnk4qFdzGtLog2exQxdbccgZrGqxyL9Ck5O+ITtq2uOx46TOfc5s
9Zno8uqf1UHkRq0p3sGNunOh+q18waWahhCXUpwDjB09a/vlK+MavSssYp5p8+8C
deZtz3D3DtwsNJj5ureQXvnN+C+7lJKBQPJFLRro+TcTk94VJMPw+XM/BCQ212s6
1idj8JQ0qqpdYyqTnW6TnmtHb20qnPkRNW1ewNWE9hmIpshzbUPI1SEmzHe8PxDP
G2JvtkEhXYPatdWB4msJCix3NMpmRZQRTOaRNDc8If3IlfplM4rUWaYAhIrCAEBt
L/uiIBkyvCwrBlEjTS71en0+D+s/vFcw8raotvEu/9cKUVfjPNGFaMQa+RMiL9TK
Vt4Oe5mUXMazFZf6q9Bnwb7yYXP3ylYc4B+ztdb3cjwGSwQpjpbhr22nSgeKRbfz
mZT5DgtZf+5xorKxHX10z3tpmhlr/byBpg52RCHUicPYDUVH84wPb+RKaAgFQ2WA
rpG+kWGzR1QZEmhlPIp1X6qCdzPHNJ7yuazBYxJyHvE1uPqS7/37GRCdh4Gu50Jo
KHRFThcIzdcxdJ7IqTVcCtxhS/KEeWry9YF/Hq6hp/QnUFAtEDau/ZQ596JYXVXI
ftm+7WBUe8IUEPaPeiOQ//AFjf4yJCLrgkSY3utUwjyrjZkf4mGT7QVbsqmBFox1
xUv54mZ0RPS6TtVMh2cLco4j4C+2kVnKeuMkVcw0IL6npRdRNAck58ivef7cIzbx
+3SYdlqdxHSb3+d9K0aoRm28Gq+DYV/QQX9jODFK3y1ihesUgZwXewPvDtVHJeA6
TvxWwZp9JqLwYM94YHLnbt9u2bFoGT/ELxxRD9dwBxD1stVmZUIqszRXZ3K9O43+
BVkfIL5evuDWiljeBWqlnP8AdKgfaGQrkiSxo2ynNyK5D1mCjttFf6SEMndn90DH
Ns8hb6fBE4A9bQuT6rimvS0991oMAnBaH0V7CLAPlscVwDrPHejNXSRPlZECw30W
pzIWfmmrxOb6fskGIiBtKff0gcLoPEwjv2SIpo8ZYzhDnlLAc6CFbdE98x0gh7+d
6UIFzEXv+HGrge+fONaRwOeiwISqFvGLC1yZxDPvmzntkgZfqd0aiaJ0wUVWzmQi
knZ662OmRRhFruvUYXEFS8pb4gr9NK7+1BKh/FP8/MNXxpKYCtndKMSb0DNkUSg6
ho0AuKXfMkn8F+dKknI8V+pH8xEW/UPrx5tVKaSl/5GvCdjiOUF+IoGV1kR9YSqQ
rCOFz/bZzFJBJgLEyLNALORx0dOTXigW3ZfqBwCIZwoA9DJ75fxrtNJOwOPfhLML
k4oPsFeUw60dtWsS3XHk/FBtghOYy0iRiwF0hFPwcr+iwxolRDd2xHdcWdg977Y7
R7PgrpL414uGZIebBte5pAQ7L0tAb1zsXwSdNFG9fuDPC09K7yc94XYLU/0XEKO6
wcPCotATXp10Mr9y/LANwepwOUZWyuk6vyo5SLUTNw9Y2mWMp3bd+hr0rSlc3gWo
CjnpFKeEtsHMnT4VmybTNrLQNHGbuB8KkxzYa0DgxxxAWP8xgYvtz5cX5D09SKj1
WOaLT7C3yZPvicA09bhGTZUJkrTKzNkqdic48+euK7SwGmNAN4akMYGBJ/NHvGBE
4VAQgZJT/xhDI4Pi8+7yYJp5pyOjkjN3Ts74CphKUZBeqXjo9k4VYyHD4IOEdmAM
Po4ycsXFgeDpErt5U+UGK0eavuqZv+Ha5oG9xWwfj8ZLzVj3U5Pfoc/sxFiyD70g
MnW0U1hh/gCExTy08FN4e9yBqkPwTNIDl3xuBxg68/BxUwKHBgevfoIghuhFYSxT
WLr3javIckIfOeoKNv84N9x+ELihpRXVKEzbeYpqU9sTB9yzr+1615DgtvB/CN/3
PME1L1Z2TvtGQmNiXOh5b7jzArgzHbkfr8c7GvWKNIxyLfCLSjkkpBdEoufPruQw
eAK3zv0vbagXWxsjp6f//3lAFt0mDFo87F+S/1Js/blgo+zxJNWgyNNMopfMfkqy
YkCkYNAB/YWKxYPpdWSx90AjqanKJgwa6fK4NXr0ABWAVOO0a0wkj8fWg4jqcGUk
Xg1KAy2k0IkiizZ0Krx4RhshMEP/P86hX6SFdzWKrtl/EX+AzUxuTM2gvGMRCdLj
4T/oPPjFqbF5pL9XWn0Om9dmDRou/Y6o5EXzcJqj+NDOa9e+Et0sUICk5MYccb/e
zJTtv6uOr6DT55B3MP7ycAFusHzNELkVrz2Fl8sJ+XffFx9voKqwNea68yWUK4td
WT3QfJiWug7v0El/hjZXOL1WHtzZefPPXxJncylolm4jaCjVQQrNRzLKbGGL20m0
t/+QlhWxH7C9AwbuJBhA2ZPzAQjGe/zMkXwJLEn1UwO0/HqfI/xY+cEzCZy6CM8L
1A29G4J7lzgFXi2CBEef+plUpyKOEbsCIUiiXBBCFWq7gM+UI9r7cfNHEHgAc3jK
4M2ZCe5rxU25tExKd0WlKbEMPfEcbQTx3mMHA4WA/ke+h7U/u0Dh5tIcgw22lHRa
0U1q6xDyqTwSoaqNmXOB39201LsUjAST4nfix7HHTA18m1tTlYNg6ApmwvWfzTbQ
xXPdz4JBfzh0JodfDEYuwKGd1WY6roBnt6oZ1rxf7+ldI14cdY03gwS35EgtoxzU
IPjJAwP15xKsPcAgZvqol//rF1hgaM4FmjDVfK1WBM/HjERv5B/AM05hZayDwrFp
IRJw9LdH+mIBO9qq5zjZZGZ9Nnuhnu56H6pKM0Tnh6nsaI2Cpuo95dNqj8BVCuKc
4R/6s/3u+3PHmF5ywCds9H32g76IGWBgAlKtVI4Bg5gVQlaYzUTBQ0Oi2bQA9bMF
2YssKEe/2FAASHariJyZIyCjqr19izxfSbdMJiqBf1VOrF26eyMg7G+z3m0rjERK
nEnKckBueQZl2D/7o2f4lz4RGVKDclFMrA9IPUnpB/DtpFuobIGM48VyMZMoLLSq
+qGl9RhfzYKYsJP1MPNOi2OO4cLUro2vbOxRHff3rlKKkvqlJjn5h1SFLzhgsIsL
WpNY8i9WX15ppCuI4kSueoizIbjgEgaftfJF578jTctCu0vPmqDZBck++7iByqtU
PBFx5YGEyxW6/R1JjwRrp5MSirR+cGsh0mKBt6wqpdK7DuSosVdKZU2F6DqhPKej
B77Ti9ul5IHUeGDETh0PPO2b2eyRpIR/qVXUuMVrDU8ng710NiSgcPTIP+ZBhNEJ
4dgEbhkOl/tldXOt6Farf8kv0j4zJ7H7dpWYjLHIfeTUvSlpJAefmwkzX0LNLXa5
7cFXHrA8fwIy4bEH/QbTARS23rIiq2U17tYbsfzpXUflPjwsZ56uVKVP4RdkL38R
Ov4Yr3cq4O9L60aBH6Fg8DDvq9Rag3xN4kV9Qd8xG6f3DWqd1Lkgl1B+0WwqLcMN
vN25NsClweAp9kvhuaWv6YJh4joPKpMvdKYNSB+R7A6SwhfEFIVSeeBxdbLbfx4U
DfOZSYHQSPXI0L/kH0pCqU6e45tG7cs3hHoet4E8kRKfiCBNapUOysMZzSyHJWTU
4ow2xN7mtzG411W35VKKKx9WR4v8SfSufnbGppZHog7uFdd9dSsryotkT+AwImxm
bQW4WPm7wImUaDjhAaY1yckwQ0aJYLclApykqtmetoukHRIsY8iC+Gq2s5N6nFG3
LUf+1BuLEhsqCw7QCpYt7F1VhNrXoXZpnyYrwu3LnV6DCrStkIPmQdRe/klZ3Qup
h1PlB9aXZIns/f+2DWPwHkuEly/T8ngO0Bi8IrirM4pWwhUnCf4m2X+R9fCgDtjL
r3lRODuJ2sy7ehYhMgGpN2xOT691Zt1UP0THRsF00VTp/selP4yXvidsqKEPB3+C
V5k2Lj09S7xUKL3OFNFHGGC8mCCF9x4J+BQIPTx21QCvejUaVgPqTUXiOvGJfNqM
lH3J2SLUb3OUSKA2A3b2UNWnMj9xYtA1GbFVIP6UFPPvqdxET9WXgGCAU7cmlHFx
2tiA4k2p4Dbe8RgNfhFTbimaEeCU3gDPMAlUCpkv29OeEL4jJreb1DhtG3W3Kcjk
rfqmFm7rll12x0XnMifla9x8PRX3IPfJP8QQe/LqbEKYDjnvJESxmZCpsRHRSRjX
/Ct0mgyL4u54BYxrS43UQpOiZYa3I2zNTKz0stawZpI1aXMohvVq3jtexGpcJzV2
ByPWhzZD8EuY6oy15FwEzSRMkfBhvmRZjOY99MK+7OBTdb1NCyARXrkPAOn5oZfq
EVrG93EP5sV8S9vC/sobsUYIHvhW/+E47EoRHhWiZ2qL6JrM94EgpUucAG14qHvO
PFwHhplvovrsIZftRplJv3r4rZopBz3cT3HlqdbfDmH7LIDDJBT/MI3ICzyr6JTT
7xGcGLDwTISSnZBeRJGQ27lTneK+tXilnBfqsE1jeW3fUHuAuw2MOsZ72fjqaKcJ
jemActTQicE8d9qdM5vpedi5hrfydXA3w9Tvk1P5iUWPeywZ/wjtaxBhqt2lgrCM
JsFRtdeZtjYbkb0hNvtFAe6/DcRoWRXh4u9pGyMjlHbmaNkIuAW27KwYimGHX7cI
yLgsotKGTpPYx13ZhU8JWeS1iF6cZXFStsjkIoTPbtRKO1UHW9Tx5pMI/dRc/gYy
p/rT0zlZ1ODhonBKp7tki+Hwf2LTezHDbKEluoJIdsoHQFtl2szjb8PCgntlr33w
vAalrEdlqsLAwfE0GmUuvaPPOP8h0ItwL4iPV8/Y5mc8du40zMiqz5m6Rq5hrH5R
i2RfgMVsrnHEwB7ctQl0M6Bc03OqV15T6/+d+AedbZ2d8rlFv1dy5C1Ok5qgw+oS
Oz5ZbCOmPfPSIg6C0MBwbwrTD1eRaoWUqgjuBB/yz8Bp+5gx52YjQ2kBfb0YqY5d
DnKapnjOMDVbm4xMPLMxWUwWXFSJCka8UtVTNYEw8vtt8fdwxjkxFHzgAcXmdi5G
E8/9wLyfJwCopE87K1J/HcJ1s2iziD/e0CTS1yzPL24Q8BC9D5hhm70+Mi3SjPDu
x3NJQeQQnJYVt1a3fJSs3VShkX72DCK/OtuGJ2dfrHTcHZOPLYUHJC2e1zchYBFB
I4KIjRelBSFKzJH3gVs+KDq/IU1OPLNCt4mhM3RR7SBm3UTTNPjxB3isFLr2SVDu
jJfyJjwHKsKj1BiiGTgU9CMU/IT8KSAZyeW5RHHO7dcAwMWL4NKAFV5p5b5v9Ube
D7QeydamkwF9icGREDOufCXnQOace1oSZEGov1r6ruAeiEcPSLQpz+hLt35sHa7U
qqnqMfVwvaSWC10rfc8NeIYo41PsBtf1MQiEs69ES7gQ+Ypk17dPCrWuRmkXkj/q
gqMrFFM22N4XHzT9+xegKHQfP9nqSzNg/zaAWVtJkETdh/1nhfLxDEtwJ88rl0j0
mhGVwb5TERJz7JDpZnWDJRw7meNq16EqS8I66Gnpx9leujK08RkJg915T5XaAwLr
E8CtvNvTRrdWRJXj/MKHZ1KKV26ax4BoSJ+kNVSY6ke8X6uMRgBhl0Av0nZoeoCX
PH13pnresOxwutb2cjvVvvNKZjR4EzDs5whuxGIJ7WZ3p2WTfA/xP18Q3dlD41FJ
v2cIwouhYGPleRPigKLYGxpHfB2Yan9hl8oqndZlsvfDghxad8QBP0pMsZCK9Rn0
bbs53MMo2RYChlMTtULrYLr4yTzQZuCJcuzZgttD3aA+nmvTgOb5EKYVxQlnK5Yc
ux2gdI6mZ1YZSj3R3l2ufDb3Obn4EnwgYFRVngMatHwvwibplQ8lDw9pnhoXeENL
IDP+y+pd7OrdPR2dlsMxP1VXGJuyjs2Roc4ZJ77atzxe/rFyDjX8kOw76G9xckfP
MDntUZCs9K8uIgXptvw7eMRjakQq8lmrpLSKs8TYgXFSqamA/NwR5vXJl4tJ6T/y
znd7w8c+XJzPWzi//giwdx3XwhuBOVTjvOWFynQlbpC3CsqaotKgLcVGR6o1wFIQ
1WIVD5WVzYUM6DaDvsblWPMVp2GVfI3pp1iASVgE7u5D5hKJULfaLjf1msbJkoTi
dLU2PpRAYaOqeytQhpgUGE21cHPu8ZDykzfA6GWpiR2cwuWl2GT65BjTQkMFgaFR
c+t7ZCffxfR4pylFzd+FCquMKd6l1AMChsT3vVbvmqg0S+8ktqPNAuUWQr5Fsy9X
cJuxWFc7pHjIjJNCtvkzSUunjt89TdJ/uwgKcSpC7pKBTJRJaMkeBHaEj9dptFpC
zd2GyHduVfXC8Jn9F4Q1X/ZfN59p6Fi+j4y+lNhNJehXQhzn+vEvw/nA6vUJwsOw
1UpFo5rGKIn0dDf7QFdsGj2Rz/rhTWx8tj/FozPjx5DjxgEAC89U6wkhhzy1ntbK
dZX1xDAf/Th5PsMkIqQwnAAIv8hxxxESHeCbRNrQVGUGcO63n4eJDtZD59l9f97W
r9kwfGJG48HQDzPMmJ7qah9eKcpmxnlPkMSYQNnHgJ8Ryjh6hffxHfgyO8HVHuw6
OzYQhq8K1H2Dr9/aS0OZ4+iRfgECv+W4cM6wQHX+9amwIJKDwFAOp0KyelK1yNMJ
ERy808q3fywdbt8pUybsvKb5YGtBt0QZ4n6UHmVBvOB8MqXvyWhLIYOlSgYfQxUC
IyUGYuduHPcpNejSxUa2VMKv07AaDV1aXcY9KdabY10HC2zgq/uFVRHWA8KKmbYr
9FriWoongNSKcFfmCbCkUV/4VJ2DQ2ejOQSD4LJFr9Kbd4l92A6cdAbcjDf/A6lA
I1jvHhuxAAtT3Nwfmk/D28jZ21yjWPR7lCFyKceZtOvRR4xhaL1bRBLE08TPeV9b
WXTP/jgqGFLignPuPM9oyx2tiR6fHKTqmthODCAQO2uwFj0rPMBvuszAABijoNeO
/0cGEtfg6j0rOiaojhFUOzd0vVB7C8jZ7ZzgfjmZx8CsVlq7NtSDvq9qDNiQjdrb
KV7Qkg1ROoOaotErqRFCdvo8b4IqPY+c4xrGcpB4V2Rhq7MwB6u1hbI5ETTeqRbi
tLW5p0x2phYGPf3SZyNgSJdsGR8O0i6syEJwU7oOgpHXFrwN5s3OjsQ52rFotE1h
Vr7RgvhTCHigoPHt87BhEYQ3DiGGNdtXWpXItG35sbvOVcY8/kW7H23PfV6L1mgs
v9Biv565//DzVO98QHKp1Ox+oiEsQvQ3aDvTvEy2upz4FafbzzGyh/DqLigXp00M
qKPjwHezM+DdDJiB2aOr4UosUXW2TLm/6XEG5xV/BN9NZ3UN9dZx8Qyj0guuIqVR
0j6EZ8a0fralE2aX+GfXeflrcgB+13LZisN74ktfeed04whokKLTAqQnMtxsgM2m
rsgr517E7BQotyTDdtGV9BocogLKkIUaxwpipSo++kmUXY3/Fsqizct4hjgBwTwJ
hZDScmL6U2OlOvygJmscS3u9XiAybw9Q1122qHtsy/IkPVU34LJF2D9fGSYSPvov
FMnfZq7E5Wjf9MlHLzcBMI87fPhaCxqHVrgv89AHYf6L6j/I0+DS7gz7TInw+4Vw
nG6W+FeypGKdnZfCcY/EpVVQDS5KRJkWf0SOmVp5p8MP/I8o5t2G84H0geAJo8/Q
vX2uEs3GY6wslMlaWkrtBJ7vawlgTIRWcgAJX8aAnuIs+m0mkiWTUPUChkjC6Fjk
PJ6ose3Nsox6x+JSiMS918bWHPRMkdcqQPyLbhqQ2UZtlpJkTuscNOjFLcEzzLtM
6BNc4NjiNtlwD9lo6jXEu4EYAXJgXB0I7baC+l/f8Dh0JF5blwuINMcT/jqYlLSr
DsvOlA9t7P5DKE9h9uipQxLc+T2O5JRImLIdHvz+sUsw92Obs76ffweU3FquHC78
UZp9557O6HLLEzgLmQiHm1TnkShheaQrz62niP3Ql+qYP1qmfZbpLLevaSgvEsKC
2lox20bbHXqlfavK8wr0hoXX3WKd4CpkX9hhNy2wfxz/keKwh69aB1XlMKFq0Jj+
sBVkQmqdDriWqWiXKe8HdZxv/Ee5VQS7fUy31Nl0fHXkbnPube3V0X2SEl2mUrDq
BJ5p6ShEESKwILomaoplOqPWZrEnpdK5494pAO4savKc3y5kyTt4Og/MfGd9bm9i
QwKzm+ksXyrwq7WWmjOaK6aWsAMJputXpqWvZiqqZRsh8CSCc9CNm1y/wqY1qBYu
Z0qKv5M3Z5RMG+24gZB9tsCnfp+vr7TgKN2GpW1XJn7WE5yiMkR24Gve0IzWXENN
3zfP9BInK1s7GDE9ch9aT1ncZSQ0hNopQrCww32Xd1IyqSZd2WPYnRxhb/6xTomT
dnH8jp2K9Ejlq1LmJNZSIHnAbBqdBNYx7Wd//HaQhpAHhfrOs184YwZqradLad97
m10iFnuP9ilr+semT3RpxfoP4ADQyYSTwaIZIHpgK/Zwk+nQERi6kVxOYK5aImIK
5Xvohs2BJMQ4+WXeJIaxrzfOzbVEY8I4tOiL878O8zpubliF7qraN9v+M4eWUTuQ
Dsq7A95hiWjsYDKHtGgG+nUSS4Qml+4Q0T7YM4qFVnLEopGtSbtTU/iV477KgYjN
4wFMZaORebuSbvwSmZ2rMeinSE9TobVxoAOWC1N8vCUbEV1va/gLc6P85ykiuD47
Uj7H71QudZuX5zFnI+Bd6jDdCGehfXZ7pN6kf8ZvYgusf3z856b6mdNoSWApa823
Sb1iI1OLKaA+ySycj6tIYRanrEON1GEOsX50p2Fwinrf8vPmKUVZFc38bDsYap74
TXowjlHMYTO3+eynAwhNvXteCUNlYoo8fY0/8V/XCQSuujq44VQ+w1PfMAjd0uOS
hjHIBeK74xeO6I4G+WG0V7ZqfBFgMp9Vs3GbVECJw1rk1iVMxK1EMnE+l4tOK9K/
Rcaju0r9bEdaQOjdUxXrSfRsSxy5dX1jWib3l+Z40XH8LZX4rRWkbqvdBaQ9vGlx
KkNOPie9156nu3giR7cEGfni4U14EecEZoz7Dzrz1kOyyn8/VYU6AeEcJaXvn2yY
6rPv3JCnCCJblMvNBUwEWVj2pvsT63l1sokW1AR/bpslObHI46jzfG+i/uNb/bI6
QOG9Qy7Jier3rtk4G1qfFXq25oJ8LyHje2fh8sv9zT/aiV/yc17Wfe6Ni9nP9eUN
7f/r18zjmQTPz8mc6D0jq4AD0ygw0/CxCTUSKmhMfn6P9JxvLjJJ0qMrlZb4xeMN
cOMuu/woMTJuBkovqpDJMctwUcnciGB05L7If2ZK1csi6AdqjSKB/8KrqNUuNkW/
JdHd1W2XQDdnVkoGMIyIj5/HlMf1ZXB7+54hGu0Oe5A9qV2LeUOYLTAT7yBbgEmA
+EI8v4oecLm2zkKEifWjapBLOv6aW3vNwLE1zYG+3LTbP27nO4oHLcJjJrJTY+71
jkfH4Bm6AFA7BQVSt+CwLp3oyNkmQaS/R9vmjOszVv7HOdWv8tS/UwZsTOaDcl7h
7kB8HWL3Zbavv5fm9GOlazNa2Z9anhJ628SfTv4ZZuFPkHr6HkrcTJ95gQwYY0CP
2T2mdDCXVGiWGu8IJfA7+Yxp6lZmkUGdIc1rK2AMC2AzjicIAVnBYXLGe4Uolqr5
7dN55empkWyIgzuxl2FE5m5xXhUeoRTq8QhRbJS/a0xLT5jWcWLuLZvzhLHeiknT
OLKKut9wVQ9w05YhLfy9eOOqB+Hz+XcQ/4OKVtsAWov4m97jhlCMJw6S6RKzvBnQ
+AKzt83tD4Dxg1wsGykfjxrgdEwxibTML/B4dA22vhJNcdcvilT96F2UTl0yRA4c
7da997eDSaUZUpIJQ4F2w8NEza8AsTeTZPaGHjPcwHDULkrJlH6dEDSYBm/Xj6N5
lTkdpcW9KBOqtDHDFZv3vt0Td+HiJlwfSjiheBfzWkVm/2o+F1Xem8egpQ3V6gr6
YNv/Fk3E/4uN3eWUPXs317kaiybP3RzZHM90+rf3f19dRBAFx3AzXX0AvhBMOd+L
qbYdeWKR7mOMiop/XPqFQFDG6r32+hdjHa0A0hYfDdDGJn2yif/wpW/54ZfmH0y7
+3D1dUs04q5Re3uF0pm9Q1G37riLJ0Tw4ruxtNrtAsS1xxDM20kV9cDG+pzSxcHO
cF0LJe3Z+GISjnJASSZSKdvuic66lq+mT8ATwwfFPIEUY4PmueLR3UXB3LYRvZza
ytra6z40ph+zfOFDhNbNKrGcDDXVDW19GAYLmLrCTu1ngC2V0Bg97qNA5cAD0ahq
/T66KNNUUkkbu88YGohQtcWR0YX4+h7tOipD184/04p8hu8pKHRtk0WtzBc1XLJG
xRFg2M9K0kXlKIuCsgMVHvK8qEaDEq8lq9KNFEX5JjM7JOCSkeor1JhSBBz+E+gO
4a84FL7b+yhak3kj7Q0IPTRzy7/GPE6Yu43JvbLKzDuTIDmEDsa+vX2fqt7QmW9I
dGw3pjzb7z+rsx7xEKw9l+6s/6Wlc24P+xP7fMBIK+Pi+vrsRt9ZgIgwPkU4wOj/
QNiTo4XWiB6giozeBlpY7GDk7+ftpahaqOosMsHwXcdYD/S3w+endT7wt+sFhIXk
VfE/mE9lZHBLnT66CVN/hfMAKIWnJgzLPObVS/VAAwaiMa+yobd2SkEI10neVEEM
LT4OVF51EtagjkQ3q8JyD87jA3R/uou25mjU/LR1MvM2aB4DLbSTQaDIFRae88aT
ukKnRph++5TyTT+Pzl73J6+F/N6DB6NWvCG2xOhlsCKduOO+8joDyO2CSKFCHoKL
uIQALR4AZyGGe3Cp88q+oEqw3uzQutQcWXLb+6L7qkipooxfRjCO0LD7kacZfrSY
HscWGJmzhcCKwjOG3wPsfbjMFTHeZKHWn4OxFR1l286+J1B8m3BwLiEh3GXuDr3q
wJ2lheC0C0QgZG2tMxq1heqKCTEF9iVgSGm5keLue3aQyBTT8WWzYQ430qxnPfGz
BY7cPoLcSU1re5vpAHDe7f83EJG0ceBkYnEDT1yRacOrmkvJ2NooT6fQ6p8uuMX1
D78y0d7bMSFmBXhzkkG2Z7Fjz1kAFY2z92JiKLlHMkFAU9jlikJbZOnqeG69QhRN
vjh9wJJ/hjYiBUSMw/qmc8rbHFjcHYHL2bDN9VXIvDFa0k+SgvjOZAzf5RSPTcku
t6QoelKQct17w6jX/w8cKG3wocL9jbbUh0GDZzUPBDw05C2ji9nczWkorrvfd7+e
TX1dDen0i3MFgFp4C+1p1IrpLtM1zsaAaSpAEJCHaGtT1BE2m5313OZ+vBjYIJmU
K5RTWPSCvIGE8FsDr/5q2om/VNO6wAAQRrwmZBVbVReuQEkUuJTdzbN5cXA9h8lf
8PbND207z0pzU3yppq+/F89MvviY19imyIhqZG2HpXG0dwNha2VxJMtPJuIWaEKL
vAmgQOJm4n7wEBgF7MC7gBvcrhWPnrbRBNzYTmTvhux2a68SQrbgO79/QRG5fNKi
sIFeHzk8kFLoNWrAJ19aEGYe87UybAOS62VYolQ7Ngs0lLS91Ef5GpNiNhmbZrRq
0eky7zFhr0L8n0eUXZg6vxktMA5SH+/zqYINme8UoKuw3LIWkih2uPjG7jvx9Q33
mDHQJ6E2Jhso44cbY0G463QMNjkP8/yUnu/35hkPcGuUDhiDUM42LCfEFOKV4XiG
fUAkxHRwbxpiDLojW4q5JaWDEHKd8cf5doXYbwhvM5R3Uoa2jR2cF7q2AIBJqwWY
0SS31ar8pdLpZKGZHMH1TAHCJKxG49KwpV+yRNSK5zcHdpb2vqAWA8tIxvoUiOvD
YTIXz3RGXze5nR5TsiNFa4pU7YoefuiEdxSsklw5i6F+edNLWqCtfO5XN0DSzzmK
o9/Q253FzYFhLsNrYi15xjr0ETtl98Z/GjolI7mBYqDiQv79gfVmAPmGDHb7T98f
uU4EPB726L5bNnqG1eqVl5RUMfepyfNwVte1y53E3d5X7EV5HoxxWAtz7wP/YdqR
IPEz9loNN5RoCZMn0uP1gy7gf7eYxxz2nMyOAjwy8a0tD4l/IxwfXZHzlnWDrk+s
2FAb527hHCwNiPznra3VHbwv+/oxHQlQpuyGG4cjL4D6BFXadEeKeyCJaugkjoSY
aZd4ztDhCplmgcyicr907VI3w2cVf5PYsDqIepmzAf5u55/MSHGAirXGwhAaYn7+
re4aGxwYP9Tp9328zSJlMHyNvOqVNkjtHEuPdxAIi0+jqBacFPNXYJrPXML4cN3W
KKvA1FYcF3kjU2+DVNm6ytNDyoH/eUGzxFwQOpUAUah68YC/x7l8P6Foj42D/cSa
hMVCe+ZumQ2am1v04a1RaYjaSkSICoqcvTgp6oVoCN0SDFLRGpMxlLF7np4R/jUv
tK7AkFM1D0LhAm3GWowAFd6pOHIMlgY2f36D5BBBIBIMQkZ5GhYzZ2CGGkBvfzOQ
rrjTzMJ6RbYTTd++MIFN99eRcj4ft5MpnIwpIM9GPwIj8fjmn+Cs2tRBl45v4Kew
uJp5xdBWYAoc7+kbfvCwCnTddzmhnTnRcqQllERTCh4xy4pCZWMssQlbTOsBOmJe
gI6eSpCYLjQXu54ndzwlMhFd0ptyzRpQLBv1GKDr54CgXYz7zTarbL/xHSbze9yE
Wn8l9hoijcBCi/CsD3nwi6rTQqt96Lp/rSHLiSMI7kYAOojEnQzCRMS3WuX/fFZU
751E4kpU3IV2SSu91G909cVFQxYs9SQLzaioQb9Z8btKYaIWlH0nf01bNWisVQUq
msA/zxbTOpYMZWWEQ+IjA0A/9M8L79IoapZGF/LY3C18GBtWea/wfR9qAA3BVpv7
k1yyJhkZrS4n0dKThxiqxgf3doaeRFsrzlDORvSTgCz0p1+iTH1kZmAKz0qisU+X
az+aEmZXRr8sG/1OpI26ihcLkE+T/m76StwvFbWFLtuw2jTlCG9Q9rzt5y6aLU9S
fUL/v8W58aoWIUoun3N4uMnXEWKy7tzww8P4Mcem4FusQ0i9ZB10uaFHTY+oKdTk
UM5LLCxPKuAoccd/OZYoEBh86TyFEw9IopC6jZgEOzaHidD8Mho4pPIsiSHgZod6
/n1JezMbjowolz8HZtMVeb5W1p2hzmLcSH7o+PCp5SYcNKsc29aREBSUsAs8kop5
F+OCwTwXugfbLgfW2rLDxbXZygjFQ7SerSBN1rKxxdKY5UPyMbXQxbhL08/w1tuw
8d64//n+5TFu3b6S+YHnrOWtonp4+9bFLn8j1smc1y/HcaBJ9Qi91fwRA530PTfM
j749K/Z4QevLFMBlzAOAFQqxddsxxEDBSgKPBrjih0wyOfsN43rJCcl5g3t9rj/W
/eKxBZ9AZu1dDYqLl2QZSFb8oS2JZr/L2IuXS93+3cXf/LiiDh6J+T32REG5cXoI
nbfDQWeFO1fVMVNm+hwxsTTP6etO0jseGBHzisEiz9Rud6N7zItqYzNzQx+dvqf3
jQcR+gCb0nyVHPnJ3okHTZiMzyRf9/L9FAuph3UFGZ0INoKFrTu/uMTt6FyoyhT1
yyrP0Din9cja55wUUhr6Xn5obV7eh17QCJjQWn7pkExDY8L8HZ9Q9McqcrqdHr26
MUNV3isjyp0dpHBLKzOMM1I6ythwciwqUMxxnUlNW7RGUYWvkMwamuIpsdztszFD
mFU93C2leD7uS9oumtypto+3rk+CtWdZu1aLbHdlZEganA4B0SOwWQO/9shAQdQj
hCL4pqttXuQiY1FWnqeaibCbopQ7DL+yVXaVSePixiaVdWpzS6PY4BN7A5O/XeF5
MVfQw8qH+vM+u6BmD22KcCgpN6t77WVF1rYr8hnacWV2yJUHDYczmtGWt8SjQUVa
mzBC5TqRSZf62Lh9J+xw+Q9X0LXuCL0Fn9nheIUlNyBcM8l66k3QCOE2glXNWhkW
BM/g/4HltRwlTFUmqa5N6h5ghWSkpXCUt7UZQkL0qK6x3dxv1mhL2AzkS7tqZIl4
ylscRdL5Y/Fyw+2btzgI4Q2MgywmIX8WPTudCHbB1MjNzkbFM4HR1X3cFf8GjQi8
JjPCLo91ykHJca2rVRNFxWD7FEjrsnstwBpwEZVjaxXg7dM4VrIytrqexP2mqwVf
vEbnqIHi7lLmcxpsqI4YKicLnIeTunlkeTpMSLZZ6Rgwl06mW9fIG8ZpXT+m4x7c
jGIye832uZxzWDonQEZQGVvmeR2z/tEIQWGF+uouK4BbK+Wc8V0/l+jhL9M+2dph
G8nVrXnc9NfsxDOOOJWwcDaVgecISuDvnO0Ac9ybmD7wSm2/5nNg07vLZRb2rfsJ
AovmMKXRgdiiF3gTEi/+I/UsQ4QamWCcF17v0WMk5H/gKTQoXMkYpbs80VSJjSP6
lEfIg/Omr620Zm7ihd8nSIbC+YrKV3ecaf20sXwljuGHPkv5LJrppISEWkkmciJw
CZPSzxtDO5CGogk/9NhXzza5/YUolddjlx/uZfhSG2kgeI5WSR6kRDBwam/yV2XI
iIRIHF0GWXNgCmxPHw3uUloTK2xDpJzvtoVJ6/auLr0t/6C9yYPyfUJo4xOhPl23
r8bHSSp+KcA0g2dflQbG8l1NPujWrZWMm7yBaU9qjpTP70byQrXuKJqICOm+VdTd
7fQlpr7JlFW1M2f6v2zdkH+XUtUhcTSQT1/GR7TtjaO5FYdhZ2XUNdYQ+hivcgex
xNwQzpa1SPmxLOCbJCmtwfEND7YbdY96glh8LHjfOIMahprHSf6XeRbuT6ytUleO
vdduhc8rR0X7x+CkgY707yRkaXctmG+RJp3QV2srOR7XOjYluPn2U2eCFjGRix3/
awMHBLR0mn+z3JevvQgfLh7nE3y6FcpeGJ7oOurawJPYME4WbO6xCYGdg0w1+AbU
vrRVtVe7XbjXWiIfOBah4LTu+FN6SZiyigc1o+4OoNrFF0gmDwKHco42/oZFqxi9
OEwK/Ag0tYvRPjoleu7uhXBfP3iihI1GeqbGYifPcVoRuiCC5E29ljW7pPLP9v+9
lgJmldcv1Kn1GsxCVFLPT2sMyXk4Yq2y0Sv5siu9TCEZWvL0O4bJWY/3PMgUK3m/
Xzw8OhKgepdFOyUB1Q8xV71FqyV70LDPbv/eZYEd4zJ1IapoeoNv7Zqbbp7LdBLb
IVhcypEy4fSes883xdXyHfF77nEG+W1ShEpfGaKuwHBiLmRLsyru6gtIWEOJ7deh
yXM7tDMajppDD9rDCKo3QwcrIR6Eu5Q8x3boV9mj1T5zJLgyYYBtTFtRaGgWhRqv
9HwIOxD5BRzei8ewPKPsBWoWdDHykpfPDbwJl/Tu0DmXykZ+WxIQDmkP0/l5mlGC
oWBaghmqQQhr8yK8FLXYddA+xzRo5t9LwKffIfrszEzi/HF3OuuAijhIXjoXolnD
1ZT1HnPIRHrDKVp+G5iqdsKQczCzgPIkI+DlNG5JxQXvjgjUydl8lKlJMVFyu27M
O48BUD9boia7P+Ps1QVZR+CHZOEENmfSPLa6Y8dF/TdwCxviScOD/IX5zJcxd2vt
3ykWt2TIUjP3RORQdQeGBH8AB18wQ/0VBX8BJtdrZ1zKTiUrDK5lVtWKlzcCtOMY
6iPtrAaCK/SH0dDXSyS1AXrxgr9u5IpYFJSjGswiTvj0WXv0qWUhcAGUD7aKtY49
SBye6nOPxTsb0lT7hULFX41cz85CaywfVk4HCnX08sHm+8Yq+9WbuxwFVnszNu7c
erUy0kUYfcQtIWg3uykwr0n00qOYEjUI5R68tcrB2BPe3JtXQQYE98xmNmv3qssZ
6W1sCV9rfKJ2kT9qPvTUDL19cPmZB1vNnnMoyTaXbA6ENo+gdz1L+XGp7Fw2dUjU
W2VUmxolty2U5oKTPzegOEKGyqng1oy00TxWP91wJn5bXV3gNWqETbSChSBRQk6+
aLpyVGCq7HSKvlvosKrb6cEeYu94r+iJSxjBfsCZTIwyuNyJS459xrn8BwwuoYJJ
5EfoZkicFjRmRCR6/nZ8AyC5VR8iRX+WRTycW026vt6YZv/KkTLVMvGIcQUFgHDb
RjhhPF1VTuHi95eZyW9R6olbynWzdRmgwiUZcz4DApwnNLgtiTtoBziKizcCEJ0T
jKh4J8TquD3KUJCpuTkfpo4rURFzf/IDq+iJEWi+ZC7snOs319d+lnDuaPriq8OK
UcYS5WgA2VHJYpKcMgKeaexQLLXeI+Xm7Zx9OOmAS2p8lYEzX9fF0qorcqTlH+4O
PCKGiAH3dFKPzGV7e5vkpLZopEKrNo3DG2KlQq3Ka9jGKCUHNmIkMPAwri6S+kjh
kGUZcouSjZ1bJBJNSCLECG7U3eNFXOvjDvFEPdOpWf2eoob9U6rgzz8KFCGgTcEl
8afpGsteMWyeVXiHygO6frJRW93oZNzIETMhWByALJDQVL89hawGEEpEwkw9E9bm
1E7QH2Pqudo0ryJcdeI5kNpWr600Vx7ai8zwh5vBl686a+QDbbLCQWOXF4nlY2Oi
kVjAKBOWh8lGqqREj7RXOJCAFIQkNaQBh1+3ENBa/qD0xwE/3HUSRfa9cXmGHskq
zT+bjLWYbK4o0px4RfO+wYrEvvJ2Rqd3L62eQ/aPPTufX0HjgCij/MOukv1M+dB3
EGqrfQziyVIxtTF0nsiYz6Ko3MuzpAixRjkwA8GBmReIddhgZHhi2X1TXIcDnEvk
q37c3qNnDstXuDWIEs20aoHCdgAvA1KLkqh4H8nkHNLzl43m5Ql6mezn5BHxNl2X
k4DTYglBlEuGoTWQ0h1UAbREI2nYJXWlRYsjY2MUKgXWPrhnard1C/8CuBcUguq9
q/3hugxedMBqe8334W5Nvqm+TTPeCiluJ4vFZLe0mI6c9Ww0lKJQwhbDyllBYJ84
qSK4Pabz55+NnmnLXz8SNbJDJpFlxO7EbdFXJiR2/078ZyHmGHKRDpeH5ryJdFhm
XwuVmCLeKLE+PDNyXCXiBL++G+GplS4s/Sr0BKQOBzHWfl/nCsMYdg93PAzGSw2Z
bPHYO61/lEC/bN2X4MeifLkqKH3QKdGrJpwwpnj0VlFdn/8FE24w1dm0Blp7IGEP
IyhAS0Jp9O7obDBxXJogNlq/SvGJnBKQxhM2DecTWjPZebrMd8NHJoYZKRwMO+wO
xUeXGww/MUOFf6HJSh1HldQ5uSSHGBw1NyJpCDeXFmHSC7h1f3JptdQ1W+16cn2V
OpIgKdcjLMkFuDI3j1H1EDVD58POOtHWYtaI+AApXGaufrLHsOMYZbdxM/z9S0pp
vEGrYxuukp36pXB4wxyN1dzaX5XI+W5Hp9M343phe10j4yTmCrbo7dPRBIcm+/rA
/TeEU9OzIM5PtSMF1UtTPQSQtpRnGIskEZQeHPOEZlCnoRm+mAC0sairgtHHfZ/b
asfnPbszQOMXfUYuCxyXIy7W4oxDvjxq/WWUvImPD5/XDHSj7my6YL4JDb6GzJ5l
/6LNQLfLINfOo98PA6J+ub+ycEUjmESQw8Q3U8DGruqCECt6sQ6N5Kgi5W3pI7Ne
0rwKHayKOPOiNsHXw3MMPGtiWGpn4mq9sI4/Z6vpMF3WvgAN2L9WCZoMP/lNoPTz
LNRPVKPzvFco9G4uTsQovn+9/akffT0Z8PsYlSBWt4twO5ESSNFCc+v1dP+wwECz
M0qn4gK/2v3T5kuqv5p5qXjyU//7W1HriPt8HL+W+1CLNnYmPiacyK4zgkVLqAG4
mc8gg8s06Hl+SWLgbp3hl4WZGKFi7pH75Gr2cPy0pYm2zhl3hMZHLsmh6T4Va40d
RoT0dmcBbYpE9OaHp0hwGih0CTB5Xt+m/VO/ZO9jTwoTyigmKd9X/EFUNrlNHu6+
b+hE/Oif4UxVZSxw1T3qH2TstD3viYiWX2Y5QNeCUJBYJXFbEQgYOtvjQvh1Ca7W
Km3el/pNVMVt/x7b33J/fCgeNvfRdfgj1nP3Cte1LJOtA2BhWxiul05Q5C726vGH
Ec2mKlew3UjrnO2Y4wjzkK5KyG30Yh9qzBxH1qIfJeYQyr9w/Uyop3vWS/4ECnfe
OIUsdQgvKZFeKCGsK8sp/TXorSeRKBOGdSjUmquijXqiBJVb0f728x8++qA9fQ+K
b9J206Q95E41+f2spqnWR9w2JpaIHX4CMeKne73aBdxJjIYqHysvQ+cDRxLbHB5D
4UxUAnm8RFGUNFewwa1zEI7Ui64CIxkDk+nFke/p/Hp/aPayKMMb8wVXw4uoFhzr
L3ghaACcEpfoTfG5IVWgSRjn35i5BWQWQFQP/rLXcheYzl8O2z/iWgIJF//Adj18
a0HxeQr0AZbDkszimqGvySEkATR6Y/xJOmqMUs5GfKcvOiKxsR5n36FcF2wcakZ8
vxda2xP3gVF4lvH87zBPjOQsiLTWdlF7KgUIL+Su1gm+U097ooiKhc6zGyR2aCGP
FRbq0kdLHek4VFwL4S02kCpmrW6bWfP3Xg0bK2nji8c8PUBXL8HeLMhNGTbOS45x
XINNjC6Tv8smsUxBihkAf7Pzw1K7nZXQ81PK/XNaoR6IcmspzZTLMePa8t7JvJ0e
GKkWif2EnK82rSkWDdBvqCPDH9spgVI613jHsy9i+0X6J7yPkuGHdr3tMKUwPvus
zaxZaVb+UHxW+uFuUqtlP4kW6OM4uP6Wbzu22tqZfu60J5sgjuTvG8OBcPcHNToa
fnF3JvbBnrnxYz1O69p6gEZrOZIijP0y+sILgGLiBj5lvNWxuklGzAUFOUgLRIha
9NEGuv5tRBNvlv9Bj7+8nZZxfO5SJ0QYYXczbKKRTU78h3A74zix7M37arlI2AEq
24rCkCeSUrAgnXwnFTcgqpkqz7uVF0HGdzZ0o0SJ0qpTzd+IqwBpKuCsjj2EbUpd
e86lzzAGIGGHKcmi7wT2LvC7yvkhkuddcvi0crtIi6qFHX+dkpk6nBZWJAkdFNKU
6SloPqIrbizpYmTz6UQul1GtwFu/o+P8NytpmB4hhAdk+YxN5vvn2UQH8TgiPEsG
kWbNnRw81CSSeqMdY9X1dQUX+nRySZRze3x0Rh4DNGRw3DcHNKtm7xoYttHBNRih
FOv1qfUCtO13lYtiokxjfRyMp3DRkS3mXffe29UV1GxV8So70saTzLHQAdNsnwXH
ld+EH81G5Xjcy3SlSLNcZolgX08585JfVCWushwLVEELNKmC9qVB1ieiMG5gycqp
k0nWgYBbklPV4jGbnANsiTvnYcP2MpHTo35uhavbg9K51MH4OhDIYRk1Jy6Odxv5
As4o11vWXMqFS8n9aLM85FOWdN1DDGyJ3gYCIrBzeDkOOlydXv4PNq/TXEwBfKGl
ASt8ioefBT7ItVfHSJVrycNGP/eBKmdVecgrk9JY/fWGBbOTbM+8HQdw+sgnS3WD
hFNG4sPLQaeCa6gXq4G9Fq2ySDj1k4KgrqpbTHC4wVrzicUzKsbfdGmOnm5Owqze
Gxw7lw4YlYp6e7o123xLYsvBT+Hr9wN/2XKn9vjTpOWoCEwGROMaCliAGZ8tbFQk
mgY/4thArDe0uSkPvYjFJ4ZN5cwFb1/eQrKKKEE20JM13PLWha/HSJV+e1sMkrdO
cfbR/x64BHmxbyORxPvYSQGVyPqIsVBQamsy2D1u3LyPJ4pQirPpX89wQWqZCmjH
P1ueTQMcnU314lA+M5zx1uFfWoIpqJxH5CG6KrDvcfCMxAVEBRWWIX1wGPn87BeF
pg7ZysWVvkf+qc3NMJa6FSQhB5+HK3xfIiaQWHAMKDURM8RGPnyob5gEt9WYtMSu
gJ10o5LVGnO2ztRy29wwZOb4Hyk2wERQI7VSBUU+R4cQYT2FbMwqFOtSEEl4PIRr
ghb8pcfHiJay9TsJKCT5+A9cZlOBPJ9cBggQlOlO6yVSCKiLbXg15bJasQepV9mz
j+OpCI0xYb5AgrRpHG2hsh2Yv+fGTPNqI9jdF4BtOVGGytdFHIObdO9E1HdoiMjr
eMM0IRR54q6ZMPxtPfzyUyvBionuowK2SSDmQYZeLEs4C6oAABAnZBOHZ6Klc+0L
lrUs+y98x6SE0HOLIllTHKsk853jPKUgC3hS86rKUQs+Jj6z3wKUOIAaj53ZQwQL
F5q5RTNESum9QSdSVL3U5/x1PSNzz0QFQKBSHEllTayMTa/XcJwM635e+Kim5wOH
anbwDrK01o7b0YKI/i6P6Fj5faGxhH4/eIbhScWIvm4lizh9ISXwPKN+yaIeIjgF
t83sVfpn7AE1p1zqmZZiwL9BYAcgpJnQ0tYTme9wowhex55bSw3y7j9ptz+qVxtK
gx5cRZK6nNFukJBtfcC3tXPR2ZavR3AobnW77QnVpOak3XuHkn5aqfFmrxmnIeMm
rpSw5sXjnYwBsX0/9WzSS7XlcKMYllsqlf6mVtZIcADPReMIyog6kVwujw8CcWZS
/Iqp4jpRU04OhjQ+X3lP3n3gR4Q9ZeL9yG40bwKzLpyLUXFj0kI2uq3RahSDpPCR
YW+o5O49E+osyKaj3geJcBZ2tR8Zy0mM4JHa0PeR3gu8xIKzJWNrtl41B1ObzZXN
FNS7DflMyIuT73HiQuPYgV0prTnO0fkErRwfXhfeawsPcwgr2lGbGmFYjheL9jUC
6Yj5yJ/DJjWZjQV7RKzGkQKQdQttN1qb7QPUtiFQ39PGiINBE9fTa/fi1fSKujXj
yda9EKBDATJe044cgV4dNwhg+j31BzsggSBUINln5Q+BgQFrk76/3nGiavXpUqiH
++IsC6mDxo5M3WBjKGEh1oaOUR2PkK7AnZFzKIkdUBk7GmNZU0zv3u+9aLy3jtVh
Tej5I2xzDs07y/W7D31qJ9qzOtKZYRtEFq7eUf0dgvYq16YnKvcfeF7P0KqVBq/T
9oluC+dy0MRzShYzZQZNoVGk7rV4iOPJn1D1Y2g6iWshYeMow6U4lJ0f2CeSySID
E/cCAFuwxTy4ZYpuTBeMLwYdluNKM3YngSocbHgkUE+3G3ztTAA0rAzxyHOKgfrX
uLGs0ny2pyfsHEdpCyjxVp11wgRkl41nVdxs1WHgOSaEwb3y/bbzBWpdoMujuQne
THFoKsZL4ZsQNXh0z8a5pWhbk0syho/VIvzsmQZuvTCq3kumy2lsa7ChxzPYUUum
e7R0EETYo4izOtPvztQbxuZ6ujRCH/3mgWNVPcOB2BovaROIUrdx9C+++4fpbfWC
QjD/j4+2Epn5Ndm2hmcFwK88xgp58ybEVHrTK9ugwZgmXBs6PuD0jpKUNjLLI063
7994aGV9iar0DVG9s3wMkS+coAoduhej/i2l6g6yvdkoFeDNo0vzhs0UiAXjNuRZ
UCHgcbXFpf7Y5vafuna3EukL+m8YR00NoYxbyUKjzLX7yfc+PqIgb2Uy0z+NLT2f
tWx6EgZd6bSJtEbBCP1qeBr9GtNBqC3tQ5CuysbrvUbbN3aAb06i7flVzkboqKVb
Lrr+tO7rAt2I7AVR+GmQqaj/QqxT8NtoEigNOyyDaLvUgBSGdFM3mE0sWNVVKafv
iPG2Cdrz97/qeH4wqajoCDXiCbRZN+ARF+gQM5upZ1MkdiKmczN6wlu8FbysPnI+
RWL9KLm0V/mLiLg1AFWx4Y8gqM1QqiIEV8OoUzCd9a5uWoQ/KTEPpK0E9JW6RAJY
krEEhNMWsMP8xNmHyBr/J7IORSjX598NvtGUPNnsMngiXxwmF3eXvb6lEseWoGne
u+l177kNQ7/TZp7/0PnoFUd/HPRvI8yq0iV725DcuaL1RFF3eoXuATa8yO1TR5qy
voGd28ek1WzvGkYbtP1Kx68stnxpj4XQajGEXAINfj9azJ3E9U6ed5vY9YRc5D1w
fx1N7GeGJRZvXZb0l9018H4GokTmEkquBw8zdHonew/5wh49n/4MY+ieTobWuJNB
2HdRo6LrEs+UWEabVAnsF891mJ0DrsSXSCu8zp4hLLd2Vqz/LtfOJXPiSB1vwdRo
7wumJT6WWLHCTjKR22fCdW5NeQG5Vx5+SpnD464n/KfU6HHD2AaowYw2InuF2qpi
stzk3Y/kkQ47J8MnR/X/YTUKmqAa3JcLSbFm/iGQP5CgnU/ZM3oRDGI7HrJ+8s5T
+kDogTgRwQYYFXwWewYVQvSQPQQddgv0qKNezTBPPJN5amdtZ8RmdPt5WDoonNp5
ZNJ1MA0kCTu+zbZ/57bIXbn3ON1GvV5d3MNy2tWqcCCkKXjZm+hjYGJq1XWjT3uy
LSd613T1nW3vW8TdbYOWKwCQQTBABIFCM/z9aJkuHoKPtE0RTvyqAkOB5/JVgsFw
skpx4h/MkjRORCJV5EGMV5l3PH6aM4IGHAndgawbkSWjuqHp5rKYPwHqNm5RbgiL
LqW9WMhZjDtm3NbxPASkqow8AGuJ1h3bz4g004DZwXNwLQeApt7iRWQP2lOwMBC6
w3oQQfelWuG7E5ZIo+cqXDbYdhrCiYU+vT/ed5kXUrtGdQsgFTkNCQdYnKHyIAdq
fIeVEUaMVbb3a8QuWuc5MrWXVALfu8LfVn5viCJibIzBDJAWEFBISSDb9K7Zf7iS
qzfmZ+7I8Kv1b8KLYjT8uqmjKHmyDU55d4jj/fvRN184JzLvBgGQiHMDo2wn2YJa
+GNeCjEVYA+oAZAW4ZTbs3iYdyWYlZ698B6bbnvC6Amf4lBg2j0+8lc0swwGqWPZ
hd1Q4elSyXtcH5nyt/NaldyMNyio28mbAetsriX0bRb6bsUEST0ZSDnj2q1IHM0U
LG34ywwk2qoWO15FOTEp49pEUyU0LAKt1VTHI2Q3iII6O9jO2QWVGw/EouHhzW+q
bRq/KG/EDNK/yhHWEihMlLqgJbj7ozSlMaFlW3+CyTLEvpBmCSoeB5dXcBrFiJe7
S8RC/gA+/wgDVwAPBiyq6SU8T7xgGQd3KP6UrPjgwrSN43Riw1Mxg6/lndEE1Lfm
w/Lvr7aPfHYdFYnjLCfABaX5BIA8PSDrc0XkRywp4r9g50ebR5tXyKGOdlhwsp1S
LBO1+4L7ZQKQWfLb77A0YyS9T5ZFzWV0VWb6bf8oX830bIydrcQz2vhMkLaP1muA
W384XASjPDbWI0NTFlOf7ZExbtMImdq9TLg/nYv1QPH1MkQpOS2PuYDIRVZ1B5Jf
hexE5nA1Eczd62nix2SnvaTlKhvHz3RkhkI22tMPk0mj5q6twWZBRHQkih3aKwls
J1qLlkEi1JX++DLLyQtwHkEbxSjVlTQlsdH6FT//c2BP7wFCL5rr8qsZh1NDkh0I
VFXy9TqmPakh5EHprmcL96eQMkmS7c/+1ROO1gEfjywI0xlj/80vALDdqUOdge8N
XoN01SYg2OXglFmagViA2o/ddZjMM2c6C7OhE+PYf6JSzKB2SdyhXskLzpVqnRan
xoVFGLjT+w4qU+YSXmIM40rx5oi2F1SxlihmLJqVn+Pjw0nDMXX1aUrsdlDDop22
LDwxLtD9czEfsj9UkKqJGI8beLlblrCsC/VJQCu60ireLm3rh3ISjdH2Q6mq6VEO
aXcdvcbesIaLD2/UyqexXUL8cJUmBzxWnswdJTp9lXrFqJg33y6gsqkI6RwRdi7N
KLsNDHsXdnzR5/7ghn4iGNrXgoGYhU1edZBISfIm7416jnJ+y+fPbIdfWmQiy/XN
9L0V+jtxDY6qGlOU0NWACJoIHUR2I96gV4954Z84O/Eh5vwqtH5yf0qd/4U8ccil
GkyiOESRIOcTPV9C8QoufvUqWLdNEcXyFAOHn+nVjc4Yof7b3lb8DRC4c6nGn4jR
QWSRha5KYglArlW1ldeGBIK+HPVKoEDBLMHyk1mHfOn/bHhLaHUsLnIYeajFKdWU
8fv3mgkal+VTblf2RxJOijetRNPO8YqXgyR0wOrs0zgJRyAAuXWVG+ukm9ekaowW
MtK0qWzVlIwSt9wgP6yYlqBGs9MqqRFXAPkglz34NCjyo7IbA6Y9Bf8koTJPaW4w
G2jNYo4XwTrXWUOx4GQ2+5FIE8OvfKO6SojHHwmcGifT9eo7c9rPfzjtOVpWQDqY
VPl45z1lasA4k8V5EX/1IjW4mXPSbb2SynswFam5ciXEIDrOGwES5mH5nxUX7G4G
8rVKBJmRhmNNdet+gYrqcEDIAFPWXpj9YARKzCP3JhCquY6ncmFdxkTrh3UlnLzT
FWLCoCD1gxvdbcjMAMvwfR99ZqDXuXQSZ9wh0iJBC5yYgNoSS3dJ2vSNl/paLD3M
S8klLzqvi+KZYKMRGTaIeQ6QfL8goPEvNV+OBn6GTpvxObgfeblWmF6OPva6KjTq
GTkii2B3W1wPT2949Jr6X8ErS40Z4EFDNcu7JBqbjn9v5igDVmOP78p90FlrCPbq
ODg+zGHcvAOfHCy6EF2JNzYiboZr4gtsFM7k9rvwFZWNiYyrQanIODoQqWD8d8De
ZFku32roblb4WJj+JP1LHm/XtvGpqSDcrOf5gPcYztxc4aRNJicPjzq42XFxKmVp
eLSYcWqOn24hZwsAMTvN7ybioueAGx/JjVE8g/rFwL06H3UoC8uhm2yjQ6R/1AuF
F+NoXPYovC7Fo9Y3lT9GnJQ4KLRWD5G7LGnmEVDaqXHfHuGxzz3RJsXvYc8bJGWh
Dgp7kpiW1YSbI3Hpjc/FwwDijsKN/OnhDCf0eTToy6EjQy9n8pskxQwm+W/N5BY8
ri6DMUO89KXVZqinPxDHEhtcYI65W9hwSXxIpGzubCPrJshn1ZxgiknrXotgBayr
adAvsmvUYVhK/jIIInX6fA3Fidd9kLOzqXmAwsenZnDnqEiXyl6JO29hIproAfrP
SBE6Ce1Qy8Inzl5NKOdNBzkr0N9Hbab69GeMqGuaSbwwmomyXxMFWMGYSKQeQENc
ZbPpX/EPOdadPNJYiUTlV69SIACHFvdrKKR7H7B1IByMVvon3zFmDISu0hCpnF8u
B47eUWVisrnc4lGMNuzxNLC1JYk8OdGllKRi5l63NvGH9UA0iCSp7StW1lKFbNs+
L165Ab9cFGkjZ1IbDWgk07yRyltDxoA0Ne1nqqiEPP/PdJdYrQum5Gbaw9fRDW7V
xnSk0KlVYKkpjXFqweErLCzALh9sf1iPulVcMyX5Mb7NWoVQ6qs/IdjUOOB+reAY
F6LuiCuhXI5GUmookNHlXL7nweHid87xWEj9u2lZmGOgXJ0rG5J9zm54Wwu/8ihf
bRXJD17X1+oKtDXFydFG3iWSUxE9nYHhwy2loR0wiK98mN3lVnTuR+0clGXJviHx
B9PSuaLWJsBUBtiBArNknOs+54zctDPBN76iqIRcZsSlJT2Nz+wF3DjU9vIPQz+8
eDLO8ZNMa2BVtv7BA5unZvK7h3/smQUgpzm8B8RPAC0WdNkNK34leoKWXisk0s5F
lNzFGO/iLC1pNqCCfU07tWUtDOF6QqZa8W7YhIGF3On/wMOOi20Iz9iOtrBvj7oK
fuaqw8FfnGm1kZMYzDnE7KYgEK30GHR1FBVG1lVCZM7gN/78f1zMgg2gu1WYX41/
tGTnt7Thn/48ZpDAB4EvyWTHCcZh/sIuctgjrldgBh2Z2JF8yWrUX2lzu90K1+/J
9NSN7XDOFrSbKu5mFKnKOgQRTeIW2/sIlwi/AOcDsmbPfoad8aL2vCSPYi7LGp3B
IMytYapP8So08gCQj8oINLyw75RHLJbP4ysNltz1Jki/nmZOX7mO+scEL3lWIXo7
VvV5GWErLQuS9MazPn/elZm+DM/Q+yzO+4HyF4bGhuHrRgsVlaHF/r/AiviHTJbw
vbV1jMxxf9lxKuDN+RAcZYmF0Kg1p51hrhgzQdS7YRzJKWTrXUBrJwJMVJYlnuZ/
hDhjYDvDFop9vEjb2vVmUZTwcMQIVNhmsIOqa1ZyYleZ5lVycml/AYQ96YZW4B4F
HuTQh93Hl0he0hYMhs5x4SUZWNTpjZPA4u0MOdV1x0nC/2/yYChKNXQFNU/iJ6Kl
nWh+MdZO68tevWTG6cbrJv1L9v7JTLZ0EPiwvmUdpKh/3Lr0TzXu8r9bW1ZhTyOO
rG4OAc9DXw8voQ5X5JOIlSOL8BsUIXMm3rKEScT0Vke2JgiZ71x83RYc0IyIdX31
Vr7SgFhJtMqzbPG18QF+3IFK1JZvFTddh28YTsyFq6SFz9q1+Bv264bz/amRr+nE
zew6JPLUZDhOiPf+BeANMRA9S6W/r3cGil7TlTuV7LGGEOyVamdI3+bAnVpD7FiD
JqDWMwmrQMlABQ4ey5y9EW06bk+Bwf6FmxAsFNHMMNSRMWlVKp3UsXESfCuOF3Nq
LaCT8uoTjkk658BIBAhXUQFIbKho20wU+KCnWaRahC2TCQ12o11uS6ZgGtJh6S8O
yg+blDAk8V5OmhrUF0Gh6iaVsebexwM4LL0tsq0ybyW9JduRpzZj77rAeYbv9+Jd
noX0Kie83Xb7OyA2ghXm9YO9hvbngEdKWhMZ+lZ/oXIEuJZR49SD2pIKc7gLynIR
SejQlaSln1nwHqMrOm/9drI26KFn+FCRT6vdPwLYax69+ACZUvTgjTRkXGTnXOE5
ZeqRgqM/EEkbVb3nyIlqC114rFI2OYd1bqpLRzjSXuJt5dt1fqzYFZA0SaIVEWUl
T0k8jTGEgJDrdO26+ilh/23Fa7/Fab14HfSC8yjAoMokpzGltEzSIbZv6TASfu2Z
o+OUvX257GfA6Alful5odgFFp6sLzTIRwnn+VQ/QcjJhjQBEHtWnaw4DrT0SzqqB
+DTsDqXyI9jDyRqTWeme5/H8mf/T7/pDau50NLo3KUDEvvoLQsW52hFR5kzeyzL5
fCE5sWZ4dffn4pcvfJaKnirLZYQM2tXMFD255HYnpTJ3fNOSWIJ3p9dger9h8iFp
R+0Nd4z0LauR/JzoQYaA3kXVEbYIbLfCcsCYR6Fg/asKB5rLEpo0HuZaBJHJviBc
YInIX0kvywnQj7gBgKGNv3I0tVtl7VaTe2mraLXatr2EG1jpY69296jZZb3i9RBs
nUkR+YgwH8p+FQJg07jXj9tDHPZT+W8XK4hnzSVlMAJljgDXB2AoVvmjfwTi1eUn
fWfRfgqoXOKcacajLlMKx8EXtTNVqgKoa38CaGzXfX30NITWd1hV3X/z3ZZB3z/+
bfgIT2Bo/ueZGE3R1raJXh5ertX76zVQGGGhTzUd5IDBB4o225cGTCwgbzz78n9e
RwS4/TK4ggyl81OdIQP0ziNwP6TcfwwvWAor5Fv61hXSShpA1ru5+Wh4VgCdiOQ2
VMpHjYQsoZY4PtMKYEhmF1Tz9uKpKaJVaMJxN2/5Ay1zKeWIw9xY9LFAriouYROq
eBKQZ+ytt4yuak+JQZmPT8YhV3eW88GJy6LgcGG8VQMokAPAb5fiy0gvBYntxXYn
TgixZODprKF3ts/r4+z1tJc5Q4mywSa9SMO6D0bSKGedX4yQbPez65IrQ01yJnkL
gpWSRg1nXDqg20+kWJugZ9/4Vc0WpXMqPxExNUy4AS0AQN/uoazt/xDJ0nyTvRrk
RlglgjUFYri6ls3BERRgzzkVhxFN15leMj9r5CbQIjBLJIrWQaFza2S0VtBTwMjn
eCyxfo34K7winv2V49CopHIeC1xwoN22jk0Qo0kE8Z9JWVG5JItWtOcFMm2hn7DB
fzL0jYG9hxtOepA3B4TVHZd/0pgVOMk2hhS0iPkwQgPHUF62TnsmkZ6oM5QeA6nG
HxQPZlhLkvtpqqMrltjDRlJi8UCgVUtbZKlv4ejA8/69yLXXIJbemHVuWoTzP90S
weHbgdu/9yEjTj48PHVwc09oDkBCzg1pNecjblz0qP5EZe0A1DPNSvFMXy9/aHrM
8lMG4paRD0NahQk1Z5RLLpWVmiV85e1tYBEjRDOfVhQWH4R4hg++vOXHOec6a+XP
T2MWSGt77TwZef9xnH4nOAUrHuzxFjazoky3pQeBc0ARpBIUUABONNjd26b7PSbO
jkze+Ed2eVtVoNRN3joZWS1fKbnWzCfsUjuiIVJNRZv3INrw543KvNXKMsvWIEZ/
pDu4IephL83DWw9LAkwfIN8OtaMAzfWVIrBiqQYQotvzzCO4iCD4dECInG+JY0qb
QBcgO47YpvYjUwr8ty7nqKu2KABN4UjfBonwML0Zjzr5TSdnaDT3UBFToY/+c5dL
rufagS4dJe7bro93BJZh6Hv2pquqIRVWTc8psoFCHTKLSB3C29s6+A5GDayFTf6n
q7iSRjkHNqT0t8FwOUdLWkejucrCheY81EKRwWNSYfK/Xr+zzY/UTYOn6NaF/gnm
9XmQ2gs4GkojxCs4hIeCDqO634QRswbSqB1PLWnuIOpwAuFSPFczuZy+fqxaYvWB
FA+s8bkY4DdsfZzM6mc2HIkq81yXY0qskffgKWs3effuJslsCafSWil/TFSFWEPH
SsAwJPkmWAT4J1OFuS6ZkfTS2jXfA2JwrDUws5qWpMuBWgpALCfEuhatXBUrg789
XKwD6Cs7KjfdWSJis6fBXYUxvPWd8eOrzPHtub4/0cBywrPHp2BCjekYFoQ8OxzZ
rHJyXKQXkUExa000s2lsiGwYPME0sTjIJlIOynr/bK595NWXcoIr6gZVff07Gme/
5Y7P21M0MDoIVd7SJ2LDBzW1hoFehPLWlRNE7tboJCez58wpdrjT+b3ZAkv6qarT
4HlamSxzIueKczmNZWipYz2QxTUd+tsgXcTfuuRaZjioazatJhYlxGJgyRlWiiVX
JEHvnxcEXHWndb1rYFyCrZcVypt0h2JTDrufem1DAAhErQD9+V5PPq2NPFOqMeY0
qzcF7tmQXb3OzubeXWaVHvvg4JxWtPM6jKUCTzktGm+tahSRod5MveAhkUSoVkhX
sBYoJybLuH9ImPKixo21kWzSZU99fbM5nyHL6BVEndm/Joi61V4IudJfBFbF9Jfh
Xcdd+Osqr7cbsBTel5syMfxqMbg75jzq7gdU/x6eYb3JYtZRGSyYyNL7d52aD36S
CgD9hrFHihciN2yQE86hhH0WfZ0S88EGToctCNaRUBz/GGaOpnDRnO319xUYkoO+
NvEBKIB1i1zIhvuBNuyqT9iOJkWHjNQ/VZuTbhW2oRCsjIrABmZoMnkkKBKGs7q5
05/4sHEMI/oTES8ehyaKKDK8Jo/ms3QbKKEEGYyxY/YS60yPr/Y7L5B8a5ijiEuw
o825BUUe8z2FiKqfFlLhcYgI2KE5HnNEr4C+YnE+vdn2E8i/iO+jOqrlKLcJtHEm
MgC+fj7MEMPDnuADVhkGXpVJro+C8kXpOSaQiS1Nd57nL7eL05wmoLtUZInO12/+
2RkxtcCuoDIQyenk2YkoKYabG4YyzEM7K9meUfsFBzvU0ua0mzctcc292purvfI7
NOcT30I8PaWkD+2P6kv7TOJV8VwtXDisFYAtJX3qxZGn8YWDqsks53BXWk/FHUNU
N46Hd8k/gOw2bJJvovoPs7aLUzpi6jBrgmdAqRyBISFFjhQ8ajQRSVeIrqL2u6W+
H6iMohrDjTnVpfrbxDdPCRtZIOI7H1Qe5ndMdUJnaHGqf+r6c0Srmov3/oFd5kF3
7V+EKX3KhFVq88JcogEBRpkO457FX9yBPMo9aG4q0jue9JCEzHyyOnXqqTx1jx0f
f6vM4LU9N6ZFfQjaavh8xLEUYTbnkkupc+77UEqNxyNWUqlmagmoafxrP8sz1Vgl
dVoJPJKp7DBdplge6QaitOL5LuURmf/0xhgSm5zxQEE+HaRkJtTQtPbCFx6O094U
NM7Tj2wZMurm3Fneip1BR/SYG+brj7M84kxiVnbKbVVqPPm2gdl88rcE8j9/Wtlw
6d1z/qjkNap6ypSS24yZmYIhKByH6HwsTBfr4dfNJ6fSNDiNtr8x2vZT3y1khBTJ
xvugAYgOlRdP6L2fIpTWSbR0VnBOzgYWvbhJ/pvYuYn5XmoYY5f9gJixpsYskWLH
vDAbltbBrEdcwssrReo+nyLAsYBVTXumekf7aBvqXmF2+B/r+1psl/XlRznriBqD
NBaKZ2U4JqtwFPKTSS7yf9Q0WtqzKGIYyDOgbegcnR1cNKq+v3EpVyhbtBf4wird
ythKeUoTppLi2v47N9xnKI7mGW3X/A2FcfXDM3GEPp9yY6718ei+y8w9er2WI8Xn
jX8fk/Itkxy0MLlHyE69NuDJP55hG5kVH36aMTBXRcT1M7ntS9MCZOzxLlLniU8O
Pxkzo186MYOgtd2verUtkcgqsfFpaaSWq4M7CF1SH8+Ajso97FCFKpRZMkNM48GB
27FkmZy5VHq6Fex4FW9YUbnGncFRBKJ8DibCZJdYKSlNCeM8wVkBXKFeNHsmLWIc
PHyo07WYa+DZpCVzP2KfC9XcnHkMOxl1qwC9Ui/Zc5k2X3iQwKoSREuOOPY05421
zlE19yoy26zwkTCcLHh3bgTN0g6WKYx5R+RdHuegT1jMzjBJ3BqU9qqfkqgu/4/p
MWx7nthGCiiOdOV6S7FMD+wP2MNiu18c8V+YgA+lSSj5n8ba6lDNqnacyUSPi/vZ
LYx7+HmcDptAtMGxfWRq8JIGThJWE4S5SjPwLmE/fsNjrrwFkwTpmpmNdV+u/7PC
W6FxT7ARHlBqBzegyOq3MGBvtWVQn30fSBQ9GeosLXOvNmxRJ/scJdVopPzbPuMq
GhMCT1UtwXF1o8wM2+yI7RMzXLkPp2dQdyUzR39fJg9YZy5+tEdUajBt6SuvYIle
um+XlBK1R0BMD9pW2fwECwQqKOEdy8KAWzYf0iRDDdQnQK3urTaTLKlD3COztO8E
RDfig+2ZatWZvyHFsX65MEPpfrMi8eyaUM/jxIbmXXYwSVWUfNj0pUmzmdNZhvcv
gsLJGQ+t24AnFD5xb2PqhwqpIjAj6+nlBsdSfkCqgMObWSk60TYaTtnvJJ8RGPK2
WoOZ6Tz40z1AaCaJccepHzkPCbovZTZl6tZ93mM6j8EzSIrKXSqBOJr+rtln4iF/
vzFARkl2xCq+5jjIr4BJiGwXNkFqDNJCGKqmTCXglDdo8ZUAEqzjTZccc1stZpQk
ngGYEhIhOteHkiVXSA/IoEv41xZxMniiXmxuM79K6FUM+lhFIFS33u7lvvAs2d5C
WSG8SgRRFbSGfxwcURZO13WE0lDpSV4cmTbJfsDOAnGemlKyemuOagSNuX+OpvYH
jhHUYusRbXJpifu5FSmYO6ChAJZ8jlHtMwbxiew7OOBrNuXUkO3J84D341H0zLMN
RLfh0kMmxVdQ6/ainvXKTAIc4w/y7UsLarp/47tfo/Aaa4htj42zoT2mkqmsZRpJ
HFp2xFgt3pDSqmmiSTZCwk8ZkQlWfItCa6Og82kcxD/pvbEGZ67WWOqsfXB1zYBP
9aOuCHuKG5QfCxrGHy6LsMeue6BkFuW2ET0R2TlTX7xmlzAGzD0fLtC+FG/PaAnN
rIhrsI0wVDzikO9bDJPwFYQlwLAo/Og0A0gGB9MVLJRedIJ3Kx3rMm+tFcvFbtui
W4I1jtp4hcafJe9qE0Ckiru14ynwoSOIThru91kBHerWAEhFGbAOrS7IKvCWBz2Q
rD1/pmjxZ4Vek+eyp4IE+y9ByecbYTCoSt3CSPnmK0cTuDO7Az/6O+dZ++s57dnT
XMrLQwfhLhWDllnVsw5t0DQERkJDW8ws7WbnZkG7VtQlCsZ+E89qC/vTWiRN2hEK
U9PUdhmcOZlKe7DoFHYzPCD8GPW1Q1jbDKlCd5UxV/5XGjdpgfZG7xTm4d/DwSR8
UPpLUPdXGJfD0xE+rdyiP7Cygw+/pBtmBUqvYDQu5Ie5b0xKqVR0LBuhI8I6Jlcx
y8B8sA9iABa+mf3djOU30xlhoMh3MecmDQQaTkQMB2yjACdoEJe7+0dsMBUop42Y
QHTxQDsgws1VlfXep7tiXg0B0CaKRlT/lkUJPvNEKLLlUIHWPtttNE1OVgRtuYXb
m6uEcCDRV3grPnM8/xkgtMrBHiC5eR3ARcQy+ThC9a4dEzB6GRfqP0eVl6X/SpbJ
cQ0knNEtKnnbCuUePz6EDCl5jBCAPsyemJQJ+aDA+4w1qr0Pt9Ge4r9KpbwMprA/
acb75tEDsleZspBPaz94Y/y7OQeEqZkTOb4JKPprkMGkamltWZkAngL60JLMjXNB
WvGcn5d7Zeu+qhvivPWMm6UZ8cITcfaB6p3OmzNK+/IJrOgZo701rVn+cZDmBWTC
O1w7CmXBHika9N35u7Y4xH+HBMQuhBTi6DTq1bHBLA48m3Etjnh057Y5UOsLGFKk
e8kXdiM8ZOueJv7LBvv6ZvcuGe+ZmE+jkh1V2oNpTUso0sJ8qH6UYO8joxP0qpNS
hghRzzf/OmfCnFSIE4DProd2MUcXNi9KoC7o8jR5BugC0rXKime8YHeaPK6IDgQo
KZTxKIyCzxBunGOpREkfUJ+YFN0MqfhKBcghCfF7Y+jr1JuFHDhHQ5qQan17/zJG
Di8vxgeVyBptC+Pn+TzIQVeOmj2t25oVHC133edNdSbUx8q6h0ki5TE7X+IdaRJG
X9xArkkhCH8i5Dm1bpB3/BydYrc8PtxUrXRwDKjsE9FG7o8Tgr19a/WUNjUIFA5L
IQ9WgVobBuEGR04vIQDTDPJ19KHK4PSqlF8wUQjwq71IHqGDYdyAnEwy0woQX0qj
6JqTT0Lr+PWjFEhHr13G+EXJjDwdoUuDTJgL8+vjR5ZDU+czisTVWMRDqlMbRivc
Og6DZ4NnE4v0mWmE7fQTQCvkhdEYAo+oI/29SeVSJSRuVOlsl156AXj85o+5ayRK
Li87ApEqObPtcGGJENuITdrvdr5stam2tFK13NB/Bhdw8G6cTE7nY3pBQhZ30/nM
hooTLaNWUQBqHfKpMAF54/CWjOGQYjsGSe473LQx7772L4K/gk6cAEmuJUMfRYdI
ogT+tLaD7Zacw+rl6j1L8K+MBaDN41QRPYHujemUuhMXm4/A1ZwJUvgu7hV86ehK
kCJr2ozz/V54jOhj98w2iO+NaL0iG1ZGoXaVFF6YT7rvpQtO00bWyzlF2YdBgd5O
tsN+gWCghn4kkI3rD3VtX6yCpuCkOEP3KARoqdCqAD8cBJDHEXb/OPT8LIu48MUy
oPHCKWGMSWsDMRnmX98I+49Zv7tyvOFuPfraFV8CfQWE8pq4IfGRDXFS//hHydyo
wa7WqnVH4rf+K/HQU/ETW+CAKxVBss3ykS6HgZCJ7Mi62khBUlCouQaOKrtlMenI
ik0V5RZa/OBr5OQPCpbVViJKnOUIWPoParzN8uP8j1TBAd/LzVTF/6OGHtlWw73D
irBVM+dVo44dYLLB0BW1n2EOm409H+m7a5BA6vR2Fo2ufxuIvHSbYJTS/636ySHg
HmScCVd8XKOj+LMVtCIrdi4+3GAo16uOMcII55TX+oieyzeRP6yDAuocVp1WTRo5
cdYA2AnRuEaye8EjgUmM2L/Ef0AqabSmXEmrzkHcuLQrg7udaaXrmfv8DAjjHMkg
Xi7uavpR1xGqBZHkyGlSBoqF8cce1SorhgY9z+hzYDJeHMipR+91B8wDMCE2spac
BAhPZWUX1qn6flH+GKE/CYryqB253ONJ4kIRnjTpVu2xozgJFpcK44Sm7VRthrp7
BqPH85Zv8rFNGxgWMpxh3b2ojp5qUuQHXZJchCIXx95W6vM+cHAVu3b4uMeCF2T3
duvoF6SzNQtypLViAs+g8N9D4Gt+JbX8Y0LLFDlISDLsVE2G42o44wqVeHAClYG0
jPm1jp9ax1bWyUigJgrUxnzKYoLvwDpe3S3bwUkTlWz7l4pQH71W4IXnaFBYfgvT
8i0TfMdmG1FMCng//Q6tAxcrvNP3khMvVJeUjCGxtNv61zSCBd6cn/+pFY0q8zEx
gDXzp5zX2WW8qyVlL9XWG0NR6RV6B/hGPau4deU7AxItB7c47fNEVXzhrJOp0uhn
GZKAkkJvB2HvlyEPcLIZogGBUuJskYihUUe6N/zUDS3lmo4/vU+hu5390LF1xk50
66yx64xRU1F081Jx2ms5aFkzJ28yU09Ir75cqfUpwZCxrQZXjEM9NR2eE8vfq9u1
mC0bVBjrXLBLxBJseJGBJCTwoA/ZEqbnka9E6EjP+cpZmoLfFclVqdzf8C99/hub
e4pFS5ofbQA+I+qrgfuQuVreqqF0beBZHdA/mAzuoAZuMJyvHJwFvdK7W4sjsQTP
4iDpmOU6v3Le0UbZKPb2wJLrnQMqtmsUXM9QEQhzcdlj7wT93NslF2MWGYugMD8X
QXbE8Wu8EOPZY9HY+BFJFO8xFANSAMqwL8Cbc6kIPC/0nxkqn4zKvnel3Oa44NwN
tEu4q6eTM2kNHwJPfv4AQuIf3RMF4FK0xdXEZCp+cvOP1yDx+z1RHsVVUxjB3FWu
0mSe0yj6rLi1E+APGhWphN7MjltdjGdekT4rcLEdBCSc0rd8QEIsbcdCxv0vIO+f
pLSTTo9Kain8ICoGzH3vopPpvk1QgLbqDS8mpQ96SKiAwqQQdHqqvxhw4ofPJa9u
lXQMhFnOnz7jvEXgeqpO+dvyW8OE8dS8u0UPFjg6ZH8VS/4adiEMgdnGqZ1zgNPV
2Pv+d9O5LY0vZCexNA1tW2tHZDpysS0cIBu2Qt4RubuJapcX4QrAmIJRbefRrAgH
RB9i0JG77+YGOS8YTTPj6e4iJa41H8CA+g7gDhTvBencJg7rudMueoYR9lpxT7HE
otitK19AYtN3nKC/yZuoevMIh+BeTEgHimv4llyX2BZLRQbbddMwGJyJga8y4jkL
9DE+JnRAljwlotEjw1QBDCnbzmHI4YTRpRMgoYCv2WCBDevKGn8sA9D7PrIFCOyS
Bw4E7PcmWl2l3nDLKGl5Clg2oAxK3EhHAEOouxn4ow1ZkwZmhm/JnxtpUP2qQD5m
Emxf0TxAy34pxAlWlWSF/uVprk4Pv1gJnXF4yaFklreKbbQym47+Nno3I/uQDjaL
T7cAHXkWtslU8AumrtNviL51iMmefN2oEx0tSj+7VG2C/PtMOVlnNfasBI4iw+Cq
be5cpncR1SzAif+wpsf1ePGyxI/hmDyvPcmAEUBV+TG6dwyOvNqYzbXCS7KjRq0y
NUmavV0r7gPQXnFZ36oe1o99W/PHZnk7n7LC1ae0uUJ2y+NbbviN6tftgujfxJ+k
h8D0eWF60R2O2GXq0OUHRHawfd87bzgdjp8rIfGktYa97RnvJa2tnPPWJY+nOaL6
eJExwHFInDEHmxN6cqxij5I7QeNE9/tEv4JEeFGzGlzNYFGhCidAwUv/rtmnScT7
IAnEl3kXxmLYN4BOhdSXdOcU2j+wfnWi4YVwzVt66HI+2tQGj1xJbf4ShaBWJ41f
zJaeHZ2ixwh0SQ9eYMKYYF7UH3ukmUzaBLpzEJa4e/3gfxIw4UgtW2RR2yT/UR3P
zUBOneN0bETrt7CVta1TYkPjfl+op8nWvESt/2iQanVLv+CKGmfb1nKu1+6rze5+
USueB0P1TcZ9o5holCYRCo4j3AY68bcOfcmhoaFeQaWliE37SPbKCawblSWOBm8E
oYYi4CaiMiGRXFQwv4GkjpCIJ3fyb97x5rCEamFtTjDrCk9RVH67eZw3BwNSfOsO
90Y38Sax9smhO5yLIAtrXrVa0Pvc4o/kpiUDlkomyqrjPvPe42Asiok5Viq7wBFw
l7S5A93szvmsBQithYDBzVL26+zRZWv/Ez1CbhqRC+NNMYUXBSe4u+Ajd2MEvalI
tKxw9BMyX0wZhv4Gp2EUT0q8XBcCCrPxZjTzqVS/+xe8sngTZ85IB4CKlkQKo+nq
Y/f+1hRv1NiSNRGNaDuoXe2SCSqAS8fYw5pnwQIAfJBeFo9AEJynBDP5yCuh+Sd3
8TiTBvmO1tSy8b9cmkOyYbpKNqbDR2hXpBiGwVgFpvLTigK+sBGS6lizFjPkSD7l
o+l7edavVPzCLCMyNlvIzgIrXA2imcdIWhiddMG/JUEt8Kpu3jQLa2FAuGfe+Pjv
Ms6xRSoJhgy6BjbT7YoReKUtZ7QbaSN9CD2v5pl5gA1OshJz/6xf8UiC1jpAqLmY
GWWM9hW8A1Nwq+OYXcoQTrb6GZE9BMy5rpNm28vnXQG4kBaMZPENFVK8urI/DGch
BeMCyN7jT8HhlhZxUaVhkUK/OePXw/kPdTqZfLYvpEfUzYN9sZBLZjloJZszZ2gj
DaqSTtQx6EJyw6DdEAddvXMj9KflD5DVvzCRlhcyHObex1vzWS8xVaRAfUr7hsQY
Y3hPc1Z9Qi/28kJM296tM74iM7mmhIQCCg9R2UbejKL/vbp3xLI4Rjd1lMuhbxsN
2cCwKVkCRb+YtoP0boOF4XyeZIlrbcIJgZbsbJSEuiosTBZdwgM9W0qmc1fm7U5V
p1RgASsg2+gvssPtc7d+d4IoSjYzwPXgCbIH8MrthMDR/272qvhuPVODYYQdBSTh
8HvFRcJqEbxgwA3+JQD2yD9oJnKtac7IerTAA1jm0EZXuphMymbNrOvvxwWt3xL1
6R7jK+eCtB8P0/nTTJJDpWJA2lfnwY6tOvUed41g8eE8RD+8bZPavxmgpS0cCkem
ZtFw5UAGbyz0y9+1+i2Jp5JmGUCd/WXKNNEFLSlwPfdOMvlOPvvKIPNbp7w3v9b5
L4v+MAeaSrqW8+WIY9Nf8/c715nFuTL4QZ6nnK/JzTTbdFeScYFwrS2ws0tqDgmE
2x9l0Q+cV/SN6S7C4y77hkYzheW0g+1Ft0y+cBpwvyDqv0jWV6rfvweFgTBQSyIi
a6zHiwo1w5Sm5EiqjFQ4hHt+0ftnuOsNbEqHm3na3xFdneO+tQAMJZmLt3Ngc6ZL
zr3iBlPapsKaWHbQOgnzpLcTJW0mcO7AAXVk0yYhVPzNSt6rI5m+Xsl2vRdisdZb
2fQAaxvwVamVKmqlkmBvgvufNkl5DkfTi1n1EpX1cEAfeI00Rlfo7TCC5mgZayTa
4A/3d78sHtUSaPLAt/RpKGiJHX5Eh8Urb8lscRorPZ2CG6OwoJCKDTQTb7ZYCVr6
jmSCRVYQ1aSZC56OmRSJrlTKxoi+Z6S9X02+9Qn5e1sB3yPekBUot79kx+ZWJgh9
D8PNpEWtJPq2HpGR7q41gGrbvHVUn4w0x4xZxbN2SN3uDVjvKSSat/NVdk1VYraj
R7sfhaadFIh/mDFhAB0jElTpjvHHwhn72YHy0JzJzWfPuS7L7HAHcvjqi1vDVDSu
sPOfe+k3dJOAmP70ZAFVbQjtjQIGoOjWGT1COMbCKYcLFpuRoSCPxJFn1g3MqGV9
tiC5YRgbtQflviYtgtH1cMp5w8lz6W2cG+TlnQLBXJtBF7PFvVSRzGQDvBAEM5XZ
7KPEMeUeF5kY70VZRO8agjdJtOG2/njpo2jA+/S+4wZUsOrO0VwyijfUxWrz4E49
gbZylZcJirVUwT7aNIqh/0qFt+J+LFwteIasgKsIvA+cj4uuibBNgwK1Swtg9Jk9
MPo1pGYttrV1Xg5EhDC2d3tf5NLaKD0kTYdkrLWpDQeEQvbXZiEPNg/qWOPu2jlL
GTKRqgBMbSmo+xkne/LUIwdx45PvSX02jt8fDVASABBQzp8DPm9K+Z68arVPRygH
hcXQvGq1pCGxJG3E8mZ8iCq8Cf0AkDGvANrsoHTu5ddnegBHSy9DJKwcaRG3mmfd
GoPh71XpvQK1iG/Ff53LlGvEBT8A/cFpz8OsppXSwzevGmXWAmKWSsbC4Hz7oZV0
wqqdygWiiJ1vJYzvRK9ru9MOyLwLyt+iTqPY/whiJ7SOVkv5mEAhlDPvpqRBQjey
m7st/8qMN8J7nT6RAIhtEFMzj3D0MDoXnP8gS2rIxWsAK6bb05lFXoa28rMbrWsh
U68c42QacqHInW1i512N0TN+jNJnsrSUUw/DfzeDyYXvaknu7Q0O6x1Yx5C9Ccvq
yY5x8vD+cQPB4Y0bV1sRgiiLWMANdMFMiQ7/mMvrDygQYZyuCGEdbjfFSo+v+4zj
jJl8fEOLItZH/SvMf9RO+7UiJg/kvcOxYEz/ADJIupuMnyGzqzo6iGrV10T7ZWFS
dv03i6IwTVtNzASPDN4by9SikJafYrQ2AtiwtqAPUCK0qV1KhuBX+iduqpZL9TK7
GdJQMv5QGTuymFtvWtGsHFac5qyXxK+FUBOSaHCP/osgQr3jGPpGOb0enJM0dtiG
ZjpwfexlNA0cKiXWAqqbiK6TnfY6UVOL4vulP/TRh5sdBfwBbjLEnn67FOFIdEqL
VUJUGEMealR8KBN+nBvdyEx4KiqXdisd3wJwZLIfZP4lOLhO0VBj14cvsYw2jskB
ItVquTbu/Z/rr6KBWDf1+M6ffvTXWUKxOHxet6fdNpuBPkLT4hsFjaLiSFsU9f6b
NTd3aWoT2iypGcz2dJoFJmYX4w9GmjJHS1+JCA1u4P2XdjQ0YcbS3F9bwcW5jYQL
7Mo9UJKnR2vU1GN1vdp6VGcMHw8RjOYmPNd5TZ/GGCEvCbxuCxWTWSsGI7jsSunY
04uwxbmtenRssOROTFjWvSMdMTcOsnXTEVT55BYIdJ4MDAy0J1KNu7wLzXXQWPXD
3tngGRlLWiPrt+lYUbAP+S3Lo2WIu2OPjB6maW9NnbQOibF+jJmefhQDyxuksVAV
M3l1+SuIpk0LjVR2NR2ILFJH+/9cZlabpzPQFsJ9+CZaOwAaxF4BMOB1B4IjAzfG
KuNoHwY9WouyoLcpe9/wsBKO3nUXXSBhRVx1yrzf+0nWaP+cJt7YweDGllwAKHVv
O7xM7plTVS5Vy/bmFtHrfqoQRUkk8L8ax9oevvIiqZbg+Pzgj+f6DBeCj+Finb0h
vczSiDIE4hQBqqKPnuE2Vs/2R7THn5SSO3wBx4l2veOsqn8WSDtCqJeyLEnOD8t/
Oik23CydYtX8u8hSbZ9ALb26MnbRZdZHPQYZjSssouanUvHs8o9SqruBqi9F48Zf
Jdr9GYlJePJU8iiF9vRRb7ltdEo1OmDp3KF6RPWv8ZSKuKPjo3mBWunGTibtjDgI
6FcEI6A04Z8ISjVi5vqu5TJWIa4bsUTxy9wJ3BYVefsbcxz5LVmbaEyiXtaeDAXh
/Q5RN2jqubdleA+D1pibfym2v/hG9TFvz9P06druiIZWQvnY4CBsBSeJ8LHQsvGO
vLGnVfsFNpoIGWd8ScTPns1JXIIozizmOvuQSVBycIAF+I/8nSEVLkE58gGtjuuv
XxkymC7iUFQMhsbMVet5GVfPxHFA8Hcp+vlCkMILfTZkhZ8g3g/CoRxBZVQEt5UJ
FGC5zZqH1SE+mS3dizvJn2hSgtCxFW8fQxz9kYAkCp0Ed8XensL4aavbia194w9Y
KX3hT6vY42qU8D0BhE9dUuwOJ7JzsNS8c1L8snhLyVaFHkkYOLQMphUfZgI+3V4g
wp5A3EG9yYI/fKzSarLpsRrEXmZsc+HUYPMm1veGZ7ZOuU80qsq3qghLD3+3BkRe
gGwPsf9ezcaJq1CbBCY4z2myPZqGlUSG5IPIuyF1ZhJ9eRk7yJkCRKzRrybh6TZU
NMEPHqVIXmnx2ZEHsNUKCIkvPHV3HCKZLJzaxheCIUJD0Ils3kt7PLkVRHdIKnVu
nvaH8g60vXuVHC3amtMgFHURhn8+hEpLXFxvjfcbbCfglCVTGJDO/2DrS4pT6Xho
iLP2IvNY9qNCI4tMXIrxmJLy1CVmn1bs8acbgfnHeNytzV0SXksyVxlCDWt+m/Kg
0VTC7y6EWrjgcwwSOsikrjNKqgc6lM6mc1ICVH88+RUw7r43oFMESniVhZbDS1Ia
aUKbW0j5IbR1kE/4I45vsctTHCj2VqT0WKcFaepttezZCRQz0E1Pj2391Nr8rCRP
s+G1cOhME21MlTDNXU2+RJ2Wd/+lKA/pil5zqVvtNEoKMePcy7XHJaNMaPAi2iDe
IijptTwmdAkYIbgqp7LybYWNoKjufffMZbEpglqO+F1arpfGz3nxBno98NBLhJfN
jKp1ZmFCkqIZCO+jfQni5k/JMxKaI6KFx0J1XrXJXIz/YDrYa9OJ60rpZArbAO4b
eZmkU4xO9xGuKpm13ioJbCzzdYUKhEeVvQcs8voNL5q6jG9DumcJ5/fnKQ7nWUus
zQ0YvnbtPSU834SjCkfiPC8NF7+zWd3md0+ufGYtP1eupUxmxiTaLA7ueRkhYWpY
gcb5jKzxfRRt4JTwGrdRVIaEZlhlkwMU8GyXbAyOd3hJUwW82j/grjSPU3tlNxEJ
nAcCMRbWHpk9gehgkyCsJnVkN7pdaOnZ+ZLtShYecZvgqsmpkj0qCTAgfeVSSYg1
aG2lWJCfVir3VucE+r2RlCODIwVXvMn7bnHU+DcoZOG5Pnjiq7zwjO5Z//lJlXU2
H+6aFfJ67ChRFdght21RoPuAdgj5vTwmO3r2VJBwlJ6AjSp7qQGN/LYSlOv/dcv5
jxn5SqfX84yq4BDPNsq0nKhODzzAuNVw8RQBgPU0FHyAas2fU8OrO0CsfM4A3PB7
7xbnIezvA6K2upm7s7he3cThPFMy05FC2WF7S2krc7GW7aodhs9yP6tcFpz+DGVu
lsqRDM1IiBfmaUNBHGSfomu4wVJeE5bAjQLddZSFosiNVvIef9uoyo3mHf8eAmHT
DuwXPvc79prQBu+lUyFFYFXOmCYw4MiFYYdIuQfrflsTupAwNb7UXc58mMk/vdHt
s0WfhHJ6PvE9tFPjnSqYczSVW2/QB7OTt6VQs3YX+JKH43seffhyG8tLPoUs9kaA
Xr4YyKb5I4ikaOIDmn8Con5fgfcJL5e3opwql5jiuXe+e2w8/3TIvH/jyl7uRhSO
yYoujmL94z8a7LwGocdcpotYN+KX0kYByR4Hoarc9Lg2A5eiQ/3ExMpZuOLi9d7+
/+Jv4iWKLPcYjAALnBnlq0fNu/a/zOn0p0jfsv6a6hyTmNzDF7+gWfXP+gTi75eF
mACR9oz1UkpPvxv4UGyksCNDcweiOgTgJP9w4Ay23N3//Ypq8nVNuMRDBgiF9cKq
yviBxXiWNtmnRn1CcRfn2HVOTL8RcSruzUZRu1ZpVdiM51/gvbzNKcyT790W+9qN
rrXP1a2a+tiYnxwkMB0UctQY2a/eSHjLMkj7mXAZsZiUOtjf/WlBaJ3W7KNe62lh
6P1prEIltaonJvaxCz3EtrrNCWI8Emt9TZxLACRix/jjekhevZJpSrj/h0JmQzpF
LYayxYZIlLgKYGQ3VyQzx+gl/tncR4jT0RCeHdnGuvZknztGiAlE2evS9984ucr+
EdthphNKWsB4lDIeAvuXCzLMskIXnpCBhdShejf3jeidkjRAMTW3rbhE5N4XuUl6
iJg0re/gIPvv5S/ymNWDB+qjleQeUrKrQhVWfdVWDejbG9yyHagaBqvGRqFEt9aY
UI/tG/nQ8gHkQlTVmliemaI0UmaNfRVOIoL9RiR7BA/Yj0i6ZnG5tbvjXAP3VQlt
ZLYBJDYHJ2vbLDwr7b5RAy9HJxUghfPBjZtbxxq4r36XjTHKgvt7OOG9JKjfgNAy
QFtAvkEEcYLuxw/ae1gfPO7FbDjy/+NwGfe7hKpwBP4T543rMeT+bmc5cAQwY2h9
XSBcMak6EE8V1TBURygFF0kHUbI5Q8fJYLtQrB+hJpnRfBLVVadN7+p+t/v8tgN2
lBpwT6BaMPCyBdQe8ZRl5hzjQr0vSFE29dxMN38lclccFMa1mUyMlF8/EDRqQJWs
oKMJY08JviXJztlG+NBw3SnL+uyLA1No9FrnKapcet9MbNvW1UH8MbaxbQUx5eDy
x9Qe/3KQ0kiqtsfF0KKWBEULauvp5RaPUv8/2PIEerI6DLKprd7idzU+vxMvOc/F
jaNLTVdpFEWJvWewMMzQ7+KGdHIj4rtxlQcKdtz/KVS2Rj/JWwQEuQRwa+TsbXJB
jeDT0ASs0OTwmSsUUq21ATjvh1g9Rnfb3pSz+i0Mh5cXeLk23V+Smxg+A+EDzeC4
5zALEIwZx2/9hYMbFqOcdCxnzNg+vLm6WBNI8R9wyKLEcrpy85lgT5Nagdaw6RmK
zf4AyVfyqBMYQHfPWnT84gvo3uib7Hbgda9uisaxJhPtafobmdYeJZm0sWpKyI4E
MaImEcHsTclp+6onCiFu2g9rF169BZvCyT+FfBtrsvO8tSryE6plQCgHRDdFZndP
0Fy55qYZGOLbuekQ9bTK7rpcBP96zLwX6sl2EHaxRPPgII0TTg6ZQn8CervJfpow
13ncOYybIXHqYpRBrLm1uVxASbnV7SP7YW/qXkNtfrMmMbi6zufA6L7ktzZxvumq
Ja/3Calz7xlg4nalGd6oHqL+ZM8kuiU6oHTX3CgEMKQatA2f1f4kyOJi0TTPA8/m
bxelXoDJxLPP6K+8IZPttvdwqDOyqak4nZlqOEQoCwJNqy+fLxVnwbgKeVR/77Fv
DOlpwEMIeVtWuewIQuT0NgpAI9sxQR0khlvmpk6JMnbSEmn2FpuLccniLLryhpoG
qN2aAzjMiayu8OoabL1qJVkknVZ+CbOo9WGy7YswRkZh6NYZrD89kARAwti/JYPt
B1QrNHTOCn/duLvwuixA5x7NXP0gnjYDw5sfPvl6B1e9DfZDVtmURHqDu2NdNbNt
x1OuUTbo2m8T8nzZbM6tiOYc285wM4O0dsu3lEGSIY+SJwYg+hFJQP+2DcuXU/Ud
0f7CHDpfxizXBDACSIIxte4QzEnduj6GyVNc8UkC5E+3Fk6OkrEoQTh2M3FcxgCa
g/xVCwZHHEoajs9DFZ2Hvculp+v9Lbtwp9dlgiZGd9vdZiFwk1t6q0mVf+EEA3QM
wZW8A/hcfLKtnMRP/FWtTFJJ8uMAwreFHh1N4RuW+CAfvw9vZKRYIxn63tkq5Gza
M57jjXYCg5r/EyQZ+/f8yQHNxo1DDkYGi4MpszA5HMeXQ4JS6OeD+WLrkSNDOwCP
Cj+Q54irlJ11mF7zCaL23GhbRnu4nJL6AmkMJI2Oluhsuqz4kICH8dQQFwgbz8R4
o+YIgOw3T+CcS3o/kVnGRdimg8RAj10nmgFLFHYYE0B4likvkOxFEs69jmt+MPn2
6HRASn5UCJU55fuv2LWHWiyNRe7loAEqdo74vJ73ikhZrkCDCXVZIN9eO78bVV81
kKIbhLpETeohP1prPattCslMfg5rXbEUDRweLdwCCde4SK0KwMib95Sb1nx5eN0V
mU6Q6oggjIuR3dR1RKE5WR0d6aelm2jexVUjP3o8MklROsD9lC4SMkSTvf8ebbi3
Y0GpNvsZvvOK0Wocmo2UpdatqXF4HVN7lWJ1335IPJmbmGL1RqUCBKpWLz+oLGir
qkIiEkSCl1X2f3jki9yI6fVUFkyjIbsj/hToSQkK4K4zeQjfdBdTLbDkabk6ClMz
VYCP3hkyG7xwZzWjOKdggLjNBc+WIUuzg7978efFEnpp8RkRscHpv/O+0J70ulNi
Sdy4hexvIiCsNbqqGUV+Pk5S+FaXFDSbaXPyydM/Kb2GmwniC5o+iyjMp/pvs11C
Z7koYIDT9/pWegmAEf7SiAjETLfCrJTJqNAc3gVhT+p4M2FmUczSgTsLEohb+UqD
m8DLMKBnB5BboURyCusS5e1mFNeaR3UW6OU9nRfX9bYDCJv2jnigB1fP7PjfF/yw
NzXc8mU6Te7HGIeUvAmjhQTQbzwIXnbF5sFFurqvaV9a+ULIzQhjFWKEAq0/8L79
+qes8VYx9o1JkKlmzpQ3ZPzArvFdymLaqTWgmrRc+BrBhbRjLztJPoffZW6ox+80
2J0EoE7qLUywC7TWCUNzZxuGNp8owjGkAkCN5CKAe+I3/0/U8+kJ9wV+W4hxz8rB
IzB33ctAxBFdVlSfnavRejvAx3ly1TTRB2FIfHuptnTd7LqRDQvkwAZYMr85Xxgc
e+yLzp/zTVXaCwqVSavJ7/QILqSXMtAD0AFRpfdbVbzFZDo1Cu4FnWkCCzbe5TPZ
5kz83ss4GskkKCF7faoKWNRt9XOGRNkFeXCEzpQm3SmVyT2Q0llwZAFleaS9ACEz
/1wsaBdvGqPo8GT3vS8CifWBsoVnJrEbe9tZRdbbP3Fwv0hJoctxwrYyO14SujnA
A1lrrEP+37f4Om3hWbE/ygk2f4bocvTpPHZdarvi9KbHYNkKwb7mNwetFbNr5TiV
e8XItzq732zPPaxI6Hqdu6KfCrxKnOhsuJI8ed8YtKb0sWLu1Kl3aXIXJTaF0/A3
4tsjjp77pXc7UDgTllMua1gQ68xlWWr4/6G0iOg9kYtCX21OUXTKZlEHwYrUeLPW
xzlrf6xdCupbOF07GXVi/6rGKk/9yiNAMdm3GGuKxEe7mptm9VwHdFpf0YDbiobd
etbJbIpor0cyTHNkWTun/bOm4z3KGJKLKjOlANq77DYKpqM4eg+1LAaxIH/4Fubt
nQMxah55DSzAVl5tyKQjATWc14dbugoPZt4MAXY0I/Vw2uqEkYP4pI3B+G0TKaN9
2ZTb8cmC9X++ExL3BzN+BoX8sbKhD3FkSCotiiKQtalbX+o0WpGzFPqyltsYPE0c
3B+hniuL0guZGY5hTek23T3JTQyoi3cqM1DkIOGMnV471a3Q5AJzoBjEoqpGKz9C
sagHgNvjcRo7aVkGcix0/duEEWs+14fOf2Ekw1NIVS0jlD0aEpvOq2K0J/mubMgz
d4yYkLEbDeoiRO1J5pVT3yDpawsQ5vNyjJBBpK0bzCvgszsIQHb8hqD+UX9yidG8
nw9wRv5lBvZjAffY+tXng60AfqRNYPnnWp63+ZMgqD02Arss/so1LiPLeajOX8Ln
pfxdeK33lAFa+PDMHO8Rk0urr6vZUo0xy220XDfowCBLcvrjdQab3ItW+8oCJDZY
IEXPGqh16XOzHbOQLE54oJBQJEg8PehGKN0guvV/MxPM8cEDIj4eD1vphrX6UwIW
RVR0iM5P6woC5N9Hy54fAC5B3f6U/naJ2vk71l94jNiPaD7WZRx7M56QiBp220fU
4khlrlRkx4rIPeo0VLzjp2v34Lync1GaNV70dp8ZIyd53LsbtifQkehS+AkK6afW
VRXnmoDuz9WFIHTSBnj3uWkv9rC5wxJhqUz1QXZsAZJ90BnweFLo8v/lCddoLgDs
Zd9i5vhYSG1ECkEDrdT84UoYTKmrJiccDWUFSjTaDzMEa1oAfEfPiwfcsBOINVTX
aRIYqsSsORL4c7Loz5nw1R0BcibsnS/kqvev+H1Cseuvztsg1llvR9QyvtVU235N
e/gSueS5Tyfxw9Af+E+7crai8Bga0+OQMz0bX4/ps+cHya3XhBYhOC6WA+RCYOWn
pIH10B+yk+qdB/SnW9cZQ8hsI+nfhpGeoIpNFOr0doHJVA5fe2MYD33Dt3uETPb8
E7/2KuFyvY0eUa68Go4S84vm53atLlYcuP+AytQM+r4LZRinzGZExSkIMK18ajvd
LNwCT6ESa4NBVM7MeZpKzHK5hUtQSlLkjRocg/VK7fqduW6aepWBFX/NczHC+RDR
D7doNXZ4SUUln9Mx4tyoTyJycQxXtPHhMXwiCGG2/cw4AU6FoVeSPgJMomQeiWGg
3qJLmOeRvIMP6MrQfFkga7jW9naw+VSt8y6F8VtdBRiSBWK7W8bPgKdifbgnjUni
g1ud3x5z48OwCUdokwq7QofuYUmW1gp/wadj+EYG8fMUmSa2PU9lD6S/+0ua2xJd
ehnzE2CaouxOUoaImXWXP5lTzEdsyVRfBVYxmaYo81nrAwEQo3d9COscwVlEyElv
5TFCVafDdo1OvAXAIfPKm9xZimyYiFrtcPcfvhQwsG8vS9uAQPxtq1niEUP1+TAH
SFoFfgTP1MkuCz05ZGKdetP7BtRThlp/kqb3E1iR/T2jYFqqxXn5DJYWlr/ZzY4L
+QKwFFcd7KgtBrDoCnJXoxRB3iDnpIyZe/aF2Dl/1vDBBcGRuDq1SgTW7pppZax8
Dc7FEFSLRe+rbRHFyACT3KtJKoY0fKpyfo7XFgZfV79ymyBJG82AQyDhtYeXaPTo
CSj18amRRj6oRR/Gien0XFVBAkSmYbsaTEWAbGYagGDJzu+J0af4lUACP/OeodhR
7Tncv3iw/yINKi8Z6nvGJAOf6ltZknJD4kENTfpW2TDwpb6Vup3lxHmyv9n/WUMn
kF3o0gaLcml3xmvnuc9IqHbq9KsLwxM+NmZXNVPhGVbZuaaLrQQyPHU75dmg5FU9
SpYTazCMRxfHGWOFG9ocjq+VXPUk0AfflZ2uDz7bV2N2i2t6ADV572XPoUdELF69
IkdUuAfk/qCMhhPlBqFR3MHbytgRW/lun15TfVbkA7b2AAoo2HhLO5OqISBflx4b
qcQsl2j+pvrmR0edY/WKybHrIbmzkMLwLJND+LcFmPb7HXZVBSIeexpjJM1pUQRs
/w2yoiW99Rf5I2oImICLoxI9jfcc2NDnWP8k/JY/Y0xXXrzAmajWNcgH+Ij047n1
bnGWxhQkkQ1sIJtzJzNEvw7QFpKklyrNuMOLArud60GoFlc7IUdfupBVSX0SC9Ix
IrNDabRvxewArF8JQUQUmpeynqtrJ7og01ISNOmnra+Van9CynJRCNEuKp4zCl7p
soWli5at7ocUxu3Dn0sv34ltmfhllHRuTgqwPnN3JECBMVxJim7iNi4g9VNXQ802
YGO3Y/+h/hL0z58fWW/YioQNQz0meGg+XwxtxXR3UwIQdYMR/7TbFE+Am5o9yGmh
q+gAcjM+hWhdK4OPricoFIPIoc/u7LfkcNNtPaFk8WR68hMSVMA3IwF77jPUErjK
R3M3Zub3JayXdZyTx9al9yb6r1mdPCwWnQ/DrVwyMn9gYigjsLuVMjYQOPHQ8nZw
+MRRy5Ere/8UGn/yZQB1ZcLoFtXnbXtZdzEDq70OFsl+ZZj5cpkwwG7ev3YSbsP9
eR7v3OGMWkLqjxjK3ZUlEF4DpIJQwKKXM5kfOj3ImYNWX99J5PdZgtdGdUkW3xdy
FQzeGzesxXAzfLhaaFJmMtqBrWOahD44LGr2rnaeIdFcYfxnzbkMJ36kWU1eJ2Gs
At5bcijdX0sje20/w9GTrgQvEXAKkx0hxmrmrRP1pjVdWrLUwWYOun4PmIcYp75s
sjpKojv1DPVzf1rt092m89XreUE/Gt6aBPCPdfJ/JRTeHFnhC+EX9Gn8VxA3jsby
EmMC0ENIyKfu0AA3LidOBfPeEMBDqAJlKeQUQV/HPOtMwAbVBrGLiZRO3gFoqZkW
MD0aOeJCNsMrDCj8ozFNXMfdpKCn8wslhcaOnADxJ905GTajfhbiuzeL8cKgP7rX
/hsb4mDHzUnunlOyDa+9hKT735yTPmvEYP8oSG1FGWTkZwj4S4q+3/ftV6peRJJs
VR5OXGcFYVzDVJzivbTVeNMNKFYRFzGqUo/N4l6GcHFBkMoAtOwxdBjSBKKU4iXR
xY8Rt6Nc6IW25t4xBPVnlVTQki9LzBGUiaf2CG5Ch9iLnYWAI8TgK/GanXlO2TPu
bw77s7M+m+G+unsfHovUUYGNWI7md8WZYT22QXpW2b0HnC/5kQb8jY1AfKNgs/JS
mTTqsEWWC4zeP01Bj/dRFjztN6QkNdMG85bJeVN6PX2lcaK6qb1kbiB4BEAWC5NE
NMCPhdVriv4TSF5FCjl/ux0WoOBVaQSjpMo7reaOB2cfBOvSAEiEY8sn+O/wIVLU
+mZoZsw3uDT3M1lRvHIDwFhuVR5w0/XKpe/KzZ/+svK774qXFfmSH/NfDX9rv9hH
6Mg5FIhxDS8oneaM92Y+T1nc6Q5sOAmM4WGcaSW//XsnZXg2TFUXRpdwMsrhlT+Q
//V5rqQMhgr1ssH6IE3dFe68dL4kComB3fdOjhw7mgqPKpWQipRnu2E1uFE3D6ka
AjjTxlBvlyG2rF3Y2E4kOYzJLaApPmBMzxKHoeyF3gNYxZSrNoiXq8bGkqFKrGa6
mEqZu17AJ92FxA9v/HeExbV71XFwwhfGFBsBzgCPJokkx1E9vrV5zG2/52SxT/Kv
zEDmvBdinXUnTg5TYQa4BWEIYpOykbl3bHs3vxRrhhTGdq5cj58WNZ1by3pah6c+
mK7wYB9Bi6zfevAjL4d2g0wI8vd+/oaKNTa8LLL8ZLb8y268VX4yesDMGNT5tnfK
HGw7oXTS6LTvvqUj94eUj1KrdRJAtnxW+LWUydML/ZSKiY8outEyKNxXU+EFD+xh
YXX9dASZhwmw13dcUqTJkUGiAq02D+acRBSj3ms/iuYXt1liA+v/2Y0Ktho0k1s8
VaZn4aS7UMfYiV4LHk5qykF1xuAu0skZqC2ZxBY8i2T9IJWHT2ekMk0Nc1p7Q6XK
NzV+XywVKAVOB+sULdjAVo+5O6S1qn1v2hTLyBQTk6rfMNHmQ5rNecZyWTF3hLdM
1yprC/KUfAVOrFDXnW+N59PcwBFkS9tdC02gotuforwNx6N3uYBB2EtPfDFkXtyJ
5kw4iGQpEKtxN2UYT8ogaXaCheQnTZcehYCelFMcMkECsxKS9xyZfQ+4ZEciQRnq
3KqNSzGsTS4zLnfAXga+YI64UmDm4blm2DSXYqywhInAIJmilHuz+HwZi5MyJabs
7Vm2fCxVufqItY7ZyyEXw0yovJnfSTrtjy0172lEsd8lkaD7JMmosGyKwJh4fzm9
ftCo3SfDpj+uF16yUVQqzW62m+UjWwrZdkFkSEjR36clSSFPOv2pZwErj1l32BFC
FCIMyHqt12tgq3j567g5oiqBWGyEIkDylx7zqlX5wdOAE+/dljE4EDYTKrtRhiIX
viqPgSA/poetNEqmI3zCLZQu+wFRDMx/jl3xFU4KzTtelxhAKYqah2+tE6z93tIx
0oSuzDjt1HUYUngjUlmYQWDQEHIHnXrWrZI8YK15gS573ZAKaUuvjq7tUHChTBjh
qxYdufZyD43yhJiJJywI0B1v8LKfzC9OxCKGWYUzqa6DrjTKGcFnyo3sMJLwmG7D
UZS7FoGr3e6bleNxobSXgS9V+BpTuTK9saRd2FIy6NwcgJg9tKbLKWdDalyXYQBc
4mI0/Lu1De8FNqBkHKg9XCn76fKAnAsqR25hHqp/nmFd5Z/24bp23z477JGxCLx0
FZ2J8PeqzD2s2y5imY7kMNGlL9oRi18PDAZqboKTb6rxM6Tf9txH40csKVHPESzU
YJt06UGrsW5GjCi/KgBNAgovl3U7uIBo+z4p/6wWwRDFEzanlrtSXkJIEmKXV3g7
F+LsEexsAy8Jbg0rpvuOHceKuJ5i4+V4BPXLPLlHZk2lqToxWqTX0tWUR91b3RTZ
4arCVHr6MiFHGLW6y68X/DZJ+beF6XBrGK0UHxwCDzL6D76rr2ZRfvGX4+twv8Cy
fAK/JDe1t26u0TvvvEfO28IS2WPWSmBujGr2bNBAjTXoWCDygcy6CS6RCWzbQX3X
SEoPIshKXz/67y7kdelYOnjWqV77Kk/2UQyrlaL3rEZWkXMPAheGvR3Dj7fpGFRF
jy2WOKfhcmi+RbiKEWV+dMhXmMoYYxS1xXPI9reOG4ZzR55DPbaeFO0ENid0e4E+
urGH3iStI8Pv9G1+tUXm9dIEo6rPuM9mchBxMVfKdS9J+j9w+36brS7goT8fN073
dYk03sraKZa8ak11TAEwsSkw+Alu+ZLkJ2J42XNqTWM/9tBdbxqEZ3/Rxraho2V6
9bNeHthnnB7PutuH2ddhDdPbDyL+oM3Pc6mcfwj8pRJk4PQ/afsHSjDfgG4ZLaJ6
7eZ6tbiisbtO6lboDExMs+doQVCP7ltI4HZrkAHaeMx7+uoC/YJqnTwKn/8bMOOe
8MAmNfSjXzI7R29pMH5JbosWULqYYySfmRPlw33coXcF+0T4hlvRx+CgBItorBpb
NAcGq98aJOAwD1Srq3UAhTwoidoKMiQYFDyjVnCqQCXTYs6V024vF3ZHwdR3jTsi
vgojxOqMpXfmMsRMHqUvZRVnK54JWK0gtRXg8vaoJF1SKC0paczRzyqUZ01M+Klh
7IKE6bGEafoMBrG1a0mVtDTBWjc0V2fI+fKUuzJ0LFRtAtESTP384CQ77nlTSBgM
7W1NtM2CfR5ezXXgaBqu/cmvOcw5w21pskIgy7EjpCjCpewspkTjoFaL4d9LrhcT
ZAKzVNkZja/JIPICC73n5Mu1ezXiHWaDNtbZaSI26dPqXkn1F/iev0LzxC1B/QVX
K2n2HmYXUbL44DXajN9TpBrF38KYXUUqD3FDtb7uk4P3pKCl3xmrnWnuk5JBtHiq
YoC0OFdWMKDRd1uqdydAxmp+uUM90v5U8hDhxn1rqpeGQAoQdhSOJxFdy9INGnq0
KVdpA2FaLxidloscBIUGyk0KTFc7qCTCZgD8oWiOkNSx70Ya8cq3Ah/Qp3l9TEB4
zfPCqlSycLR+TCInWPC1ZkdcyQeTsXGmx+VzHrMEHZIl+b+5uWtsCG8Vh59HvHFj
OheFhut4tnV7Xfik9iXXql1EdTcT3q+mWUFl0UajJdfugTDkyQ+P8ajjyun63U2f
u3j1NzVkyCEFK592wuc3hEDy1xDQxFYHFKpI9WRoqCecJDEI3zcb/NHGMRSY1Sdt
FmxAHTy7HqkGcB+o32qURBdUohTyn2zhwuCPiUwiGmOZH/W2JIRlyaiStkQq0uJI
7SXaQvZ2+rtEKHK8hbpj1To0ehk7cKF6dCKhqm0SZ4xn9qRv1oKRrAwELzMH2yP8
0lKL8U68eUe2WwwGX8GHdnzlk5W39sd9qLJTj6HOovx+T81vzEEfWHDSoXs0i2ww
5u5P75Yg3TG5h/gAvvFKxd+sIOojKQL93lyhG8gowZOVOgqck/VZjKVZ+A618e/l
oNq7j4w1HiOFrmzo8X5olR+M3r2geoPU/J2c6CYK3UW8SGYUB7+4jVFtgpOYJTcK
shVAKnRU4GJUmCc01cecQPOdbNLQnYwkEqwA41XxfEXJ0EvHyfxo4XU38gAkCUtM
V0cmyThJlMm+ryLKyC+Wa1B5FV2VK+DE32pcBBpqdAoUgJu2IV0fcFjhUkKTjU8c
Mk1QrAS30PaUr1HI6AGHtMm8sGQCgeWhNTYxOLTpzwp0lUqWg49Yajyw9ojQIZme
EEXsOwpr2jwf3xxZ1CTEARmRtS3o+iWwcmv+f4BAd3dfE8RtQ360Dh7SG7g2gPBD
jcuU0Q1eTbrFOpEkuD2fEQf2MdQx2AG6w31lC6iAS13aLNuoLn2TJwqfA7jZrswW
mNqrw6jLFM/fF1PU55SyVnGIj18xxDNByfKlD5aSzAf/fUCPugACpwZtI7nkc6EB
APc/NDFZOIe3oDf/hVZ4fHaZxaPvTsZlRKQikiFOrqo0orqb1InjoF0TwbiSx4NB
vcwRapfxBWzFNYliZUym5ColExeVi3rGaZl3+jLAzzTPQcIMcfLW1Wm4EspPKQ2m
sxXCRR/KhZxhyZ0EpHbK92DAKnTP2imXz9LLm3JzqIG97Wunec2D4SaUIxfr0ul0
UWDorbM2CUPjS8i4+g6KNsO2GJot1377GvLYHw5d6iwM5EryanFF7Pd3tzUBvL3u
jOZXB9Pq+ORPqlzzt6Xkcg+zTDfZaz5fPdTz5ovZRpwwbKE61FAvyOqSlEYPqLW/
fANnmIi3SfYo/Fa0dIS34Hgi1GSE+oDTAp15Am2bbo7NE2BSpm3Ik8SE/7p0y5wU
LkLDfOqFhEESO1/TnnVNUzTlueoW/ltKe3kRP4z1+AEeprQM+zTMRllrIn52KWhO
0HXQg3PczoPMfvJjEsm8OlgoNOkelnCkIRWioSXLtNqW5x8YIbIxXpLGtr6//xuF
2n+VrRjdMNA8PEUm1sM2j+2+quUIgU/z33SpVgk5QGpHhmXHYKLSKoc1rTl9IxPP
rCs7V4AkV7Zr9Hr8ocCzhL+TqBGXMrPlhfrT2U2JhiFW7t2RNbdileb3WjfAETwy
ra+a2TizpKF7zTubfmFnzA0bB1PUHB3LvvzqgkNLpaLHp1gxYjHShq+5wM3ATm4G
UmEtd9rYIPW/f8PKVO8AXAphxzfwH7vTiSOVUghY7Ts70iFWN0v5rKOj+eoLQYuB
LLZwgNERY212I7HVfUItOTWTMK3ReR9s2PT6Bl5XiqCpYH3Q2xbWvC7DOcYc5OT3
F+1Mxi1nDCJ3dY7WqsBcO3dIaMp0WfAnQuURumJ0mV2qmj4PEgOFy9VBhNBfSKTw
4qd6Z0ojImB46sHfqEcT7LpBxQUaDnl/JcICbBNyglcz6e4QqfJL4Rou6Hnsnx7m
bowvVz+/gdenOmOiODLsYeKxVA3JzpBsL2Jn8HbsP2pXF1oHLpPegoltOc5rhGDN
zgWmw6scYxg0d/6KhTtX8qcF5oSTUvlGKS7AZZ5fpebY4SKMy040hwTJySqETl20
xWP23KE5eE3oBbm85DQ40jwFXypMVbSb681OO4fN1UtlPDHWE7ysY+b2fyOkIhpK
+9wcYFLQpMjn+qpG1rnM7Qo/d0gBS+tak4MkZ+NSh1xosy2Y3c72H8uaw9T6y65y
SmupoN4HbxNzxw0PZMpM0kXGAci2I7h1t9bstmlMpOsZ9VE7m0yFW1LDwui3XZzI
ytxLiCpouXxmLKr6612nM4Ncy4EVzxAijL43B6+jvBbXhzrOz5VuiyellHKCkws8
Etf/CRbZXHagqeof1qXcDLvUaJXOTxBKUIuoPSuepOlqnbXRNxsmyNjbrAzP+JCA
OVVW65uyWe80HuuAjhTDQgGDzJiY923koXYET0lqO1Bl+iHWFqtKQMtIahtQjvGv
VT5yK6zYrzVsQLNijeyvyFl90UBRPcU6iyuYHIDiCdQNmBvCCbRRHGTosFHfteGM
Mcj5JJlkneV+F3EW+lFbDedE5XZW9uPynMdkhWEw+dN7lDYtYAiJUHj7Z9ijKTEm
FqMNirOfGt2nJpalf/KpaVRzgcqzntEqRGB7e2UymntQfC4rT3Wu4DpWidOw+TkN
PBOxrrZxj0fuJGdyBMxhiWewn7XWRku9calhAEnq7X9No+DR1HMH64U0zXM9+QRl
6zu7iYbvaI2kdczSaXpeJN2jExRZiZr/9NqYTIzm+9BYIVqvK1Y+n2D/H1XhKq1+
8TYRVvdHhdnFiMsMc8eGNLtl1D+5Tb8d+8oVV7K1Q8cHoG8mkplxj+7wD1pW1wnP
WI0DqFJDwgKzLxAiS+DT15BXjemiBydCv9JREP0wct7pNuYr8ziXrD3CDLpgvQvD
lB9lxbZ2M29MuE5KidPZBdjyTpAv7xOXiOeE2U6XA+lDUNiqG4UdO0hhin4Zs70H
1ocNp306oyANlUza6+NAci7mHHDzxlXnmSgjayV3FIHSxw5XxrCoIjvgGZwE1yHw
RM59ACo2BnaC4+o8Ehp1yG6Hb1QRqMYCLdlmE4o1DCPi9gLEq6DxtCk11RMecTRo
ab6bIfF6Y6FPPbYsIBCj4kGuHvi4l+fkhNJq7ygJuVYkxCfu29R9uLjeSxGkEOGd
WvmXPmau54o5b1vGRTP/dTUS2ky3qDwRaJAjd6o0P9fSnZ5s4v6YYJiqWW4GIchE
L4BBowoxU34GzlURfoE3tsXvDr1Fc7m4X8VFmLgWQlAoriVfKq1+udgd/ARP4CRh
tc4ZW8UzYfCJZOGyGP0MpDsrqjjsd9pqaLJt4QdhFhGfFexNKTFEA24Izz+g/R3b
ZT0fyPVhBYv+oQsyhYR0M2RIEnm1ZHfUJ5LDmRUM6shASLLm9HrrsawJPNs8NM8t
K+W8Hcr/UL/lIVVFiTbq0pilK/dhuv1AaIVrWC7lbqtfSrxc9eeiHbqB+nKi1glq
TxlQrKnpflle9o4qv0SwwZLCSehDsc9R5HX1rjGkfHHKpVTW/leduiu1oJ2ALrNq
3Cct1qFebPn0iFrlGXDEZAr/dAeJNgTlr7BpxhjJZU/HhF1vh14esOv/yY258EuB
OZgS+5CCOnT16rxrHaTTsfGBMLlekk0I6JbpcS8gyMgf0GGGzz8VQxJKUkaGLZL9
Vxy4grO9XyvqCCXj1RIhqiahbMsTd6bM22SiIqqknyrcuL2NcSgNwi2sLkrPQ+0f
wlBOf/n2kjCSgL+ERI9ctg6/xBktty3m0TJJbtI1sxIpeeqXeVk0k/0wEe0z8pBz
HmsiuqmEZn0+ncwhDD878pQj1c9341sts2nJkUmOhjeRl67pamnnQ2BrFHzRCpKC
IGGxONhBXFyo4p8GSmSv6SCMLPrSoktO8TAvnGqZWVvjXouF866IZGIv6LO5ubHC
E52ogtL1hntUUs8BwmkQWa/+9pjVl7CpRUsplYgvU4QA0TIYzTisMu9fcaSoIGVb
NTBe04seUFj80BPjLNPD96vvSiXUyLVkkGMdD1obmahTndM1FNoUI6E7IWPQ1yEA
FW/7c3n/Nf/COeze62erOtHZhheYW8Ap6WlvQXmgguleVcws9MF6UlGqOxN+x+XS
tqMfSBc0Pph4/SxijzXV+9qV9eY4jPbKSL4NX2ndkbqllnMXTtRd8VcQJOhosO4u
nPVXfNfEw2pvxkZlO/v7seE9ZPf9I2Y0uLcyxOxj9Ss7zOjNYSZfeMjbbhuIKp88
BZGfFLfDjhEok5pk2kV4bC39/mI5mrIQHVNDQkU5P/t3DXRrYCpzx7uoKiv2bnfO
CS/gc4xG3FBZM6DG5FlhgG0sE0LZOoXgavbz1cFbPWqvdB6hXwbG79hadZ+jpXS6
PQxoSFCDbnTeNe0C9zLzMDN/eQ0j/DqMM2oIuBvvfZYvF2Zh72dlWKeQQHOLVyYz
OiPSlbFlq98awVpqc0/ZoX/yt8kvAn8BZ8OtmGFasd8GZs/0KLBVtwk5zIuZ484q
LEQfxGMp3aYHw2bGKiO1Hq3eCzUuost50VMWwbTJglN203GUcAksb7FvH84JQ9c+
7nDEtF8zbuDVH0CkmfhXS8ASaKLU6BO5sL/OfAr+F2R/muhuFgcgO6HD4byJIj94
avuk00Na8S7wBngubJRenUubOWe6vCZ1PpwUlH1Yr3CTCL+Avca+MY5zlX/DsCiS
jOKIwRiW7//TKDc/vKwkbrLpUY3WV2xqcHJKhjhqcmHuIrRDQ5AsStzBAS6fufgW
k3TEulnoRwLu0+TzpfomkoGGGrtYJKLhJwzJoaoka854oD0bwFORw0PuNxImgU0/
+MGvOW3ZZaCslJPeAcP+nH8rwmFfn40+pPDz3J1ew99bit4MOP957lvIk6jSA1FK
nEM/5GDmmp6u6wLQSwABDgNVX99PnOQwtUhNXQyX1DBKiIjcKNBq0Y2MRHS/2/dc
KwfEL8itGKElCGMlpIXcmxAaojkD6H3Gim7oa80DnhMYuNFlKShiOGm0F2J4GQcu
ze8WFhuYqYnZOVI4QJEwSAKIy8Q5X/Qz0sMeDAoAqlwmo2QDK7pT+cldpr0NeQNm
/0GvpHGARuJJg1JQJMLTkr2LsT4qQkiKGgMusdhtiuSDLyUJCb2TEn8nqg3yr49Z
ym+YiO8WnPfFN7g50qUnJ8hCWKKk9D3zRLCZH9lb6fp5ce7qZ/c9XlP3PffP/EIN
Gvsxrj2Axm1NfEYpbIMzPHCvAvrBphRaanJu5IcKMahj8NLrwwTcP/moBtAFrTxc
SyGvs9jvbhnb/OrSkjyn8IiCOFNLWfTMAWK28Xk07Y4ez2wgAFBq22KXw475wcuJ
12lt/EPBJCr1Zb//R+dToKHSXguyyQWdrbe7j9ErpXLQquSMIxWcenrpXf/FVa77
vOP+Af2QCQTxMw4IwMctgcyzD59szQFD8OhHS1580RvftB0vFACgZa/r3Aqw2rX4
UdbQ3v70iaAi9ps0PKibboK4a/+iExC1rjxo2/R2Oc0k6ojK5iGVyP7FeHXoxb3M
KbCCU08XHEfSsyRiu/4jjeNxYf01DAnETfHxxOzrtMCCMT6Nccs4AtMJLJGJrHuM
KwyqcjY3PF9OVBObLffkmC5pFsOENi1Sv2A9KJzKJbVI/MfYermKu5IKm97/t+P0
YQWH4/RPy8Yqhe944KWhbLwbFrQK8WysPMLmg2z4GkBMW4DtjHCcwOdjBS+16te2
Xo2mEtElZQFyFQlNj5ve9wmDc53OzwRgX2aedyXQ8PwdEsxCgX10YHRiucpQVAyD
StRkqsvK3V1/SGfnas7RXpSlc6u70U9gZBV+YbbhtOeAWO0BKV7jcAK+8O0YOkNT
FGDUMYpO7kxwlJnOdnu7d1X4x74KGo/0XZDRDRW4b9Kxf925B9rjYMq2s0Qw4JZm
kBBIvr9Gwr3IaSMuetazkNM83kkn4kSKXaTpJcrcb9nbHZ3w/Lv/lqAbzFvkrMFQ
/JhuLW3YmWB6WssrLo7ZkAs+OfYrgz0u2ttXgswEPnyRwOUAiHDVDaxQllZlkMXT
72iUHkxs5dVHKFBM6WA1s61cTFff9dr+sSyqAcLEnvxnisLf8Ds3wBN1FW1mXQN8
VmVBN0kBQsBG+vFYO/0CFhxp0l5jHjk/t08jC6O/C3QxGZdO0UpCGCcfPIXhNE+G
7fR+SP57by/Ff4Xom1NMSSYWMtYVkKSo1h7/HnfPw8IuAvaDC0NowPLRz+QCPewR
YkRxfEr7O2NxQRCX5UQ9etg/UMFzEN3CzweW8CuEiI08lHZ/mCTeSYKG12lstwu4
vKP58lR+pS3mrNkDGQWR+7CBtCOxDbmgbSS7iLDCX9nqci5zBeI73PLFjwXFjS3X
fDIsNlIlCaDPyjWOSx6tk1TarjXqZhDlkK2nHvbHaEX7g6iMViVOIomBhD6ynI9V
qNuEzdpAkDtXT5ybNSqO8OwhKhnjOxYG9KD+v6uD0/hW6E5FCUeuTYwwqedIj2VQ
rGVPYICFC+P+o328Xo66Hq6bIINgQSfviUNL2E4KS7bdeZdbG5tWl46M+pK/FkPH
toPcUyWZMEGKbklEMIfCFG3kH8ZoZna2/NxRQFWQA50r9ZRk4plwe3XcEuJVeyiy
QRmRL/YwP9QqliGB8mZttCnB01KVbpqbU31qjOX8/9W/gweaptMvw3UUwtDRyP25
5Zq8QGbiS554u/Ir8VyrACpBLvstAcb1QnVnHhqNmKcbxtIbBvmxBqfsi6kZt/uL
Ciy1/bsHXhUsCPo52QJ7PyyEmnULjZYV8IVO4QPJTiOzH6ORM8tD/cN7r5DAhbyf
rhz+/EqokoSkgNfS0yjH2BZmojv6m8P3+jYYIYrfpRpCYGPS/MOI41gXEpQTwMEk
XrNtgIN83fBVEVMuhYMMK+AZuc+zdOhTaiyCCl/TmhXsiAOOdxEsSG3S7GjApKM3
sNfKlE0dHBdIbvl0UBB8dY9rPIsGCkiubSCTJ/L3wrM5opPZRIUgoQiPsh5Gkx4r
v79THbKcSVppEYS2qyQ5/0R6LOBhg7bcUUT9/qQFbyDv2yzuUf10dRLJD6DzTOo5
WNUpzXzR71/NIwxG/HKC6wFdxqrLEHWkwnmyk1IXqcSEmQd/rTkAZ322eRaKlmsg
Od/Zz0sJ28vPCaOtfV6+xsFtZJIyhSNVl8AU/cD9Hvn/F9711Rd6UZ47+DCXuud8
G83y324L7elY0m5fy4bZetj1OuwEZBRyLA49ugyylmUtQ9ShTnIUM9RBptpOqWtF
OOOlu8QPPZf/0C5FiF7Afn18F4q9zevoNDw0RRy3Sq0ITpO3bmPXyL/gRK3lnoZm
4cCJle6QiYcO/s/a6FPUCtYPumBg7j1jA83qXEUJi9iQXPvhN52pAyZKfR33LQhU
itGoe93VVXDF4A6kY/mUmaZlDzDD/nY8stDJ/fihNlg+kPctBj9onDfw/MSM3lJm
V4v2UHCBs1MnrdCJkm6J1/4oKIF4MQmb3szWBbrrtYTkfMI/q0FvtE4PRqZ92rsI
fhlPV0AgJGIisYQD1oAOfl2FaR59dPQtFBUtVfxlAYeY+nI2nOQAWyrveyfeBxpU
BVjIFU6x0kSXVnEdAdAHEZlKbiuiMcoJdClY5+mMy2wZNf1Ya320dKunoLFFwkl6
48plHnsf9usT7/etirTawE8eaFsSKibyweCxwmlJS2Jp1W9cEsnBEd09A5TMsBAO
0O576aIJZ3ODnqlSL3pzyaTSt8MxPt9KHCPbocXk41Y6udLNMnO7PsoqZl5/YqTg
EcYXX9JPUk5ohBAVHZQ+BcyE+HdJwzPe15mkky1j+WiRoqrR5ViZ9yS6CobnjDQg
U2qNOJ6xbm06ZDPOjj8xrbtC4+GM+K5sqyCcHtM/kkrpUo1H8GzwAaJ8Df8BVVzQ
FkqLQyRDgsD+L5aZZjVyQmIHUAMWRZsRyV7PvuHwRArJ9EtpuCYoSZMfMVS2/06+
ardZ7sD7i5j0HCwF+ZIkpCNSA/lxrSV8+I6Vp/6DLbwqAQeb6OFL/ehRz2BrXzDW
TjGAUJA2vYppPTEpjkMGY5EIzUkLJFW4HWV9LQFjsVfM1rvCN8c0SVzvu802WEFC
FORJqAC4uL9F8wsMtDkCUCQn6CYQtwZYv5A6Znd9K+uuEIdD+7lv7FUmK1EPlxH3
zxPWEKHhFUqMJnYZcnRysnyg+86MJ0cozTbeRLxbjmbwrJ6Cli3u6eplBBMfsxb9
+p72I1aD3i1+VmI8HxNLbMQLVT75DPImQ6c55iGwq9/RsYvq4xkqaQzWyNKocRRr
4e+S13CK/VfGg/fWSSFjOoNhM0AcvnlTh+Svlerdxg3uOrheVA9yhrB6WzGlopUV
lzxh9jgqob/8m+lb1rH2ifsaJNzVBZ5QvWiE5IMU2OLeaP7n3ENgf9kIomYfyxEk
6Uu4us9a0gE1l0QvRitiyyqmhATtcKbG6eDx8k/xckXaUn5dKzP9HAz+Ba3MZmfH
RWnP49yn1XmmNArmFf1AXT+m3pOPjgEXkMElYVF2x/L0p1wchwwC75wZljOjWhjj
gquUPd51eVt+5A/fSy9S/M7x58isuQmABvHKpjgdRUkshBLkXrM4ew4ebSPb+i8U
UGJQsVxdoOXyf0TwaS/sl9WHKUr5Yl/X1nLTthU93KoMHLts33RL4xtym39dOaQJ
YIEEpEzZEwxDIo4g02Lkq0LZHU/7cZrpqWk96Hs5taPLbWAWAOY/jHTL2qmMoVuw
XiBpQ4fmrOVIRn7YhiNxu+7pgm9Nwf4tYNT1kv/zWmGTOu+l1vgj36WvPk02Pelq
VIgXCIkt6gLS3ZHib7Y8ayuTGDQM2hkfihy7T8W8vnro9q1KVu/NOLlXbQm2FPLK
Hj0IRJT0thbSdR6YqA+8AuV3Pi0oY0kdBOzlCObloXNNP2VWwF51yoKdyoUvaBPT
NruKqzqqiKpEtwvg8JGb2IcAKdtajFkGikr/FndXK7Zxygr2Gj0HSS3qBtgt8RFi
gjM0EatrdLUV/fTsxYsRPBo2s2CVu8w2fuQgpbG4MPFZYZAgWB1seFDqzQV3cCsd
DaE8SX7K8hD6w3q5Wv8Kgg9IIQomKKeWv0K4o9dSB/y47Ifj9RiJaBZYg94G5pM7
dfI6gZKE9U8EklwC1vbsegvnd3DPtA/r3AY0p7n/gm4KfJJ528HK/rDU667wvalU
pDxrC3fz1D42/1KZnwjxgFksSD3zCl6RGHvoDI1aL+JaVE7vPiJ0/W+97+g8XXMs
Xv6IQZix9WLLvDNFUhdIJV3zpcROpbWbw1LVZzRYv2BB5q7XEMe5Hp1L2yTDPb+d
C7peVfqIPzC1eq2AkzfDeglEidbs7tw2sYISEaU/FutecxVWRrwra4voQFHDNxcT
OacsqLC2ma0rV0Gnvb7SBhmkrCK0I121ep6eHOIT4jRgRx5VaiVKz3bexNpvm0zr
owkoqtSZzY6SnmpJcXdHgWJbglcYjgi+Mj+whMbxiwgOCiIcD+ujPNKmMV1dh31G
pxpWXDhWKha9yQiqLOxCcUNGFhcDzaw5dp08BXY/hbMSrZIg50KNWmQma1vHqzL5
ErUPTAZW2Ts1iBw0gzd/3/WNW0H10D3Q/JHTkoBdAfunIzMqErXd6vJcr1gNBZzC
V2relYghpgCr7ERuJp5OIS8EcgJcWldLK5WBTI6S0HfD0vgMfvAAJSz/yh+p0Sok
s3kIXMjJbji1CNIFP9F9r0lm8OwDGyy+GeKZDl0P+fRM/0tOUj8gIoP7LmWai9mH
X8KdxaYcRS2+4wNsC8fzkwVnOs+XVmzZf59Apn6tvXurBI/P/J9UActJInFF3OXj
WDB4O+ypwvdDbm1AcYEJGmscoj1pipK3/pVzR2vFNEEoK0rHPNHU7dpHg9wOQJaZ
AcP4uugzDmieYP9IKlWVYXkCmX3oWT5M5boG6yCQQqXlCoIju+OTYpIiqgnNP4S3
+1w6DaOnnzofuf5nlQ8AGvBOvv9pGavrgKNuitEGGQYzmbYcP9/zVeXTzzrnJJ4k
HFipK0nZc+kwQmPWRKqrDOC6XxH0Jq74iPnLWfLVmRUSabAlveqF/awZMI1bhoix
wGL40HJIs3fOfDUvSHKxNt8b73qOdIIe2MsYkE19TU2KHgBELSw12flneklyt7tt
yg4oYXBpRzZh3FKib8tAw77KL5JFFkJvdPM/ytnzPc4PoBBgXIMHJugXSyEdCutJ
TC4ZWhKNFa3xZBpJrAX/LXk1RaQ7G7qunl6JLDV5gErLnA0TUdAMACKBaDbJ4Fup
VxFC++qO1u0lKEbvlX8lGLS6wQnde8YhmjzOv8MSjVt5r7Pi0Pg1GNSbr0Heo+Sr
ygCwWFHCK1wgKLFYHgnC9T46AjPK3KAQ5lkMEtt+SzgPWS73EZh532qQn3P49HJA
7+oRBnNSpjOdYI1E+YcxshoZXo3xgWtopMD1LiyDxJuXsgTplF57eJAmXbbzwyo8
2zlXCuMl1+JLJzWYmg8VPA5tilR4owpqkqYE4+MYH1NPPBDZ5bVdw7b76xBgCVfL
3XXWGa/B95x5sfBR8qaCR58lKoJiXB2XW8BlxqwXTRkK4UOH/WPaq5SfNss7oGtH
UoCvZ/9P9X8svFN64q9tffb16uSjzgj3Pl86Ibj7P6gif/AWjC3/X5kl2du2YAHc
/rAfKt3F+uPhAjHiC3slA/NU7YPrxWzY3iPwY18kRSoXfXlguLcXk6KK/NJEggqG
tZUCZuCt5b/o4YXhLxMjctrLRxy4FYY3Od8Qhm/Lh8aZGWgEnsU/ZBJeqPv0G4NH
EpAK3k5wET82Ib0yv7QF8QQVjeHQAkKqmUyVwzRnETCI5Z86dih12DrvJvN46m+u
KQTrqonocWhHFYin+P0j4zdRsAwAhq6zURrT1VpEHk6PfJL/MsvEnreqTNMLmkYi
YcMlnKBAy3tyPIlkBoYeEcAQzzXjDAZUXNm0g9nCGjkU2sxk+bjzVj3l0lMIWNA8
YdabIcs9E1yYoWmV3fp7DqeYBHzofpKvHzacVCNvSMT66U1YOPM+pxjRLa1sbq5C
UKHTqmQ6PvPWImux5gs1TnM18207lbAOJErKyYwQcwcJkvnqubs9ncXPNXOK9jOL
9l6kCzxxl+RIqMTScQ0WgmA9FxqBBq0O3qITnZvJVfzyES5/BvUihnIF7Ti8rbi0
W2j5W8lywF9jtC7XnAUafmtFZ72N48wvpPXM/dpnFSULx+t8D6UgIR4J8SUwtbTz
J3FP8GG2hU5Wvqz0wmZ4r+ZQHr4ImlJJAhX5j4nREhy+3nMjTl6m/mgHemi5mB4x
ORx0Q1murXZes5thQBu33Y8PdlqIDooUBOIImQ9nTNR/ziAhtLdeNOV5FEbWF+UC
OIqkDoGrg2GpwM5XfoP9gxFaseERDNaZgDnHtgD5sZ7iPNyTWOnp5jJgsC7Im9vJ
l49E+GnUfAJSxW1dtl9kN3wJTrTXVeL+46nrn7GGzije8j7eGDjLErSxxz3GEUv6
N3l+vEgNXIdTors+GHPu77lk9alIyJaOxkLGKpNwdn44D9V3Rkcc4IW3eTLSHXEr
fw3w6UOX9KwhiYMPYWfTv0JqStiYw9WlEwkuoHxLY6DcYtaZhR7n+uuVvfmw0cgU
ET72fF7B0ltemm/k1JbwzLPgxFgz217wGBVETicTZLTm471sAopZE6DT4Lklhd4b
WgRJIedCsMURpEs3+eaVZ7PW+PZv/EWnJwzeJix5LLH0WonUTVZJSshc2v8yVETC
rvSs+C5ebviX+fxChsf7EuhoayvimQWmfBf4/RSmy26eFB46Evrg17LczDAXFI7x
J2CgOxDcc2Tp8//Jk5YA/E9ets5zgty1pNemaV5Houef9wQ2WEYW+cBefVAtbCfZ
OfFTSIzZO1c6mcbWV2Py17TKabq/2fH5JisS1SUcP6RYOPmtmcXNqcGIYhsHNvav
cavw5g1mjBFjVB/oDQVO3NRaQWiJv49mU1PQQ4+ecEkua0cDKuZSNONoNCAeXaF6
YfHkc61taMP0Z/vn8d/q5OqB+Fo5R0+7EkrJM9kGlVHwx2k2UvkhVK/ygsf3pa/y
brKWjtGjkCUcCK9NCXvj8P0Okg6UphsyZ/CGM6ppbj0o+9mrMDKqstlpOphW2NMN
nVJH97D8//W100gI+T8RefZCrTZWU9O8j5c6/plShztSHaHHi2JIZEJ3MFcSS4WL
KL6BKN7jMU5f87xpI50NA5aCHiC+qeYWaoIc19f54w/u1dpQdx9PVu5N4wMxkIEA
1Llcaat6xnAQNiNvGS/KyK5SKPQZL//SM3XgA6QN2Z9fQlO99ugo+kq6uWJbejDO
5akbU7rrjbeaOk35bZUo/YGkDar5d2UJ66pz/Joz3Z5O1ydqPeOTAWpR7+gGK+9l
1xdlvNJfYsYsIgLAnR4+ENJygI6BYFcCDgXvr0995CFooN5iGLgQ4ngR1atkjQ9F
Lls/FFmCFRbQ53txpDL5p4pTl/+nlY3tT3m/g0SzgOvJ17zd9v4la176Gh1RiiJf
9tVB7znSGKm7ekWEZ9UdG99s2VgTh0FiqjzAGjIWvQYB1Nejxb9jz2Xs6plGBtvC
9p6e0/s/SvDjqrllDg4DDEvtqdn+Q1ZqNiAsJoziI9W50GM3lUTq129Q1xVntl8C
34d3TULUWQg8XDnSW2+3qne4GEZGFJwk8IcI5bdCs7m/zN4mgIsx2+ATfnUwiCz2
HmAo7FbERfIM3vHe6iIT28CrU3tYcdXI1YEsdq56LIXGBCle0udd4DP/O5GqDgk1
hvwGfD9a+84F65vqd1BGl6Srj6CxRwjLf6hM3k6fv/e30P672syNZdbayWnWMqHM
PPeLHMiib1V3Bsna/yWV6++d/bXdPM2BCuC6XSlISEumLEtWpXI4XKqpBU1CYVbT
NN8WwOlNlt47fdHfqPqeHROPTwoNHC0Yu+Yq4fLSEkRut5T/Gmak6NYn8QhnocrF
WnrB/+Oim8ybP7nV/1F5M3+0Pm0dyHPXbH0/zHz9Sf2rYTtIJJxR8XaXJpvfDIt0
fF4ScH1BgzIUEiWSt87lZecVmdY6JTD43JgAtsBXXC0u1nLlJTAg9JrYQ3rUnq8F
32CxXOoxoGwdQdjeYVCUTsjrUJ9WYFp3byp9W9wWPO0e79mDIs4hL0HWHd+O5zVt
ikCnUAF93KRKu6f9O9zEMxhkm+Kb5Viq5cXZIfraGJgi5Eskr/VeIGEFMeQOOo5t
DX/lWth3wOYYDA4v9ta9wf9Fl127ucDiU2BJBr3QF+PMQH67SgRi992qTymLBr0I
ImeC96Fwvsc+z99FACVJrEaZuAS3fPpD1R+OGJU3oU7TCyeN/EPT86PQ+YUFlqfo
nGSumCZIylac5AZMd9Y3wSGmJCkDNR9+MOsddTlgdM+Lv/yR3GKW33sZ4uKk3TQr
vZC2rqL+xRgGEs22JGnQkqctSeM2dple13JzuQDlY5WEZI1K2SZ8XHaUmLij7aE5
rw6IEXxsz5Wa9T7WOIfdBqsHvhUX8Ig41gildT34D5VlHpL9udc+KDPbYmgXA0mv
ugqCYtc44CVNDfphV0mERq3hHUKxhAsfdjlHiViP4+3UH589m9GHgxnKUCDsRJ22
0SNxruUrzrN07w2KuOSZBMi6Jo4rlC3boylxo48x0cV1yBaB3Nh3fv2P+ml70oFU
UPJSyOhhlJDhbRuR8akm0jCeLJFBl4bakpxBM4RwoU31vMCOjsnPJbrmy36UQ5sC
1dBwr+TTnvjHr6lMxCaH0K7wbtRuuIudkhAPSESEU53Kbcksgffcvyo78tGaE6h0
cFt6DBG309yDSWLNKBVA8hfA3qjZ0C94nLaTo3kXnYHlqFBKsXIcE8eaIXP31zuG
8HpKj1T8Yw01U2SN+VhEYgOVKybXDT6/CSjOgJUXIuoN5WWzB2/wl0jx/APOXnnX
et7tCLitlOJmkWtLcvEkuLIF3TXLEfyBfDxppKRsTJ1pC1kzT2FAiCAFDwDjyyto
ApTwLSO0o20nnOeX0fboWNlylMx4ZG9ZhzMPEX3GRBV5DdJft2ZzNmPs4zfBB61K
FTiux0k4IJ9/YJH0j7dHdOKm7MVN5EPvJ8RKvYtwxJrD+Qqk3qc9r3XFajWRGeNz
7B2dwnuWDbS+vVTMlh1YiNMTP44oW1qqel32w7bQk5eHQvgLN+JgPn145FWNwOTL
AQTjPXY8ZDjt6c3dU2zxYCfhQhzNZh5vtMVhaKnjOOqLk5L2sqwvRHbLzJpKSXwF
rV6HCh4vJbNxCnCbRr6dh77Fpnd3rPQOa9I0y752nFMR6aGKEX/dgVJ7lDjSjkZ0
CjqmTL2fLRdhzndZe0En2NMNd8y+8kA5zI4o5QeQQLnB2QpOASXrcvzbGgHj/st4
75F0fXsXIqxr7sCwqP6xfhj47kLhnj1IdV5y2hpVLd4KscH9FfWo2SIYOAFFYm/s
d/iZYpzlGNFcBLWmFRrqHB6hn48PvHpbivio2mxexsF6oDa79eGrCi09i+m9rMUx
rMRSjfrusMHK4uiRqrf2LJfypsfAXwY4XRsG9q9/mO2bSOVvoccNEUPWKZDoXOsW
VTA+lb6xzpfFU2iQOm5+arN4tg71hMEEjI1doU80zNkKFndbqeK53Nqas7cOgd9G
PHTLhYFm5fz5sq5jEQ72sqJo4+05YJOXEo3GJnep4qqbamgHXZY0WIkmyYbn1aVT
VdfUjFvclQV7VsCWxIKtCy4fONz3js182XXssy/EW69b45i2jbIc8c6Q0HkryCbu
pXYwCRgs8b6vbxcACWsye6ohRLNnnAjs+eoYs53CDbeWQi/jLryq0QCTg8+Jo615
HfcU7vwY4coiPjeQj1/3eZ2H7pSTZt6Ccn8LB1R+aCSiF9kWHOjbRvB/wUMMMFlh
ei0AQvOucBI25tQL6SH2rgZUD39DgJKR90tb4WHZXoAdZG3SE8ejQIV6xj8wGYsJ
4H/qL3XrpCHqgAV7oHRbmhxwZX3Gt7L3JAoeoFcN9iQc+sFfwjfGshgRn0AYqWX5
5auIuJEbZC6YD7bpUNReTRt0T12YiM9xAm8eDtBVFrbbbL1kBH7tCyuZ+k0lstdT
x1EnI669B6BBADILhDGmEA77hlO8IEA8pLCqifxxd/oEGT15YGR2k8ObvHuHAI1n
9cP5NDrtdlG2y9pFtVPCvL1EK59vM4lB5h5MQbJFvq+G3r0jXmgMxEaMQOiBOPF4
lnbz4eQK4oxO/juITFrStliB7JLhFamv3weNLx60DdgTC6U8SE86shOvsyz3OO10
x8JmLeK+sHYXD96Sad7mgGORi6A6ZD5yDNApSPQFwmC9Xxozeqf0Yf7PcwZDAoDv
NJN5I8rl6Wz6qzTS1QkjSnT6KckW4MlGMSfdIPyTIxotYNOERXNwz8NfXB5Nfqke
WXoH+Sed1wShFmAIwkgPYslSgwSZ4Lb8YdLAtdz7cknb9feesTZnSC9YFop+e6Vk
NGRFtwymLoscGDKZQNm1DBTCH24N0S7/iL8e3m/XaZWdxm4r7DOc9nfm7eLzKCuJ
cexIRTUkk1tMy8FbH7zo3IoO7Hf0CUHpxhYBerFl4EcgpTit3wTSgF+giYqowtxe
1FD0UNR9SvtC6CZnBSkd8eeApG7xdqmTOsUHxQY/IbSIoeQ3+1ef6vjjC9i+Ha+f
RDAcWJ9n1dM9puwp7TzpcObPZRGj0v9l0p78wZU3eM8jSILfzEN7ttXqzMMBlQDl
Ic4z3rORhh68xGApyYWQ12u8TALuFxwdQ3gsO8JYmjbmdegDxN/4AiJZIyFiuREs
nXagsouNKBMsFK+db0eLzqwG5/kyx8cInr4Z1mFf065wmd+S7cuy3BVByh/5Schr
xhvUQCZHUHch4qBtRHaakLvA5Nv7nQCDMCpBp+JGMEv62bsrGdTAngi7XeKmoY28
mfdLPgdDbyRi+FgNi56SIHQR5h9Eye1BlfYa8YpeUcF9XTSBCA+xaQLwIAvfhuxg
7XknT409EbX64o3EiOU3GOVHsQ4xIOrwr2tq+w45ztsZnGFDzTzIiIz9qAwA1vwR
MlCApwAqFp/KxZZZ8wZnMqAHUnD+NAcb6tSgntDWwtwMVtelCoopI9UpTDOIbjXv
6h3tJuxvYcJ14tYOm6IvyIK1xAwenFjkc/AxszjlmSlv4EV+xhe/lq0h09jzhtAo
kVYuvludsBBngiKR1V9q5Z2GtB2/+sHr6DLcmTZUfQ3P34BZ916wuUB190xIP6jq
1X+BUmjri/L42tdCJ2hFK3yt4YjjB8LACVwoLF74dhUCbbwXY75WzPgnymEWOOM8
p+lVbi003OSVepoCwHDWYpfT1S5Fg5XlsfcdpSE9JNpSMbjzoAnbJfxf+t+6vcCD
DqGDRlPHLWxTPtbZbjzIA8iDp2S/FrhyUO9ullc4zl2GwnNbxuaDOTT7aq0LO8sg
iOrUG7nZoVa7v/VGfE2JOnlfLmWaxoxMESjbZvp2RzF9f6F/RnswHWXm3UGTSdjt
FoxUEmKfCOhU8i7bCxfg+bO3hcgTJplyBHTPhMYi/H3dlS0nJBb+oAIOBvAUUsoS
ssexMauoasI/5cDL6CUQ8w4ydEopQnDEi/ZAU5DKkeEEiymg4Z61D69gvW1ytYUw
DczUFuAphqXBHOep+OavDGn4Wtx9ik7//3aKJtoCObLatHZqegO+JnZM2mw55PYh
xWgGYkJzyPuzUCZunuaT9FulbofwGUhZ0cCB/iYjLJrJKhExAphN1MYnVoQt/AO3
Jqx42C8xU7ENxx6H0SadmHcNTTYOB04lVkPkrnbOdYCcu+KVzZLfUrHsWy4N6ROu
l/+mmd+wT8YOercxhYbsteSvLfwgdia8uzRN0SQUWPEtJGU1SQaCJCY+NXSlorU7
kDZ6KrAjvgxwM5A4lfLCJ9NK9eccqty10TvZz36avK0rA51z5PvIdlyyJSYtJZIx
4WPFnyIVDwa/IFJn6hXTNqsKXPWURmWU+Ea9WE1FSaRIkU+mN/kVqTsU55SwUzhH
sacM5CJomhrsTWRfMbDuCBdvTZjXz8I0zme6Jz9cyoMClTISTyPHkVw3GBaWhvCb
yI57ZpAKbn8mL6Ach+f/nD+ZJX+buHZjQy6bgS8Mm3S8BgkPBiO7p6XZmVeQLQ8W
zsLTNHJq/YHF5uvq45ToAiv3/gSene94TuTtta3caztPfMyDbZDbo5UGPhSE7Zy+
rbqoxxoi3y1g+1P/6Qd5zk7b9mdLFcmIZkVxdq3rXIPLFnaKpMCYj8aYFeE3N7vl
uU8ToQl0QTOSrl/WjzNb/caBtRBjiPf6BZJN3OH6Y2NT7kRwPURK5kBRIavZjYgv
VHL+HNoIaCFgSvJqxioPpTjaQNE0baoatqkQEhefjSXV+jFdYu18hRIhSws9YJgN
lAED4uu4jTwhDHRRwLmfVlBmuT15sDmSr+oyqfYHKKI2UV4WUV5SiHKhmwwF523u
Qv5v1NGKL7QNoTuM2XILvwrRYFm7D62UwNDUXyIoZtJjnx9yeKQw7E7JQqlX6m9O
niHqHGA7c5OU8WRvJYrPZSma68pR6oKehBGyEHpw64+yCBOMTT5QrIW7aD+f6rAM
y7zESs5H8GDIAUMC7ZUAr/e4jRRaI9l9VarLQ7VP2x8JqTeuUHuiREdAom/TQgd2
U2+ocao3uqXikSy9oYkfAiYd8dzvS0tZRYRAm7IlZc+UxoXKyiByVTg1tK6TAGlx
CaJ9mNMdMtNVomc+Qiy9s5PpkpIVud1+tDH3Uj40j8L6+bM3JT5B0gU7aW1ik1cL
h2I3d5zBtawFvh7EkQSdtOGyb+8QPsTnGWTAcR+bvog5NCB1Q/uLmsSl0myKx+mD
Sual3XtZIRT+JaClO9uZNIufjDbAeoSjrAD59jqUnexiPZos1rFwOY64x26zcH/l
EeZXDGfDkghdX7SaXtRpMPoeoXhVN3FmmeyHihRVzVZxIVPqvw5QRT3+3bGbU8Xp
f4PAEwkVHVpz5iBsObmnDlNylKG8ia3OdC3MGr45smKKARZ8aL9n9J3BsoYG4VIr
40kf1W/QKh9JAGFTlIgfnMuOxhlWriAP0h9mPihL8oVHxRmkulC7Okttn/VK5ay8
U/0pRRXSiMItumKN+5CdHes7hhqRB5dGm0sB4r++V2CntoqdSYak3kUiqMzp+FQ7
XMfC22RP5MzD3iIWyQCiSZWCcYY/vQjjcbS0WD8q1VjAxjtaoNU5JrLTFAOdr6ah
qdwPS/JDgBtZ5agv2HxZML+Zj9gfGzi0UYg1W5q2fVNUiw3QZ67GNRX3jZ4v4TcJ
HwyeH2lk84Ku2u31rUjIIWcqm1a7RykNz+Au9gK3X3k4WaIaNZ6OrYXl/SB3cSCa
RaV3hIDYkknPxAQ3xtebGHYXz0whj4XaSkxlWydFAu017mO1I2dStTQi5FY6U/4i
wvvJc+M3N0cOgFLaxVKfYX+ZyZbxRmknUowgWYXxSXb5hqrk+fhdUF3QwWbXBfVO
rcF4XCsGj6rDWmqAzXKSPAnQnrdLDKnS+LQJciQOaf0=
`protect end_protected