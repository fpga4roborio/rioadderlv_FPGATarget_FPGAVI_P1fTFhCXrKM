`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
ddtXksX2+yylW5zu6QL2Lhnb2d1sD00763mmSITNX595NcHTEkwn0zB1Dry37fOW
FufOhVzEJp80NC5qZ/+F0Vk7Ik02dIR0elf3clrjeJRK85K4e3Hoo4xn7YbFUIms
l/8VZSb14+JVGURjfswrIyCUotIzlzVYZ6gzoZwDXIi5gQIBf/gI+KxNXPaKV+PQ
Ufys/12rjO6aI/pPlqSm0hCvftmBcnezN2hk1UeXgOIuKZnogjOsf0iJVX2aOOWE
6pD/psybjbnsNB6kH5uFTA5frkzIzkzl5d9+YDm9OyC+k84E83I/7/j+rk4L2dah
QJOvksSIzN867/4Qt8qYTQ==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="MvBXkzurAa5VTw+1JJ70nePUfoQXBvZOku/SMmg4TwQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
oRtzZL4VJ4iwysPsC8SXYCzXS8Fw2gtZTOskLcDV+1B9Nzn1zTyNtlo6lNICRmmK
ZRVu2BmCc2G+fmzynYlNTnSa7C0Cuel6FYpxCBlOuk3OF2tzAmLAuDyOH3Z1Yjzk
a0aHuoCdIRKv7BrZCdALt03JeUmXKPdOmIlkVGFl8yw=
`protect rights_digest_method = "sha256"
`protect end_toolblock="Jn9CQpRhJt4rnzZPRk+dOpzAubz7omckX1MrFd4p81o="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 24064 )
`protect data_block
gD6l00tciPUa6pDNTk/+t0OO0nC/UTtBwLB41d4inuAUA3i/ALrNyoJVcBnAmEQW
ptbcNp5fxEUJjnOxnedyZEuEBxWRieZFQnkRdF269oMMtEnxiUgqgoYfZI3dOVHz
jRzosq4mkO2ywXtp3CV6gIZA/O+xtnqoO0vm9uiXQIGfaNnL33o5flaDMiKFIcU3
qBDrTJipME4W1gyrbbkbXOEUzMJ3pD5A/6cdZzoaFXrBaaha9tmM3CpTBMnoWDdo
dDIRVQKjuPe5cQySo0XpsRZT/jf65PHoyLMSNIAEXSHdAkqwj/Nyw6OSXvNPbbYR
kHwYRiqZ84K0Nju51auScEJ49SHQ24r8O8dOP/KPI9/5+NRWSoC4/fo2Kaq5Ajmr
xKXmpjVPGMHwWrm4oYi7a6ESdCQxS8nIUQErdOS5PC9t+pb95wwdsm9qSylmTuXR
355lX9ZM4hlIdg03f1ae9+uMdM929LHyvimKGqJmsn7c5UrBPxZ7p5hxHGM+1uYJ
cqpPsY1aTcrlWHc6+lQOCzlIggqAfi0KLMr32CuVj/4VQagqVS9Gs7EY5l9kkSIf
rVg/bfWABebFZJVoi7JAOTDdNg4oQdruvvtRR7DvjntsVp/0xCoTTajap3fod6Cf
0SBQ2HC+S12aEl6ASvXOHzSyX3hnkdTr+Giy7hozQ/XRoukIr7JeWjutHxMZ54d9
ft77Hj8pFbhQBWGtfFPaRANjH0MQJD5FpQUl2ubgVceWPDorFPwheUn9Iq1bDcKp
DVmb9ju5ZJ2Ikbv6sFELEaqxirb4ezo4RKHjPfI4mYjqW6PowmIgCauUO7fIB01M
s/47pTr6XYOTRVBJcF7LkNLuOuWzEl+P1n/pa7AHI9FNBtFXifkWFuio22ijvf45
lE3QA15UyTUqUs73F+SpmYTZYYkA0wZJZZw12iVKq5XB8SEGoP9oEI1gzijJCQ+m
UZdw07mx/mLWtQZ0IuYydPI3bn5ub9zil7lpSJ5AIxv+iyIo05JvMPZSin+9Q2yj
5sFNe5/gPud90gy3mryHI/K2FlBDgMe6dGrCA+nQe8p375xVN5mmA8Gx3MxIYtr+
3qz95mXlXYOsDlB91x6HR5diVU8fzZcH+HI6YWq0A6T3hH22N5DPQuE2U2J5mwjG
aOeY6y78dkWHHBuYPQoQ8eN/HegP6rt5dEUBBPsyb9if+UsHflEpgRIRdVNrw3aq
GuYNvQO+AcaCHsdvj2VtSU4FCEDpoEDtGDTkbi0y+xVPSsrJosg4H1q4kGycOQwr
Et8a0oyFlFhOZhHEenkGb29FEvf/5KjSQh1eCmQABMvNFAxrbsu5QBfatkKCT0IR
/s1Hz4VXmpAr93qZkK1zXwaRyJBhgqkJVkeptE4CcjqHs+oET01pnpsdReH3/UZN
CV77p0ehyhlY0zgmNw43SUPAQ9tcEEgKzK9NbXvqvhreJykr6Va4H6DBwWGY5uNN
Nq5YWZ6h25DrAiH+Cwqao0+ot7FcUnMeR4ktcKhSP71f/WCWhUHUtig7QvM2ty1s
K4uWC5UzDjyZRvBZjB11XXSe7bxpd/JcBVjhYpNpfIcoDNi+O/5bMXSHDItVuJKg
YvYY7sD4+8HcT5wmG7LBiiID7RlNr9iUsnC5PJ2m1FaaXk+pFZmS5ZsA5U5LtVlj
FKQ4f3Xx97zLPJqRGcyhHSo0nwYtyGhiEQOPBnKjzJ8yxe52RL36E5lcfySUbmy1
7jiMzr/n4HmN9+j5U+Ow/dO5gZzfTxPd3yVaS8439yr8PlMvbDSauA9QPIWO9Z2/
jByp3qnvKOh2dKYyh3EB7erH+c3wAD9xE8JhzVcx/Uyt0a5NBm7QhdoZiXdzwjk/
OhjEAT4uL8X2ERO/2g7PrA0m3jOk3fcD4XXNZclkP7a646DPM87qBbuKENAmna4e
mKJ0jmzDLUFZC/Hn97kIfcHdEibykDTnkQ6DylwHYObKem8VG+inR8KL8mE1B/iO
HMdS8gjBM7dlg180mr76A4yJmoBR50nZWL09XqFXtLqISgQk8nPi9nOgslYjX9+a
R1m0so3eMXxVNvEHQzpzZH44DITqyGfUHKb8rpNmyCUm+r0l1HgvL7LOMV2g51/1
aJhScQD6/kQq63/OyHK51gx46quUpAGplbizdhJQWCkcKavYSqnUNJ19xspAs48G
hXWPuViCkJ7PCoWYrbpn2LNbo87JYDDoPHMJw7oGOOJG1LKrSXztbkdv5JSxygm1
ciKD/2o96WVI4RPhHfudujtJJB6gA3J802/cJcGb3iVtL+pjdf0MXWsxeG+WctjK
uyIzCHJf4LtG7Cyf5pDaPewZcaKCIVdKQhJoo+tQEvKZpB97E4UMBSUrIGPM9BIK
JajqPtOSz1oaZFiKD2HeScNaf/CWO04BHmOyIuNnjzyoha+e1dpwGSqL+5E4aGw+
TJgKV4jbCn/+YJYPDjSY6pXGADugH5qhLxsSdVKvIytYxE/wbHIroGfQPYG0ccdR
yhWfPEGuBSAN2s4cN7hUGC0pcG5DH/RaS9I0S/I6Hx1S+kQbsfYiWr/e8KM6mPft
74c5qpqi7gB1SohUXty6qToZb0DhtSajlAwEyvYJvnKuXhV1jS6EcVPy+sumSs1D
yqb7gJhaVaVB0W6VglOT2CU3tl8NM4qt5t3JSKNpcIEJGwoVMIlJ+Le74WlyxMyS
hKXJ5auhBcDJPZapSdP2q2aTyihaamb6U5AvMO8i0RE/CbC5ba0wTBV9Gzo6goFR
pkcnXyQNe2AkHWAmZVVEfgMlTeDwdKDm0a9jXt3YjuVXvwqCXiaaYdgIcjc7Iumn
rfVpO4h6b3D20+3VI1DkQ6niBJ0AmO7WTz/RV4rASn6+fK1nUizuDTwbThsF3fDz
c2L1kM9B9WQYK1RXnj309hRz+PTTpjBLV5iQsei0JvF/Bpt2EYflNZGTRdwY5aBN
z1UomhKTwVAOH8cfG3L5bGJwafvRl6I5OCdaQ9YDACv9NbM3mEZpVI2wYtkqjhRY
J9qM/RhxKevg61Fe11rXT/RSCW8R7TToEpMYJ5Keq0paF1lkQEi6NSRFQwEFXrdG
EzOOQeR2QDv+kEiC6UxC+touhS6WSq7Db6j3+UEOZRElrVNdu4V4iy0U9AjBRr8W
id5ehtp0D/eNmUEq8Xp6TolPh7auXcIF3qhQ4x7BbUrLGbd/zQJ2Lia1NrUu66Zx
DhjlxbvoY/aZB2YPhVI2Mvtr0ALU/Fu6zr340ZzMsOlWCqn69N4DP6VQlzc40QGW
WtTBunrZUevDHp5g6hlkyBEUU9e4/aYTQPJ8gtfs63c/fUTt5ZUqdxeUI62oFXh7
KFSH4g92z0nL1ZOGAHcNJriqGoJE6VhTovVlvdt9ngUpMUkXVqT040wB2T7IaqFB
jpnZ6lG+H0XPnY8HXrnDIxNdVgxSamgW9UfHfKHltYMD5jeUJIm23oxLf6ZRu786
V7ErK7We4+qEKEyxDeTJ0NoelvO5jaBL8RWhuyAHaTSMw2OLGHY/po9PZXoJNeHg
nd2coilwNDSslTzyw5e+2H0IiBU+lKj3Ziwr6mt2CZx30T896135uLO/CVvwZ/8q
hgNaPZ1eVILYPCTu6Skq33HJwGImTnJ8Nd0dyHrzarvIZsF+XK0wi3SO+LjSkqGz
PK6JYUznTuJYcKGdMR01Q4m/8E4YvoEidoTcIN9zCMvkkg8QiA6BCiRpkvmYX3QS
OhY0FzAgLg7CMPHT70Ln3xv+Ogr+iQM0LM8PlKYWYjOPmHsjcmCN2+fr/YaZj4Bz
O8s0NCF2S9r4SBIc5h3ALFPYxQcEahXdXvPplJNRZaPu0RobTRzGtyq7fMTRp1fE
HyifaxPtYA4cz8l3fucWs1p4Le/UjKRIZy4/imWaG3s7D/6TY0osxVCc/XOQLvf5
xP1KlxGSP6TnxENEAo2QxYPLuZCwadfEmbazrK8/DJD9s+jeCNOQuGvkeCKHPnec
G0BKtFq1Y+ycJ0Mq8grnPTIlql+rbsjvtoyCmctprsl0THFSafLOqEBSO0sODcDz
7YwUr/9PJqXvbLlwq4F1MY19xEhdDuxuXWACDzMfEg/Ndn9LsuqnF2VQCtoD7XJw
+8Ggedw5FtIBCSoUcy0wvkXSmEzSsHtTtndxqD/ooyaChUxyXoJuAMW0MU5sTjbe
n6j4cjK2b9ox/7Xp3v0h4VMkQvLlVYsaF6qYN6zFRZuyuHDTCrycepmAEKdGErLM
94bRyCb2K/t1lWragOn6S/KBEnMsizQRjCaxf9RT4c/yMtRbEbki3vDhJ4TUwEuj
HCTQFfPBIYFVCkucrH0KelsSqeKZ418VgiWEt73gyEQTGMMkwSa09sId14J8cD5r
7/QhkXyRhVXFWQnfmBCSBhGAhdGQZP9M7TYZDX/Y/lwnOmElGKVsBwYZsNPlqS7o
E5YJXWTDsGh4BGaoN1LVStrNycfa0SGiCPl/fBVw9C2z1LBxskQqXCE4seUBQ47Z
TqyoOfaIoSzCYA+b8BaGbdHbXEJ14MQa0FkHpdt2BOTRPxJC93oqKJTZKX+zTNFs
Z6v3MVaMHzHaTkxxRU/UGNFv5iJkcdVU3dp0xx9dGB9ZqwRk3o67r4etSt6yl5n0
czsYJbUvPbst/KXK9648Ug37rC8MuvsHFdBKSKiCi74s2h1rutMLPVRO1pzw9NAq
bsAjLO0d6vwlIBqW/pQ6wlVTYQbhYv1MNyCbb4xNG7CU3s8k4C4i2FKUMcNhnRIU
qjX2Zs8V3h9JIc1lL5LjhBT1R7qNL1YEF8+akc7oDyy5kYtYv1QrlkdUJPqqTjZ/
42klZpoVgd6qfmO1fapfgUndxpU0rXZlPBGePk7szuttv2xCgM7LUJP5u0KKHJHA
td1d9W8gvXWnL4tWUOM+HTAt6n/8EL+lFlq2echgKbflBQ33EMC0p7okJM4i82Y5
bFJ6ylOxVdS79MrZftE1oJOOdBfkVUy86KfC17httMbZ+GOkhmm3LsWPM6d67ch8
eTk8hpkgKzfhcNMWWLuPtkCzbO6rhHAtHfOIoknhRR/GsCF2bfrSh3BLRJ+1MPg1
hDTL+FXifbRbHa+4IqjC9AHBcITUNP9wGVzT18CZmrcCQ0PKOxlyD3pIalwA5tYY
n5BjqawnhbqNyEXayBvgJ43RSevuCBOgn/FOalsT9imx78QwYE3z7zzju/yD+hAt
ZfDpShUYBASm1kt/93TIbsnf2XknIAskVFI26rCodERsKa+SdnJAM6nne0Dvc/ZB
AymIWj3oQMTFGnZQVbJ7JthoVLjRqj5j5sx5Le9Gx89QpLX44xK1O52rYCD31DgC
kML3Km8NSx/uJISa2nqM1SpzOL7reRyaGTHVQL0wJ/ebsVc7r3cQMHGs7AfoaFzf
4aqbPfgw2V4QQOIxRj0zw5EOOcO3Bm2ftip2CeZUx/qzHQvC2Q3QoZgaeL1QmaMy
17Z4/ZaZi+JfO7uuwyT7FowmWdDLMKPLCmGczCRBiWM9zQmDYgGE/U8HJmP8pIxp
7YFrUshHuUWqOftf5fs3YuhYzvKhYAfrX4C42VfJTQ2GNMNgoCK/7vdyrTUbRgnq
y6XYC1T/LUHIsF84OHyleu8GqMkSnckDf7Exs/V3xUnNhgq9ZmxJ9nfGNivu6mgL
HfthRB8aWjVvlTGaOxX92lP/a33b+vvavA3LMylnd8YkXLVTYL6lvV9U71cm7sDt
7480d2CKKduVXgWUwk0ZgzixyqR+ZcdMsJ4lB5eRuiEHaEuR7CctS/zmD33KrmsI
3fu59Bkm91qjY1LA0dp7YtSaYt8t0LJIKpxwng2MIDh7TW8Puws0A4tkUF7oI67B
zcKEbdvSIQ/2pSPyR7oSAu6k6IAPEkmomnI5yox9FSFzZz//lE/9L3ggV237+AEF
a05/D1d+3xcfWemOrOoPnJD5yclMSqStFjGC6IfEggb2hattuJ+PHyR1AnrXMObf
1D0ZqHIvwI31DnnkG9GRBi7Oz3BAasstBGXhYDB9WMkpltvDEy8Gf7LP/ZbP8KCf
5fVG1Xwd+cLT0b50kMg+PlF0vPf+9BlkGFc1pQmlb1E26tPdmzSgUEA46xZSDx8B
6xv0+fCcVu1fTfuciR8PIdYedyAGLNDCHXnJq9AkJpewjvyAlTEuLvF745Z5GTuw
R4yTLX4c2JM8PZ+hE2oTr5ZDqJl63gUDZuPYL8Lr1V4E5XtBinBSCAfC7WZqUNTp
Gduwz5pLLlI7/0Cd2S2n7kQ7+viDIVhpaXfnJ2kCw8l+FzznN/s00nKbWDDZ+S2U
y5pHs+um3j/FOHXPQWjffdIVeNERhLgxXvlROq4YUzNjDMCS2pO/dwk4DyEkNG1K
jGd7k3bSgnK1fM94qMDGkya5FuWW2UHCUPhIHRHE0or/unHV7h+QCyXHY0BhJ9A1
vegOYnl6s+8xQNHGhqRpZ63iHqUY/6gLtWIKZs/3zo8LyqGD5JpIzCh1uOiSDRvp
Y1WghER2l6RIzVULjnMMgUdBQVEVYRV8G8lgISiJ1GgYsqnTDgm9HSSqAk0x/80z
16B8MKFEuKSlKgvccT5Ke9VzIJ0Ytm5VDcmUjBOBd2DgBULp9Ze7WMuCCQPeP43/
xsemb3Q6v2RX1SnqH9G84u6xejDaTfsE4FQ4OPE+M03eelLklbEiAO0eYcGLEaQQ
t3GHA+se8tcsXe3JJqVjma/upU8DB8r6ymzbQ2mVUu8nVA6+YcQzqUOjzFRLN07m
H6B9wmrNqz2DgPwfKWBbHSepogJndw6H8chbJz4EDubYyotWNSxF76BJHI+nmZAK
oXploGrcniPUCmL4/oxaMFtSNAtA4TwRbozZ9gsYq/YqyG7qUdHir3sUXj8APySb
zRV4cn165Z5qmaOSkEQBZ6NRWNOguxsXViE8omO1JxrhqXxkVAAR0EDn4uZPuBEB
aIdD6jGmZdqfswrcmjm2JXYs3DDCcO3TypQuNdbF91zbS75alFo7DeUmf0U87tUo
Q6WmJiI9ne+rDefyjaMX/eJMbBCdf/jfqmXkFAveX/EW+1Sgtn/gYUsgzgotpc2r
G875VxegshB6OXBEw2UTntWdyiC9yu9sD13aCAN2IbRU4b4mVpn0pGcVlanKT8dI
KxHxzONTMsrjqo9wyCDeOVFPHB/OFH/G/cqGJy+fexTcl4ova7H5chGSMpxVG/i9
6t1wgWwqret5thqSrAs3qH/3P3WMLwvTo63//Nhxhqc8kC36lgKUur9MqP2SKnFX
M2zXtuQ/CXLUisq6w4P/Hau3p+eeQpA2Nlb8NjIHnjqNvgeN7ynMbKtBjeJ11E/w
mNpwoSPxRNkOhJKB9ajmDV8WqcCdzi9N0jzzoaHlLp4K8BB9VAH5seDNTe4bhYJ7
AbcA3NxMJkP7N9k+n2gBSQOaPDVBXpRCyyK9ijzN0dhrTvkV5pUGf4Xr+7XS/Jpn
t3mEz8/0cqU/xLCO4Z1mQy6+ZcrSNZpXQ/SW00F6a0VrCa1Dj90PvTpnQoIwDsSw
5V3jThXPDXRzNzy71SYK7Ty3CginVYW3XxttMo2mAYsODCYgybTDhx0dvh5vM3hD
Hxa4VpNVsFNaZddapVRUz/jwDLSyPTWYHYfKqWqNT3QOmhqcjwsv/iU4jJ/7z0D1
TQvZrMoh4U//hshUfpsvfq7zEXjTNOtYQ4YMyDvMBLtXwEusWrTyaHIbMmKnLZmY
MGUkDJwvjKONLFr4+hJNyH7CZL7whXaPjfgzk3NX4iND5647KZcaNqE2DsWdwJCo
NnOFJV2AqmwjkM7gwAul9QPFk8/BvG6iVlrpvYSgWwgze0reDF9F4C1e+atow/2a
w+iNX8p39Af3V0nAYF3hIf6fiOTM4hHaMPFJeU20KCEDzBNQOMO45yGP/tdzox1/
Zk8yOCkT1sAP9jl6bEHbAo9VWm91h9rqJPhBzvUScBTuacv7ruagh6pKNRPMZRGX
zxAERihXQ+NyemxOSV3fCnZxdz+J8GCkyOQBFlz0aX64yyDqUb2y6RYoWfRRTQJj
E05wRI4mW69jdtpXl40W9NSsxe48QRK+LZD8moILw0OEQx0RtQSauDrKiPxNO1ab
GcHZSchh1hNxy+mjKX22/5xG0XhBtdiVUeapGeri3/2vE/13U2YlnOOFInTxBjLe
7z9qLo8vzCsUI9Y9Z0v3wtJJXIfLhlMDxgsWY0qaSo1Iymon2CplThJqwFULfpYm
DB/+krz+NhSMSW0i9HURsD8XepuD+6OQwV++n1kvhftfrlIdG8p8iFhyaOf8gvt3
LQukB4fn9k3Ih9jXAeXg+U0MGfy/omoyz1Aq6D+Wm3SjjBIcOYN8N5UJ8YbfHYOo
Pp1BXYFGpioEu9AkQDxnmcS9qZLWINvUsPjlowX0ppYRGnD4tbd5sYzQaoTjVyS9
Ws3nvsVR56HIJPDh4EBg/0Q6czX1NorR4DU7YwklGpJyZ52P6Tw+bu3qoK0I2tYs
xve2TqUbStrWVdo8PT+gTZKBHNpwQQAUH9vWaz77hCZUFT2eMxxHbPCOmOgZ4jnW
AXV0zxP6zL6cr4wnmE27Pz/GakNLfvp+TjX6yfyNxKYFPU5zj7ZCljx0iDrMLcWE
GPSXaji9EnG2MDFJXJPzF+eqFRc9442xM2qJl3ieDLF5H2UfjEr65NjnnY48tUpO
A/n9gfJPAWnAGSB5/ylY9g5Y9/GNKXMMXZ4goPQsXoA7/1eD+JloGrCKpiCw45bB
bUi+meGUzHwp/jMFriJt38gZ4og9+zjffLr8pMWYNrum66gCVY1pWbxy8AMyHSF1
X48eK8tPFehvb8PwW+gMDCqhKFEp37jh6QZrUHCOi39bNBgSta2Gv1QHqElUXcxx
pH362mXgrEwPR8WLd15/18jy1t8/vNxqAakL6+uVxv16/IIQhVSp55t6QN+dapwQ
Rgaaxit/feLK9mdYj5r6hotu2Su+t2qsZvi6ybPxrpGGCvTdtGiqBA7pm55lHm1h
Yu0WR9RbAvTpSbPA43KKCRmAuQ+IfaWtpmT9ew/HuaVdxOioA74VhtAevy5dq+hB
NpRRPS6ENs0H2yKTW0ftVf08Pi5/Au8UiGBvPPnRIkBv2TUuUi3JACLDmHV7hESw
BjM5klSmRviv65Soe58RxzWvFw8pCWV4GWLnKaW0ceIpc6IqUoVkQjIEmAThfh6f
dj6OzI2dTs4NJ75GcqZ2lQ5YlwUVOc6ZRU/Wb6smTTg4LNFVY8ebIm2WsvInEyrD
kmsFoxkHe9UGBrqlU8X7MwHpqou8qWfsru1KLPMUOlt5gsCHLXaBm/ogPW94sS5y
Mw68Y/rsNTatR1O7opaLWYojg5PvcCupL41gnbZfLfFspUdb1pd/Lwe/RW/sXJeo
McBAsnF6LaboMlG7uIuX/QL5AxTLIf+wqnQGGTHZT9ep18afZohiN9qVYcxy5VRj
P6XxZoOFUxJPVjnSPeSDw3LGybkKUauuXHX2+8joA0EKYWA2sp1EtwpEYkNfSmFL
lAmSW2s/hq6hGvrtiJgrAqkeUzaKFLVypCYrKUpXH4/Etslb7ftMrz+FcAEnnuN0
O1b6efntOtW8emR/h+mmbFpVh3IsHhcE1FaNJDECwyVQSAM02wjc8dvScDebkzjO
GBeORjV30fzqDZlyTbmPKwzmfmYwpxA2tsHnjcdtVNU74c3xuCyFn51/34krB5JT
lpvfM+6jDBYprSVQWU5ae8RLhtox1qbgg3jYM2zD5KddrYbg8Rc+u6UpBRZNLXLI
PqXJJ2jWbRASzM65wETFTMEWIWdPX2j1YAFzfD6Ze4izUykKBF68hOd+uOCSiAzu
7JsD2x2Ect/OSFDp3O6EpcuYjo/MR4p+Gkt11tVqgudepqzqPpSdz+tqxFLTM073
dvv9kQ75ubfXQHyVv2NPsdUxo0p9kzi2S789N9M/OAhxpZ3B34OhtriZfrdfWnlZ
Mk4JTeR85N4k1K46igUpymuzsF9Ku3jft28lM9sgy79AA8nI+eM5Qji4ctcw+6GU
n2CjW/U26j1yZyUdBNfa/4DKZ1IMmlHhrSWnc+MgHCMaaxcHSl8J2X3STjzDpggH
bRPW0ZO/lP4phZZDPPbv3ofUiINc5WWkQzHlGwLXwCbnnfIQLzXd2XztI/2NtWMt
r9A05BYwX1q5Fgzks8oI5XnLQO4G+mn21a/FzjbZS41qsvWAWPc9hgLkVtGS6Ehm
rKDCgaKPKknu248PpQJyvKamzcDpdBnF8sM6v04Ia59M9yKvQcXnUgbJx0bN1ztM
2d7aqZ5onLbpBYfIHEWbvuOjrogVfnz+Xa3f5mJxPhEZ4xVk08L84nWGg9CR1BjD
/jEdZIwPDdQgAwlM5OFijPMZSEe7OrmcvFEY76Enox/R02KsH6dytZID6yZqQhJF
Gdt5O1B988T5anwHK268M5RZ3jryHKJ703Mer9eZRU03TT2EbJTOS6cUDE2bL2SG
sqBkcvxq7QF19WCjiGXgmABSWyhifyfqt9jQJieciP5umc7S1HJqrtQXQAZuZnOX
Qa8yDVxU55hV0acDRGKEcsT1MYlMGfBLx42j470DRfUsezHPhVBGHjPWXhjrka4R
A0qupq6SB1RWMH7/SPuGTWyk71NRHK7K1p5BYf4W3V5ya4xbtNaFzs+oaLVnlI47
38EJHLtulSnkbelcz8sOH8zbhYxEWJLx35FFyrBnJ579zPp0V2XZosmnTj+tI59l
BLGpSmSoa8WBttGveYAQ3wioTeTEebyCld8epuPOVbZ+M3lTr7wuZMgMysR6CFdN
nFjoYFhdR8BD+lckRTcWL6+Ku4NImYu8n6Jncstj62PfTdmu+uI3FUQpLR5NbUQz
ARUC2I5lLEcktCSLelsNcBlz8I5+SnUmLDxbk9O+xGp1h0XO12BSb2XzsfQiABmB
sqYhWQFJA91D4QxCfn4WLL/3hyOB5tmcws49ZbgSTnORSoevqU0Oe3tVjvRm1mes
qEDEcYuEpFyJ3woW7QVVuo1bgUWHplC8H5Km7QNAG/U2IJkE8y/5MV7Dw7/t1ZTV
mm8Pk2hm+ZLamPhAvczUmsoUjQ1Xs6raNw/jxPJ0T1MRrP1T4W+MI578VPlvYeAX
lHnYIO7VLiG8oz9rcZ5MvRbCXZ82+YqOC1erXKWlPxqsqTTM1bTSTYzRejhFYyDb
weXnx2PFz4ZAEdXcPrQAb8hN9/pxxsjSoGRiPIhFrsI5QZsAzTxjwO3fPjb30avE
ESg6fYUo5JGQC53dEgPFbc+h3vWqbI32L3JXLGMl5eqvSE/emz4RBrKJOA/v2tqR
6fQ//Ph9H8Y/r2pMpIe5fquYGYKGLGOjBjquUvaCvmjPzPCRyihUtjnxbfK3rSY+
D12IGeDxHTSxBzglRE72eLTypWJyZG3ALrr62jJD54BQloBm5xd2xufTJC4Cg3Bo
SgQnnHYPqD6Y3F2JVjJkMIn5oNPxJABEHTxbRgKxJZ8jEI+IQDC2lHSLpfjk57vH
1I7p60Sh6t2rWNHF8ZVpsBmvG63ORyjk0suW7mZEbPz/P3QynwmYbETX0X6qAHT7
AYVKnEc/3tyYxFNfr3gW6UCsTqH6ABZulElmCa7SQ4Df0OayD7si0mTGhNW0Qxur
W5ASrSDHQTQwTFxqtLhn2lkHQUHrD/p5q3Rw+sNv3NwxnwxKdpgR7FUrXygxfOSq
sYf/kuWIF8uw9ClUoIpnES7GNnN8NPpLZyFrPck7tNShkq+W55ihDpAAi5Fa3mU9
THbMv+VkNcrrdezQ0+6fNqRpzhaI5+CTsiizkQYY8hQeJT+v4MRtjt5sLMJnYBvY
XeBF0ZOCUmmSuoGPoBk/kUFo/TwSH/ntWFzkigYAuZ/wwzFLELsUiL15ozGKdnJT
wgUOfLHiBSRBOJnv678KDY2/uCDgrD+cKTkcLfZyiqxOXMFDLTv0+E+IYaJh8kxt
aBSKZfSIOaa2ai+Rq/ZyYVdywfKRQR1Sftf7rsqClZoi3SIb7jJVY3XUg67Gr/XO
XSw/IBTADJW6b1R5d/mc3Ljpuiwq31iDrN43zGnoRWGnLs7051geUEG6nwfyDVe6
3Yv1HDeiZw4EmhlZuKTaeyki+e2bRaixRoQfTZx/sxT9xHhNJl1MxpGUfJ0i6JeQ
fuySBaVjXs6+j2M9pEdThwUp5SCs2lhMY7KZvihq+wjE4AZyLa/mXDVInMGnNDLG
BKFD3RZoNdAyY5qz45sJ9Ns4BaXzbGZz2HD/lUMMzWzl508+g6ZtZvCS1XMk6EQI
BJQVCsNIfrix0pEiMwf7qci2J+ockSAOgRO1wCZVEMqtOz+ee3AQ8Je6c3+m1hA2
WlPJwZfSdehFSY6U2YHzswDAA2Cs9fRXaBwR6H/tJKmAZ8uZ+cs7KtlLzZ48Bb3v
ozpkj/QZ0ugPHwJgmVlDojOUBtV3oyDEIjr3AwmBm0Vdk6fuvTyw1nVFd1WW6Mjk
Q0RdrGr6D6fsU2gAByvJkJNJpjeXDNfrWq5pQZj7Kwwgn/+PKaClR0/T/iQ3BsWR
MHrHC1c0Bab6ApmMVeJ/xkzXbEnBMu8qlJWKSoQdGCWM0bc5DnqQhTI20NvxUmcp
hCrXJUzTMdceeaFr0dWDVmX4UGauCVHJzgSkgfLR85VTT9rJqWuWlTJ52OvTEj9U
zOigGTdg5CtCt+uPwwjD0Ch94lfazzvEvlqILJoeQl+HBI7K8PWQMhUGaTkwFSlg
h8NnazDr6M2WDo1t9xpqoAIkiAeCav0kq58xlExZGgPZbirYTL/z90jym/NmlFr/
rKOXzrX/Za5Wegsoqc7q/er7Td/qKSUniFVQBUla+Y306F0aHqiyCTd5TUbFkYRW
/3ubXxkzSZDKZMgxNRpcEFXsxrmfUUwc+eRgWMpgfKtfhZ0QGbI2Z1OvgHO9H28B
C4f9Wi3UwxhUGIzAr5K6t4vEWOQfpXylCqU7f5smMcpYZUk8dXB4md4KmpWoW1XA
uz4Oc6f/F591IXhcUZ4Kfl33jrK/9t+XAD9hXYYNjxX9wcMF+fKj8lQ8A0FUBNsj
qvohiViw6MV9cMgaWn6NXh7s3HGClyy6D2POjdDeDCk6bfa4bXf4MKAjD02ARv0q
JfKpj0Zvq/cAwYZZ75HWwIX4c3CoRuhKKEYF3Oo3q1iI5sXWjO6HZoSfRoQ4N8V8
acLHRV8hoarzlXhLJEcdtVrQC/bT6Y3Vj/j5aoGb8JFaMTyD+4T8CAPZZpF1Unkl
FAOj5sIW3hIz+l5m8KBomX4oVYu3IMFK+ijFA0NWk5TDBhtuDcNo/69O8zFgtmnf
20K0AyAkPE6Uv9lPOz8pf6XIok34jsTgdwOoZy5kYIO+TNwSL84Ju3+zc3DgcZsd
tYFv9IdbbvL5OzAMPhs4coyDbDpMJElob/fEdTKXHNiBiXyirmcoKZBwYdQguUnL
pqmJ28cdu5nB2QVwSIBe1EZ/coHq6+ksuxZnsaDPX8PyReGzaFpYbAqcHO2lNvC5
MSIgHNCZec+sGfzXokD9OsoiHSr1ZsgFHiwoRsA55U8lFyP0t+/eP5jLyVUwVUur
y3eLI/5nSFKdH4j54H72fuQDNEGqRQJUcDyEv04L7kg6Vq6Ee8xiBgK/Ovezrd5d
dYG7FC4QxFJv7rrLEIfMDlYYOrhtMRw+hZmaF2er0VDe5dd1xeM/QpdFzrj64MFe
oF71qZZv+cDZPLnOBlzv+aB8/3WeGpAFr0OG4k6kLcIzz2F7TuiFLDOUKm9A5lJf
BjQf8doF+qZWdXLzzBSVG+I/ecWBPADcklEnLokZjPXDv9Ed9QUG5sjMuKfpZfAm
r6K0yd1LAkDlSRXDbOzjJrUQWCzw+6nia2/VrikR8x8WQjcEBjE0Rc4u/S3U/qxT
5eGldIRVhHgjl21uiRMAv4SLWUothqe8VkroteQVN6ncQzN7OZxy30zZ2iB7iOCy
313EcwMMq0E1uETpiDw/ERS5KCHBMagJwNH1bY0QgPhRoHnMIZGkjXMXMbynLwQB
mi5EfpVv8zsJyNTm6NQsbuKe9KBGDm148X+ZFcxOxWWFNk/ug7FQMNS2OIueocdK
VyL2WgEVTIBIRJD6JSaCFfqaQA/G/kc19gZAu27xEq8w8C1S5O0ZbPIsVjcitpLN
mDNHYx0zmJje3GxyCoK4OXQqfg0wi3rG60f+QkgXjq4IYb53vdyBbb+Q0P4e2Krs
TNZjt7MRlyV2ISc/TbcZmTkSYzj0IvWnhYo0o7DTjkAVtmb/JHLg2MIiwXMzsI4L
8iLFvWbkqxJszNrKcsrGnb8czY+J4uN+ocWmhWRoHj63BInkSPKjiv/FnSMK87rx
W+QG65s0V04HoLfvUrM3IhoHZgV65U5gaAE1Q70qFrz5Sozy0qQHzfE4HK5n/drp
8QVomZRlFbnU97XngA0B2mNlYxy2ncddioBQ0wU1Jy+UdznqJD70TwgV6HpHWtfx
Oaj4nHQW5/oqb8vUDB1l2XMH1YVCnrV0JL/rfLUzLg/ioC1h2yFUbUdVDpamv67u
BDuKSP72EDCU7ub54VbjjdavUIGJCvYTN24G3qxXw+6KCgUudMopFidfIUVVWU5l
4kUkIkPJJzt8sHEZB5s5U8ORKcbtJ6L+++fxsf38PC1HZ7w9AhTzGjLZeZMHscv1
oLgv6i5KVcPJWqzf85+ScSSrX/aR2DOX01gCC+rDjJqyUsXaXjC1rUXJbRgOOURf
2KlPRpMB7QuGkYf0nWMFHIWnvkzhhXs4xCZqVT2u5o57eEjN7gdLCGuvVzuNX08V
6QKXmssHyWBgoSP4xYyAV9onU58CZ9o86Jo3T56o2ZAW4npSgWgSRJtNfkIYUdla
BLP1Q6Noui8vKhh0MCprxdgNCQnDAHujs6s/+wB8uyFIujFp56Rmx8JvwGGEXKhL
XO6hbPQMoVq9cyOGRWYnkmX7iBNnACkpL393QWNtFO60fJ934inm7crx+OAFy1dx
oZG9hwvbIAAy+sxiNejiUHdqJfyjHa4kPFoUP8naUYQKWZFekLAAoeHLylWo/n6S
rs1TQ4g8b1lCaD5FJraXW5mcxCbU4tMnG53OpMP7rvMzK+YHugCBwm6FzsqzNOLp
f28hCUSj1AuJ7AaG3TspuJgKG3AuUgdDiisGiNz0X/950Ql3Y0dmNWgZCByTTVYh
lXFmnr7+UY7wu3/6hY0/XBQs9vF3n52G50vJMS07/9w75GG+k5oFzzNWIFamPtHd
CNiTVRvnjwPWkCt3Yej2ObgP7RYiGh4OqcHLIUl0GOdJTUYAVieEpHsQyBesjiJM
jQ0RWJHA9X7R993FYkSqHTZxQiLysqpwjP76m3yyqoTvPjRWI0Na+nc34iuWlDbB
MaA0/kZuSyCYxU/bAiLdd6e1XB3wOlO5K6Qzy5lI0uerEGjqOmXylfDtg6Nr+2KR
l/11c4Vt/GyuQJy8cb2h22IsDpfj+wLqn9qp08134sXaphF4y3bfElwZr4rr0VQP
Rd+fsJJ1r+zRzVipxROz+vl22a76v57g62QRhoIYrL3z0SEj9CF1BWQrGauZ+QAl
IwDYF1pyXVnQeawqk2UauC0a5a4HLQgpTO9XUKYJiYd+zPMZFAnvggypIp7nSu6A
vvdWXCO409dLIDxQPmSUDft+f6OWRPJIPMivJJYl5zFct0zQ+ZGlQHFyhQFXkrDs
1NEDIz6R/2eAoJjfRQzAf9yocIF4I+jObfTJImozd9MVYUpTictLrbzz9Ya5ALzk
YSXhZW+zppL/okoxSBJBNyL3K7D/Y3Tfb1ZNjDbJISAN1NXkIluVp4ijxrEIGccn
qeJPSoVy8lXlAmYcwszH96ZsTUvNNbduDmL5kmlv8gYqjRksGuEv3lvPE+JUbImE
NTvL76sf9PdWaksIBddmsOJkrtlIGFKqtki+lVtaL/vHKfhOdSPVc4xIDTuICMvI
ScgjJoaPyygiRkSxfnt3BgYq7QrIyCyOqWvTVNPbCCcqsEebHNnzCNktwvZcHkDn
tuMSa7RBblDnkbj9xYy3cSN/hJKdJssjKCQRPJGy0ajOh5eYMfe2PFLku17TzICs
j2/1P88q+REgs37JC5bXzTlS8m2mWOaArxk1xm6OCePJseJWVyzIfTPsfAdOhczl
w/cfdQfrDiyIYF0qmHHU4Ia/D584nA9Me1Jsaz1tfBJ+kh/J7uh3gijANoWqjlbT
nuRQ61C3b+FCBtjKtPS2vSv3Ye7cclKJ8j/clVsM1+fnBk3IgfLK8bq38+zd+cj7
vWne4LuioEKOyHNhrkQ20lkRfDUiT5iDPaWXY6kZymd8R46DeZ4xS2zuZQUtl2Oc
iF+2mcxhuiT9b59PKQM4199xJFkLfAlN0LijWNjsdrcKOWY0Xv/KvLszD3+4QKGM
zh5cTSZHjiMmsQzgOwjpnnN/iGo8wW7JQhHnol1WKZo/9XvYEnACu3Hqs1GqbxRo
PCAZ03wQHbxchRETCJoN/uu1M2mPIMYRCgzpYtEn1/YELBQtt0LeeUODhFVs7sqq
qqQG0J1LJwVhAOs2txkS87MGB+k54V1SmoX19w5r4eCvtorwFpoh/RahDY6OxNLn
ym3jKdTF7CySBnI5NvxpA0Yuh245Vd6vhlhjrd4a8HQA22GC8PjQfwq/Jx5QVeQn
p8uVEdPcR3WP/AP9BeB2LTQ+cV2XY4sk4D7Xh+uo7va0JR96or+DL3HD3/jIWmKN
InQ1haejZDD+qcXN1wiBQPhz3UFgyTr+oWKf5kW1CDPQu9d7X5l9MtXmWnwtfBAK
v7ERfuJ1+fLysHQhQXr+5xy3/WlmUcRPL0gaLWWUVCOX2s9GC5AwZPTvtlWn/i2q
lRlO0KIyTEJ5xsxjKC3FqbgzBO/lBQF7AbnBbyYxQh+kfdlo5myDy8z1WvJP0cnc
PyLo8OptAPfsZAx+r1wLhCJUIRAJ6v1+ibHUguNdGb+jYbdH+gGfkzrRP2drLcms
ZNl8+lM+nW6O0rjyzI5oVr32eE9quHrfBjTjj1m5ROFE4B1QFCu2+sguwk7bkpbT
DgePWvqhxjyWsmx6GFgcUoTC5Oi7WG3Ll+kajggIO05hnBHwl1fxhd0Js4/GpZ1w
6HrMIUmk522ZdcjAhl1Ju4uOVG6eus5wnxOKQN9h5HWidTRknZemGu7rEwjnXdyN
bf4eX2R6YZcno9djLElfzbskqsxDTg2wVKodki0ScBXKyS3o6T52jEz4I2LFrnSK
vYqU0+jYYQDcL6wWmLoLS32eUe50ZmUUR8KcbGjxGD+IBhwcsLXM5cXeD9QOW+Md
2doP79OEiuYZgQZ3zdon1Nx6dveu+NsciQE9UBH+GTCOS4SwGcVlzEs1zqx4NE/K
hfKdguM5LkkqBI02ccxfuaQDkhEy7vgQb3UC2Ys50peywUYbfGkgJWw9Vnm77OM6
fiRkjbweAF3fS5YxmJjHCM3QpIiBCRr9vq9K8abLYa4vbEXx/I0MvXNDXMTaKvsD
/4B2EF6rUFPD2gRi53fWyGwcWRMNQYDkuo1JM5Rq5cYjIWMM+IX51ClrES1M8Tj9
MAxSZEJYedNOiYf7xJ9YYYCggNruvhl6IFYcgFyoCY4MxytQ0vw9qUEWTyBUYh9Y
sIxP7/fhfN1ngxqL5VPUv3mnPnOnr0KGv2IbOhpen5FrQQ+KZ3IQ+u5gz/fOngE0
XZhhQ3r12zw1NNj0yqjFj4aHwBo2p1tDJqLC9WdwDsHFz/UYVBNMdoNKQfzU+VeE
WO6zLhDxesmCwu/4fnB8AZjKgegnkrSnkAwBAlyYGhhuTBIxF7nONRu2d7a+Tdlc
c8Rv+1RTKBihbW2rFTpGtmi0g8q70LUaBNLRiGPKtXksFqKcoYlUQbjpvnd2zs4x
MjZoSw4NhFoUI4RGIv6zFiFAnStSxoUo+Qe5kX9t2n1IIfvuSobAUEOeY6ND7reG
7hcV3udQMM7jMY8zdgyknY0N+6sR+F4lYAkw1Y0pjWc59YH8UJM0BhaoCZwRhLRo
hyyiSzdKP7iErUE47evV5qVSxgmGBvJnffoVWMcQ5wFEMZo2jHtklMN4NmncVffY
v7s92bW/OAOAkcaxdpdBYgFCoFtYJlKZf2JTy1q54P3p1FtZ/gFCz65mHYzYQiPd
EawhYKPbFiTOlgXm+T6sNI0kkWfCAJ7A67roEqm0mA0kH7DTfYjdaMnNZFzWk6PN
TP5khPwemp6ui34kmVABfjizm+MZpM94nOhNlGWEkBZi6p3cUcJImNTsp3cYW2e1
XpMHD1g2EOIUbHDLlpCIWvfyy02KL2FXJY83YVZ4UKRe6lp4dYeVc68lESlP6mNn
r01dAOTQ8aAmQORVSUdRktF5BuUzw7R1g7tkjL/D2N2TxZaUWAUBgMvk3Wy6tSAs
OP6VmCethFhFBGxmgfbretbhf7ShJjuFiQzsVwsb8ajj1HGPetlGvKzvPCtcM+Ri
r+ApIg/vQenak7Leq/qzZrKDvj8ztFFs15knphuHA0Cq2aprnX8WgZB1F4Jh/fv7
eeD05yAKXGVOPFuI1S2OzHQG1UZMNdiX6U5eHbbb8SPoFw6k8O0KUyENQArYZZKL
w/mrY6H5b0PwhER/xz8Bb9sU1rw19gJmZlP2xL3fR/oxaFA6VuNyNpMpyIIo7w+K
vamfzlWym4ws5UR/9dRDYKQjeDxV2gZNlzF0VOkbILJHjFGJA6mv1gbS+ENRHdto
fiYAf6Vx0mlZk86iRZAZlnXKE7WuHcIOTls9uYYamz3XnFgiYjiGJUWQvP7chZbT
gyktBHwH9mSummNfMr0aZ34lBnU3rlgS1Jjl+rBjmhM37Mc33VAhoyJL9NYO+15O
kIj8xKL5d9KdQQxylFUVf1N+7pOaqMMRRFawl/5FWWhO1hUeqSIAtLuz4FsFI0lM
RBspAKrbIX0Zg65TkOnNRbNuRFFKfrL/t7cC8W9dqYuMz0B8dZNyn91Z7V5jDXmn
dBJbEI9pEVX/CqOj42UiR/kV4NfOwetzCI04nhm+Ld4+yXOe0+K7hi8Di2KRR4eF
JufvCJJpkU72Wg1yaCzaiv443Yr79afG61PgxFvhyof1Sb7FwHBYKr3QHGXn96fN
ObZnM2QOZODJdp9O/ZR68v4S3yrd6n8O2+8XZH+NePZ2e9Y+BbPwwwObCYfvNcrQ
MERCL0bh6gkWeyhb2ykzay1M8GFgPigwPZWXDAmfUmf496Bi5eF5bh3Mw3lHeOY4
WM5n1Mb2elzT55pAOnokl4m8sS1oAiXkhCsKrbvCPTTYlGsV/aEAj0GlfS7AH1G5
vQu++8PHGkcFXoH/yoDn6dXDa4LdWJh+l9Yka9Zo0Sc1EvWiV8hdDG6AY6XzCa4a
kTf+HJv6yvX5R+CL3J1X5CwlnrqxqZCuYJ1JYNQNwpoVR0ts5hl4IRLeMW9jJxqe
JQ9cCC4cP2Oe8iSPcJglAgueZtyM9U4dMh1uPeQJigx6zNOnp1ywoYYQKQtUlMAT
fBelIrWFbzncdDq3WwSIk/xt9AqjU1gnShNs90715ClwhuaKGWDRAa/rGoO6KzYC
SyPMPxbk0q3PxeQt0YA98SA7OnPBe7GO+l8udLliqr6ITo32/dAVm+qectWljVsM
gKMhfFPDkTIBc0ljzXWA1ztja8nBBdoCFTW/Wq2GZwWkcl6f9zNorKUv1Xun+gxi
oiSDo82X2tIz4X/BVwK550K6HRnmm//BjuNVyPm6Mj0B5hnv0G0IEp7ktvRK1NZj
0AXOwG5rq6y0F/mWEqLkNZ8a+3NPTFWSyzaM8UaGKpuKy9/E8kS4L7VDqh+1Yfat
W/qKuCaopXO2MtO1A0nPmIkPzu0UzUMKGBmxfxbSeS0GGitQrYaGyNZkbJMXcP+U
17ILFnZUucPoXsVy5HuEiOpN4OU4OblmZIjqKr9WlMUrNhXpih2JzsxDhqLkqEvP
5IpXhmvbMtaCpRhB2rnT9PYQHryQnDfP9nr2TtR5QD2yo6OFCV6Nxp4DUOIFe5SZ
crXvax4z3UBPJtNI2KA/K/s0vxC9uyWdljexLOfMDGPaGubwGunsAktUuZ0Lw/Sq
e1VlQ72b1QaqLfTb1EWMshcD6Qcu9+yZUhcY1ZW+YrZiz+7RJKNcdxply16k+VZy
chGf3lCznu1/M3hgAbk8Wnh6vT6x5bdnfxCm9fM9Vqt7By1CaY5N7ngA6uABiPwJ
hvi1/nRiIbB++/AVz2sVcaQHgCnWwakO+SLwS19B+lTig+3KgVN12axfiYyaCLlX
EakFvBQBSFMUQIxJeueXdkBacvszmO+h34hoC3gxoaWqY5Ac02KCPkA4rMi5LBbH
XwjUs+TSdGktvcRgjwMcOtlD2hCSoMkklaUZQGr3AB/n2Oebyj21wV6fy670y4q9
smEeoIOuSpZZ3a6+YWUeL1LUUxEQ4TnzGz7RtB4OswWgVkRKAx78sA8C82D9fyM8
DkejZmSr21x3TZ/hCpN/czU//8C5z0nPAN140JuWC5a2pqaLaln65137SZg9txJx
GfG6a4ZpSxYsm4AQr3yzf7+7/WY/Iz5qbUE2pnSY0rV8J8NsmFyJ3je8me1rJgQm
Mj2M3nNm7sH2nCHMYrqlEtVBoXHlp+7NiGLehl2ARva9vdmxdDIu3Bv6NNiIi17e
/K6w9eb0Go+KANtDzKP3rz37rW+JPsfii4+V/+eNIvTQekszk1rFtcItirjIZfT8
G00pxUdX0EsZC2+Iv65ctBn/Y2j0vbK7a5R3RM1TX7qEfWtt9RBbhke1396ISQ8t
9qQEt23rdDOilPqzqcj+VbYlXOoD9nz/LUGtKZp4W1gsTJcRo5FtxUNhqybOjWIj
LLOkOwNHxHS3G1S+H/TitBZnyPmwaj2bssNvkbDsheba0EO/z8EMU+aTOQ4VKSTP
/+cBXcOJ+1mtzV9CT3Wr0gPi2NqS022/Zd6RyJawWGfeJlWUNFOn7BYn5dfM4WE2
HxBdjvya3mhrZFGsxCFDKytMArTu5IaEf9pKcE6YWQqaKgNBwrKe19e5EF2/GsZD
VCxOj7guozXwifQkDmAXU2xcXsksptJFhf7wZF85G9rzO8TyW9V2s0wgIbp5z9ZQ
ATeGbUvZCCyfX+bdsf7HIsysfmpRtpQ7rlneXeVE0TyhprVy7228Ru+X3+4NIqcz
FogMRSDthr7G46jexwrwec/zelFpNKiaFwRPjVn8fUWimPTV8A0LuJyeyaGBIvGT
JvasTexkRIJiOMEF3tFwAoAwFtWAbPZhLnUUknd1n7F8aGghBB/tqNGxq/CrS5yS
vSf+Q2jmTz3s1VceblsWvyaftz+EHZnmNPUABkWgSgXzTRe6mvxc89FwU1v2e9EB
y7TdsDjCCZVKPkOIHeIdFlk5r+Z5T0OM6cIdwYZcaF/lIsapG9ivAeXgmdm5elXH
Vrp5bxeZNywTNtlr/Y6wlCk8nag9ajm1UYqL/SI1l4lz7p7XfR2lpeWwIapaHaSS
TAQ7iJq3RfMv++RSCwknUc7UVZGJBZJvgnhWfpT7fWACU1O4B/VNow7ErDCU1p0u
+jmZ5qHxRG9iJ1fKzjUBOn5I1to/MqS/AelhnJA97Y6GbbKyw91NT3fZsWkhugZI
AO3qbhZlwI2+FDlcH1ln2x2ikbzTyF2Zrv1aHZI/jn/0m+p5zvSnptgz2+WmEIxf
F2oHnepACXmvunrrR8hQtU5hTrrVVmtjO/E+OWuJpbHeGcPAMzqUDX2umUMDG0N0
GGtXRRt2eJzk6UUGl38DZpWlyHT3LF+ClMLaIOZ1RmDaYE+eNdl7OqrpEgi1Xix2
b1aT3Sds+HYJlgctunVyuB3wiL7TASqq+Q17hBHnPjS+ZAw0rDZ9M4Uik0Ij5egA
cEEODGz6ChfPCmhfztyxcHyV2ZyeA97B91U5FyuQV/k4skq5L8PWNXEcCMRqnESP
OIxsPeHg7LLC9RnZMTe39HOdd2eLD7PEmrotU4/33WHFUg+BMxuURsvGVVnSpeLE
jWcrE0pM6Jp4jd1vlRr9ghjZcnVNJaGuXLs6FQyck+U3anljhi1gWFfJSylkP1aN
16svp80iZD1EBTt6GvyQCtq8AT3ziWC7saTzSYOmdgtfuJbqQpIEPSgBHkmW+dE1
XnaT4WdoL6V6jDw6kulx19mp4577shcWwN5pf6W7FHfOvr3JU/3jG6GxU+2tyDwm
L1UpPUvfHZ0m9Y6NWFWch5GS3lrXRtVTl3fBQbnlTL5QOSqIQ7YvOMEWigZx7peT
BE5m/I1F1evkdUmsMAfBxapb2/9rP3IKMqhgRryEGJeabIFTmc23mwKKbd9fNwSZ
cFmGhD2Hh3ZS8CmnTtJsS+7DqleApb25eavPaQhj8Y7CLpRSThVRd8HCzHukOUTh
w6vRFEtCvmY9GHUI+7UPC24CPAzswzAleXqp9GI3wpsztzKNyMUwWoq7ZmIsEGk0
7zCeH+px7bWXl67uye30KZhRxc+EB0aA/1OOfLyv5SpFy8EX75T9U+Ufq/soyY/h
aKegZCVJBAnSB4HnNxLgKql0LovZ/OnRLJTv501JWfuLI+QM1tGC+tD5sONaWVLp
tTr/lgi2FhsI2vuj1cmG1YjH9ve1Ya4RTdkL6sVsAXNBOgipEzmStHWo+JQPSrxg
qLrvi3JWE0KlSrfaR1CWpUSRXPdCfPcjaSN1Oj9i4hRpO3Pw3lKKeT50gkq5tA8N
puCAMUInv4cxmPVqoXVrONODCygCi3XGHQu5PTXnwrvhpMq/6xJkrk3DgtM/sBoN
ZHl7GvItpnSRo2b8Bvq1PFJIpWFLu6jNxsOCebpY6Nq1fUKbtY6qJ8QcT99UaJ8Y
3r2a35QIOY+tF0jaZdGlTdvmIou3vYrKlLdJYYENWsFN2G4J0V6fiYjCAi02zxRX
4w+pS80FsaopQEFt51AvQK8COcXm6rVFNu4hdkx2LBCikyzfkpSH4F4uTwF5FCfL
eL2kbFo8HWQz8FEuHilYCjTSZCe0ylW3qJ6uEW3ahvb1tpgruYBSxpKjOZlXJzOC
YoySQ7/jOvEMXdkJAmH2qGI4H4fpsqXtIqiTnlMtjDxrkLjpgHnqoqxrVXyzMXWz
vMQvUqQz/OFjlTeX12nqZOw4kxbxJxRGKG/Rihe+CFPQ5AMgVZ7kw79ghVlehE9v
IKRKx21NGPVSPqZcBEfpQgKWGUQsv7YNXnIJnfgaXI3rQJIycthvdPGL/BHDgi4J
ZniypyEZtiSsR2u6USNynkuUpyj+79AESW645w+xqhKGNeFwA8qwJb/iG0ex4iHw
Xf8o7kNBA7Y5k7n/gDXLv/tkSAfSXDbmZZFgyz4Yrblfkm+LYf8iOPDXEt8mkBF/
dAXtgXVLC66F6cyyyg+Bk22mq1fovoA7Gw2aA7Vz7YnzglTxQiSzaH/W2VRRPHdu
3eg3FU7l7EwDIMf1dZfIskzEgHQVc4tf8aqZQE2+hxOrg30oanHQYd1IlKNtv/fF
6NrPWnSNh0ts4EelSoTwcRfHk4v7frmZEKXK0whcfc/qi0dLjCh1aRUtqOK5OGrj
HL71X9yY4LNJLo0DsvA8O3MN4oPB65oNlS1t5pROywZzgTnKOJuDxr2Bo/OxdnP9
lSBpM50VXCn92mF0izpolLxLMAnOZeOvk16UFbLbkMK5xx4v5vNeo9Ketbcvgen+
toreFUP4OWfmjJeIyttRewHGIi+YAMG0k/xsLwVDUlyaF08LFrtR6n9OO8qvcBC9
/aBblLWzLxrXA0cL3fTQqji9gdslaQNt82v9zY0ARWaOCzxJXcdJmyPDw7+1yGkA
DwNc1xGdRdOrD2vfk/aUIc/EGX2EPZMHZdQZJkB1MwOzMIhY1js4t3syLR00sx03
JyEigCtqDMu4TU4jz7ElQ9oIvUnj9VBqFo7byiuC0UGqfHH6PBVFzNBVrB44wGLL
OtKXtM+4+VNf21BS0nnPAF7hxGRTQpUgRyKj+rLeIbsxXDJjUkwj6kopLsN70ufX
SRhmRHaW9MzKz3VVRrR8La2TvUG8LMPBbOUsoxeUUW2pr/qn2AMxX9xvglT99GRq
1MHCjVbSeZAZBouyvLFDY13eYzLVXyOHzrRuebFBePSocupq0j9AFtyKDD7mJ7Rf
ydwOJBpglo3fwvV7NhRo6jiJJORih2uTVvgN2RZIySmhgK6v/1nSrcMTJVBvAOJE
nFSaBzM5BVtcU611a3z0Zh7llZiIceJNYpFHvypTTaUU8uWmNm/DRL1DsigyDW1R
myUuIj0AKhgPjs1gwtjt6WRMYrh93OVdcvur8S9gVFFJJ95rgK4F05/n9LCReOm5
tlhj7EOEvHZN57y3cM9/14FCQtKK/Zsg3f6D2BuLFCJ5u0oGzyAZuhnV/9Zhs1MQ
Zq4Lb0Xjezq7oO74cqy8K/bv3HQVtyaBm/5kPJW6jXfsYv/F8CafOFUmm3/olIsn
g/XuZXysfP0NsnsAZSUobISnoIp3wqbwQL2dQvzqlhJPiCQrcb3JvZnrLYrGQngv
zRXD19gYQYKRa8TYvEUOQN63p9xJX+FUEsAZ0qY/dq6inOMH/P9FSIkaIDFEWC85
OzIPsPWWaIJ0hnnJjRnnulxvbcWErVUe+WzK/++OZqekSze9BJHcjqXvCJm1rOOr
IL12cnBYK99EyvZm3bOSO7mhoZCysSWlh5ChhqKZG6k16ligyUfzq3sTGK+FUKX2
sn26zvF3vE6KjC9v1zw4mbWINCXW7aQCp8xKfZ3uBw+roecdxLGCndmhFMcK+WG9
t6HSCaZl2dsGaskHFmgFr17Pw7MDcV4eQBO4JhhosME8wwK+kXLQgUwOvbtP0bh/
3lFcx4sA/bwJiu0XfzmcpXiqXr8hq8LI97Sz+E6zYxaYUPrkkI4AaRNRwAgB/lSq
0YmPX8fAe0TEOLppYXOdvKVc7upCq+9Q4HtGCDrre9TldB7dNzHEi/4sypD5nmfe
ypvnGrI6uM/7/Bhqk+4MSmqOJIgp4iyOYQqSJOoYTej5wbyBzJgF82SMeM/MDQ4o
ahw8ukBCxe9vJ9lcq+Xq0pCm+ALLJ00jOGf7VbxKzsGZnOFoxhxQ+15vg0sCDIFT
CMY7Ggh4pDA3KWFUXRvbsEavWEgdNR5DUBN/zLfVV08Iiy5npPw+rz0Mo3kPS6xJ
G1QJFPR0Ej1bIYD8CbK0e+VEpSllhKObGEfrwfJUIj49zYznBfeX2VnnaBg+avUr
JaCEKX9qWlQz/WXNshKeKFmA97TDtHhyhgffK6sb8O67lzQ/zH62EAErTXvCMDnF
5o1qvSCYCb1IEix/I74wXL1J1fver4oCFSS3pT+tBiQUZSAe70YYD0y/X79Ev7LK
KUuPq37FpMZGrr6exPFMcD0e/cP5xlDB9d/oWMXqNmS4H2Awu2qxKfurgQgCLy8X
7hL6/+W5jT8BdQGiYQ5r+CR3Wt8yn3cMdzDlD1zjjM38w6ZrahljG4h1Z24DFwsY
jWdbUXar336m1B231vgLa6sIn+yFPLvBOZt//gK/QnfSTAhde88yK+udPqHOlM2A
7dPnexZJBOxlxYN0W1Rppm7S1wgww+hnOo2bBW1AbUZBFc6pv7WQmFlvKv+mLkTQ
BpeZC4U3lRh3kJhacHPOP751l4UVJyezAikxO2BVWAhblBWnOs7mHLTNmV/7Wl7/
QDHZdQYIWPzWtgnhMqbSC+txPcoOShqzds4YCVGgbnX26aiFnOrGt5sOECCRWO3L
0NiFmSzGHHddZtQa4RosimPP8f+VAhJ2h7mvnyONxFF6mET7l9KisU8BoZbe2bYb
arAi4IxH+PoDmmTvk5heWxUVf8EJ65oZ7cy7Ko2dT3aaNpiE1kDJlZOFLh2hOz1c
xHoOXXjp0eq167IFVXdWtj8OkCMdCU/1jtGW3RHGC8KEG/Z8GbyNUjLShY5JAAtA
xpqwy7vF09uuPzer4GU3kslp9WXmuVu3hn87UniNj+oE0gBngo1o1q2bfP7ZNMOA
gtb5HgHclcxnCV6p+QaIk3aubfoKlwjNM1RLcwBz3m4TIAYWBCav5pAlL+0uoQnA
XLBz9KcnUEyLyI/zeJrn5WH5dHaiNTs7LHdCM999RdcR3ZwluZjozj0pBKYDVpsh
IzzZhr6zUL73mcr4SZeMcsmPrzg1QQOpJ1+85xTVbWIkJgpBYBJkckBoaWtFT+Xz
0o0eiVvuQszE7/h3jjgCJIPxkMr6/Uc4Eg1FR51QOX8FpkrRnbP7qlc1jYXNai4S
e7EjxUfhHCqa4qBzs6BGiiY3e4Q/UBVqqS3CHJdzQhwo25008rk4R+yYHeW2PQR4
aexA/HKC157BPJI7xCtRVx2kLlNtmh419t4fTh7VcSubADl2lCv9R4tappAQT910
E8X5oxWGLnobeoM0Hxem0e08e2+69+Gayj7aGDMhN+HKRZiRjA9wG6TJNQq/BSgm
aLxtkCzZgAYGyQJ0rH6ofbsJtRpX/ReNOGTvlp29yOwfEFc6NjUL/TgNtOo/DTeB
FK34CwsAv5yovUqzWK6/dJpUIKPPW4Gu2s7pjXODfN3cyEVfbEcHcaD0F1AOR5t6
b6EIGZkksvVzDmHnfxxcCeQzr3XvA5H+XMoXo9Za+L0OotxwVEyrCpxoTlXYHm8Y
1sDh/dGmmTJCvLrNqVeSeGKbNMmi6xdPM3ossYSt8gipMxcMp/EYoqALEqu6q9PT
rv4Dz2rM3a/NC8NQhpNuTbk7OCX+/m4sQz9l0cUaaO/cX97VnTCtW8PRipwSJhyB
eEBVKriu2L/66TLvsE5qpv2Ns6oLCPJ74d+R1ki9a5zRMT6L1M7EN63tkfuXas4V
M0QLHmh9S9fl0JC9Tz3/77u8hiHCxMCvtvkSzYspOrosiHd/gsdcbfjJDnjBWwrd
zNmQe2Diz5VBTU9avmzgJsZw2oZETN/vNL6DBP5ZE36UJc/ZPl6V3zDPPNunWWib
N37iEb0Q+ZBGT+z9feXB2SK8v088hF9lxw/Z9u5HLkKftZzthCe4QYz+4wgzBEFO
6LmbfSc4Nd2+X22oXOGEC7CwqxxFgDQ+eXlCIt/UgZOrBhcVEG9cZtUedlaq5YRk
CDC81E3Hbi93mxyfitBxTEa0E3huUYzpqYf0Q89oglUGh3LicNRV1b6cCi3swRt6
IH9BTidrdi26UZzPh0Czr/2OYykneR93+KRvu4oL2ELz/IrvmmGqDdXXzha5XemK
eziS/3TTV1NwRloAqAgsdwep7DaFe6pJWuUCicN2pVjR3+nqqjPJtBPSxIQ/sxZ6
5lOsw7RMmbJRd/YaPYZOx5LMeXmjY7POi7ds3binSHfa0il7IzeeKDhy5X1z4JuN
M/VPPgZse5qdyIuTNALLiIYrCCxX2iK0fxR1tGKbNguMPT2L3vMr6YE/tLCO+l3E
Kki5SuCEa4vqClmW84i7L799WpO8QFcCrfzxtNzdXsfuAON1gqGJuTMp1etiJKOz
QyIg8jkHEDmMmXYiJQTD+wWL5i1UmiuOeCY1jYZZcw4OusyEJnpDUxMHkjQMomp1
+DEuGaB9ESpUxqqu74f782h3++4PNUXcHuuxdHvH5td7DZkLbi272jfLu3Q3vniv
0saUvrZNOGa89ek0VP/5Jn9Yjd/4bMV8mYrctVtVfOimWV3UP2bxXeIWMV2DnxZR
bYY8UWk8xZDpquEuexPY0XDFnU3LIhuPBX3J37s9vBWyCpeSNSLJnlpy7OS3J7zA
V2etb0kM2wNJAtbuWPmfywtYOA5pfU3pR4NquYQzLEUyMpQHCTb+S/DlOyiX4S89
Ce631x5BKpYLBhjaCpA4n1FKKR4lxJnXnueNpcPjOZjwZ6xqlKorknBtTmlnWgvb
TvS4KjP0Bwvqk79cYRK3LmolS8z5NoKSxeGJ9R9K64G/wsq0Sftc8xoUs6tN+mTJ
IlZbz8hG3VLP4pjZIsz0gqN8gP2sLAGNTdJt3cAHEmPR0KUjRaBq2qNLVE8PHp4h
gYAGL385+1PmDCH9I1i+D4oj6q+5mDkiAEbE3eoQoFjfblrj1Rgp2nnZq9a5nReO
KveqJbGqqd/SNm2VTZIO/cwd4Oz/KGzjBE1lXV38eHux80cT6ofDLDcAIk4J1GJ6
t0bVlrhej/IIWgT8IH82lrp4CPYkL69l1uYpWYfY+pL5zoYOHlQXegIHp1m4Qacl
mdkn2ZOXRKdZx9pbdcCwNw5nfQlIgOhZ25t/T2bQh8RQVjfNIG3Z8wmqnHvRCRnM
6hT0mSCrgcocm3uZKUPIpPVPxtRjDuCIAAN/WybixQ0cnNV6kgXri+Eqe8DLCnoq
0lLDHQYiOq5H/3XEDS2/KfnKKOStfg5qLRdQldjC5diM/42vV9A0Kc9bz321YvAX
A5GhHZdo/kizactVrDgLmUPfRpXDLTrnNgyPBWzfgtXI403MddTZaPw6Q0UiGmGU
NF6qvvqwjrJ3rMvPxoqNCVpHXNhicM0rAVgxrbX6xe7S2YUSC7AQS1J5ERZDz/56
+q+TcNbZ9RsXKshp/j9wRelukcK4mdLVtcfDWSgo5l+LOcIXQa9hTl4lnxEgIJ+Z
NieLqOWUTqPZaxBLyLGU0HO5SJstY55zRGmawoHDv3+dUEc2lHqqRWd4G6PHR4yL
22yTmthM2ljG8S2cQHX3QekN6nMSCIY9VAXlA5gnIiQQuNxNGHD9e+UdJ50EiQwV
RORuUy00uzR4YSXBfpr3CODCXHtb9nEPPl/h+hdl0SCh9dN4dq25TVepUlFkiPxF
xth1vZZUvjPrguKB6waneI+dVIFe+xeBppzAiZO8EHL1hkrq7k4yIqm6s9eWu+XX
7ADPtzKeE9z3zmko30xOad40uBQrgPWCm5v3O9yf7M7avxmsd7tf3ovkAp7OdlIq
eCzztNHHuAD/RbYxXImKYXlN3zSDrg9KS2tpwcIdcvs2Bru7UFF6RImNShRVgj1X
E4E9uL+qpandgduYO+pkGHcm+kwpK8cO1UrzeG7uk3g1y2i8kgs9sFjQ286EZAEt
ymZrpIpE/lWl3RFG4DRok6aJLODhwzQCnRFY5C1Kf6cXc0HR48EvqVGRHtiFEfjJ
1Kz1OpeMk/7dgB7JuZNBgSwHCQ694uN/KqV2JpqaQkI4w5RCHvvavLQeZwXLVI2d
OeIj20oPXUktB/qUITJh5sVvhmOGlOHTghULZTZx/vv34fiB/ZAL1Ihbv0MQMLML
uBAkbyjOASYTiT1YcLTEajHkaYB3rRQtNNPcoI5ZdQGiAkhoue7ZASRVEBM52B4w
ySECjhEc1s6367zromXMpA5jSCQpQ874O9Pz8awAFOKbyedHJ0Rnh4d+yuFxDh9U
F0tcLRbZ82pJJ6hVAAm58Ykd6FESbnIWKtMuyyCU0UUvtabmP1BH0LnI3h9hGxGi
Er+k/eWU+R/7MsWDtMkLqKVDTC9VmQXpVFpUzJIc+HyQSNTVHkPDAlrH+jIGjs/A
NfkoFUr4H67aFun5aaCOsgMAON1+urJec1UsdcATzFWuBuVUi8CXNoq531eCS335
PGT2KotsHJhmcOKITuhuFBS1g5Ku89H/2HpR7J5+amKsgas5EWsbQvw+nnwka6DU
LpYkGJTX9NtRsIGNcHP0NJfShaPVMnd9m4/4aSBCmJQg8FAlbRjMX4rw4QS2T6no
l7+bLlasD1LVBQ8PdM5j5FIE53sZ0Z4F4gBbxN3Wo/0YuvYebSVE6b4Y0n8RRPE4
vQe/XWYvvrihIWQdyiL2HQBdw8nOtBDsSipDNp1hlSD1f1Ow1g9Xb6BYqBNiApei
sUWEN9jW6St8QBBcW97tsy0HdR7KKreI82dUTnil6CMymrDPt/KOFcdOb2bbdYxC
VAqNBQIOEnpGU3Hb/1WccWd2RdIKwZhILKS73zvFmmdgaduEOb/V3dKxf4Qpstew
Hvb867AUizFsAwuMgZLzFI/5uSvgXAeMsqpJOaC1g1NuP1uJw0bpydNYZQTWqVW6
4MvaL+utn+nnI9J6kB6u/CJdXCzEVM/ag1kV4vG2sA1XV5jOsyk6qSb7hnf01kdR
a6vmk7mUHdfmU07XNcxfFEnjnT9wT3c07oXc9mtu3gA1VeJeIFu4976YNCfs/KDn
nI4hhYUhioR6ucJRzc3rrKCeSnIffm6YIm6HqzaPHk1inJPST6AfKXxNie0rM722
c72IeWkQ1mfBP9wCknNwxfn46SaP++KD83DmC6ngdj8KLdf1pt+ZmqCFJbOdjmYT
zdVq8ZFzL5AKuukhFuBrDOznrRFQwtP9AOJBkbBrv32ImDr9C96gEZrq6WjYjPo8
+9q9AWmoAgsBNc2mGanlgo5h84sMyyt+dmW8Hi+mB6jV1IGGOvmqE3SaFr7YNrWZ
PwOVzFlhibbg7YqFVrexHDWdGZMINL1/wkQ+ImWCH3J9sFWdT/0a90dWffTK6GzB
9sEsv8xwWvasy83puH4FS4fNzbfutjVSHx/SC6oljDlrVZjRpAhxNN2WgdVc17lc
bE/4j+0md9pO/t6BMxagWlXNCTpacy5JkVyfStauvPFi5WgN1cxJ+LlBewnKcszB
9w99emG4APjTYylz/Dh+ORkDyQ80yJn7hTZjNU5Il4zGVdTUkIrd/YwJj2sv7iym
2A9QHlurOf2etmvHwa5BmI1ha96AxApMDTBAuN62PHxG/ieBjROhujn0WxbacZj0
ut8PE26jMfvBuYbFNPjtiaL17w9KFycATMOtMBDcdAbMm7r4MU1dlO6FaDX3z+1b
t+gB5Cjrzcroy94+T8oTpOYVMsG7X3TXQdm0LrQOm+Mb6c7Fwie7Cm3NKYlTsmJw
2RU7tf/wZcGb/KfIjz2HPGZqEgZtWNZeoLarhciBwJ1V/OwLU77MgX6EhG8PX1Dg
pVuoVDhQ9Gg5FSG0kwkPEch6HHeer7y/qpQgIK78tiTg8EBSheILt4Xqrt0IgGtT
I8HlcpiuBKiAz4ZbV8akjn6mGzTjKbHRp/YZAICJ2X1+cDKqqSqv/u0j6LyX2kJf
1MLT8Olk4csve2GBwMS+KmKvO1aMUXqTlu1oEnfRYdHh/kPb5KFkBEQ2iMga0POh
25HXoOpk8hUCqoF8/rddvBtavBRwBqQXX6HuKW/Dl3tK0DmIwUbje9GfBSjHguIb
g+45fvofNJOBLvP41W1HpDslPrl1s2t4X4aqN8HAAibgTDhdRqrJMucilfttuaCb
rDRkYSDBQ68n32DisqhW4UMrzLm+ilL8S9KUBZHFfAxTi9WvDPH++Z2BSYg+Ip6U
aawZtCEXsKHdy8+1NIvgLYkgax3JBwavxbag/AIcpxO3RAK/UONcDiZj8BMyAyVn
4gtMsk8ARzbZfOTkmGT7czu3iVWGuHlSzgZQbGhRIedrC0h2WL/BBnftR57HPQoW
blTUJszZWG8xhnLh6PGS9+uv088nmA+5Tba08RyJAvSZ63BzLKVgy4VZye88oEqf
IXSU2viX6U2mFgKk7FTYv5LQRsAInuCukD8Wl66I8BxJgyQUEe+yfhNnXYBH5wtP
smAFPfDgkip66QI+0BhpRZeuxVlIuekJqCDP6BKvcNHePfDzOSs3ujACf05DGKc7
kXLW2k8Kw9aM1lqJeE+jfqHX7lqrCzBsmQE6pxD9F8ji2BWr130r6GSriRDW9yhS
HVRZBoyfbh1Mqbew6JzzpUPnke8j9yPuxDx8LhVmGwW3CldXKxW+ISKoHrBj076Q
8Y2W/sDPt5n5FKJmKfoTq/ugsYUKu2e3JDC3ksAyoNM9JFhVwY2KNssiq7YPrxGj
SlS3OCEvpHjQcXLOYnasDlOfJ2LMwXuFH2tXhczweCfXJbw7FNu4e3UiabT02IW5
IVLnoMe4baP4aRv8Nw4/s6CQXyqbysQMd747Pj+jfWq6Gu+NLXSn2N/D8ofrjqLx
7bS/F+a2z+PcCw96+sr3gWpSQCI1jHZ9+iRWGVFa8jeFHFUivVbYTG+nT9IlkyPf
fRId2keL58kaHy/01GmsFrqpTO0kUGUYtva/xRCsMyt1P4v2jaQhCYZeHREBzAd3
CXY7krO9tNVEDFptWOr1twsZw2f6H4Md4KUdzXJrklMMSee1+e0yAd3FOVbQloJp
e6YxZITX/4nMP6qeJALYAC3Tp7HYa3+gmevgZQAVR8bjVesFTcFVoDIshPFH6JyV
8PakEq9bgyS9acts9MC71egxoTPZi0fa6thMA3QJ6gkmceyHhXuwNnXo9q9EX1UT
gJzW/hMnAXScN49B64BREg==
`protect end_protected