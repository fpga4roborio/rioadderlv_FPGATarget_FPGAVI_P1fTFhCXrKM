`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
ddtXksX2+yylW5zu6QL2Lhnb2d1sD00763mmSITNX595NcHTEkwn0zB1Dry37fOW
FufOhVzEJp80NC5qZ/+F0Vk7Ik02dIR0elf3clrjeJRK85K4e3Hoo4xn7YbFUIms
l/8VZSb14+JVGURjfswrIyCUotIzlzVYZ6gzoZwDXIi5gQIBf/gI+KxNXPaKV+PQ
Ufys/12rjO6aI/pPlqSm0hCvftmBcnezN2hk1UeXgOIuKZnogjOsf0iJVX2aOOWE
6pD/psybjbnsNB6kH5uFTA5frkzIzkzl5d9+YDm9OyC+k84E83I/7/j+rk4L2dah
QJOvksSIzN867/4Qt8qYTQ==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="MvBXkzurAa5VTw+1JJ70nePUfoQXBvZOku/SMmg4TwQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
oRtzZL4VJ4iwysPsC8SXYCzXS8Fw2gtZTOskLcDV+1B9Nzn1zTyNtlo6lNICRmmK
ZRVu2BmCc2G+fmzynYlNTnSa7C0Cuel6FYpxCBlOuk3OF2tzAmLAuDyOH3Z1Yjzk
a0aHuoCdIRKv7BrZCdALt03JeUmXKPdOmIlkVGFl8yw=
`protect rights_digest_method = "sha256"
`protect end_toolblock="Jn9CQpRhJt4rnzZPRk+dOpzAubz7omckX1MrFd4p81o="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 44064 )
`protect data_block
gD6l00tciPUa6pDNTk/+t0OO0nC/UTtBwLB41d4inuAUA3i/ALrNyoJVcBnAmEQW
ptbcNp5fxEUJjnOxnedyZEuEBxWRieZFQnkRdF269oOiu52QN60nM1awZHUGppCN
sNqz6razEfzV49bDMOtBuyRD1Zj10imdc5fLMeeVIEeDeUrqNEacZ81S/1BByoXw
CMQ+/WXkEiXW60YIlO6nAGaIeBf2SHZ/zD5pt/1HKZCmDDQK9jV5Vsg/6YRXKByw
y5rWIQZNmadkSNc2UKO+9OzbcNEF+7yR8JW2f3Mvxl4nPoMZWGZmivWFMGp9YHFu
8L4O3fvXazeW6ETgLHZf3qjiboa7Si9gmjlWCcKutqTPaUbiRUPsIOhMAbSF5Gqk
Hn5lmytFeco+YYBe8zD/4/8wBPqKCEhNs4/kZntDtOwDBCjeS1Q4e3wmvblwAjYq
ZpoZge/8oQOHBpKoetoydsP5ixkN7Zpdroji93az50euWPA55k65pmtC22WB0nkB
pZz8VMrVWg5SKfmRfQl7IWpho5XFf5nJnUuVeg/ysOyAzZBAXRSBzjbHZ+0U2vVq
6YLPBm8tGT/1ds5kp1VZxkwIkV56CxYWZAgiokIp50nzEnnAcDnuQ2HBptyIsiV7
AuHqzaxn9DEfZo2O/qRXjmCvCzuijQWemQIq8YtQPaJIsGGKc2akSzsW6iqjCDNA
EKkcQYl+Pxj/LqVg5SktvfudAt+kaRAVSVh1aZaqZMgy589y63atIdaDZQiWQLr4
JKOMtN2accfGOdsrfqTocAEAe9ZEBWABWW+M87VIa/hchA8CHTTGdZ8bCUtpACh3
9lzUEfJ2IFxlR7RtTKrXcaPADNd9cm/JH+xZjdnv9mEQbjFVBcfC+1j+yM0qMEBZ
GWep1ssyWYgwug9ikhb759dgcBrvrcciYZqErq51/xoLnjBBcRS802dNAFF58vsv
Ehg/dt911Q3S6FpZ/6YPI5WTuLooAiMzoRGRng6VPknWHScbkoMlrCbYnzT3Hg5B
MpJhOLPa8LovpjbkHR7vqeCwfdtcEtvnpFUaWHfdfXFxBUFajRm1tJ8/F7KcaD3d
SGs3u7e1bofbV5cPtOD4kGsnh63eOYmy+m8Z4x0zB3XjCSOZNmKtNx7FKYdxUsG+
BOT/iEDGz9hZ/PY5Oia5m/04ENt3W/yx+D+u0T8Y9tt/p7mKyYEgci91AoOPjSWQ
SIzhPxZroWhnoUaxn5QSP8xqCZ9B3ydzQD4Pk4UWACEPYYw27TX0D3TMGEwI2kss
l/rtGjAAOkFj1diLSIlJLYrQG12lqRS0QJkzT0ZMVyVI5L7uhprhQ0tGHgfWZeTD
OmKxzuPosNpEtzV+fm0REC8fBeRwlRiBeW0UVvtBAOHZk1vx0iaHVWCEhQoLozeF
zbFIdBovX5y2IfVX3KTRnG8vFlJT/vI0xaxNRgsaB7E/Zewz95+MWEeNpYQnMEa4
XBtcQurFIS3lVRVt84AYhB2S4JKZxExM03KAspqYCM/D7az6xBDbBiZMr1le0gxh
rjFGPZLKWJ+vSUt7e3RkUKzZqt2r7PPQQ9Fi0/mXOm6AV+ESd/h7UxK+suwgMiv8
luYrr4guS9lLovwCZD2E7kn3hVixZsD35TVKFadgz6v64NMVuXAJqFf27yedX5o/
Q/IXTmhu0EyrTDHWRNqaqrCZvNJKbUf21nVTjbsEt/4F5i9xwJxJb5rTHyxbozbD
4HN0xQt9O2Sw9gIrdShKijXwk6AWj/iYaHkrcj7oK0wc9MyLYxZd9tzJIKMnTYSO
70KtjhXKrHMD07ghll39KvAMSzHxmbONXQ3iS+KJByUHwSAXYqvBWv7lzteG5vQL
VzayH/NQ5Hi2ZEWtRrJvwzcLhPCJJ6hiZrqEScGOjCp3xH/9H4IdgTeKfNsAa6vv
ozet4p2OlGAB+SzExDrnaeQgfoger6RLKGMDxzAS+pZkyIcR3T6wCsSbOIPLIoaV
roc7cTSsae7kjN2oKuIEJu2H5WJUAp7//rAi+I9uZcmvRY+d5T7j6g38yuidKhI4
gwWXzdwRl+LMhK0NkLhvURHJV8MNjbK+55O/BtRIg7UPZD5sk4VPWuJfTZ7wUTG6
zFGOWs4BHB7nshpHrJI7IIzT7aZ/Wv4/tJcjcwl24jhS1AuDuUVBj5qNm/z8xwK1
KMF+X+oyd4UKo00WH1GF3Y9OetDc3gGNDWn8T3+t6ZGOAeN075GmN0zigFT82j9a
8hBucDEFgKDfj7owbLsESEQG3l4GeGAdUYcK3FEju+rIZEFTkailqvhnneysTpmZ
FkJXJNu4HdouevG6Pi6En1+8G55Fww8Ih7kw5reZnczBdD8plXvqmeum4b68tzE+
ILPlDFg9H9lO86v6zC+ahrSZv4Ku+09+1BoQpEoj1mQvyCaH0014wkkJyLwqej6h
OK8PjvUz7GmQfBWiZu2jXyJhsN2TE5GaYyT0WZKr7vTUa8ma1Scqulvvh747ln92
Dq9E+w97T8g51Rnc3oDHDhFtbZag0ICMm9jVZaryiwNfmnDE5CLJrCEv5GSMoryp
TT0NEdHlLMSUznfrLkgIP7dzt9GlVbo8FrlHJCAljAkQu0H5nLBy4uSzZrT6yaqa
V3JV/LjA7jmsvgfg6qr6iJtdgdKWQ5LAQTDh07CbM4JuhodrvrMTI3Q7extx97AG
4tRE7364T7kwRYarf5ec5mfwpx0UcmIBnTqGhAx2ORAvMeaoWhiMPCmnpUQRHL4c
u2hgBP2IM+udW7aDLUdjbk+MQrZ5TsWF9DVdcwXq0xD7lh3AjLvbhJG+v7OfRGEl
3TDW4xDkXfWyWG2vykDUzaspCU7wKmbDPL1D4+85TR3r801k2NDxoVTlaIQsE+PU
Lu1pGrP8dWUR9sNOtE9cSylPHTiioxNpDGiuIhCgHr5ymtqcz6ywpt/X76H9eie7
cafm/WuS3cWIHly5aoCuzfYxLVKHvyl0+PIbYYBpDc0FHz/pZhGMv0j2vnfawphX
JJCkUv15vePTh4Nsf0ZmxzbnDO9IikEBCR3nLCVfijtlvCjebZBY2+Vf+jMRdDUU
TtR2FU1EyzUoKHNNErL2+mO9sPpF42RmF8BigTKzLgA/rmW1LSj0x5NCB6bFRDYA
Uc/jMit6LF9H/3Bci0oxoWN6VvarxiCUUpMHhzwfIXkuNuiENsiVuAF/4zhVXxH/
B00CD+s0pRIGeRBES6MrpsBGm6Dep8uw5zG/H7k89aygunwU9lD4E6/cq3D6fEUx
Lr5TeTMjuM7jdVJGHVzwIKcZmu2RVcnZJ/g6LhAYt2XlA7aC6v8Onr8dZEE5eMdh
MOWbJsTZ0Vs4KHKamOg3BTpx2o+rW4V/Vr2O9CeVw87O9JZOuzKAzA6PID33bJ7O
0MYs9LQZFSxOeOmWkoAeJd+759XugJcAxHdHLxC8QHNw9/YdO9EukVo7NwyOJZ2f
shL6nB8dtuSUc+LUIcSD0O3WqWj2YyOPhfZitn+7fBTn5aAVMVINtXRdwG2j9tRL
+oPx0A5sw2D+JZDUeQyvKwGsbq5o23lw2JbUJ05B3ON/uRy3vbp+AY0aL6hAMsb/
5lKc48omjSvKPKIcgAClD3p52pM/9itQsdC8LMajvE19yH58g41c/g8uruZ1ttmA
3mEoURuvz4o6zpoImwiGRssLGUAbT/XUj7HYKrr0G/ABa2A9vpBf2KLpPtL9jVZh
Db9pG+5z4oBYV+wAw4+bUQape13T1+0Q3jtDKu8GXPJH+x6BXBUNMZ8dedNdLjnT
+pJhyJ1EVg7J5DUvMAP82FtSL3UI9S6JURoEaymjt2fXRgmHmFzvnWCgo3bKR4Q4
e0X+LIc07nkvGqaqUVQmHO0ttguzANoF0nnMERRYTi+ZIHEXod3No/d+VBkJ29yE
N8TFjDoi4AfqQhJLUdeCE6gbm5+UVUb8QLE7sO9Ry/OEjNWl4JDpKQw1cALmxmHR
RLu59wCYugBm0f9DY9PrN/SWKkITWBK1T65cFcbYHpGzKCG55SDwH7h5ZkWhxrgO
AXFOQDXiCcFYCXxlgrTLnC5j3AFrpAvDs73tHq3ptE4E8SAewgArl4oJ2BHJyWTz
dVIR5E7TjjSnYfNugUN+fTtPQ8R6a/Liyl34rBBvhSxG3xeWbnOULmZHoOi8i727
Mjq/SUMfB4kXr6NmoDxBxGJfRPqPYA101WphX03QkkMUj1tMSo7FMlsjE6r3bK4+
3yECToVbEgJYx7TN0eSSTl3Qh9bN6c2t8mq8LFyRNiLVSunmUMWtdI5RD/hVk+/o
S7usEBxpaMZSlrgDKcIWctDUz99bO7k+a0J804bqgzB0isfoxS4S04u6lfEtMMFV
73V2qr9esWcgho5sLsbwSt9YsY0B/UlWXuySXpAdpNQCLFNMnZw2iAPua32WbxMu
eghCFgyU4hNaQDdtEftOYFJRbYfwgVttrDWLdo2tve0MpIQl0iL4Hpom92xSCs7k
wRVNuP9O5l3HKKWY113XS0XOvVrCNfxe0M/DNySYyefiI+0RQyvlxWxapjY8nyc7
++KvRUeYqj9n3U+gl7k4h38kuaRU6bWk403SBtkqhY4KWDQmdRq9Vy6KQj8LVb3p
p/s6+/cc+/L/E5P7FamqOnf5oZlAV5XhgMsH0Vtj/rsTyUbs2wggRUnwoyRRhgaw
3pUiA6gwNgPHHIp8Skqo3TAFoy0k5fi8d7m0b86VqQn4sRkn1Y95XYoYbSMR1pOe
oRrmhMXS5CGwhFkmphW18/Xv9AjCTZFqhxz35+DYl1376fFNje29E1oIdp3j0dzv
zWDO0iQgEtSdU+m4TtZ9DhRbO3YOyVKCha6ksHFYXzHVjdV1F+fSOjyBY757q6Pf
MZpZklauVijz9LqGAo4WX/qDlanBnwXig/cQrzO3WyB/P7wo9bR5oz2N2XZpinmp
xk3RTNPkmD0aBwiGVsssM0MRwdnZX2ezyBR5OmxAMCPssSsJTmMPql5fiT1tCFK4
eHsb7eYrUg10SYNawaWcgqQEIYh4Vho5e4QLxRI2B+bjW2swdo3/CvK66TpwV8Yg
30aNEvn+I8nONOloQDq6L6hKZIHcNO6yPfCjes5cXa+Lhhk/DuQm6ELhNEOtrQ4k
wiW4dDo8wKXSqD58qvLOweg8e/TpaPifKP6J60Kbwm22kU7cwjH9bEgS3lTljmU4
R9xz6mjv/mhlb8VwPG0UFGINcodY9k7/MpTrWhiKqBf+4php84RXzaCCnmda6Roq
/7eKDbOFErONCvm0NbrHiCp7nEwZHfwIXX8WeEmGqq8ziMAd6JDglZJf59MIkRV/
CfWMREOEx+/KiKvb3ffrONeTiQ9nSd/Oqw2NEPYo+jCFGx37e7OiGDZhedTkAr3u
WmJwrhCEYw5pl8uCoi+W1J+yxi9swQiGU6mY43dCyKVzyf4Ml+PO+LbXInBlwhx/
ceGQavzc4gkQlCIqxEm0s8KGv6UxtQBtUEt49VfikkLVBJ1JGERrfqCv9kowklud
pQ38qDwf6QKbNGC9q9vMe7nxgFpqApMJ482WWiONe4vf9dSEFWPWHq0LR5Y30lSH
Sy9iJi0fF0NId1SgCxxPIwLnBg8Jgv0J0xDirNoHBMDwhHURXqtXLVwHspYNdLdq
cOVT9C5daIfUXvqKZSsrV4yJzYbdt9Ge8b7JOOyQfqAR1BKHLCzS1Yngk7E01hxY
Hv4I9yQ7/2Xuxim1OwxkCyuNeO1C0qtuJ9R36MzT/g+pG263Z/D/vOAS9/h3hnzu
35wTUCy2VY0qmdGqlNfXWksJg17oJVz3oopIHcK565ijOUiH+QqZO14924X9i7qT
DFkTlbzmYAqq7ms1PJ9OqB13uvHNe1KdCuBrrZs0vbNqQ4TPIcLCdcedRT/5tcuk
SDfNTkwQPoHjIkGJSyZsqPfuCHZa2ftwn/EIkKUWbn6SOUPK0u7S2h07t0VHJiod
MMkGWnQhzCFNgmujIamrVq2fbDI64cNx0q9Kv+UzSdCe/e8qGGQHwrUtuq1kntYl
Sai2usO4tLvFM4TmYlzjSBtndQPau0z13FY0EB28AUhgbFNtbagHnwBzDJZ1apU+
pdDUxcd6L1Wh07quds7mULZmSzyH/G8UKar7fmWLZonR2XS1W6jFAwvtsaESb2oH
VE+fAQCXdtGw31aPx4LfzO1MZhXt1XWLTtbYRxSKiY3F0S8GitdBUqsYyv19D7Or
uPiHMEnjx7/QnEHSnr8+GyQD0TZe9SHJ1IInasrzliKUDOAI1j05OdPlLTp0BKSX
3qC5SJlryrmiG3PD6cf1TTjwO3sYwFuPDIuQZNAhuLOvGbntUd6Of6J9mp9Pk4Og
D5YEfOwseQn0R+pw0k5YZmT39kiEAKe7+l8cyRjjf3kaTrsY+g+BW3v6Zt/56sLP
ShPv595h+575xvz0+J5EEtrIEBPB0QN67yPl46r3Hn5qVBA9Txg+ja8Z5sruyrRi
NVXF3QD6lYaHan7+p2UxDDxvwFEFS4qRyAozRgek7se3R/mgnKIGyF6i8qPnExDh
/aLXosAHoaj8/I6ZcwTQp8auNzpvh80Su3OtLhut+Yb6IZRGDoeIkdcO05DqT6Bi
WsD+jP4nt1x7NtORgMfmKLysHc5Lk43x1sgxvdZxXiOlDXRkM2qVQnWJF5wJn4dA
n5lLweLgi8gkqNepfOzUIfgbpTTp8oKUBDAMVU86Wd2Aqycz9NYTVFGOScHzVqhj
ssVnij4+QukKiJTWB1ry/8byxnUN1NuhNnOf1my3ln3zXCa2MYhLct1AEu9jxUj1
cAFARU1vj4ExfEH/5fEgm5Od5ziHneVch/Rq50G2sWUAupxvwfAmI7f0djMFCyN/
211h9/uKkv12QPvyEaFYyGGWccWGqR/9XZM0GeM3HYiLnzRqaesCULlZWEzxnzHo
9sbWS4LCUL1uw6eHCdimiDiz13N+OSyVuaxG9MLz6qxWtNMfj2vmSIvtei08vZL6
kmJNTwRpM7/J57xOdRoClpS0GR6CQkCqq68KH7odb0pUOUDckHZJdza2fLhKs7+Z
bdhsod+YOXB/4ADfHcpZ30+jgAcOsd0Xb8N78TMaFnuTconAvSB+1VbqdK70khzo
d3ooXokdy6cubxsSqtN3WaHXdpY5P34M3bjYUhtNoHxyvbethESjmF5UyO0LggMD
A45QlN7ew8BuRf1Ahf9U6C9OXutTOOmkzLXWSMgZqciSCa18uO/FsC9cRhGXImlc
PtrIL9SchlJps+eW/iXfYjmP00dnRmdbtiFQu89N/wJB8j8k0hHzTaIHxmzU5OYV
cxN/Jn5hzBI+mxUWXWHK2d8W1w2eZAHKH/y6Pu0+qRog49I7h05kkI/ONoEJYZHC
TF+BeKi3W/lYteordnOv/vhXmthnOHC/5wDaF0+jSFbLJNTX3EyXKZiPjKvvJmDl
ytaaYS09BVfefNKvvvkru7phzMhsjRi7d4Zq72KrzBwjfKYsPFJzmDqAlcldA6DD
oM9kZwfupPqFgiVUoDsc2aSOMryAIzl87Ct3U6D6CLtZqnKEtCPtBT1p5DhfwtbR
LFgIsPC6mstHjBMBbV3dI1ytFL6VuGrcNWKrKiqRLmws3czF87Q9eDEpPQBPm3s1
Lwc84e3Hf6t6uaE8UDuVUd50ZACso8I87Z9OIQa9ZV8p4Zm/QJYwQ3zelCZ+hw29
eo7tqHh77oIeR7uykCiccM06rT74tqX0vcq6WyTRWxnsMufVFCz4QnKTDX7djNZg
ABbWHRFTWlXI+a7IJPTfV51egXf2vmFvaeDZSp/LvofRF2MeiGSOQrq2kjtMhFst
luvXFAbYgM132Z25xaAJDv6+iUQ1/MYF11GNeLhk9RDIyhSZvhjXnCsi6YxRmphS
CXCL0BGICy7kdse6WZAvmhk6sa7dodnL6QG8APTETgWmkv76qwlFLdx87kkmrfMF
DxGZq+jBaOF0Ey1ni0DProZXQfo0LPZDyPyFpvSmbdZMwFJHH3A+GkO4eHBVwRlv
LFKFzMFe4EjCDQEwdS3s2k9dNqQqRtNu2WcfMwpbON61V3/Lfje0j8Q+yFiC19Qb
cC6yuANHzjNEV95ksfg+j3eK8T2ZA+Xok1rmHlQuozRcutEN6WagnOlITB2ycBYR
MZ8971jMj0x++aMAA/A0Knt4K/MWEa64PqjrAKJTyzGtI+BmBLmlyR7I9/fDGHrp
ImN0gENMfROxM7t9DhZoAxnznK4yjgbvcRp2LsnJ5TH6MDVLKOJqRVfptxWVDcRc
1cEQHiZQPktM8Su90tomJt3jEj+bMtRG8Op/7BLKQKIA5x2XsniOrZEQ9SDQc+PA
Vo0JpOlYXUe6tP9rgbIOWzGiP9WC4Q1NRtTd1Frr5uRzdO7X119781sAcDgFB1hi
98/1pobYD9qfjvEsa0w7DAi3E9EYbsm1R7hoNp0IPNAScjmgcg7kB8wDDwvoBSAY
c86PMGIbtqmfiEJ9mTGzGgoArFN5Vdpum+tbAmQanNaZ3GYXeYlas4NNa9B+FPkw
NdSDPv/2JPYUupDOH+UCNOmxPdGf0zWFtmgM5nLIEnwdfA8f8b/ZCw0TXPbhM8Ii
3YwK95yTEsRVoQaaUHMBdSTqtBzvWwsnxXwQGzs93P6IcRw93ByIBVrYLd6a4l4K
IG3CRDETGPeaYQSbLiApdwzwT+9UUm0No52j2iyebVshwJ1PVMg977kVBQyvfocD
8FxZVxOcvpbvE1S15zO6uvqeRGHMhlX7idc3VZ7dbVeMJYpqILCmNzgKBQ4VXkl0
yyUHqRRAsvUmQ3ATj2OlVC6FRiBkSgV2CHaLyxiAdom32fAfjN8jPh7eMqkpu3uq
HV/zsCEYIOxJcRw4SDUk8F83AEoObrEPPnSC0/QSbCn/XYiEbnsskTeI0QMHObzc
3TWuQuSqGyUGa8H1Zh8dZrsgla5t4gnAG/xej+DfQ/ISnHdagA0X+BsiVQbTBnmz
SJz66CfYvc9I7YojHVjBX7VQrWpWw10XBhZKUeWY4S+h0pIN0vbnY+aIGjQ2a8Pk
Le6hqtAWHwnZUp6YZK2DgcpXt6yVIEKnGtnQZ+yJQl91v8KbqRdn06Rn+emzCAjl
rh8nntJtoWc0LYthnceGCJ+c1+y7RlJNPLnmfccsZeTMwjLzuhCHUDpocb4vFZgU
2eOX8KE01XajndAkgWoqGcFxW/CWKEghO8vO9INNN62opabtZsUNgrSX6acSX0QC
RqhbM4u2XRCiROrv0qm8OY1ZHC9VMku60UnasL57CzMax9HN4gO5OxpaILLV7G6z
Zi6k0wrrsvJn4qVMxbPt8bG0qVXr42vr+7Hg5/SSIghRnvLfgQ+8IFRxItW/3ixF
1e+WDrah3u2q3z+wxK80uR3MlEHmnJ9DiW3BhoeM81EtdjHrmopZBXSOa16KCOEl
/i9aNUr4vH9DMccj+zZoTwxxSZ+rIMqZyz86nw6/yz9MB2HdnJHzjRui1hT2aZDg
G53Z7syaFv2VxYzYfZTJfuxG0HWmA8luBk2eeqIAWGIDLQ89KxeHOIDh7XQQMUFm
EroEuHsmuTcvxWW9Rprp7VCbmLBRZ1VD269s6rq50QyWS9SHoPo0cbArLa04ABCZ
q6BCMGJ18C+vkvU3WjSRtsANgXqTOJsxHr0vmAy/Mect5S0vf1hcz9mBEr7daUJj
/ai4p9lLA3oe2A5wCVWR7EK0ETPVYv7IQLbk26cLf9q4VQrxSCeC5t5umyllUrTS
Y1dBlC7kZI4Nuz9WybQ5Eebh/BeteabMEiNeJtq6SWkgelVYyApfzrOF+vtUJ+iB
+Ck/OkFmFkQjQAArhSRY+rdhzQvG+ilbnnd94IlwIsE2Y+4HZ/uvdljOzkDkBhJX
tcjg6wbrBF5rVcRqTY36rzVopppZRO7mWztKrsGn1LswJjz89v9MQR1YV+lT/26X
c+q45EMgAFJ1f6Sa4TAC/IVnvw8uFmk+Y/uNktgQPmmaM4YoBwoN8CPiq+21Sq1B
r+HenoOJXwZKGH/odIUMMtbDVY8QlW17HLeeOI2GrWpUIbWofKAK85OJiPe4KAMy
V0vSqo5dMY/utIQ2JzEid/293h4us61lrlaal8j8J104zL5gJm7sFQLYcTg5sTEH
qTxzVyHFvfaotZwZyscQkZHseZ+lzaxo1zmOvkxoBi01B/W5aRw+DA5C1ynjdtu0
FUd9W1559TrT6lPfbi2154rQZkW2vmrYD0aK0cbR0X3SD9hEj7Kz+IPHGr88UKRu
L2THoSL35vhe6IvaQ1NEApE+dLOFSX59jslUlmVPSi7TDnScJN+BO7P9z8IsruP3
Dfa1g1wSMDIkdkm2qFgugGi3M6vX+aKLUq4QO5Rrj3NNR270lZ3tq99p5cZM2wzt
LjTVQXnMbARQ4115A0eYJkCuuDI/AzxNgdgVGwg97uDKxjlcyXIjBk/VDEKqAQro
kxnquCIfLhZjQEwSo++qBjtE9gasEtx0TNHBHDMh8l4dNCLN9r+4VDE///oZeuGy
i7F/bIFgY2TssJu+CIF4+SD1DzpMwCBghUQNOz8Q4Tb9aRoprmM6pNjWaF+Gql9W
GdKUiMlKYx/lS8mbqCUgULO8NDDfpyudYUPOp/bD0yv+9WfOzO7kn23hRIeomRLv
01oYWSwATotbKjVyknkVkhWAikDrgcSgwsV1yU4VC/b78JZAA07umQQ3KSekcMlc
RFTZfxXSfxTMOijYFNY48MA66pdsIEyA++8uWkD8is79Vglza/TnVNhUEYxfS1MQ
ISfW3BTXLoc1t3B6tHB72AUVYYVy/aZa6Cn6+Of7OhU/RpPgXbytoX2qu3Ek5QSE
a5gQxm+2nlkrrTHwdkRjNVIH9WQtIdGfmeblaFE5PIk98pFibH6cCO04qKcBIdzO
+QDAqFSZCG86kRhHM+/cqPn/BNj3wQNc3cRX2JIgA5/5rKwwxVyLXprDtKnYPXIw
JLJQglxgD9LCie+UNTDM/e37QdQ/8h2+TcZrKnlXRSNl23OSuzJGRBFuf158jmSS
Iv+osj11HIr1orjSt8Xptwm3ZvnjtzEWGBmVuCkr/nTswHk8ApquSRWXG18px2zY
M5FFSKFZ4ikf8yo7DzBh618wDAPMtM5yx94h10K5CTiof4HZ+MdD69DpB+XML2Ht
LkWmLDtPvwHfh6XQTT89tB62o8ZpEo9dZXep+0wCIbNNePbAMGaC+jHEgAEygfcz
yAFa/9XAYwK0lmhC1h4l/Q1r/e/Yr2+h6jvpCUfwUv79gEl4WZWZz3+Mrpc47gt4
uW2D2D1t4SLPy+Y7/ErdEoabw7XIjWlO4rw5lW2EzYWD57kST9OzMiBrq/JifTsn
u75McWLGhniUDdbvbqUeczp1MCUamIkMPAIPeaYWs+XPwfN1c9nWqkvAJG7O3srB
J7wuHJXlKZ8OK59Fu1proM1wB5ir667Zjyr/27jzK/wxZzYiINO+TUZ74HZLVlCG
mv4zRCr5Q7WTCCyjNgk1vic2WKn+KNmkP/C5/XkN1HZ8S/D9zJaC9mVFIFkG+Wag
IV+uRbmkhMoNSYwoGuebwmYADUV7Mh+dNfE7GDWtRAvOrreVrIUPaHFBU+H6TrUI
QChJmDNtLqw8dGoVFREjKYfn9gsNVRSTd8tBqaovNVlG7b/DI7XBXMivXRRZiHZ0
jbkdQA3nv/fJxJfei/4vrOCyr3eBTCwtyH6YCYxmZBiZ6TwpAGCYwdoXQVAwBvcE
hO9XsmhKmJqiRVSCWdqoerHV8wEbT+ET+rIWnTHm0m13QTw5NvRKxtKBQNCKvNvH
mMuqQJFMGGIxAsq3531kSQCRwENlRgqWQZ+ABdqSZFOeJTB8LAwdxEHWtlJtmNAQ
IUIF6SbY05FZ0AJECAmMEcUA09+jld0Dx3rdFXZaeynI7do2ELaX93Z4MLvz2JGJ
0cDBJrVRa0+zZoMyYafd1Y9I3fj248k14nMbpHqPPK8qEQ3DC0aogT6DQLRB7pBt
6YoI/foXlm1iwMrsUgDcgarz/R45i+AvQ4IBij6UtIZBVGpbuIcITotE/xSI/Nqf
37lP9ffLsF9E60vRu67PZe7f8jWM08peVwDSOdr15CgYcZdt6UWqUcsXa6iNM9W2
F20mc1WYK1ZkDpScEi5YBY+EQOq6wyuTLmVPkY5ib4vmqhqfHydxpytWndyTRJFh
y8sDvS3FsYfGg+xVqIkVUTsd7F8CrUqBNFcW10eFQ7eNRj9ZqH/E0kmKqC11j2dU
3roOCBHIGsAf8Crw0PvW/IilkcZY6LBBWarbfFxA5lRqmo9JeidwPEyLjERGkHhp
MBKSVE0/K5ua99gpVLeaMbUl+FeUDYHXQ/1qubpEljAXcE5RcZuRnCazl6aRtaIA
yqOj++gIOAdlauU/OdiwpSDwUwr59BJIP7G7c9adqHW9y9UfiVVJJr4yHw1dK6ec
9syoAQyMuvP6OxiKK6t1IQHiNJVwYJi+psR7yTUcwOWVEUAgimsYmvYXiqu+lZ4G
UAZ7+YsLWR6Yl4JNneMKQHIEBJ5Lamh/q3VRqgUSxFJAojkgj7xLqqkPh2ljPQvZ
cKq/AVDdC/JsqAk288W0sLTuUar/549QZre4empMogoZSn2/8Msd2AFwJSnwu0YY
zhyODFwjRG4InTbU/bZJumr+etF0WNcTER6ACcFGMRYH8CBJLjsSIDzaaYvK53JR
8r53fBLbl1pExH8HX0rRyCWuY8r53x+wWYs3EODBeNX8MqWmi//wJfN142w/r4vG
dF2O2lBqY8CvA9nnRs8TSRAHCzteQsaJtJoGV2GSqbtN12wgvY6ZluV6wepKYK44
JVPBOsrGwoBHSogwVSx34yagAHt0fcq6jjJyMoWHTdBgf5Ps8U/dKtGnJvLHx8Y/
rn8DoOQRWsw50O1BDd1DJ9x/2zcP9+efm9YsAxEp4/JSMLZF6tBEWRfGTN1Y/6Kk
eQPxHPM0aFnxlfG5vSHj1qESDBLUZIGcd7M5nnKi6p/lTBfqA7FrtCGdxj1v9lRJ
zgtwG+cpXxCnu4u7a39WQk+/LTLI+y7EdklWqZBrAUI0bp5mMHn8YsKM7Pkb5yWy
GbVQokPCuNXaRsEm1uhpCdmHncxH1psP5B00JMdfyTd/UNPOI9kwb5Sjkd4mEIZe
D45f4GZW+nCME8/B7CVS+lvIJOAEI7sRmZMnczLKdNtOvEh6LUWxFLkTf7TJrQog
Ye8HHrAmbZBPqtmW7DNsS2MVBGTcSnEu2/JtmtRlHy2LxScokepOcYbGd5RiPFl1
FFIr/51cjnffOVVAkVbCTesqSQtx89ZczHEVfadud9DVvJMsup7w/RhcQwf5fEE2
CLAuI2uEtf/ktryS+8ASWla9v8fYMMy18CoQYgLKWZEXsetL1dO51kqUOks2xyD+
mMumeTBnjEBuwuXMqL5asWr5qN1oQIX5F7d4dt8hcJAfINqX+lnyU1z4UZF6xtSZ
ktC3af8hZqAc7DW8wpyM1Dh2YcRJdEnKsvDbvIHuwsWVPFS3lCiwWpMvh2HRYBWg
jeO4e6PbJi1LrXY1LDJHzDa7Z46Z4EkCqSS9bhEWFKhgEehcsiDxyis6eghhDBNJ
Hy3sann477X0c+LnTO8FzZrgTv1wJ8dKL8eBB+3XE6sDELmo3d4Cy3ivDHSXJwCm
h8ia9lG4FikLe8k0IOIePBrj4d9Rz8O5DoMw0TcewCDvQCmWj0crL+fA7blwtKUA
gwSEFwEOqKR65mcbI2yeTq/0Mym8QoBHiOVp6juDX6X0LLJJq5TCC8tADR+sNa1z
hWqaJO2sPTvguXw8xd8fw0qtPIH5CqE49wggnWD1Nwa/+tw60ggtowhv6BwM0k4g
KdcuUs5W4an5NCR9XL4INIu3GAO1bxiZuLSCBDdpUe3i6z09dKyctTI7Gp6+F24s
5AEV9A7trWgNWEArqc+8IYXA1drBzZCxbw0TXfWj7JlHeVQsMsyHvoR1TGVBGjZ6
lut3Olk8nEIw5VadQQ12Aiy9BLA0iWasUxh2L1J9NdEodgzVucJz7kIOg7Gio1FB
AlFeRjwSR5czRMpF5X+MGDHKRmtOHez3TNtcLIA4X8z6Eo24W4QkhTZDTE/nddv0
MqSj8ydQrzv50LZit2WaczDIvhlteo5z9B5Shlp2OJ478+B6ygovNPkdL54LVG6E
Eg0dl32oknPL1JwFXK37rTIF3nxi6FiqgJ/DmRxwVDAtkbMNgjw2cVr5oSrAJ/Zo
zmG7+SmbHB2E1dpSjR8OX/ncoXdPKZheBHb8SPY283jkXaiV1lDMJEOGdK3MbyCP
hlQp4DCEE5/IPoV0VUuJ0JP37/nETMmV0zsDNBZAbZqMgZAGQIEpYdtFvQk+lxPS
gJc+JnYELiU3BKveFWcQlyta/WuU+eTehBvCVc7PT9fVVjL15Qy5ezwfwGtxUagb
RfWXq0zdwFLhrzAMD3LI3Gdc6Xp/jtGHsB2encgJK6NYgEFQyBtV1VQyujWGODsy
PqVbRq+J+12PO9m3LG+DInsvfHY4MbGa6Qe5dz5dG73UzxMQhq2JfJGObt2STGg1
2ityNNUzVCiJxjRYaiZJhXoGtq2uvqf8o0qlightV+cRGe142i6hHqdivUMTw46Q
sH7aCK3wV5KUr3x32NriRRPkPvSrEzzEAZXYZjkp2v/BHFR/avJG4kzw+hsMm/vZ
36oGAi4RgEYLmEg9qymSmhBi6NNlejoB+CCHW8YlTCqoaeI1tJrzV4pXXUorSSOK
Vc4Pj9OK1jFtIj1sVSJsmayGAgSvJQkPsUxPHCFm/ydDzpmxhoJ6xadhTTpiuU9S
TmOagcS49j2OwJp4f6BkS5PzyvAzhf193sDCKaPrTaBZM47wxgjp1HHlrMiZXM/6
eGj7o54RBrB+uwpKDlQcWnL3TkgUSNa+DaK13Cx7dEGFXE7HprKM8n24H4Jo4hbb
E08j9KTgoaccKEHRJ7GR9A/2nJ/riH+OLuuuUWCFFCJCfZt7UHsz+2St7Zcb1Q/t
5Jumk0rLNfyWkoyyqIDmW7HjkGBi3osJtZVg+/cI2Uh/M0KvjoTo9Obz74NkWZKl
JoRrMWlXs7TnYjc5L6GjdxZrXiuchIxLu8N60/y65xoSZw+/GE76y8OfW+8Ks9D2
MqQjfefGGuSuSngfj1rLK4i2XK4lA6EZEoFfnnOmU2kOdOaTJJs1dmu8hG/teLI7
SFiikK7V/iMkgMNYPKIXty3wWnGZqf1CalRvUqUmD8TQ2TLbVwNGpCKcysr4IKsp
u9YBoAkYLUftPQXSlWBYI+exsMZwstnNkI32HEEXWYq8HFmd6++U6hQgGTDUKfci
vxM6U/1zEEaxGCmYf2wSvFOicxOWLAiu9WRJetOy3/oAeMkFH2JW2fHIeY9Qu6wF
zNIlDXyrKSM9ZOkNlQwzrwwCK0qjUYb8kIz3tar57IU6EIUogtHSF9a5tuyOok8G
OBuQThojj+qdrMDjJg+3QHedGLE5cr1eBJHKIxoQrmRwfpYev6Nr2/aLOqGw3vVr
+r+24u19wAARh5Eu9tx+Stuvm+ZsLOvb8xoaw+Gvn1NzbmSPKUNUec7RokO7YYtg
VO9EVvAB7BMgpVxsw2fh8HATFWjMWFwYRycJYriIDi2L30XAJyBpwE0yNNi7igS0
hUocpAmTS5eLv4RyFV05mLKysXV1dkpk8NN+DKMlR92SbUw9DE7TB9fNCetwbqFD
APxfS2/3/JDhYXPziNGXPQ1tXXxOeXmt6o6ghN7ddSDD7h/cQoTk6NAtAqUXI5Bv
imIuHzLIUqiP37QueLqENaCLfTmqWD/o9+mL5tLthxOy/e5ValVc5mLa5FGDi27Z
a7k4BpAYjhJg744ahXrNOrU7DHnspBL0/0n14xzeOgJ/hMCUCvIrOFzNFtk1YM0T
S9QTP/oD1uxp6QiDL/EOjgqISuDcPQPJWsU8oun9RxlfJrQR7dYn2qoykH4NMaYY
ffqN5B1x/qh9feWgMxW/CoQ9DpQuOZhXRau0bTFrqwu0KfJ9u8W8JOe6x8Wgfhxx
ym4zDs+2hCYeDl7dgGRb3miaDFsOkdAge6+6E4RYRwnMGjH/kqacpxKKz2mkPmt2
F2kFxdNjLLjAqE1o96eyTmiFwzh2aI1zYR5OdWEKZMPwMnc08eHWQhbkl6ekFT8w
EztPTGZMDzQ3g9f0uQr9dlGYnup9MAgzTEp7MNaRPGqYos3+kU5vPPWJDbcCq69s
+iNQgM0slKCIX6V0Zlxp41ydAFlS2XJIgxeNrSmnf9mzjUeg4K9DEpxw/UG5jaUb
z5vodAmvY+Xk1735D6v7UAVarrS+qVOYxfm2uEZpA+7p9PpB2YEgrNohN1v0Lpjh
ysSF8w+16KrcOJa7m7JXB4Dyn4/nJb9ctbc17eMgUIMT3wfsDhd54C8EQuUZWxRi
uCJ7uqCj5t1oajuGeX8Ia9UukeLbq2+kTF36xOl7TsVqBMlE6hwO/8d+vdziPSzR
GrOwZaH/z3DQp00/la1tChfGa9Yds7HgQNrhdVN1uCs3WMRMqCoJoQPPUqw2xmCF
fnSL4jw1rvSxuJasveo2mBAQsIFf/azZOAK9rqJXrg5oEjDatDef+rLFWVyBZJ0W
K7B3manSlSAwcW3m4LcjUIlkc/ODn7gu2V+BN4qxRc1HvRt2h8psiyHsDwSPGMpP
6dCKQaO/CM/n/x+N1PGcZwo9HE5gTy8Xw2L28eQJfuUFI58+M3PMqdeUiXIvofnl
ItTMj5SoVSTK43zCsO7gNvyxlUWjDcxltr4wu6I98exqkM09mp6hbcDx1JoIHMx3
UisD19bqxPiBkRM9ttE3UpS4OfWy2UehI2jD6BrjATgo0W0Ra5MvEd1+7lXdpL/4
DvVkwQRFG6nzOxkl1yz/w8VJssbKrAwdO2J5hnJzV/b+Ka/u4880I3JrUc0wz4FA
RYtNyIpMCx+kMzIHB231AZ3RD19b+yrGefRXA8M0Ov7/aN0TN55OzRiG4MN2Q675
vtcoy4aCnskcvnIMHJxtP0WE1Y6+Lalu6uRbg2EmQwJLKsKxWlzNPMR3HTIBgwif
Jt5o6rYa0/Uco4rqcHfiJRuiekChP5002pgtoGjuKJdaTAvuiZmz1LIbuwy2o1tY
sH8dpn54VaQiwCLP1HaDudxh3eJbW+hWr8n+A7fIUCnNSX2IWQZOXyuDaSYiZQmP
JdnLBBCOksPwwl6VkwdPZuFqzzfW795ItWE5XWtWkE/fCuM29gUeHT/zUhoTdAFl
4OGm3dU+XFntfHowSfKiFXLbp3E5yepcl6jEiZB57+HSHqN8N19gQJTAmFZ43810
RZmTWVLtUIBfFrEQ5+KyxAxepaTn7b8qkvdP7beGR4TlGYXJAYrpJE5VZBR9CGz0
Ng6wmzRDBhSO/MDaPN0neFHKlzQSj/idmMbASEZYprxg4gL7tMpeaDYSXtFWiTnx
Z0uKJRYzl2p4ybNRS5VVHWFwkIiPNmxCCLTgPQI6njcCdmdnoj+caEbULPA8Y4CA
iRdpuuD/B1bL34yC79X9h9hC6tftW7SH95fmpUoX+5uXTHF5xq6U87nYaONXoG+x
rjJopCeLUZFR1KEzxcGVuH4DZlaNx/zH3JJ/Pp5ZTZdJkXW5c+C6hPQ5nN8H7LAv
xvpvbYRf8IQJ+aQ/Dfuzv81hRNISk8jZ7vk6ong3tSczBS9HKpHDzLCbyyymoqbk
3PKMnPxUND4tpc8329lzxN2M1k0UZk2ImSQdFKZbIUb1j135pn7Ii9TMuTvWHmgS
Y9bOzSit3lDdNFgxFOxqG5UJDz5CBFKW/68Ad2zSSu88I+4WFxRreHTR/rlrLDo6
tygrHp5nbLB57cP0M/Of8PagBFYXu0K7o/Kg1i9HsHzSEl9i+mRMyro6kfFU5G62
hEVCoIQAmVOuon3OovRVp7JRYo9OCR+BS1WEA/cGFlWu5N8EjYQ54snoJdxBEM4b
idkdAoeK3FjbitVQBXbWtEUVaxzw+cnzsSvFrFtK0ymEiZuP/PGUFloSmUuhkktZ
I5yVgzQvcVfqJsqozz3iOlfsNZkFjNWdgnsZHJmp9o/ihi+8VNBDVkMjVQEvqqfi
m6N8qB5pPxvqrzzbkDK3kZqwZ+ZOgFENUwRYtB5AQENs2HPTUzyLN00j9UB0KaTk
eqQ2/s+P7lZEDsNaq339YiXu2AmD3f6O67sRqHvieITb12Pm+xoHoACv7k7tkgaU
UJvUhgesJu0ZGbnv+MInYe7NpIpT9bHru5clXWx4FQTjwfi2XIbBuLjmcKeX2AzA
kqwuvLsz+CpIodDNIyDnSW1wWKggPlta9N1qfAWTVA9x4lQk3AHM+EsXf0NlF6Sq
JzUjLiCq5jLohGmIEV/AmtYJ20iTvhI3FaEquo6wA/TBBuxNvFL1T33ttB9qzthQ
6+SmFQfgBR+bf1tviBXMAigtu58FoPSuayhgJUABNsDJq2hpMbww3pX9d9P7ikiI
W3TdiiutLG5hgLd3PaqgMJnTIb0mQtjnfFPaHQqKuwFD3pZjka+Q6xUfzWz4qwai
5h0e3gAuxe+spRjdFbpDKtQvPpvKQR41Bj0jY++y3u1UWpKz4fVRrl818HVsT7WT
/NHTIkeILUk8J7y85S6Z9Bas5jPCZpgGXqz1VLeYIabOJcBxHRxUzp5aoXAvwxfX
uRJJuEqipjtnhFgCHxZzHEDvhQl2NYd7aAJUZSX12PSZ/3Y5OdLFcvmujMuvkSQ4
gjgTapy4ZB+H+y7FKb2PdwflmJ8gM9cdZSPu94J6o9P8iPz7sFglZsxg9CJ7cApN
VPZQxP6akhzkvOC/9feFeyvSuIOlO9PWv1XbFx5drGsIPfalsJa0+6eQfMnMQLtt
TyRRadOw/DelGuwskKJ2iOU+K95FQ0bHgFY/s5sE61isyM2SP/xBiytXmvj0+3Fm
XMjENHnOXv7OQvWDpFJeWHLUpD65N6QVfYTf8TavztDO7XORrUz2hb6CxId1jabT
FBdJwP/6VwktMN+NGQ/wRD4Ec6JFFoKoHqOOYOcYG2UuKUKkdx4HvnaaAHZRCP4h
XlUEr1wKhY3WuJm8JNBHeXq3RscnG/mGfwoED5FcSGU066kZg/u+eegVFdY7JvFW
j6jsqX3Dyio6UijayqjRjBd1wCYNthqjawFpsByhxuRrH0IhukE7NumIuHW+rIPO
HbtctFQtYfB12W6iwyEJSx/4iL/srtsLvqd1n/0FizztgkE3zIMamNFWOW1JjL1y
LvIjYLk1abi0Ti5rMULgGsU3qq1kWeRTgev3yWtChMsj2F6FDOApYuvZriQRgRZm
8gxNw/cclaj1P1qul6edk7yrfL5/S0V5IM9xfKkWNpbGK+AjkYXOv7fs9U01P7tk
UeRGz6HPYQnPGgHbQz257/uvmhSVHUaLlCaaOV4j9LCby7m971FKRXM+7lZDiMkW
y9S92p0MeGqVWP4JoYXM2DaQvfGRKNJHnAbENJUEOqHEi399zP07On/EtCDEp/9w
W++WmZkEircWMNI1McU47CxWe48gzyOd6VIXWS2nfwyJ+KHoLAp4wH2+erDwQ5gF
4TA/J9VigQMFNAqkwUlmrpKrWaQkRZDck2VZpEDIbKmpZ20FOKqxL2VLfmNRCrYF
B/ewNhZTqTaIoVH4fHxyeTDjcz6VlfrZgnBTHF3bvkhryNKWjQY6lYzaNZs2U+fF
gdZPW3TKhNdFmSC0eXnH74u3psHwLkxPhpMNcvEUYotzxOAAP9eK3j8yK3BLRw30
Wd205mm7OCV3GnmtKJerIBrOsS8AzUZjkyedwMTGKVD7u5nPOeDqJHowXP0z1hiR
JAYm9SMcAEhxRS0AxHaS7ZfIFSJ/tgxV5a5JLZo4su1NJfp4yAL//muejUVOa7L7
7tEP0im6erilzhQYqnKg9KTyqsbrt1OtOmROIFNmF6KRKAVOyERQ2ilNiecNXyP2
moTf8lKo/gH8hvLwzPJF6OoM5cQAJDFamNkIiRpHg06NhqH7v1GCeP8aNo952TLU
CPUGwi11H12hcII5B7uohTEzqvut+TPVep3jT8Lb+QZg+EA77z0KTzllPjSfQFJi
qo1U0LAZWt13eOW0pC/3/Cy+Pn8fgNiaEGih+g1ACgcQMPXlDeP3Ct3CEW57A+ug
qjjbp7r/NawbZ8x3/Es42YeFdTUwdifeueqTsMZeQv80kL/6PBcRhjRPT8cDFs5s
VwuTrnxds1rJUbnc/+h09A5HS+xYVqGNuTNuYpTORYeWyY4rsxKYnOh+vBNwOo6i
qi4HXIcMEDxhfz7CmJ2C5orxF9snED/DIGLK9yumFBnRBKwD1gPRZ57Cjo3KA7S/
gRnz40D5Ju4fcPbMZ2x9Qa/Flaf/6FJAZmi8Bj9oqC/SqchG7Y2LEDbhr4P+BEUn
7ssr2YJVAbiHoD3/MDjmXvQvfsETiV7pOKwnutJakJJJVyefl7vOnDN2LQftY8IT
Hxj7Syf2RoZdxg+7WKPe6q9B3v6IfXCU+eF/US/LGHZfK7yJoQ+RNO/6oSYy+GfN
TtEJr4gTuv4yWiC1k2Uc1kjZJnO/91UPU7xk5C9PEFQvt/2cfZDKvVd64OlzigY4
ie4k7PMSVcMkegoGPxcSl3v2IBepP4aGXlJfQ6MPHUQFWcTrHFGU1nDGOxdh9bK9
V75YjB+qnoqX62XA6XXA2uW0v76JOhuaEgQoA8hK4J0X26hHOr9ppTplGbNF4BmG
n1Z6ojI2L3yhpFDI90CrMt/kHiHvliXkj7aNC7yB8iB8mnnBIiHQVunI5ZZQpHEf
SM1aEuvM9RPEBAKAU191TDLtZAkIMxCuu+RjxNkAyP/4mbiWvVnqwbntCLqRX2Jx
/H53G3MFuUPeSiFyU8pitdO917wWmH2UZx1zAPtTgkEbxjh9wEL2+/+oSpd2YV0N
ELMTaAdQB//5QUrFCmkbKlH7OxdszWMcF8bjXdI7CLBI8oqwzDiaO+x+5xgYXTGz
l0oKm1i+ElNCI9PTJSE+X0o2Vs3AjqY2pi/Dc/Tsy2MFaPQf0/GtdETyWBr3CMf1
twn9ZwtHh2Hu+gk/aBP7DlCMisDieDZSugGfxXLq4uUZkTC5QjIScnhamK58vKw/
WpFZ5+O6hrd0capa0k0l3QtnvmRS+41CtmSVsE03A+9p5VJGdEhu1B2UQ5kggeBu
IEKBEOSujwxv6UHdu3X5q9jNhkelW6N3IuB7ja8DYd3xdfF6DV6E/FV+gHuZEtgr
JYaKQ6ea96qszzfHHJKVTqF4zNOU+N7mkgEAR9ScPFKBbVfoazjA8Wf5Klhi3f+6
PT+w5f1HvrhjPMznJCVaoUkdQfUMD1azdFsoq/faj9wA0kzVPiJo5I09SBMO++5Y
AtX4GGofaxMbZ0B3FGye+RRvJ7ly9f/ErwmIU4/A7KmxMLShy+BjxJlTQvdai5wL
iSFDknCfz0kQXfj1KXoLk/0Un8pfyHwqCF6f0aro9YkPq4m4m55eE0jRqQdDzVK7
uQw17r7BrsiSR5cY2oBFjfwyvzmChpZlMB8j/VZ/mNUxhv6QIHSAql+fnmPWhjLU
OFoBynYgazIEaEcMMF/bMDv5GRGt/R3v4kf5trJoLNLhnca7AK/WN8eEuJpkdv9m
2FnAqbfkQBgWdfv7kwIb8GWSItsz3GT3nGeg3YjVBaeziU1198aJiV/LsnwaShLc
9ibR6ApzzaSK5WllPsKWmtm1JCdm1toJxdiIb4c5W6ez06dd4rI/cV6F/8veBVL7
6l1ue6IPRA3XP4H8DbtZBCrDjdp9soWZ2FezBMYzPkpNRfvMnjB6kA379eNmhx5o
I6ID/vFv4BSOcz89tx5mbYURmdpmtcFXaRsU2d1hScKAW1Z7s1Q1nc06C/YniOZ2
UdSN6PpfCR1SWQOCGKn2J+Tx17DSTW523PoLRj+/Qwlh6XzO4jq49YbN14z8X/Qn
HS2kt/6Ey++/9gjqzcs0ywD8J87KZx3EoybEi/api05KirthFAFzKmwx5eANANfP
Rpna/9ddSUwe0Q6KOQi7HtAqINrL5O8CmifC+MXnEexTA2PruS1lEk+CjSDvBq7L
fPaIIzC7JerEMPc4Soyd9YLuQp+sv27d52G/JTRpHCkFV7R0MXqDbaiKQCOSyX3q
ZqKjDeJvUHjFwdOhkS/PXe4C9EpOTXhqOPeGPAoWYCRnxuA3sS7mg/+xaER28rzB
htDfYVm2u+T6FAsYQh8furaUJvAQqOqy8oEMWly0HC+X0oIIYPtyQt/pY7/N1tEj
vy9MoObU34YsAwyx4GYPKQK8XJ+a1kNs++hT4ifg5qp6e0/0fao0mr9tgq8grObr
aVdjBhju3SDoi4KTwyihB5yN3n5QGwrF0OTv5jiVB2L9YrpgJG4Tob0UZWlOaeZb
rzp5vDf+J0WL1yVd4OUouwfqvcQ48qeaTtGB6otfkHwgOw5ZfiidPS5o/mt+PMXc
qgFpEjwlKwJe66C1tpvf6m2Wxi/EXpG0TMyixNiB0Ium2XIgkiPuFq3vpzksc9T9
TM3hojHQPcsAiaTczWnStdFtr51UlVg0hdaa6dz+QA30Rtcl5leAAUWaWYkqvaa5
MOYLx6mdiSRuST6uXnsvq5zLHFw9a4yAVkBbqsEclkNPP4e1lQgsray5Lou3NXg2
jONI/m+hBV0tDbEzZh/Sb8v4CPJVNWq6Xa1zF2OdnZ1g7IspYpLUj+sCIGMX1fQn
U2nOpfYilZ2FMNsEXunkV/wBG4ATY807NLXQZuDqPFngI+7ymQESZKZGNgcD1/Ji
CxXoGvtPozqxFvvqp6tGSsW/JmRljBKU4gXikWINc91lBoPkLjwlMoaNTbIU7YgR
rc38uRBR8Rlu0WuJ5qNlC0kpAeUC6drXc7GGJhZPYG0mmkJyxzFXAT/jnXIt47+K
TJwQGe9gArBYs48MEWHr2+RzMDKZxcVH/RmYQK61+UaixeNGRsqsmW8FIzbrLwZQ
R+uhFTCNTE9aHUvyT9AKzXbjDl35+W72fJkjpiQ2ndz7IfIDgitA+YFC2HcA0K27
dgmYYUOb0PUI8Tbd3SxhpOm8ziRgg4xtumi+I28trgzX3pp7QwNYtxqofMxcCDF7
qBc4iaZwkLn+8cORDWVExARYx/eEzB8e8PaH8cw6sPv+FqmPLCsCbPfCHo3NJzPo
A0BQqNTbA4k6V5oUNG0M+iP0uKAJ/KwgVV51MPJuvMhUKEi+fpcx9ytrI+e7+RsY
PhOdEjGr68rGe05mnBqszx6S64nO3pOx2KqjbCYp9bfath9ULES1Usnwv4B7g7Ub
IpnKlmeo6so6Gw4zsaI/rkPzIc/zJ9Cw4a6bd+JU3Shn/E4Ov5ha9z6qHjJSuEx/
motIFGnitD/FTfzkbGg4vkZzfwLEQXipT6QqCVqZIjTur3Tciuj9BcoMlXXEDOIE
DUyYw3F346KTYihLH0GPIqk04Gkt9FL7soS5gSLR57IJYqNEWN30pxknhBIGTPF9
RjRp7hOcnVw58xiN8xwf3K6QBlPLzUZlSibSiFdKSwAtzC3sxk8ZFeARDCabmNrl
YJC2gj5a0sjRkpnqPamwE9S5goxg0GfoiXXgbI/1LDFFOC+WGMquUEpVycWbUVSD
JxMFDoI/grnxVH8nFtyQ2YBzpsyUn4N3Z5qwk/+HHTZ+ByJ6jw0Zx1Q4WlTNfWOi
fOm43NJpJtPVx3NQjLk5EUfmS02SJHNvI00TUU2GVuJ30Az3K3tQom5efGGHs4IJ
VDAky7vZF+UcBTFqpfE/mm+pR16HWQH+121+JvZGze+qLAGS2rSkthLc6SBZ10Wa
05tqGuHm6P6lHd7YtWYDy44e2wBbO/FEBfGOAaipqcSIbkKIzXcu7XovzM2MGqSz
KklSMbACjny/sMasdpjhAKUFJXVcLNFregnzg1s2a27Mo2fxvWF1laOyANZTjnw3
abIJdzE9VK0597xxqbzjRbWgz98xyIAeQ4fjYeyKQieHJTU2/tPfVka5xDWp0p/t
PAQYXTrGk7qRmRQJV1Gb8tiOMgra7/fY8QM3+Jsnk6jAHu+D6o7rVPffRMxGZ8yL
V+xwJgNrJD2PzWVC1yWz8cWXhl5tMeIwMLWf7cE2sa0yuZJRIudbcddNH6JCNgbY
BQQcRhZ8VHuCOn+FLGvXDpS99C6NO10D70BjlogOWKwNn6BSuTqG7Fq2zq95/kgj
5lpWtDuLCXcZk/b5YvuJDxaYeJybd0t/mpqCBtS3DbXcmUd2EEHHXh/iSNKP+TO0
IxO33DRiz5ZUKsVXGDZE+vfvr9B6b9x/MJO1wL3NGLXcwZ4o/jW3+xjI0PmRlNPa
oT6Qo+mA8xR9evSegWUQhGUoL0Omlko62CPepZwyKUucaKwX/H/7wPbzBBpD7b3/
1EO+AFgeBKp/m/oRviTS0D+jCSFB0BgBV8nytVRjt73whueIX1gTi4h9+QrVuem5
jy8weN7GR/xT33zetbRtqXDoPxQ2MjS++WWQM5qdKnVseFY1JOwPH0pwjKjslaA2
HhD6umFtXcLS5LXBU0fhyrpOwUwYuBrBHHTP/uKjarlH0K56UeDffVmjGGtXRbYj
tTlT6S52Pmf2vmVYb5ZuR5lrAxSeaVda7gPUFFHL+bof3q8yNk9v20eBa9j5yZ1r
tO/RmmSYD+a7V3hMcgo4p0DFZR2UoaEud64yDpW4VR9FuDI0qLUgrIwogCDLT9e+
A+deyTKEt1I+4uDYdIJsLS/BlZEz2mKk/7ox3wLOWihC10dCp/FW+FqujX4yW0RY
6RdnByxS1CGOnheNOkosKH/uFiFBZxrc4dmCMP+8+wRgBMmo56hhtXWLm/Afggqm
AqvGvjm0cDs85DYb3Em5U2iayUyEwdL/Pp/bz5XF4xq+V/juOLmfm1GfDr1eDBvr
e6PyDbfvRQRydlMXg2DuCLrjAt5b+c6Iy23LU6T556OfcRBZGKwhBn0Ga20jUzV7
2Uom4tCzf0I8jrYeyCcK+a/58nY07nULoksVNxuP+mWnoGbcXal5H+e1shKf4wdT
1wVfrF2a6VeslmxGwtmEhRDPUFgVKzFHgMbjAmjR5D7L4XFEM5S2FMiRKXZcf5jp
Zml9oBhZ/9JaBj1WWLgtNIHlD5o5I/ZWl3r/JPL8TINSBGLzaWjD7zzIYPuKMJli
zZ3j6auFEmAHyzvrbCVbPmhxR3ljjejlERfGdRkVsQTgTzhe/xmMnxr1GD1TImKC
dilXkduMR68VoWdiVbtm40cAXBDtLG0GStafral/yE55zk00R0PuerHQyP7rMlQo
U8U7MgkcPqH4wirk/KyO1EWNjd7d7hd9JErcGScRQaon5MtjP1/p+Ibq22B62Oz6
6NMc4ATJKiRy5+iiYpd0bVeYueVoCD1o/Y7XZ62fDyahxTCAKNGkVU3F73J/DPN0
taoJWUqxKz4z00NEhE+Z/qJOX2cugwRndmT9aqF1/hHtYZVh52eYJ6D/dQXFFXyW
ElNNwaIyCh/cJ7YfPh2Rb8PLeTzyP9XKkvBi4WLaaurxzr8a5gSwwYl5LlWcTMUF
F149Dt6CgCuGsadOLlYHITj0XkyS5eicNqrNYAiMR1OAK7moYDqq5TQAKgSNysBp
RkV/VPtrm+hDWOjz49WncSLeDd4qLz4P9qtHyxY63jn6PJj2ZHesuhkDWyzQ6Pm5
xJWR4fxERojfeEEqG/hRic63Ikt+qvAAwycbpmgfWZna+40NkFHtGsAsBiDv+uW+
og/fimwMoKbLt4w9nQJLnhEdh3I0DXPVIKpC9gIlXMvklrRctYeajxcGrSLtXLKg
QpWadys522EL7GNl58UGPoa/4tbJDIdXJC3N/iN3STibapoqYF7ClludK31Pgs2Z
TYOY6WaXws9+XQ5xji56aOPMKIGu3tLpZwmWwl0DfzSRPN33KcLSu+zFQPUIWse3
vD1I4rqdlWV5Q4WM9RbH8dS+TApM3g6ck4YNdA7ELwFlRjmfhlU6YqXvwiMFTBh7
p92RjmeRF6z2b0G4Qd550eoSCE1UbWk9N04oClilux3ac+dGcB0YKPgYB8bu0tUR
P6tB8NTisP/pE8YM+s8siM3rW5emHg+bERKGo4vRJ2BX0dCCo51B9Vv974vxj4OG
se31zljYDTgcZRMDAVCkN1YCfYhbEfLkyf2egq9pi02tAmjr0bLKWu+XCtUMh5Nu
+/f+p/uZihvW50JOL7P9JqNT98gYwLM9fTFilpgqbVSGfROyDp23X55inumT786u
gAVLrliun3/w68+LfiNOPKEnYKVpJe083le5agUMivx+U7ObEI6frTpsc9pf+aME
XUNPS4kx1yJ7XNY9OV9YHGDZgq/4dQtysBGmO6tJisPO2g58jj9Tf16qVv3D8yic
EBtJr093mK68PHvSSNPErD8hQc20Naa+p3zeLbnlbBCUKsB+CWn/4fEeq8acc+j2
pYk19SKmEFO2IBqhUOx6CN4GupKStTY0L2lU9LbNFzyKIKyDYTwq4Alc2d4ISZfd
4M5it323YHgTUCqfXw0eL7Ad6nO3bQCtchJhECthPvkxVfEqZfXKTDnXB89Ng7Wd
ysle+BSrW8npOzugSyrXJS9w4uOiSO2AHA8Lhdv//mPCcqqOvqg188rErkZUga1B
vxzk2ubv40E1Beh9Uf+VxXpti4kgHxrCdha8GLa8kcckjVu/6DTchyG8l/WOUbv4
FlAbBHbUzmDTbgSpp+p/hrNG6wd+Re2bnp7VUGXR1tvt0W7rOi+reCSJ8EVA7kyW
Gb8NlId3EqSUaUkQd0kgbx4H5qkR4S1+7czFPwlMCpnvmVrF0s50NMGEcqrVLaAY
kbsT4y8Gsa74AcoSBxRnOjvzF2AiqGqQVFmOEkHse/DzV98HzdJPnD1CH3auDDCL
+8WeZGhNj2qYJqq2yjzNhd6kYAehbbZ5NiQlVleTNALBgIOW+LdthesfS0HtL+fh
BZilZ262Srb+QTrc6F6+tToS9zJ8PaFknFip2O3mgpUbeWp3/7Gg/+5GHLfdebm4
XvnuqOAVBZcG/DDDURyx1J9z3TiMVYyBsDuYPK38P4vB3Xax9veeoJyhgzjNLSxC
x+vFT16A+i2XN9AGBz2M3PEMqXcZP++ZMq6HQMyVHJiW+wrvfCGdD04/LIZB9gbQ
qdn+dNjujTEPj+hQWgDIbzVIHKfB0byyu3uf2wxoOA0e4syvwlv+BJLt+6nIfoLl
hSvj4tE7tktzFVNclCFGHzadiTLZb/F0BBAE/XRbaYRaOrkHStC+TXqPqS08GCbu
yk8M2tFEqCBAN+tbBircecz3doSkub2l5wyqQ+Q56LObxWXVoJxR/9Kpi9SOFRJw
4QXrdTY/Ci/xyX6cALISYltfLjp5Y82vQviATFeYzuDm211kl8HpJo6d9EJv5j2T
vALDRCUoXQFCYsYzd9nf6hN7r0q+VKv4BN0SL85ayZuE+Rnvf5nl3kXBKke32gwq
py9DhuN6b3uaLnirSa3no4Uci1GiYrZ3rrZkY1f4kyhR9eE25JAw8z5L7z93JURw
cyjWwjDYhFDO/X1lWyUPEiqS5B9PK1fCsZp57mXqY+K6vdukyZ8w7NF4t9qeDNQm
F4R8zEtj8IwVTlAhWh7zC6G6q1iyUJLpiLiJgTlnnbQn42FDn0ztVaEj63Klsehk
IXHUY/ATs0USf2S/k7raciFe1+D9YjjPoOp6BP/Na7QAPrZ9wjE5jD68I3Aeyoob
fzSwG3wbTxQLzLYCi4a/tM1Z9qLCedkahXUO+16G8OKpWEL8B4W7r6eSc4ccXkTo
owZQlfkfbDqK5wmP4efJ4HF1EFL7HaLU8iTOesCtIuEwUdRxqUsUsgJBWv0pMHMv
92+CB86A2bmQH7Z3Z6DMFHOecMtj7SldgpG8U7Ko3a+iXgHWzsnJL3OmZCnI30OY
JhodOMzTHRRrIj+jEAIljr6B06B/8bC3ABs4H3YJW0HOzFqaFE0kzMHpEH7g1TDc
jaEo5UCELmb8q4S6yNfOcvU/U7CTqras1Q3lOI/Z4XoYrr0IsONSYG7kGWWDHnZT
EMnLNhMAVp8MzL+dt3Xga/QzSZb+aAqgBScMQE366l1xEaSdySb+lWEpohyiBnfZ
/4XnolQJdmeKj5uMiP8I+wd5APl53CisTiljJjgxtIvsX1sdc2pPNqIFOtCd2hIZ
GayQ3Ly7E500lF4uwPU0AZglr0fmaMZP2LwSfu4qwRrOHxQFLXIpAJ1jLIq+2/ou
OJwX+IuJ6oxae4WVQMPnWreu0fPU7eadGmw6orNbyLBPhg40SfH6W+F4G8LjllOx
nYdvGGqleKvGB1OatoJ8ZZGJ7utcT05UMvQpf+l8/jNDcd7S4oMTkP+AzBcGPPwy
oz1QG2G/dJFcYWyLpXNjdIfk6LVMIx0cUG54tR19efGR2TucQQzO7kYnlf5x1Mtq
WqY98Fk6Tv5ZLuc+FEkgcXUz+OvaUQHr07k90oeeO+rPcXnf75nuQDGW83bKCGEs
0467nDej8aEYAML1EysAPDI7qETz9LbmgI2S8r75aN3MRhpQaRTvtzB94I52ldwS
UNnYldhu1rDlEOrJgraLm8RKdinyalj9QwfBpix2Mxx1dO0HHRk/Anul/7l+AiRN
7EFIz1qHcr7YYNUWn+KjJ9xCV3N51gdsabvm5+ltMPgo2myqcGdKLGr8LtWEtZr+
BsZbUbh7ZEG++vN9SC3BT+Vq+VBdr1+KrZkZBVy92G96I5PnTBcokB9bW7o3x/hW
dLpECt1qb8NUKiP5d7R1tnpPRqzWnr20k5CEElCMbNw/C7t5NkGwtHppCFmBTi4+
stIFtKqvhMHK0wOA8dpR3fRYYvmeuz7Ff6tynW+uQCnGa+rw1BEf5tcsAzhQ/pCH
NREl3HPXmxh5RbbwzrqHbBu7xHbOtJSGsAENumNfxXU+R+cVUt9WT5breF23O9zf
lxlhAQ2rqBK21+HZnc31MobXIv5XtiLXsP/Mc+5V/Rruky8I14LcCE6drjXqTy32
uE0oJgEhDiLJ2MBfH5N4+3U06KPJjc9AC9eDGL1Qe8waophijQe1EprRv5Ncycgt
9sqFXI1Op9CT/7SB19oIMiynjoATY3/OSVrOaXoSMqkD2UaPJ+ltqmnkLLBnxoHq
2aMWcuSDlJWQyL/6EumjGDEhgeKV9KV7pMYPthForIGUrgDInZaXwgDq3rxjNSnD
BU6LJ+tFSUlr9sG+3KlCvGetAW0nDe/HX09NPtylO8ZviVw2kKEZujxufO+2k5Bw
9bUL2Ol4ic/JKyT4znn7RGT2gDXtvE+/6wp74Bnh0TNb04SZomc2//0CzWHZHAKK
ilFYjPXqtL+xnmTiJM5tfsVGoW07LD+pUelcnWxwMcQMZp47eG/55YEVLvlNjQLx
zX02yB9xsIGx/0HydC5ToDNk42YQLPJ9fs5KvONLFx+3i7BjSBVx8zAVr2UXXM1m
IL4PlBScVDgSIbkd6i53DfQnvO+OedGXGf46lx2vVijDaD4/eFRoJEEQ2/YA9NCU
dC32hqLfY9VWs7PMwID/mV9q6iZDrG9tXAB4lbp0Ffk4fItD6HucqfBFtL1H1fKJ
oFuw1d4UdOR/hY2cRzUn6IH8uM03qYSQWMY8wYZeNGHgOzQlk82iyIrRuOLBVHbp
TaCz4KuZJRYrl+s73LREcQx2jcgV8CPRi0F2dv3iv+bmJfBmBtm2S16QI22oQ9PA
lPWAxOQRbtgdC0+BBsEk55eTVdk61zYzDkI75Yf9izi3txukj+L6VAWYZQjlRURw
W8SnrWYhBHg4D8Neb65BvBk8pixp/AldPHMtsAJx9pIzvD1cO9q2eAGcmP4UeOYg
KneoQI2QYTEtKavS4A0kcYKtuG1xyMUKioikb4Jo/rDhMCPk6lEuu6ZNxx4tMA27
zTNGMbEyiXtmfyBT2ceIEsOx0us+cixDOzRYZGM0azbp3C7l/VQTx+K/CH/Ju61L
v17pUeD454/AHfYj86jQQT5CM3zOGJmhJCB5QYGJWZVxYA74dUowDHfk1RO4b17O
8rkDtc1K3/h8H3dAi+jXi19uidyHO1XCh7QVMRbA5Gnqb8UIkCX4zlVat4qG1rLn
l0A2K0E2/rIXT1GnDsuEp8rd+fW1u/kFHuOZanymPxJKhZJMDCXoKIk4tJqHIAyy
ds6nzbdyQOIA8B76JQ3ey+mjHrRQxf0WowoFNyI3gEr/snYCqjnBI3FqPt7YfY7Q
VS8z33qO64q4u/sLWGVQ07sQMGZiVbpnpBg8DMSoyCqAygt2K9skGtHnNk0+sm6t
3p0mbFazWBqmxNdmmJGm2p++6OOSqPJn3h4zuZ1qTFo2o/PcXZzcsxTqvZLE7iP0
77cgeLef4tP5NTHctKOtF6xAUWjmiLcXBdimBwH0yYBTxmHc5MRhhRwn0GT5tux1
BFw2a8kYfp/wPwhbDWY3JzRIBhpX/bjomnGpYN5ow0p4evsCg8eguPm/DpBrQzNF
IV63mZFb8GsBEkoRdx9MIyscQWiYN9J8UDNOoM+hK/9Q+AZXUWTqWIBEGc6C597T
sISDejm0IAPkTmHpkjvkZ1Toz+9miF2SHquYGIAWJxfCwKJc/sEtdWigKTOBCa+Y
7dKaldSUn93fAefOL2ZPf5L8G1J6k2Cm3QcTQkhzzUQXrVhUmvEvBYnNIv5jbvws
byX5SeRnoRN1YSbOHxSyKo0rCjessI5c94+JMD33AYAqlGQgU4omMHYc0g+hx4u5
eDFGyjT9KzJCB/CywI7KxcfH8N0HDNg/r3+xBp8BQsCzULz4VZE669MqbIQzLphV
ldgKNMdoJvtfwtjsgGKKsWqP7ADk2DrdvFlaHnqphbKYvomaDaKfE/62QzqrZMnK
911cCg2X4+JE1tJ9gBiLbnoCBBdlbFSLCJtuea9qCXJZ4ppT6Wcr3/UAvqqJiSL5
lJ0fyCd1U/6isxx6W/QUltyWU/EPdRq6gWvFuBwalGOpWsquT0FmFffQlSStrRMR
sVrdRLn1CtGfTfSQwkcnTVZ6gT8mW9HC54UFa3dpzw1XW2EAKFN+K3wRghg5Hs0B
q4DNZ5dbPkcdR30xiEFp1XDsNm6ZU4jUnuGKvR+ra/Bj0T4OsfHBAyoGTnta9xdR
dZhfCNr0fX3/WGSfmXjF7ehQrqOVY5lynj2crTapEx/XpQPZPzOPNLA30IDAm/Su
B7XFQF1R/ua0XaYFpvG1dAo9bUb54u361CEK69UZ2wLuzR7Nm6/52r4qF2BGal/V
2FGA9E6FrpWAutyCo7tvPrLNapZe+pd1Lm1Xn6kK6bPn/vZW4d069CdO+nP30d7E
5ueCNk+0GER/+yPzqa5ZNDOppY0Xq3g55CXs8EdxwDuauIqUa5p3zujxfGN9kxTX
ZYdtAFfnvIuDGqHStEOsJLhtMCQX0f+qxTNKQrFtoLUD2FmTiT3R+XL1u+QKBgJP
IS184e5Avge2zmSdPdTfA6kXYBeUFWzG4KjKU7XLd4g0HjmVHooZjQ4I2OOGIHZC
jIecy5C6V+9bgGfR4b3LuHUIm4NUBkYZAG39fwSivKfFeE86iSQyf+GclH8bVaxC
KderqIW9L0sX9bNvzDfxknqATkMuBPJ69W+JWovsYyoBwxuUI2WKtVooy0JVqk5O
agdb4O9lNBsmTw7gBBs5OAKXqj2gD3oFKRPy07PhX6XxasbpR5Nuo/RgC51kzAYT
IuF8rjAsMNw6YCbWC2b/gsUETJDYFGYVXoqkAIE80QbSF7hDfZ3nf3eiJ0u6Nj+y
zI3M3hX43l1QNSdM9s6lPYlDJsLjI51eDbuYNzuMCZSvtD7bdnMDCecpIxF+W6xp
ySXFxFYQ33wdtvWy35hfCTfwVKHpI8693KKwCfPKEuMZ1+bZAzNLEEgNOw0J3Svg
gfwXBekc8yuqTVrmfadaSyq9mn2/Pdtbf6tckjlJpFAnr7h/Y3v17WAW+Jl6+ISG
N7a9Ua4ouC/HzYp/GaETc/tkEt9YvRmzTuu3xU8ouNf9mzCPaHhBClsAD4l/CVpw
QJZ51u36wHubTcyw08eGBw3174XQoI2JyB0yFh+hHD8zoGvSsLLl3v3HwBul1fvt
8n9P+6H0JPPhwjw9Dzx9w4NDL3qmuoOzp89UWmuKiV4TrIhEihGuLvlR8Ka55Yr3
7MUm6r4QpzZFUQK3iVpyaZiBdNSoKOqBi/P+gNutke3T/7T/Xl7Ird3UgK9RzWTE
tnom1x0IaHSrZnbirGbH6+WYxDpYSzFFpuGhZdaDv3Qh9yJZFwuwrFgCKnHirQJj
8oABWipTMaJJMuUXYVY+348kaJ97Hzo2oLOjtmj7vwqQ/h2JxxVAb4PbNoO87+SX
WPPugC3cg7O8+qRtWXaY0V19lirqhrCk3bdfyPKjukFMfkzVUX8pBPrMhhMyQ/MY
AXcV1Mtz8X7ziB4rLm8BHSC+wF613rbx4KtKejM2LGGpGRC/ofIAwQWfBnGPGfXH
MTU6TsAHh/+94Wvjb0ioG0Jrty/pVMN3YOjp8q1U0rt7Io3LGWScFkEZjPHDMiNH
fSGIjb3y7pgJg+poRvOOPFr6scBu3MIQvxWOHBSifftotnpZWFpJ7ZNQTbpWElqN
QxOxGPVb8fqNBnSk2sJ+olXYUvxlD5mAWIp9vlXOlCygwzOV+GyH/lq47vl4HOsO
3gsKfizuO1NwjpfKxuY/pvMmgP933qiS8rWkADgO3ZIc8fcq54QTZniS/uBojjxO
F+ER9ivALTVo2KateQrKCuBMQtISXpijAEFMiWGlt9GTGvv6/hCbF4DBO6BNj8Ei
IC/CU2a3sxfbby8n24OlbO/+6Gp2BIPgydJyYkyu0GP6dv+XQDkSPGAr5n8k+XAx
SmkmLGxvHYvvq6pfrPENLbv9VS+H9AgJnQRx/io2emFBVWyuC20rhZCpk7AytjDO
+Gw+Zmu78wTs9x09PNJ1wfZeL6dZN72tPbUpmoNuEnei553ic3V4NvsmgODmo4VM
tjqYe3R+NIifkJx5QIWmLLfL6BoWiiC5L9nKGpaKV6kXTt/oSaeA6mhclfYPaWxj
AaM9CaMmWdjJENnrQnh3X85RJTQgvKJlf1EEzSz9RlGROhIs0+qcmvFsuuJmAN4X
WVcLPciC0y1TNImewdVVDZshoJiRAbY3D+woPu4QhYwEYL7YE2FZYnIZuk2JD06Y
IffElvTagk+yWNaQ17dIAbhClFHjjY2qjBbjQf5R47nPa0LyJdNj++gcm3P9jpJV
s+BVq0NtQf3nLx5jgriXVWYpQQ+O8Vg8mJN6fuOdbF6dtgM6i6n6oraOSX94g+B4
7t2chr5OrViWiWlR+CL+1XRbqRPE+7ZZHZiKAPWtgr+JRUvRpYsazSoVYEjgO/4O
hrzAWTGBdGlpUTIrEbFNObdhhcvon9BZaFFdP6Vn5JFN32+JsiGR4l4xlhHThgw0
mWmUC8yxlCMR3iAYJLB4Nn/45kgeLl6KBClmYZlp651nFA+fl2LiRxH19BUT5xKq
jL/KjaAgqv84KctajBdqUKkIrfvSjzMhoAv3GfyJarlN/DYw5O3gKmu/cwb8krhH
Yy0Kf9xTX3PW8W6Qic9l25F9Ph7gPzmPN3vlkHINjrIQLlX8rMNqaD/snh6TUNMm
o9WpXRitNI1dzFI/g3b+utSRZCoqkcrClA3zVXvlyjVJKhR2OBw9wqc5yqATUcOd
W1PBVie26u9mNveLxrU2EKAg7G282HvWb6vXfZH3fPOkoLZWi2gchPcgwRe0VyvN
axd4nKz1fuDO6DjOI8LO0ZL2LGK/gPuJilvLSICcTjwKRkgc5rDnZ1tX2yflqyGz
8Rh2we2heYZAhssePQPKy9jQNZjHBrF4Ji6G6UWVrmRdKCPoTXuqTZpflw9+eDWS
/RMi1NGMGzOm0hLUhN2ZwlrUPTho77t8Fw8qNVf/DKAViRGTD6kTSdKA93SdFicQ
02f0UOQXDVpC1wJiAWpp+6qmvo2ZBfx4b0k6DlqE72wKy/4ctBH8V8DLxGwfjZhJ
aV4UOov3v1Pm2QW4ZISNB2McLQfutVMXs1E7oYtMa5NoQexGnCiZi8mk70krh2aZ
C1ks78eYkKju/PBkBxs9jOK83wTxlX6bJ1oLznNSBZuHKMR7mEuMvFJux/ATkOSW
YxSC1PSiTBPwbPgdZPvx3vRfBsh59mowsPfMovzC7yteFzqJ4aZcDIvJrADTF8KL
BlZGnnOWLC3RJOaFH0O+5xAwhRV8w/U2b4vv/8HcWijaccyw5oFMYzQYwtEtx9Ud
tuDGl1k1vMfG5bXb+pIL+/Qe56aVJzlZga2ACsE4Ng87/ViwEo1FJTBIJExvsS+Q
fG/Ny3KSh28IiyjK2ddHQeY6DFeO9NEiEBffReKtiwyvx694lGrC1JYryQhhSsW1
QMllCZ/YPP5/n4jfuF1IFIwGpSTQ8bW1+AgwnXo8WmRH7zYVhAgQbc/tckBJW6Vv
NZytBXXon+q7T+H2zIhGR5HSGBuA75zvrMz1P4eYBtZLCEV+8wAY0HqJUXwZx6Hm
BphQIWH9nyOWK9sFFgPc4w4JhNNvvZd2sL35I6Y4x0y9o9EdYXOJfe8GJC27P43S
UBloo1cC66J7fTuqxv9WeCdmVfxs9EnGQYZ6b5WaDrGFf7Tw4WQsNnFVJr4Y5Okd
SYMEIT53z6fj28c2mSYv7LqLYdSGpArGDWRlw1TKYwWQGTkIrtC1erf1ts7I07H9
THBmFISGqS69w4NHgllwkRzzYkejgjIqsJplh7GLh7fyxgVCczOim2X1MRTRS3cW
LXM1H4UTKeC2mvuvKqwO65yTQ8OQt4xZITomWV3NO9LKLCugC/hn1LZmkxEerrIb
aGX3EwOZjEMJaF27BbpYqO2BPq86hugShDOt2eALYw23t5ZoNFLQmgkxEk2eDjN2
WGDrJbTqsxjIUWXFalH5taEza+1/W50rtWDBRKN5eUuvX4tizSAnDDnSTbBvOK/J
nwvbq9wDbkEYin3p+YAi7JqtfgMhLwOzkQXhTfhf6wSnhmSWbGyur+OMPqE7zvu5
DAYoTaV6M8LF8dNypaZz1vDM5cCOGR+C4l+HZbzCUD1gV7zo5OGioxBwj9KjJ+Rn
xnny1uxEak9J1gLC/TCASpQ31mwcC5v2vdbfgdaqhvQCMiFzsOVEI1fPxTdOLlEJ
6QtXhNY/syr8WdhCNXpmuBHZ0ZiMgEkCA+CqEuyw08dfeOBID/HckTvUxnd3LoT3
VHInKfFB+CA/9IVpwAXqz7rn1itZpCYd+Ay4ndffTydVEX73F810OFn2/DJZf9/p
2ocwQw1ZI8qozdddss0RyRSzC6cy8MKIX0hD5i/Hh+dl2yzjBDV0aa53PEARWNBI
7dYzwSz4lH3B1JOMPrPXEX0jMtdrMhd8kYlNvy0B4UwmV9JKBz5EYc5o6J83K3A2
pB7ktGVFV93wfOifyhAA2iJycRFnjeIYLylHOQC6nWzgBI9hNDSwKWRC7ANY9Ttn
uOP4MAHpCNS6qZRtNxdfq77wyepeWr0kKK9P8FhgHZGMwVIIL2LWmvb1eZmY0AUM
llG/4BjDlrJhG7uvRgo/zNKxY8y1L8Js4K+6RpbyFwM3LX0LLIH4WmGfvdxNmIb5
fga/mM9MDRYrj46C6FKIrXW4BShm4o0jKl5oMPKS2m9wcTGsbq21V+2b7PiqFE3P
i+wcbmmxLIx1jbsqEHu+kULdBUC6r3aNKjByfp1wLhMYjx1YVIDVUDWzYj3kiDAk
4ZgubRDvdWaH1cfwb6owgW2TtVMKw6twGyjBlkutZs5RWIuUvBIVZOn1vq5Q8HUf
0oITgAq/XPD1t6cCu+cSdGIIqbLC0rm23EUru3vRFozu/ePqyytIVD/A01i8VV0O
b1hkgYDZm6BQKgyqcEdTsjhGcIybAAlC9gATd3i43G7SNgQYabyudFgoxT2k98Qk
D4f8t4QgCCPJTmiKVcrU4ID5xx9TBP0Inltmb3lVjsHI2AIEdVHywqj5gZf45XF9
HcDTJBpjx0OFWLYjSvDQttQA1E1QfvZ/9UiJLRoAuGv/2dLxOmoDpG+XaJKouqP+
Hewz5wfZWBW3lq25sua3C1SvpIUINOlpu55v0rCUgVvaH9bg0HilL+0aPc+QAuUv
oYMtXN4I5ft34K8kksddyxbOZ0YbFubWJQSxfyE1JMElJMMm21qLu7a7s2pd3+Tt
R9UmuzOYDpg9aLunDF5ZfVZ4eKlHR/PBTWxooeHBdbkoebcwTrZRhVlgKBr7CtBW
M+o/hzWlogWNeNsIq5MzLcqP88hysVwV43MIYAZJPqn15LyXf8ar/p91o55DEDNm
lpU4NcEYpTq+zyo8Db+YvMrWAvj0k80+4L7o4WRyxFh2EP986hpa3+a0jzhzvBeM
43MYNczjvftYg24STSSGd7a88SvpecWIbk/ittrQh8+HI/0r/d4nnz3Abta49qs6
tZkbmSwvrH3N+jWqSJVF5FjojeRmb4q2Sw7rsMYLvapB9lnZVf9XUc4UyGSQ7qPA
zMsnnXe6RRefPRvGaazRtG5Z3eq2ckVVIn4+gaKc/8nF81gRm5RsIqxH0mfj69Ik
kRXseueZVVyKKSG/KvmZMRDYbOvgKAbFzRwsvpH7HxjwGyzt5JmWd2GqTtQ4YmPp
Rp5MlGSKtIUA+xYFQIZFVpJuMNrU3MYWRQzDha1DI4YAL4w8PBPjgHU1Z8LRyTT4
3N4E/lFocPuglQNFQySz183S8fePP74tl+JEIWNmEzk09SX0ARM2+BXZAnrEt5Z0
1gPfIIKFWjVWOxyHKtu4dkmOl5Abee3i70ySnO9Yz1OJYWvkj7IeYcwGQoL7PoKF
TX0T2hZcRnpVXMfLLlPvHq4cMhFYrIdTMAYBt5LDq2Hxf1SQwssX3JedhPL52SJ/
oC+BuF+oazQCGVvX+XVX7zbzmBz2+Fdo4+Zc2pPl8Y4SgVuIRgCLi6WWqzv2KcY3
7MjcRIa24187WsNwAoDYUBgOaYzAqn4F3ABgr8gKKaOIkxukMqYtzI2I+mlWgF2B
kFfG7CopRtKeFQ3eTlayivICqEBTZltuACySU0MHu0jwQLvMfMlwvpUDVi+3Bl90
bEBpUj1QW/sTPRF6lcvC16MdRPSrEArWZwCpBAVX2lpQEKM05IZMxleEAu5Qc+0n
chiVkCC88aW4wHfQoK89OxjZvINRYKVv1jPVLkkehxfsPneJ/VNPcd8EKuULH2+C
jtXt9dIM2Rqr2fmq6d5QgDUt8TSmHNy0kzpMImabD3YPgCJwMGufmWJZF36LvNfa
ORfW0f0ZbRNuzlTUV02Oze3sNzEYW0L56ZkKs7ZuE6iUuEwIcVBBpgJtZeLXq4bs
bqTKffDPpGKpUOgPljbmR26lkBPbntOslFVHodGf66dWTeFETDC372u88pxm+Qu0
zJwWUzGoGXmcUHlR6d5tQ06ZfckunEu6qmTmKbdhRdWu+hQxQp7knD1AD3KPdC4b
oj+IOrORY2IrD6j6sNiJCtPbUBL7wRtMNginxcavvobPy6dUsWWCxg7DZutCoNQV
BVtg+FfkWfRnNPO39qGDtnOihaA4YVPCS9fu8YV5gwSHIgZlsAe7hbtzimF3GuEb
a+1qoF2c9Uw6ZkvgIuiIbKHlQRDZ9bwtafItRdbvM09WzpmYFHgVm+z7k1QIfrzQ
07huGJ0Va49tiwAGhynIdPY/2XwZ3DrW8BAA/jER4QmoTmLyXNMScLbkAdB6wNGc
5dpMewgxcImA92Gpj9zwSIBE7qh6oYAotnp12gxrAYZmkKRdo/H00M0zA8l+6bm8
ef4t2DTMImBNm1LQ40FQWUYAo51nqFz/ABsIBZY6P2aA/JLhLBKqZ99P7hDwEGgf
3H+ZodbqSPK7YPF9MK5Hzd/XBL+UVG7wRWyPPFVEEkCjJRy49ld0aF7S7/cIAW+N
bwM+/26sNObYn77+XDIK9cShEFbDjw6A6kM1iITXBhRlkQloiL3yIjdzEmwwO/kF
mchecLq9ARiNDcAfZCcG8o7PzgSPuVOwa7j0dc3QbMTu7Ah4BZYKwhdlaCVDGbwZ
et0JYmtNESjqc1fIEtgmG8K6m3C/UU/fvQUoIXZW55Uzz99NLPRhT0wB+skqozBM
IrvK2jpv1/9GQKpUUx/qGcG7w4fcc9D+7jTQBP1KTUz1ajjOX1Ra89KBdG2jNdLI
4vacBpeoOAYPV3v9Zntl0pCy0zk4FZsuBjWcDJ/8q91ANtNNw1GkaY9nrAfrnpun
WGzjen/5ueT3xZU2/FNz7hqdFpyThUADC/xhmkPUy1wsWaxH7zZ1Y0hPtBzUfIch
gRvz+jDdP3DTWa0R4WkAqXjv010jgBfKqnJyJ6+8m2XE39U64EUczHfMtJKU4pSM
SZi61OgIrhhBljfQpqb74xpmqv6MNR362wwClGF6pvxKfEW6E37hLNjNW6DhVWY1
m/u6dk93coO4Sb8edZ6AtKirRzpHdG7SV1KvbjjCz/bSeRljsqNUlD5JX81HnExU
jICgzWzi95f3tB9HabOyA2JA+w8h4vMrUcbDi4pAa3wQwDk9WK0IqNII/qxzNCCw
XZWCyRtSQFOIvks5QZ9bGiPWR2TlmbrZUvOtgUeEU51JXd5ZH+Hvr6yJIbXmQsUI
JSa2q+XzFzQGRkFQ1DdV6fU1jPmn5YXmrgpeQ0YfRWgaLQNYza0okGAzeA1HQ9MQ
C6Qhsso3XIlaubqfFGN/06+PszR7m2g80cL7BYTWAjoX8rAp9ea8W6ncz657+2bU
lw4f1zgdHufd6pqX43cNQYsUTtgfr3TkraTQJibhvUBKZtfLreeTmaNvg6sBv7wm
AQuUEMukB25sqnTYexbizgrBqoeQ0dcXi7bSTxPkiDe6SymwOh0xfumpPR1L6m6W
CxCopVtFd/M1yn+Q2X/37lRXIJQGZeLDlz8mg+6CXp/2CPR+zshXrgyBfH4ClSX0
WY2Ohse4AV3btnvu87HWr+M87IcRkzMVbP4XjK++DRXVQmwALliOCZl7bamHWR51
p67rsJNtwwhlruWp8pUog6ezN+cueXnOkJCfTfZs9TeMomvQVND27/xdUkYi6wRm
mLz/85lIj8Ih4rnhepfUaKKXow7ZUfCGT44KoMZBdpOaQOPxYU9H38NHYMaOdhmG
lj5Rv45NUb/JI2gnkehqLcvjHg40YRuHgBLIr0POy1rgzbxJ+wm/RBlgrrR+/BKd
wwYjXB7w0no7o4jaUAMb42P5AtiP6e3DhkO2Zh+qFOW9NyZw3xc1d4lKtaxqzRN1
YeFnNlwTshPzvW7CQ+sY6yAPx0ceeY7+ZMUGbCmYBE483uJA0v2wIeHl+Qmn359O
iczrBdvfy9nOxR/j3K1fbOJS4SsGH884TxPR+vR1gylaLuzd5kIWhS2DBeJa/uOP
h5CSdKElL2vQMGPiUFyibdlSYceqbyQaBZkISHLuj+kfH1UL6uMzOMxpMSnfel/k
nUovx9gU/JRiP4eX6x3s62KfxOosXPINkivxVsIllR0TPVqJhnQGhSzTV1qaPKAM
/C3tYFcpuBYeX7PizFyiX4IW0ErsO6gAKQwEUFwU0yx/pAoRfti/xCq45ueGCWWa
/IZ8/MatdhjHaoDx0N0WNlGH1acldyH2/2E5hoNNcNVc+yuLA+ipsS4rDgSveDE8
71IEf1XtCqlJxekOX/OwPwx0opG6CxLmLpI6VQlKpP4AJb7ldtvpot/R2s/66Fls
qkmvgYS6kxXvIzP9ZUxS77TrDas8jcfXeS5ziGZmdN1LkMfI5MYnioDb5Yo10YWt
DLJfXeaLEBj59jNPW0GZW3EERulKOHgHUindc+ExnIxO72t99Z+WgITREljGjhnB
0FM3t+T9ewNT6cIq4lKvjPu2dLbQQyxM5sgylrKd1ajeN4rz16NK2Sp9ULBJpLSN
Jdi84Cyg3VxM4rUU2e4pNo6wQeGK/OD8NObzThAFWuFaOjg2uJ6AXo1boeKe3tOM
FBElaqLWfKjGJxAkwvY+jdgQdaPfeDuVZY4ZlPXhYbJvMmaT0TOLAE2jZ7Zytji+
WwiNIfR+xNWFm3+7g8GEsRPPhTeAPzrUBwBsr1Efj9sJPqn4OujBLYNM/ZIvTsBV
V/AoArQjqFxL/BJpexho46tS41DYfd+0Uv1J4fxFW88Y15xjDqDavgDTpBpj89Et
E5/nmqGBVA2p2vuJpEzEOA5RVSAKDPI/KKDxpanEqyJhZi4WTnJKBAEsDTOpz1kg
qFyspZPeW2Q9ycKVe+r6OyP2Rfnan7EzkwHh5a070iB1qufJWZz0eGmbWxy5sA0Z
JJujBKH6jh5FNOSxMwjspeRWjjxWz/yiFwptKsVqoeOaAATlAmoYAdIYN3SgVchv
udpgtT74jFf/0StZCX+10yftxUmGBGAc7kqafc2lkN/SWJAmaGz+ylDw/V3Xy8Xy
ZFHL22iqLfujlri/mSmPiLr6WhVbtWexFHbNxEOQBZV1FDbdNIn8mBS9LiUtlqpO
JADbt18WKdOMY+ge4pLMmTN5UzBfeXwS0Az2cykn8c/6+mv/vJLUDuPrSJb2W0Fr
1XnRVTPtdoQhPZOFUGrHYET1H7DYJAQzzNBDzbSByufMIM6DnLq0PrMRxgyUimjk
SDAskYzmoymZeBvkWe68BnFBGZVWZh8bgfVfD1ZyKHjdSPwTV2+UE+Enf4xw0esb
tasFHIHPgq04rkB65oJWtsH8z+IfnJFktZAai0g26hIdFw3k1xjgdiPjUGEXZXAw
ZltQltdotBMVK0j21qtaPwbTsp/NtICmmoWHBugxPD5Wxq4vHijVQnQ9kU/jGVPH
2+a09Uscqz8liDpbTXLPJuJGd3e6Rw6R0KTRJp+v50do2YI1K5rr72LI8i+F2LSF
aNulL4XP15hQvTMp7GYR+2cdFKOsSmXrbDe5CVwAc4PttxJjZcyV9Khmh0KaEU8N
aXsqNTFzBGatVFUJUlM3hJZe8olzgyt0ZQCHdpIwxPhtuPfmB7jv7zuVRGnEGl+W
ckR59MvhDrp4OgEKGJ6NU4vMh3YPWuW2wIaCE48T2e203cg1HkEGQ4tGPzLz1veF
sRJgH3DqkDON8QY2ygaR4KsdMzIT3TSH5SF+y7L0chmrJcq6VQrp+FWDRCjOJOme
MNuqnNEl5aRvkm2AUyq3TK/+ryLKOFHPAcLBK/mQTDiVs+4Go5US77iRnoh5A3Ra
hsYYDoZEW13C5QhDx9xN8VtuWkdruAdhsnrwR59NEMbQ+gda+28DiF2MGDbDbLJR
xnTkuIgqrY+g+9fa9jYsWKyCknG2N/dZzH+BATPRtrzpssEN3hof5Jgv1c0n4jcm
V2AzRKhxijgtKhPsg7vA+fo8X9ay55Q06v/8t4oP/2EpOnWKY9DDSA2LQhSjSojO
O/0nOIXTIQJUWI1XmkombTKLDvmvUMa2t5Ezn9BcGJA7MlJgu3Mqh0+2p5C1Yd/b
m4OnVoj4oqHt5Y95tQq69Gl/IqECPP5P0PHYa/ISTlm2QSnN7pNd19Hlp0sVscZu
OCbX3uQIJEGySxV0+NvDz0Gq3o1ykhZlEtt2ChfgUasHLI2cEwtvY7z0etscnKpq
hUXcMhva8mfg8JOf+Ym1Uzra9+G+gjKTYJBuVpzDaEvZt+7UV4RXcopvNmw67OZ8
jwguqcabKWxaQf/2ESZP7ghzSeUpp7m+8C02Qkqp6CbldPyk0Rn4j5aV+eCTV1+r
5/XEUyuiYQJ5lj/ea/q9HovHnEjzrQy/c7P/GjBDVQCC8BQtXo1Aggt7f8vNtaPL
Bt4+ZOWoa91QrbqdkHDtuiBBztE1ihc4Ugp6JezOYv2ww4xnnwxILVTaLzQNv2YU
yuFxtKWMnjlTafSDqgK+TgjfQ+I2yQR0mUvAMAH5yNqVyGfez9RUMq1mRskV1zVl
iQCflw0iFQB12zdISWfsd2lsuJDTj1j6dx+QW4vn4PqhLupYWPqBSaTM712mJ5bF
lB0Lnyg+KDaPE7LHO8/H0CFYGgnJnbBPfBNikFCac6HMrJxojqDeZtXUkjDkOFga
3eWk8Td+i9K/KA5JYaq40LZAm7tbwO1QGX2scnww7eFtFgCByEyxYbggYwFOSOWa
vXOwid3NL2xKO8PVoCzm03bf3wzqzmGbIoOJOE2dgXqCcKxV6XUZbay97NWW0Plr
G0gayN+yqtGi7qXnXvUKXgLETrjTUhFjJ/JXmQLIFZ/748MMA3Hol/K2Lx4QOSHm
/qzdETinEOJUuI2Vf1TA1YBmIYcpfnAvqY0gG6P6Drn7SSHR3Hq+fM/geuDp7mow
R8HR9xc093rScTkS0PLnsNSif/32kNiA0d+lcvdaMkcngOAwAPS28dtDw8tlaJXB
XvPcPExTfvDTB34eSLtCy83X4AWNynvbWgwF2WYX2CGPushUHU0ndYKToKVex0Eq
0Kzh9+2+QdHHUUgPgA4HOJcKRV8RXhA0cTvemKR3hf3kE932glet1OPOQbWR4/NO
19h2ZTFKQyRRIUKfU2IRuXo9LtGAgzzmlQk71u2MioyqkHiZq0s/6BsA30hdGBZX
XE5rPhK8VrXb4v1XLpvaz7LscyUFy4NlqgBYq2/ut+6jwNxzW9swaDljKwu3ihqF
kdVpHMXJVG+9QcaIW+lk6DrkZ1zjsfLS1j/tZvuCwnsUoUJgqUapAUtWp44zezM7
YLhP388eBxm3XoCMIj459JAcLv9wWNDWZpzRDB+RDYulM6+Z55BEPu0m/V0dkLWf
dp0Q385Q9COt3wHVJ6atFTCGCTprUzh/d2/8TxKHNxGlICSa/jueTGIzpRn9mBag
FkBC6lrup5RnMs0eMF84bsyDOGWblAHD5qvN03UdCyhlk7Cp7o0MwMMuiNI/hwFV
gvEvchM0kgSKwZ4XIEWMG8iRCMTq5oOhXB7Rbmycpykv5+KolEsnUozIbRm/Uc92
qwRK4VafyxoatwA1humqIQaLwqFiDoQy6vfnw1xm0+L/oYXEJ8z9Fm56GsDfB+7m
MmrUlynSFMbT/Uil2WxQLlX3PtC27XoVUfzAL03oyysdg+F/5GG5gppybBBUJIzO
ptCkClnq4YOTD0Zd/G0PH5SYhSmV77b2WOvZHYIfl1yrXrIRuamX0Ti4WoJOZqWp
RTpKQY8SvbNiIaaJrNQk6xN/oeiKORnsLyVKSWcy4Qi91EN2yX1JZEUkt7D21zkB
tzXv8aONAHcOTFbz+fb9AY0jRu1Sn9W1f8TxNV3VJzJrwnm/osekQI+lKKvuSvAI
iGAhzhdTG8FXVhT5xz0sIYPWJ2x04krjgNKcHE0ag3TVxhOnVW1nAOBolRfMoNN2
ZJmkJOTCZr7M8gvQ/e1OUGPSL2aDfH7JMkWtc1MOYawn1JZ62WqHSkmJwVmac/9q
Jys0wMLXDTymSBgypu4CF5W00PV4ReO7ta1eacrBzwQfkxRnKQo4l/wc9V8KA2rz
jATFv/keki7WdRoleKKWl722tYGB7WsSH/t+gq4T1OmnzsobqgvZIcd2KoAdo/Sj
4GfLZsn43mC+vpTRs134fMdUunL/Z21xcNZxJu/9W1fyoJWS77JZOzTAWumWbtYv
cE865GDEBQ0cWZgHc2Zya7CxJTzqAR1yUnuscMYWysSUX6wjR2IYxa6lFd8MomM2
FsneRS8Kv85+3bvy+v26PhKgI/Sc5HlqCbsc7WOP5QqoT1pok4+smGExUwHMgP81
n+Mnzog2uFYiJ7n7GoWbZjyCY1lYIw6AbNCfk4gOcgSoho/0TvAIW08EptKPBOE/
jby8kIIhQEFoJoRZZ7u/dKdoQuYapovDuAiKInJXWUtXcTEsVqRJsjRSlBTUYWJC
83wo9bvAyLg5CQAOtHc4y4ib8b9hAM/VCfSarAbroBYNFMKqU5B9fogriLV9bzdF
CmLrjApd6QtX/BckiaDCFEzPZKO00aLs4NE3Jn5P1SehjgOCocZDYdSzaL9559qt
FiQjSBtYrLWGcLYWlZinY3o6eaBqVCfG3Fzyv7T9jjYJp5UCLcbqES7ujEA8vqBC
GSjcSFPci0cKY1nPKGVDDP+SmR0v479bbHzYGK1dSHt8rJooHBgKWTtFIA7t/B0i
iAOsnpolqk3lh8bc5Ew930To5qQXHRHvFDexuzZnqgYN6fvf30DtOx3LUb+PqJUm
XjncTtqFXrFnQISyfd+fXa2+cuL2s5siBV4BZuu6HG+Fk2TvUNpoL+sp7AGujwhE
3htRe2O5yaCSIK33eZSOuGJ67pfbojaDVC9RA9ymKpPCvEB3wAlXhOnVXc+xI7Tr
w1TZwP8I9CCTl78xf7WivDwVRd+kmokLsWysbksaQTnWVOBemJzB803PX0DigRll
4UYcjJQu0MXRsmk6TcXy4xg2A3FCu9UWF6SPDkZqdIU5UAEhI/0erqi66vgtmKEH
gTCDuFsuXMi9QbyZPf63YJNGYX+HwuMhGEN7+CGIjfPV7ngTrksko9l+oikH1Rmx
B3qb3cJPw3r+Qj+JE7y+DdaiZvbvDHvjdzDc1oOB5wQZ3px6lRkr/YKEzeGxzsg7
UAJG3IE8M0XS5Rqj0qkXF2Hi1FypIHtbDheRUkRB4KuGBxA115qwcRxE2y83bGF0
H/co8OUc8u9JnsH710SQhPblJpZygf0DLaKbahSpIJgYcA6NQNvQkoIQJbjf/ZGj
FsBtwn/M2zhdGZO4NcCz2EFzBEngVsZaXOMzZ/whGXk+ms19jpTZh0oVRS3dyUNu
ULPoyd7xVK8yx3FKb3yWpy/fx67Ua1TXtKgQHSMAI7Iya5EaACCDbLHX9tLdo4SS
hVye9nenIzZ3QhOd4jEnTcmpNoh6Y/yizhfP5iPoGRwfQhCgZS+lyxHSTW/jicWM
Q1gn1J76E1xDmiNJ/OWdmb6QOjUCS+95hsYuVcHnVDOBPUbgKKjXXD5mxxY55IwT
bNAFlCfR4vMKTfaezn55dtAF2Nd7RAYBkLmaSB6kaMc4BPycpEZGAxCdm249Ao+U
/a1i80oHZdgwsQvlTno0Z7O3/diivPK4Qn/5dNoXNta9V5IRuqHMSIJmLdRT7GX5
RFEZ19vSh7my6IMYnQ7Tm4gNa3pNOBu2y4ZTvQm2bf+R0NQVdNOtgsHA0V1l0BN+
UFHuc9ZvTzValEUjnUnwgzo/K4DCehdV7z4UQaXu0tMITdRXTYSU3Hz512qlwzCi
xNkjUZHq7yPe2CDizLfGX8EIAA8c1b7wjcVhW/gsHvxx1fSiD5Q2UUnlarHPF2Gc
VS2XUZpa6eTpvWhaqa0JOgFJJHGLMHx2cyGIRl0wWjxnuirJWLV7cE6CwKOIU8GD
7RHZFBAzrVNKgZSVrfF/8nQdIFD11PLrGVmtDjTXhO4ZAuL4NDaJHrYhDM6o3z4b
EjFifiP1kqPBbrI0pKkwnANukdvSmHIrLQRIviAxTehOIoeXCS8Uz2yON/TarHyV
CFaWkiBiRyO9T/HQqFd9yB3xOOsGQ+pPl1G5TXJXW3bVcxt4Bumb3WtRJvrWjYq/
kKMGKiDLx1ZBjhX2Yfb9yrlwLaPJsvjEnrUCrtIelEsUtD3TUp+Uu8tZ4gjsA3GH
7l9JX8GoijvsqGbchyUhq3N5TUN7BbkUgzp3CxsJ+UlriCUvFep+YOEipCOrBOIM
5hKjHRwl6bJh2roDF2kMJC9C7kPUe2x3x60bJARky6Q3SZZTYIh511hTPeisx2/4
sGfw3Kl3DWWsTKnV0dU6HT3zmjB+IVOdSlOH+NgvBvpGgvQdZ5H+X090b6cuYEgT
kEINjjckXCiZIGtWg7Tq1Sq31cdxHl9ewbllALAxi7CeHTR3iYai1KFMBoNksfXc
WI76Q5JQpZ2roLf5AfKtP18vqbTmE7eui7P5ObTvypyYkm9f771NIhp3lVLFjXsS
KGMz2smloXvwCG1bzfVEUSMpwEIx+elsYYo/Tx+SbLRJoL1se+E+yidN353TmQ2l
eXk82W/DjrZQfejzsmggK/rZcADsj2Oz6tYuvANbsGfwYFdb5BxrrmWpgq2KMz8h
F7LZLVHw8+CNZRNBra0X8KtybL+eCN7kCOnlTpnBuZmP5KW8v2XLf2FOUzs0Pjg7
Cn7bDdkU6LfMUnlQGkMucNMhMpEBFNC8HkYCbWefO0vlF2zVp32t+VWyP6WHGN/3
i73EkOYXJDZC1jtZlzNfe4OXWSGmj1xW5RdZdM3BpleDJqS06JKZ3SBFgbZKLNnF
o4FmxkrvPxVxz1JnzK89nI9PiXLQvlb9Cw/VJzUPMwAjR5yMGeHsXnsE5ZEmHh+F
blmYG2d8fTJwHsggy4uo9alXwc3V2PQzP9ZGJ8PTyw43vPI8WPtuV2ndPSI1Lmui
mmnQn75YRH21dlX3ZaT1LNxNU8WPm4OR5FjwMXPTQ8KOFUvKx4+6wmHlJZQ0Y6hb
3nTyfTO+aSXOB4ng19lfIaqTGQf0RPcAsXq+wu/W/I2QMmWxWXKwoKnZTsFkPnL1
6o5O+XL33T7XqElO4PESfoC3SmXgMg7amL1U25khK5WM563+va5cwR3qU/cVNjRw
h70Cau0huVzhUuxUl8VwFEogASoud2n7n+GmQSJrLLllYx4RhlXSUOIX7V0X+r3a
wvHHvNDek+RdCf9nbdfrj1wdJPSJ9SiY/n6pb1uyoQSVcepr71BpXgTFjZFbr6R5
ZJkbAS0zlvHlkllV1T/GgX2UmIW00ZDufE5ip03wOse2U+CTKEY6Jcg/JJQwSnjL
FCx5X3yQ2w4PpWcQACIj1ArsJ1WVc3r+S82YD7KhSpxxEVWM+NFbgDxtkoEVWfSD
cs/14eqZZpeH23Uwm12wULsKKD7a9e93sQ8b2HtoVUzvCnOc5JmZfrTcuWg/wz/w
zsWxgZIZM7kckcc2UOtC+xO9/iMW7sU4u/zIyY9rfSqQUwYs9qH3yVgLmL8z8rDV
LtDt9cD0h866mgrzQbrc7nArXoRKbuBZUC9QJ8Io0H5jqa7NpS3LZLYWSEnGqC1u
JVn5FiAsdsKV0VjW4yT7X9/Mz/SYC3d1FwBYH6U3y150GGKcWXeiGGneFvh+yHhq
QrqXTX4O34K6Hs5FY/DsEN5FJiLlXGepGsL/znJHdrzRUpu+/Drbryy9g0gPSdqe
r9ITOa6RiED1j+lO6D5q0jlQkFBA8sYTrSonE5IDQJL1Gskf2up6Kw+iGErbwMVE
lVBW/acJvNwPRMpdla5CBMuOh/xZWR8wkRjEI3q40gsnihNPno89yDysv/06NKIE
0EdNRadoxTEuxkzf1xXSrazSMz5ESV5gW9PfWvXMt9QtxEsjrrJx5/SqIjE0Nl5f
JAZuKb/FMyNOHPiMT6x/P8sST+R2fiMu744S3HuIGscaBKQknmiKwMTKiUI7J/A9
k5oiae6Jzd8dwAI464D5+YmdjPqI5hK6TCZ+Tu4lbIrPuiZVYkbgHGhI5GEVn+3z
EwajT6/7+4Nk2ZdSSMMKLeGTWhvYpJh2DSc+xl+kf/s7TBjzM+CyOfF8kHP7rUdK
Jhpo7D/mmj1ioGPWB7ZgEN4yxVLLey95COD2Q0atQCo3OEKX4kGjtjsdQIeizBa4
AxaVJH0GF6DjjPgHE4lqlUg3OYToK0fy7VoZ4IZclakqUOSyHODtBL3RZLgSGyHE
WGavXz46/SoxuOB6+siLnNhPElvMAr/clGZb7uBAvqAYn7vEp92atHguipGF3fyx
5BZPN04XbUYR5GPc3W0gQ+psEuluqNsr/mmNZV3+FDFrDnvNW6aPm4BnuqVw0W7e
8wEU8G1gEJzYch0arpa32AT36SjI7MHpVGgHMwAUmZu4lj/s4BT2IAW9FCs+Xcxt
sg67GV4A+hJeAl4ZfI5t8ezMgwiIGYmE232rmjVRK+elFgDVq2kq2hMejDHyHddM
MP9e6LiNJt274yGPLvtUcSFe1KYftMY1QeW4XW4urb6FhhlW8fr3sD8O6XSlWMhH
VOaKtzv4dpNfnkyTKeoUMcGOeSlLMqEHXX1qFH5J4rqza2QsA0fbzvg6c0Je7PON
11ld3xHVuaKim/5u01MvX+3ANh0I3ZS3sOz9H+LrAHmAJOt0/iiTnyKBwrGZUZtn
zENghG4q4uYS+u6pLfo7qyFrxADpurxANso/inaIsqcASbQUhx8kCmFZBl8eLuuB
dnpwL4u9DzyDCiTwj8O7zdjMAmnQeDxZcZGdmFAM20PKgGW3jdl3Ab68i/m5lEEP
vKhaPsYAOFgNAgnwOl1dwKiF+rWTXD9y2mQVuHEEk0F19D5Q8CmJ03/YfXeuoE5U
z6UePuFWIea+jxD1hiT57boQnVDJSMdaShQX6xaQ8E3B2xLmiqmvpwkCD75FknGb
Sy+8wstsoUT7RJoUhVH+KmgssQ8YidIyQVRvSaVSRYf4GpyaJJtEo15qjOobHUw+
3LUVONSy0g655naFBentkhnH29qbnxQhAfzvCiFtju2dWq3dhvl/mgQ0w5rKes7X
Kk40XaxRatbTqk0GAhmKQ86141PQ5YHn8J8+3NTA2dDs8ZAC/L2gZetyCY5YQwQW
RajipBjTUvwuH3oTGVyjGCiyiEHoAIb+LEewAIAp5ZMpU23xwnqJJPwekb6Eie1T
EenKzhb9JDV/x0i+agdRSzhWL/2HDBEbMhm7fKn+OgRYJl6YgwEEvJfXFpzhtlsp
39f37eRP1yqLvWHAD0367z+Wch0SFVQfDYFB5NlHzmSig2OTogbN4POFP0r5Y+kO
Fvk0Y94xVLv9aVPacqLlUZBvozgH1fdiwtE0nVBRuokTWGWqTehbalgxk3guX3al
f7/x5Lf0W26Uxk+vuIDV0beBsx920e2U5mZ45QnYDgYgJT9u3ERUJVH6+F3tOeSk
FHK4yhfmzSMlrmvIc765ebbKNTkm+kcYL1axp5OudzoFC+Nb7qe4Y282w5IahLJ+
JO+5eMfKKwB9WbmXVMbb159GWT1BlbxctDAXOM0st0ziZTGsukUbkC/2Lwh2ZgVs
sPxgpkEh/qHDy0wRGN10eR2EyhDUt2D8wd+V8Ym5jW+g4St/UL2+wGEb3en7/lpe
rWxA0ObeH36GxehkJVJegCcMr6sDl+KuoZq0YuZu1rfpqNe+me76PZheXQq0nSoR
5Z2p86HFU6o3d8Kw2vge/TIhDuV7bi021dyI0GFmIPCKtKofkR1q9cGVemIo1p9x
abyEoHIod+r7ODd295sh54vsx/6AeC741bd9XqrkqZuDzOXiOGCcYCBkWAjUuSag
GRZYLlluo8P8t4C9b7fgMXGcyOeWoBHu/qB1cRKbY4kaU0sC4fv/bjKHnaQtGdPW
PxQkVjBtELHApTUW0TkeQA3xYiET/7RXGPIoRTH9qrEmNnkk/eG4fmraZGukRiJ0
RY8VUknqGIv0OSgAVu2h1MWJvt4tyicRyHbpi/RhR9LWflwKsbs5HN9vrRQ+zyYB
huCCoGEThCj8oM65yzILzdcEwuZ+ZfAqobW6XROrxoDCIcdCUpYbRK2/Wy+PPnC+
WiQeuiDyOVI8dAkw/+g9ckYgFvbhzRNBXYFwkh3mGbdssNjFJLQ383b8tW/GxyWc
VCLLZRrp+9/GLppNnaocFq/eQfqaOeUiHehOl6KNZFwp6TVRNr4+yLb1e3CYUlxS
loCUkUDH3tgjEXEz2+Xm5sBgAftMDI7x1k0j17VsZoubDSAhcXL0a+kYa+wayZPv
GN+TwM2ThFYkiwXZYZgbxpHL/5tzSBBh0bAjpBeuMEBibYHad0JQ8aj+Zpbg2VFX
xACXtcE3PVeTAe8Ora9c5YCzCxkpT0KXUdinhOCJni/753rVtAC4rTcHVFgEuWc6
7apXIVLOoSAQbQlUUlJhdgJ3+0QSfm9GU297UXiIKoutglrtguvfCe0vKYMANZIp
sGA9RarxpkpmGs6O5zakbyAcvENyfpVWtthfPjVtv7vp1MfquCXR9EgZnrWCwp/Q
C2z4IKA4NcITMG4UtL0CEIfiTip1owkkqR404dFmt6bI8IM74FBV7rTCU2Im3elO
BszUx89v4msJZCLiLnFpNiy1YM3PzzlWYKJRjtoHtkYg6hnhnneUyga7TX0Dugk1
mb2w742RKBphM6ScdWFx0mQGHm4eyXZ5GaUWwsdyVyAQTKkHXEK0O+xvSCgbDlt8
er95llIvGvNYImqkhSRlBvQSfybP4I1ktBkWs7Zn7C6ERIZP3DZNHt2J3XUjAYK7
aM1r7KjZRalN6IdqXAu5cYUEJDStFMGsWggHwU+ckBAMkMrALZ9HkXFx4Vg4FyKy
6FHYAHvG/GsczZ9bhcMjfsisQaBDwNrlqjiFHyik4/IVX5OvDNHzYpHMdmodLE/Y
byW8YVECYDHVTiy4WJSjydcf9X9iE90OUUqCN+lUG7YJbG36ixFHntwKlhq5Rby3
OFAXG/3ylWujcxY9QCYTpTkarKNgbiNP9zvvltn+DcfJ0nOmHGzw2ZC5+ouNXQND
uDrGCb+lBAqbXvntEqvW4Racy3yWbp6EuMVkws6K6/VyyoJLWl5D5wGXI63xhL+o
zwKoDqSzP8L2QVNzHcTAMmSnnnPlbRnQGHk5EQvh+ALj/kmjBGQ1ei073scaAjTl
I1sfwFv8KlI6aY8dNcG9nYwAGWMYWeRgyeeTO9HMczNIyhMzr9HDI1g318ikyyMl
U1z9jXoVARfqOPTp358rNnMopU1Ewi419SKF2q6pOjAId7OsEs8qj7fNrx68tqC8
V/3vVbYsdx7WWqSWk9GwYt2DIZTymLvhLlhqOJGVWxwv+4xBoZk1JOIFXtRdfpzY
CmhQ0srhXk9aMklvoR6PyAAGTmQ0x/nX2CEBjNdNW6Bd+gqWXyLgaaauplkznKQX
0H3+UbiBS+l+fox/Mk6lIe2+pIhf3AUkj3c4DU6LdpjAS/GJ2i2veX8+gzOjvy3X
SkIYirQ1+DRi7nSZ5SKdC9UEAouNo0hsCGfPKKV31hnQCxAIQQwxY5SYsCNDPirk
N+fr9QFPJr4WFvbrPb+dU0anWBbI3Klnn7q06yjRp9m0YeGIjydLstXrUWggpEon
1tyH2HiRnYNo7puo1UMveBK0KMmHE+HJBDrqsdp+SjSewCr7fZ84shntEjQByYwV
fo6p+Fn+16CE7OLswLq9xbEBPai+VJRdyAWcq4V0HEwS6WaepgA+jkLBbWo/xt0a
f92X+6QI5i+Yhk8knZL3k7jAuihCLurEyUmbZXDEBi51thk+a3/kCYQXg0lLBLLY
dvgIUQaEx0aJSrtzBUK1DLAXJdfufB8g6TMRqeTbVioohdXDoslsmjJt1VdVfRVl
rjApabHyHCjouWdLhxdKCx4rXuPpZzyRw5Bw6QUlVc077RIp4ierUiTAHa4OCyBu
Uo+ik4riYHe8P5M/E02jnsT/DQaiw4UVTnDdyDdDgXuKuGuhwXRB1VbacRSGHF3t
QDJjqB16K+PE9VBHVfLZ2G65s7DC95Fr80OFc1Dsek9lEY7wg8aSK2M0XS2zFIN9
vmgQNYznsTpMEjC5+P3FLGpwfnZVJw64KYJDccGyADYVPaaChwCGKp0BGezjPIU9
Sod9m/bV2amdzNCtvmVr8Pq5LQ4U+E6KKPtrvOevRuplpwUUr2sUy8edL0YlL+qt
NWqDSvOy5O5/hfhLoAV8uhzbNJpxNZnvn+lnAzfejWunBpJPHC+GNkjPl7xpRrSu
V52gMfRIyTOp5g6Z6txrshbq+/scBk1dk14KhDG4n4A+khEM7NVFeZ+1TDCz4ehg
oP6Avlwq5n5KNdsgzarF75vbC5zSfdNJeJ3bFsL8lHLCPiah1o5D8ULphsjUblJM
EPXJXrjWcQWoYItIMxud9vU5lBfaPLkmSpFqC/loIh+oTpYbVTYCB59W2csbh4Va
educSkjL5FsYAS7p+yZbqp2L8EBbLN1+b1MDisePm8p6WqXMcKGFyNOVV3I1jbxY
eujNXFSxLKl98rNJfWaJl4Tn+6MGBHe6A6BZdkiE4ZDr+Wh/kAE6zOBhIZQrB8qp
06l52rvKj+V3SJspjY3CQhU80BlJwCto74xPKQj4IlooKFfxfInvNEBz8vxxg2cW
IWfRijhwozNFDzxRPaBgvb/IaJTPH8byjjymD3gAmwwV8eXFfn5/gJ+Tpd6McYHi
yBR4d87rmm3wW/g2dDFBta/UVw84HLz46kiZnwSgMAAouYft18D/1erwVzGACjWk
dQZkTWOycNVJLgqxzUVUDYyhaDYPaJaRQ5w7IW+87etY/vUekYaJnjx8k9847kJb
QncWKt2Wq+UUQLTPSQ3XyeA5cm+8LUIbXx1OY6JrCMk4DdtqTZSuDMObHJzwoFDh
nj3ShdHNSctoi35gnbdjndoM3XW6YUqcj3gxGNGmMQPHO9GwDn4zL82GFCKsx8qq
dJUG3NqBnuyXr7FOOz53CyhurltgvW1Eh2GOtu7H/lZvtxtMHcBqhEGQbFWRwsZC
aMMQ5PMmizDklJn/Z1sFnGNO3YdT1bz8MxDl918ngfX++QsYGCKSJK52UOBEjq85
X8mNhOSSLJiH/OQEP0QW9shDVNaU3qitSGlawdcntSiYV+NzwQElVCUClHPJbL9S
EOk6EknIWmo/YeIvmIw59h2aIW5dwX80ePaNr2wOeCie6KyA0NOeV8HeW/iMhRhk
MLSpuNOz/9NDwAEw1KvSKhzHvmlu0++JuncnIHZ6kCr0VhT5d9Sl7qH6zeyhD8Xt
wo+RJa7IcGcLwb9lkNgjYfhYxZQiAEAY9cTJpwFXzA2S4fZ5Q7YF9EeGpva/D/s9
yiqrjyE8Ztyv4LuJkMFFMG1Wxo/3sHRZCyZ1qAQMkgsTvMCl4/DNmkmXBW4dEqGf
Xch+dFv6gWNfFwuuUa0tyGfankwoAZHcNzSL4B0U2h7ZlUJuHfasPY1xr+aPnjA/
ZK3VEro/yRWRr0t3D3SKJmZARKni4lSXUPW4ZtZE2i/1ftCvM5HJWi1MrvD035ZT
4Zkequ7pxgVNzI4PFGNtYcgL/mTKSXC/AXWaLBvgbzWrYQSsHl/U470RYqsZ493n
cpUxxOw+lzV//u2pPY2tHJOWyLUG6xOzGMFnCmV+4leIGmc5/LdlYiFSrcrQGb+k
tEmbnogijUdycXwUjHb7ST4IiesTshnX5UZKTJriQq8cAb5KC0WQyurx6R4q8rHV
bs2DDtqB2XP44UUmj0hy+QlZFXnHoBbVXKJ2VIG3KDku03GftdN9BzbI8LxW233n
isU8lUVcXZ7GWuxE6RrUMsWusaXlcshIrUbEJHgiNftO5snlII4wZuecIC5iYSfX
Zyyf1933KEFuq1mnN/4zxm3w2g6vay/W1xvKYmR7tyqXyauDiKAYxMRHFsxaaEl0
13vqdwz09XBFkrv7np4QUkZAb/WnP3CFk77mwtbPDG94pGfYTlC7i8LFGto9vdzL
SEClrOzoX5xwMyt7Uafmt1NnUSxg+3h9uYudPibfQt8ubkEMgNtN7aIJcKbaPdpI
ue5n0Y4hLmuonmd1WHttWxdefEN3zf9oHbz8EghuuNnthCd8sDRHLfIviYkBFpgO
V5mAKl98vBRhVXCOt/spSJxSmEbni7LxOaZ1VsN99mduJkFsrXdKaA1+lOJ68uqk
/WR4EBu3/aCqLPfXlxH8B4EsrEqPRNpAYUDXpz1iLU6aw+q9sOrfWrA00B3HmwIm
5BLcHQEUFoKCMCy7iIzHwHr2A80Keg0QKL72ZcI+saITDIU3/Xq9j/2PiMyNTotX
j0La1d9PgzsSgoAHXCtGM6YIyQfE27bsqF8DJcLfHMGEUo6WfraOL8OlCM/C9N+0
GrVJg0EApfRzKzv+WoJqrfY2nBrxjR6ME5bgn2WVs27r4iCuSHz88xDC6vQiMfD2
ZtzFpb+42b4o+YRlRn7UNipyjAn0qv+fMQ0+dGP5yZ+P1ThRedelUMGNQmk917qY
uiOlypauxBo1ok5Sf68h/eQiyJFDMv+h3g3UYtQNVwolJilC55JXgRtX71ATKGTw
iYMRFGKdVdAPCWKlmPBV9z1j86ty+plZP2mJ0Q2nVGh4f3RdaPkh7a6wLpnX/zxV
7Rw0rrfxExqGZRdAEeXzKnbSL9IIFQ19oWs7oXLqR9pWc4JwWqPYmUqSuYG92ROs
G+OA3fPnryNHUiyL+vYYI76aTU5nDTAm6qSdmkcA7M+MfU0PTp6VV+ZUNwhYnX6+
216KrOL1dp/50Cxp/0JfJGYRjMjgZ0yZZt3S3FnwPe6RdkHgKttr91skShOfgXur
nWVyYcUCu9qc+Ox4dDWqQRHQ/49OFM3X32yAbEZoQbnI5nQz3gH2oOWzsVH4t5HE
u3U1ALabyF/+wuvTgthSZbTslnl/OosMcE5c3IUTXeZk10wufLgo8ZA0cKsWvf+d
61KBxrrrXNwdG3x5kR2rMwymo1YgL9nzzccct07qCeb3J1Urn//mqxaxDhXje2WR
8PZCsM4frTtJmpMwAHdXtG7s1+bV083HB4wr1Rf4wt8hJDjUpqGzpJGX/NKRjX6c
phyHFxDE0SULEb3VJzVbCgeSuEmaSopcO9iApXF+FKHa75rXayXwOxeoZy7ERyWJ
MaAlvGtfXiIvGb4Wo9mL2E/bY7Jb9xE0C+IVUY4xZDKYLCv+I/qqvzWmtL8pGlhU
le0yUu9ZLvK21nWew21QYGCBdOllNYP4CnUvNXV13KZXZP6Hy9UZgo9+EolLqvVU
V+c36uoBmsovQOFdbwPBgQN3k5646G+Kj020w5+WuP8k7RGOThnsr6GxQtmBUr33
cgsPp/m694/RQZpKXrTMTAzonaCFF/njDhkLRbLSFn6DE+fBtXf7qpAjoHk6HhHU
NWxee2s7NusAx5Ln4QoMGhD1IelSmFy0lEQjp9RwoStjDH8GxTwou7yuOK+xHXGR
yv8GOxUYY7PgNL/peMuO/uTHCsbQptWNbbf0gB/Ehn/972OFQNKMIDTZGILP/QMb
fOxCpgdiMWB2hItyHUHWsFbjjqglsaKhIoxoZK/DA9176qIQJ0vod6FKtL3IBz3/
yxULmr5frdFS54LO/SyLAg0qTgMx1GHYZnq6IRHZ11i1rQsyVbbGThInj6+7LpaL
CNd8uqid0x/DKcSO632wnj3XIi9TggXMzcAe5neiub7qgWRDLnXk6BSvIam34OfU
hDL0eO7nuFFS+WmuNu0A3Ql9WKKJqQ66NPpUcHPBbJv5er9b1nMqXhwsqZKz4R8M
cInxhnFJskuTISCLro8zFcybjJYk6EXeXL0KiY7HBF8QKXICqSQtKYsPxEMMptlC
1u4L98kXQPqJMKPP1UXPy+PXaCBX5lvY0D+Hd6vKfSKDucuRpaTNtOPZ5G6n6gqn
ORnWiGRfFQ95d9mAeQTIrLnKwk5sfEe2LbCm9rh0Hg9gRt/jFpLuejuwft9JMQ77
RTlgXPpoSq+9sQ69iUGfqFiXvx88lNvvGcxAgwgMmRB1O1OL4aVkBukdlwzR5Aar
Xi0u55kPVcGoSao/wDEkS6iGqJVvGOiW6M58XrSHi3DHRP+A56UvkxJR8ewrMLjt
KgzSqIGC6GUahE68uOx5Et8vyvYadb5WnOiJR0SqKqwERDmXvahzXai+i9gHVFKm
y2T8yzFDlFhaKkrybvihqJQvyQFro1GYO0mfnp3WTquovzLaQlyK20C2NmVJjFrk
Dqxlw65pWBPYxiWv4AxKJdERNHhMDfLzpsneLg03r5IRo5ZkqQJZ4V8VKTDHxOdW
yOpmFFj/IwAPZ3ncbqCZbri2e2dX+lAqmaY6eN5hfSGamJsybNRv/DTTOnLIkfzm
OdOTaGQuDifog6dFEsshAwLQKmP293nOsm/p280/nVwLwNcjUAFnFxObxMgJUuFJ
6xv7x0rPV6xwg5NWWyuvXS+fUbCNCincCoq0QV+92M4oh2iNLHt3lPLAQZEjkBF6
xcCewZn6OS6zjBXHEYGGrTYQaBFiPpHvkCPJSgiZ3r40ErXTY/poELrdvk8jZkMH
q1mFqVAfvWBb/YCHzRYBesrt/EKgLxos2e7mXVh0GdO/3qsZKU4TkfTO5YnkiHrC
ZVpSH1zXIPOnRWlAe88U0CZdwudl34fbAa8Hp7oN9wKfLM301Iy690IFGlpsE9eN
IAZvDDJK/9k2T7pUpumSU0wNAmSGOczBpgzQrAZ9Mg6/2EdRbjt9MigeSlYXVICq
4p2NwAZ/pgGeqGp9qoOoTXbBVqx0CxTL30acJVacZNv1LPvF/fPvE0h7oj3IGkPG
e3GdCVSPhE4DFqNoHJlJ9ynuvxsLorSiyGzJV55VGbqVv45st9JPXtFLwpG0DREa
hYJ4/+IsZ8pUZnzL9PblkaUjsq+G+HZzvtZy1q45PnI+/dQXAQFRbYK3Q3KVmJ2d
N+UGU73cqoeMh71gH41U9Yc6+jM9kpRfpjp5rEQ8KN8A6w19wy2PddI4xghHinAj
pVuvpTrP4L/nhrIpgP3Etn88HfrkCCcIZVeiwyc5q4VtsSobBXbAB2H3cdCizY+W
IXboJ2/0WSlSAfYuSERoXgVoOHT8S+4996hNZQFb7eBpqvVovCfW3deS2LL/CqT+
lfCemS8uNsSiA4fkeAGbRHbsmChgW9DLiI53fDUIVd3wVzLyr05Pca/QJ2aFk5hl
LZzLcfOv4FnywqKwB/eGy44iPT0+dn6q68qF1xe9ITx3vPSA5TpDzLruEs5asbud
NfOvmihgZX1GpOEjT+soaD5rA0pC3g1Xer4QChjFIODjQtdbG7Nfwrmv3CcuISQC
ZUu20mCQPBnjpGm2WVB7lHS6XAiGbcPbPmZptD+fu72w+XWrTRwVYooaXTYJWkfc
K+DKJrbYJMQE27TuhaoxDsGaXDZYb7gVxYNPrtcgCGuA5TFIcBR4vYt+4LL/tRSw
J9uKJF2bKQT+/7x//BgxxBY1OreOBgxhNyLowg7RLQSszDOCOKCtqDFAhie7xBHO
LDGs1EtM1RMEVujC5pC1ZhMc8H1Xk1QX70ITiHIxRGt06UHNANqRTKE31+IqXE0I
hd7hLtTrYizL8erg8e+5vL6OcYWT3yV6lXPjyrz/D8IQ6mVUmdoM4DHLjHbChw6Z
05d2xWxShwuk6zZFf3iilqYKjf2vyYKtJ0M/PvwJaIg3Pd+0IfNbf9LZb66QJLY7
qaRbbyVdRGyBXlxHclaNNYhe6LTFwBDmop2AnxTCfu+k65geNB/lDVZAJSAmvMqK
Yh7CW5HqluXS7bncVvyu86m1YsNd7as1kKCBy2D/3XtCQozijG6o/PwH5vX/D63F
BNF+z5sdqItrq8WWZsP31mCob5ZhKcPv02w6oxvKbCKMV2O0nTQRoXJzm+48S3Nd
8tJ50pmM1MzO3w4iC8cWbL8dPlw2UiSgk7YFSVe7z2gOzQesmkFp1zwVj9vTR6Ai
14ERtCJQQQth8plw0Pb1njUaS8e41Z7uFRBd0gUyhsUcRPa2oUaZeHrMHkuI15kc
8w4IMavt8sot3xrNw1wiO8/YafBn4fy/x5CfJaVt/LXSIOqobIe+ATq4/hWP3tlE
0CDMOvyJMe6an84yiorZzXupQdcTKxqhxedLDtnJbmf1Qczctlu/N6vK7dGQYdmi
pbVZLzERES0gZFFwK5hVQdpwNZayH44eNLo/5iIPwSvI79sbp5SHawSDcAXnWr+Q
Xv/FS43hOaevfv+1FNpN9AIPYHe/pewfqwN2Aa9zPh88a9nrlyKn+gzQgQkI25dY
812C4SWPJi4FOANrYQWAl3yMaAGtWFASUMbxlE6WyvPLorrOet0WqWcxi0VjW4wt
RAX1KSAUo6/C/tO+8Qgg1L2nI6GiHcsmXg39r75jf1mWKY/fhlaA6Z8fzaYS15CA
R5YpXdJppWFxFCeykn2pJeMfHtlpve+mONmgLKuZm4vNGa3t+7gCpSw45obQs0Y3
+78yiKU/kr33/VqTESqUlmO/wOoKrtXZXq99S34sMNDbCup+DZLZVuv6e+72gVeY
0mKbZQRp0hrfAuYGsoEFRtrnsovItpysgprhiSdxIXMI3yJF4r6VgMTm3iJOjsWL
yPZyvDN5c622bxMFGOB39gEuzdcAd+3wVczibPPimZS51S32/6zn8t/TnCLaClrd
R0rcFypi6GsPtllDScGPFyd54y3WuOUzIOjSZJAdlyaBFaaxcbEZfcWpL9zmMrJv
8hUa582zgOc17Z54U/1AQ9whcnS1lrYzneEUfXvZXxT1Ei6Yiqx0wueOmfrpUVYC
17Iss5mHBGhbIlBYVbkXJgGvIx5dnfja7zlTKRwtUVC1RBslzZk30HZPRpOPWSMF
Rio/4P1EiY8tgJdB7bPLpJ4nGiwgbeLp2b3KzL2gLoVSASl50RfUX5R8iyJbRP74
p1/YKpKbFVg92n8U8me8XWyJoNR6hWzV+5Jj6klhgG8dbC6ggj5TS4vJfpdaEqrk
eJDxJkPWXSr3cooTcqqsJBXzmgZAR11MSxEk8BPF28kT2pIDBFtVyqDnsJvQzciZ
gNUYbl3PQKoJBZNLl+DkGZm90nO/2IaQbsi5D+O4dP6j5z6XCJcEhph7mOJrf/fC
jMU4fM38wFZ1FJsKlyZB5p4+uQfan0i8u+5lrh5jYsJ87Qc9H+bmsVYaX2JgSyb4
bIHQqDB2Vtv/FJodiEvoaeJ77tVDh6AIHhGWoG6mx74QQmBrQ+zDBJaxM4mduTh1
GrIrk4W3b1WhWo5E4owMoVO1liDf+zkQOrDtCJ8gp/9pODW/8opuQMiVEbkyyWqT
2VGswG55XPkDtIBXZd/hUFoU0Tk+7wqoU22I+Ih06U+cmtnX2cIjoxOXFLThqLvH
fb4Ikmdgg3PrzyFeAgMUaPzVNmKOtaeMp6mSlSsbCbrXqjcWynppSuvHmMPjWXW0
Y3eWPJJ2UCEweo7MxU/ZOUs1gKrJxcT8hQw1Sp5O+xWay5BXrJ8tscH9b8U/vsuY
`protect end_protected