`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
ddtXksX2+yylW5zu6QL2Lhnb2d1sD00763mmSITNX595NcHTEkwn0zB1Dry37fOW
FufOhVzEJp80NC5qZ/+F0Vk7Ik02dIR0elf3clrjeJRK85K4e3Hoo4xn7YbFUIms
l/8VZSb14+JVGURjfswrIyCUotIzlzVYZ6gzoZwDXIi5gQIBf/gI+KxNXPaKV+PQ
Ufys/12rjO6aI/pPlqSm0hCvftmBcnezN2hk1UeXgOIuKZnogjOsf0iJVX2aOOWE
6pD/psybjbnsNB6kH5uFTA5frkzIzkzl5d9+YDm9OyC+k84E83I/7/j+rk4L2dah
QJOvksSIzN867/4Qt8qYTQ==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="MvBXkzurAa5VTw+1JJ70nePUfoQXBvZOku/SMmg4TwQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
oRtzZL4VJ4iwysPsC8SXYCzXS8Fw2gtZTOskLcDV+1B9Nzn1zTyNtlo6lNICRmmK
ZRVu2BmCc2G+fmzynYlNTnSa7C0Cuel6FYpxCBlOuk3OF2tzAmLAuDyOH3Z1Yjzk
a0aHuoCdIRKv7BrZCdALt03JeUmXKPdOmIlkVGFl8yw=
`protect rights_digest_method = "sha256"
`protect end_toolblock="Jn9CQpRhJt4rnzZPRk+dOpzAubz7omckX1MrFd4p81o="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 6176 )
`protect data_block
gD6l00tciPUa6pDNTk/+t0OO0nC/UTtBwLB41d4inuAUA3i/ALrNyoJVcBnAmEQW
ptbcNp5fxEUJjnOxnedyZEuEBxWRieZFQnkRdF269oNhQQeU20GgSwA0LULFJX6C
BggG7x2+2aJxt5f2k9uKWCPsYj2Z4xl/ZWSEoTOHOuAMD42AhJSeu2ANEzfKoLtz
HJuCCGcHwOmwRab3dHBXXk4XuDjaeCr5nfQ/156SRGh0fLNFGnp7OprbjneRHl6t
hmCqvMoVewIpgIeq9VP0M4KvSuJgcegWyHxYD2PHmRhlzrsCNw7S/LTjrZ3SdQnE
3UX/N+Nvb0q9uowZ/ry9EjluEQwGHZiTlD2/jIIr8ttssbIWJ98NnqCbz/eLoVal
2Qgv2s3W4FwsJPCPY4iI4yZgQRwxqkhmier7diYJA47pGxDgOC0NpzFE2lvJJdvZ
0QPYmnz3GBXoBHlsedVxjYUw0xTA8n+uZwTzdZSYJKxeYdqsa6qUHPcAmdu4ZXKA
LQllSdOXFbK+9uVHr9KfKJ+QGqnV7IytXC/B8Tue5Wto0zCYdFobT/t8dlny1oEc
8IaMADR5sKVCBTi4GmMuD0WD42GbaIoxXhjsNXw6WrcAYI75znlJm6vqynItSEVu
3y0cWHve5uWsE6YJInYqzYIOA59Ubv8DnP8TzPKzx3/5QKZAR4ygPWPqCeWDMGve
5hf6BpLfWoiulZNQXq0b4hEAkSF1m/cM5WzbdiW6J1jlI003R6y8bYcVNDqFG5la
nveV/6vMgfVXlJWKESFjtymcVvZg1gE4ikYdnMAw42X/QUvl6HeqgtMZBLVnh7ZV
KtW16S2fEpUeQr8+AHTzHKYv2OsKqQ3V0zIOQ8S22yknEuf2dsNcRdATGLC2lL22
Ht3l7RSh1urqTK3C2tymfXZ2Zh6l8vK+aIGaOfAYqAs7+9PsBROKpNR+aFHnXPQa
NOwtknsUVo2M0coLDlepnj2V+4DYEWblXNMUm/DV+TGW0CUbjcyZxw7QWX+2lWo0
gxN2Csq2G0//HCLOR1X5wNehkCbKmgRajLIMiHPbIedjbUeiJ6WVH6O6fYoXDP+Q
hnsw85czftS8C9L70txFLwz5DeXM9tuX8nEBGNGK94PxuDvXPoz7rc+uNbS6U7Tn
fGT/ndKpjsn9LWhEjDhdlLrWOqfr41RipdKvL+6Sn8E58MJK+okdDpAz8OZ508BT
wnAaLbiMSkKILAllG3bxsU6VL0iJSSuZ6k0Y+QpzmXjWuGYfJyoBr5fF2MMhc6nr
tmujKM2OqkX6PDKc7wB1N1tQNoXzvp1k4kNpDZFh0vmliT/Xr8ML6pjUttn9phuM
kf6kXm/sCVhLP5gohokccwhM7CU6h9jZTQBUV0YjA7OCXtO8zvi5x1vSAoQEvzh/
upiBPcD1h4BwU+uVpfVRYVBE+2czri5rOCKNEpiBQuWTJMtxgD+7tKob63W+TO0G
76eQB1v6qdCi5xyEr19rNaGIlUn9Mwb93x97tYQSKrSxijDyRUC9t44rMIsRm6sW
/ImbYvAMZQn+qGPNaAP/MA6NhHhQEs4rqTVB6Wwtxnh1MZzDwdbEryZD9fp5DCXP
ia+YDlsFyI4w7BI3mA15OuF6W0gN6aVN5Z7SVhYjyhRzBEGmkT5D2B9pB0tTehLI
Qj2djLThwHJKZ2IGrmMpS+q1jIE8nfZLtetbtWiCwqwvdCCiJCXil0PnPxxft9lO
WDuXVmNx6qkgZdsXaiKDY3ONkdm/2PAzRxQ4023tZst5XErKOZht0yK3egW6ylUi
vboe+MfNxgX5C7SgRihhdPYUv+i4cicEliGDcm9aW2s1wscdspKagI44Co7+xwto
hveMUP00WF88/p9roYS0IoV298j1GZsRnYpkGOA42moBlHZsSEGX0oFeXqs/+f4y
vpbNRj8IPcih67c3fjJx45aks4BRTTEVb5lbBQT2dfdgxBlWFT3UH8u+UHJ7ThHN
zAobXSKQToH9weIbHHWYtJkdRayEPMFFzSbI8e5pQget0C6kRfACE79ebkRCucIf
Sa13LORG7PXneWVM0Qro1L8xhSdCLxP+E8RKr8hppmYraFaY1qQOwdyB9s3bXa1p
7tzwOht7zYKUkA+oDLHPzQ7z/Su/5kRfyGzcpppaf29A15zc75aP2X8D714ADpNG
klmxxsd56FocF1vO+BxV4irgPHYqTAdS7ZtF3fNScA//0FlzTM3t+ft/OFw5jH7R
is2qhLWTlsC6bd0vjyqB8qSVoGanIHMH3Pw9r5ObUJENqOLPkKg2kQuDKeM+jZmQ
n6WLUwnNEt4Y70I7T/lUQ+d+QwWeooLc+BKUQldqINkWDWZ4ZLSJodl4ORoleG54
PL/9NhT5mT5tcyIimiLgB6ZotW9JM9R8ZVmMl0izdiJkZ2sMTFGVL80IzIgEYi39
h4rLbu8nfcx/s7QQoAeqiKD2ZF8geUnqED5kTxxEOINHNP9jtGNv8U9SnajR0VCt
Xg9t7w4dEKOTPJxIz/itvht2IBdzRWQ4l7gmoanaH+qZAsioGrBXAADbTbYaJqEH
VM64vVnjAZecqkvoSKmEanzw2AfZXvB7wCv000TNC4DgNYMXZ8yjyclHqYCeV3c3
ZOUqVvSF4NMXyzCb5hsfUakzDkstz8jBn4g61NkIfKbUu+61ucXq4RUqHV7KH/LR
/k1yA8cR4vIJOd/A6Ji2s/U5M/7wJoDAxmI6fisuK2X1kMyHMDrFw8ZjpKnYs5dg
8peNuhWKtOKn/puk/8G2cUKp7zruKGkkAKwwox/+msyoZQOjHA8Dp4bvifN2mskS
0JxFi6VpF4wfp637T4nV36siCZAMF9mdaCkP9nO62VNoYLmkEXyWbLsex/biZBQb
tWVkMeDxLmBqcFy12F5RjwO/kObOrJKikg4KmNgXj8mEq6VJYVJvWuhWikcMYoqy
3J966N9R8mYYWxI1w4zAy33XKsuB/Xc6tdHrcY7Y9pw2fu7saNxzpaR5UT2iCS6b
8pdZIfuFn/TT4ybwzhtPhawFFW0BmFobqdJ/2CIvcEXNt/jsTYYH/4J4iS/WUq9w
TVDAuUV6PREFmx10escvWT0BtCoAxqrmaRrkP1gb6HwAVwbCWIcwLknJtBpQsR4R
jqgR0TObvUlMpKjczpgVkUsWeqaDmdWbcc4b/KylWpU2cGP4XIhg/H5e4ypWGXFI
muEcpb7AlWOSnBvjjVFs56Q9tds82oYozwVzzzsEp/nqqJ5Ou1ku2ON1nf3VsLXC
rbp1kCku1BCOHe97+bddDQZYOIH8gD9xUcWomLtwHMyovcSSA3Aj78PovHv5PQuS
rBNrGl4gpoymKvLKPVL3gH6ZFtDmdbuOWULEGlITZOaOFRrzHhd2tEaSX/XVdPv1
1WpdKj4jxAv9Dz2dps2pqbvUIAiIRmHEQQ6Iz2N8h7JjArQ81JCNoQ3r8VATcsSE
3HYwrSwmvFC3UAR47P7oaZkg0ZtjrXHQ9eA4SdmkikjKBlQD7tNiiZWugkGEuMhD
CihA8dWR/y0rOB/Km5DJwU1bitKjZrTlrS5CKjzaQt2hMn9v25aU7xZ6DJdhjaCt
GGZYb2UOewvuqTjeq8WrwirIPbVRSRD2lldeEP4y7sS56AZQ8gdjeqTeCBgh5qUO
UUEoeFXc3mUfkLoXbuQDp7sB4WlcmrpTN1QQ2HnRGCFIyYbuMvfBWrR18jxZ6+vq
5MfCP77Y0547adhF9BmWcgBhLxB6dXDkFFgJ2hd7J/U/iq9ZEP0QAGg09SQkkGQw
Z65AYGgCfwK9DTutq2VtiIrIEyyScDwyogKWpQE5XTyWlLs7/ER3voKgYiz6s9Hm
mXGTQWC2KxuYHQyUjg7+7rnZjdHbSi2Ed/zCV3TTjxCEC0jyl9ODQZT/DxUKSa0t
UzS0UN8j60/eiE6WLr+cWVTmGtqEEFLbTknX43yjzdmEigD+HSyuxjL7VictWeQo
I2TyEGrgzIjR5ZuviGqSTRIklN7k6vMNPtWRBZQm98q0bFspuRWJcHRlkcilFCyw
Vh8NnQ/i3kRwinYaOb3WPVMQjkdwZkWUjLDMlAfmD9PtvaCLKWycudaF662n12CL
zMipXMGgLqhnWP3Pqm7PSaeXo9v7xe4Ns881eyCWr3qh/JnXdOmhkKMKCoe8ubaO
ElBuaQL7VemKYbIqWGECpi47U1p+sU5Ya1//wZcFgf5vXTXeOiOIdjLsvNjp7p2v
L0g0gRzcxiTObXygBRJM1O+0t8BHRS92GOiyyGt+p4SaMiIMjrqwHHACDKyscyrN
7e0zDPNLIvDRMvuQ4j5M3lTIu0MZWnoxP4lWwZ7BuFvXSv0PX7xY2K4GHP9Ae21z
xUFqYVSKQcfnLujmqScnMT3c7aJ8qh69R/ddyUMPPLXgnN7EAXzrVIdD6vrwlTXt
X8qI7OwLJB+fdJwkGDWcVXN7vx8ABfdYy4Em3A8x8WL9uUBTmG656KBaGfRApSYI
PsgIcATsaW9Sa+9o04+aJM97qC9tGT6/Og9jhFztf0+IILyB88/gjnXDKvsEsIST
aXy2/uuVwyQvgDa1w4NDP3B9a3tCEsNIADur2FhJBIYhw9YTziSV0jDRgjt7xKGx
TL7kC5Sn+AnvkkE2H8zJc6HsXvo7JCYC3yx9iROQeQURhX10S1zHVlS56qds888Z
FNDl2+IYECMJUcYQjBq+a73xFSjHlMInoPUx001YHbYvWY3jxhQ6VOckNND9s3mX
LCsH0KjeYLiNCZLajhH5LJZu/1mzMBy8+O3Utg0TWX3jK90uTDju4POFnslIClt+
w9vct4Sw9Sb6VCKRAt71/J9QPAc3igYbwHkb+XlQ9BsnWc95ZffbOFeVmrVrIoGL
GO8w3dywbCV1t2LrEWhECmY/T6Ja/hIA3JoeQmGsZJVxKnwhzz3XzsD1718FQ7Jy
SXOvZXaAk1ZLWE2ipfMeTRzVOSDO7986/aUeoVgAxWiVVvvUVAEOTwV3PGgy7x6U
FMFbuZN4s7ovabeM+/1mHnZy5P/Vu/dlRj2OV5mnNSMnSzF7/Vkce22ZwrBhy87S
PIRhLHm5Fd5Jwxhf0kAVF/kcomSlSYT/k24zW9E8DVCF9pvXOiDUDgreUr9EOxOJ
Fo3ruKyMB0YecWUQ1fyXeiICOweK4Ummzu/5fSMV/jDbdM0qJWXVqIpKifYNdPsN
w0LkbcFfCu5TG7Zvq0Qq/LPWZn9PpskJK0+8cTv22b2VSjsMdrw20ktT+3yVO3je
Pih3LAONXYFESu3njg16z0O98KsS7Z72fQm/HnCIw+/ZYvm0dz7gj3ePVK2dq90Z
Z9FGbfQSU2UjfsoKHvH5FIgtGiUSnH5maeOVkTXB9MtXLRXCUYv9hiRMuoZzUj2C
dJXC/PBY8uuQYQ5uCyajaikXWyXHK3W69r2ugOnQptBA1rqFBcDF51lo++zpxooT
SgJ3ZM7Iz+UwFmRSS8ZcKg/N/JX0EREwNwwzMFNAiWstqvLX4KcdwoBe+vNG0cY8
mpHsyAjC8ihwWzLV00sxrueWoQFpA9fA/HtAB8l6jiZH0zNdgloK62XxY81danFr
C9CpmUv7yBjLwmOIn4tuoN3WG0Ua+3qaLpUeO8s9QYzYnR7RSABCCL4DOAdPCGgO
6Eil121v0eTUm1l5CfAbwOQnI1sSQAOF5V6zQh4EZCle7NHgRwgxzXY7DSSx2rqm
ljdVNYNiu1dx89TMPUBtfRzFGcec8RAZP0SE/tQ+4M/8jJQSxtqXHFAu/JyGr/sk
WVAa1d/e4kVptO/h62arvbkrF572TvG0Q1Gl7s7EJCLX/uJzHtCAlZ3PeDQMiQsQ
QzcAEArHhKBPoV4j2eb+FfISFiKUbA4dNBFfW9NEf+2j1QENBl6MqX1lIP3vzUqI
IbdJpXwMZjNhEuycPneVZQNprrRhLO70L2q3DpzbhWNgyP1HQtt9EGS1MWyPT0GQ
NJ1KY0ycFWJZGtksY5zSj/lXvytAr2iEWVasOXTN9zMtV316ms+Lj+n7eKUdBKny
IApFgaONnf8Fh3C64vQQNIzNxFHnNyRqqWlxTJ0CcnrOlPXSKEnr8AfkAjzq+m3J
hLFcw3k8HdbpreE1yB4Hh/p68TwgpNcpTWNDglhanrm1s9pFlJvlP4zGnBlj6/Wk
dI64HuLsvzWgerG72hglfBhz3zcE4qkZMNBplrWURSvSRoIBtFb5JEzqTeib5ZEa
4cHPRWMmBzLOPV+gAjjTkEjXS9xiOdTxM/lOK/Hk7r4viyi7/i4v+pbopOMpe+QU
RYKbhL9uOfJzeDnckXtYhBltF64ibMqBZ9+2ccaZ+SaiCp7BlOYELmK79DAv4luG
+paWvsndbUvIBQLjM9jMrRnKwb132Gp+BVjZnWv1wO22ipJYh5KAcMSk3ItEQYjK
cbuP3fpvEE1/EOT51nGRxqZC9kKwMdi+ZG26WdOK58Ky1cfqPqV9A8HjvDGIsyB7
aljRoT4g6v/8HS8Qiv3B/WWkIYPdpTydZlr2RBRrJSicWFobuh2EZbQVGyuXtKnc
sg3Ji9w0OjUJXfyc4bh6y9OJ21C3lTcMkNdqPitNmR5QyDOZi2vueg6eFhqRqPjk
KpcuUAjkiMiCpib++EA68hjlqDp2tCHFIE2OFChc3SSc4XyFHlhmRwT4mfGu9q5i
D/1B/bB/WzFvqu22xhFW+qp85T/r+IIPAT5em9rOg2vA4nPmB7LnHn8tW3Epb/Kb
X86HeC91Qje6mWfkxkjI9PFqP4s0Tz4WcdiZIsNyySj/ot1YsQYPt1BAixV3WaXC
KjLTrhQ1AZZWParLNLmrpoUOAUQSwR21/10Y8U8lzOMlR5zo3MVOuiZME6QAl9Uv
b4V6Mq/+M5C15ewJZirvPgix90DNRzphvMMn6zPhT8XJ5P3L+ofab8FxKAYkD9Bn
ZJFHYl1ihGVI39E1R0+rVM81NZJEwCu3YMbHNubDQvAc0ggsPcfQKRkL+NhxS9rc
KqJGKMRfvwR3sK4Tc96qiOjEMF7vJrolHO2xj4MDuroXKXdcLZ2lZOuoAGKUpG/1
TIe0adPz1rPpvGtBCY+7NDT/593VtKJUQziPxwDuURAbd1OvZ85anF3d9BCOPF9J
FkQ5uOa2FIUM1p+fO9sWglGjM4EgW1i0VKWkM1jpbvXW8WYLNUPLkWZ1xXM+uGHJ
xTEqvd04rL5EH2naeArxidXPbmxIgNpqm/fsSYmLXPiU+nnZBl64g3GLPV7UYS89
6U7Xu+qhceJaC1Hmz02XX5UOvB5Dr2EuANlFX//pIw+T3H5WdCLjHJUzPhlqEMVY
idDaKXMsb84VzHJ7rZumDzkFLZt8LMM9CS9gNjbVSfJvKrB+y735Bodl2CadsquJ
5vodEwnCdusCttuY5YU2tuckCbKkXVLghTFc3gGqvhNDMbRsJ7yDrXE4kIfdRDdy
PPDfKOONcK9eDEliWVKf0/6ZKRwG3tkEWKGfNF7hE6mR2MDsGZzm6nqtNLC5GAZI
ZR+7gszd+3mzpAWKS3vsesoDp18c+OXdaLaWiue/4DGaL+i1nRIXlAkIvAF0mBhL
bjtkURQEg8hnAU4GgGr6TrVlzRj2ii1U9vHB19OOGufD3KzOhuLZptpijWip0B0s
B72YJLOOW/g9F6Yj8pJaIPGBTQnsvQrkJkk2DU4mHg/UOfKtQeFfcaOAqtC6h7yt
TdbKmRYq7Hkw+JDd1uvl7/xONVE+ga8TCajkzYfVzgceRpdWO1fOjC9jKFYV8Vkk
0FwCWChbjegufJoSAg0juzL60IA9P4EXVxOsA7ZMAozY0eiBEv+OZr/UDVSJEFro
ekR1MXP0cLvo5Mrd33yULX1EmGpoTa7njsE4iNLJXOmZhevopRyCWqKGmdoO9l7z
tWMJw2vWaCHYdCJPUSkmXgIyjeHgtBESxUiP8xGzhptsABSe7flZjZ4VuBfmRzMo
tvOZkHchof5r5QiJaYXYsKDpdVcj9gLLfcePgKz/Yd7yzgNyIRbfSWb3m/JLA1Qr
lKe6gDrbxSACu84NkBjFlzraiPjSNJoDVQbjW1ADJZgq9lF5ArooLwVnUS5I9fey
4uLRGKM7j4gftimqFPLfOZdEgimY2bS9ivjWBIyFKFEBiMw8D/8T1UXxU0cQCLdV
ZyouOom0wB3dW++4JBYY8Y2BjY1uu4TW0zBBXB+7JlhNsgzegSKg0YnceKomLi//
OOp/dAWp/F/vw+x0godScmKpBy4H86LCVn55tl/Z86s=
`protect end_protected