`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
ddtXksX2+yylW5zu6QL2Lhnb2d1sD00763mmSITNX595NcHTEkwn0zB1Dry37fOW
FufOhVzEJp80NC5qZ/+F0Vk7Ik02dIR0elf3clrjeJRK85K4e3Hoo4xn7YbFUIms
l/8VZSb14+JVGURjfswrIyCUotIzlzVYZ6gzoZwDXIi5gQIBf/gI+KxNXPaKV+PQ
Ufys/12rjO6aI/pPlqSm0hCvftmBcnezN2hk1UeXgOIuKZnogjOsf0iJVX2aOOWE
6pD/psybjbnsNB6kH5uFTA5frkzIzkzl5d9+YDm9OyC+k84E83I/7/j+rk4L2dah
QJOvksSIzN867/4Qt8qYTQ==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="MvBXkzurAa5VTw+1JJ70nePUfoQXBvZOku/SMmg4TwQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
oRtzZL4VJ4iwysPsC8SXYCzXS8Fw2gtZTOskLcDV+1B9Nzn1zTyNtlo6lNICRmmK
ZRVu2BmCc2G+fmzynYlNTnSa7C0Cuel6FYpxCBlOuk3OF2tzAmLAuDyOH3Z1Yjzk
a0aHuoCdIRKv7BrZCdALt03JeUmXKPdOmIlkVGFl8yw=
`protect rights_digest_method = "sha256"
`protect end_toolblock="Jn9CQpRhJt4rnzZPRk+dOpzAubz7omckX1MrFd4p81o="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 4400 )
`protect data_block
gD6l00tciPUa6pDNTk/+t0OO0nC/UTtBwLB41d4inuAUA3i/ALrNyoJVcBnAmEQW
ptbcNp5fxEUJjnOxnedyZEuEBxWRieZFQnkRdF269oNhD6j6njB5TMCIBTGRoOu0
cYX0FG5A5/rgTiv6/NEJOwOBGovPclbe994zCJVxVKT1zFWJkppcEK8kFaUyDvWN
vH71Lpw29mZZfk13t/pgM7GbfYCfZtQYRwbGxvsl8Nb6iN9k14NBuAVLwkUS8xVV
O7cKjHnbyYmsUDika8iDl7/qrWAPcY9fB5xKsmf0SiE6Ai0FznOXfGd5zRYaJu0R
aw08Uw3CWsbRdFM9DPr9lYZImSiDB9DtxvfykBoaLvx+gSZnPDAhXzZZO8mVmOBy
CN6jmbfCXKtTfomu1rywonKA2K2G0RUZxNQZx6JDBLei9S4C9tnyKH7VEqLWxP8A
MlOSBqq4B9cEkzHBQFfWXDw257TbpPFJ/GR0qjs62dxjhjeWYDun3w/IbuCgRG5/
uR0YeFb87TAqdL3eV+mLOsGbW/Q+n8qDC88t1MZdbXRaqUWPUNwIzOCJPzXlL3ty
dChCo5z1qe1NMPDtNJnB7y1VeNBCYmJYP8BPhTfcr+GkkXfwiqhny99Qx/CoaEzl
Q9ht7z2lsW4Ms7hnV90gHJisBBXUugpkcFE+lQU8P41GL9ZTaWmWvPEAMlAiJ1Y2
nYWisKz4Z1iMQGViNk/3jDLdXdPsgmPdAmIE5er7b1ehs94o0OXuF0CipAmmozNU
OM4HwkXMYQ/ngGEs6YGV+jZ11kU9JxwDoEumrWiGiGYUauY/3zT0Ass0nmhHZAD7
qrTDWz41x/ICgCR5r44oWxdquFxllAgzoV+y7ewmSQ9Yk378Z1agqKnvcX56NaP+
XKZywEaz2BoHfKRjSS5OpXVrmwNHDb0/iM7bM3yLpOTFs90ftI41WSJCdCT0nxS9
yXx20K9RE+/FF925hFmGwlZSPXobFT9vpI1fQjrTL+qiVO0NEJ51eV77zFJls5nA
h/ZbeubwcZSsoi2nOwkoMdmmMH005MhCw5c/gfmdjHP2GI3W/c8c5+Av2PZP6Pf2
n2l4c5PfuRSTfPy+T+BZ4SGdDd1AwjoB8S+1+9rZqdT5/xdznbElLVgIZFn5OVKm
U+qk5wzRhkLfzqmORRDhEglVLoBCHKZm7d3B0zL+NtDG+24vcDoYUKzbsxxQcn0n
wmhf11+bkVzNrBslvyG3lUyah+k/PJV1W9Lb6CnJSTzJx8cR87ObHsUH2rVPgIuK
SleLC+qdlb8s6eISZuYtn0iHjOuc3PC5Il/gMimgS4r98JrKDSsf0X7mCY+uOzGZ
DwErRaidT9qXoiEbv/YaBT+Viebgy1TGDnDOGaFuljcsliSg4Jhzl517fDbYALq5
I9FKDlNfSAo5Nm+iK08TyWIHKgoe4lOI6yTK9OMjb1Lv/QwtooafPzBpC726Ahx4
eyoknfOM9JH6V8GUtOdCe/R/EIgCaw9jwVZg1ncGGlgZAuyRNpZby4IBjkF394J6
jsA/bJ7TNllnFPZNhJ5dtlFtilBxn+ESfCZDoMAshNEbzy3TtwIYjrfFzPKHLuAt
q04OdbEycxeXLPMgm4QtcVmaP618IxlQLZACF1xJ9wyL4HqhqlsbmYmwq8nz47Xh
UAbkdBgQZ3svVccwCfm71amVTncIbarF1TSmFl9A3uVYOmI+23nq6FPY8v3Q1av8
N6gYJ+xKsgmS8w16yES5kExMXrjOJvgsXU4/vhYoHpKDFigtweU9nz1hTuO182RN
Cf/XSOkXDTiF6/ezxB32NDK60UwCWLISNk9jFtveVFsPNuTxsn9+GO68v0eefPEH
8zfppS4QI0gnE1RBss/Zj2UUDmiMb52V47IhjKLVhFmclG+aZVpuodz33dtUowy9
vE4b/OQm/1fkOrn7oU2olKXnvxKKlY8kBiMzE0Nz79JvbSFrMdkbVYLSwZ9o2brp
pK1cINaQ3XVb+KPQeT2qFCNYQXc+k+rpTgHRZI+Yos2xmS409my199QdfSbK4BHR
RNSiY+i5Or4zoiKZNcYURIMqstP42p7BAQYzzhuqKbgn1WAicIToYtEBX7Ed/63k
j1d8jfv4pAA66HlTv/oMUeh04IfkFzQZA0ZXm4+xY+PAJmYHOP/HJjqN8AlNoJJn
5TWVntgaqGVdFHNO7MH4UnMitja4yAQaGtlFVsho0WhRunGnowyqdAG2KN5vVQ41
kdOM5DP28EvuMYj8Vm6RhIsXJaiwP4jKSKotuG2HBjwtwxTSCBwWTCB16lWgepa+
8tjZ72k7WLPXOJVs3neoX4h6gr+tL46mCwEYZDIEx5NfytuZJ1F6g41HBuGIaxz0
USPUioWEAwTE/E0NufZ26AEIEV/HcKjcBIhNdcySs534kUzi26vM6qr4Ah9mgs/L
G/5MB6CwX408aecX8pmNVS4t5VBdgPGwkGJNvre0qCgFtrD0iLbJ54YIJAX/rMUw
83cXghoSSyjDWBBOB5tY/RKvtku+0PP1Z0Cn0EQNjriQ6uEIuNSNwTkGR84azTun
KUxmGJIVnnPbf57VJboB+ekfdH1rU3gmffhH4l8zPeScf/yQxPoMXH4BO2+RP+6k
idX9BGrzeQVjoTn1bAKjAZfBnUqWn6+F1rAa5u/gl4D3Cs1//vb3RS7IcZi8hn/Q
2djAv7LnAnUgaD4LkDxIScvq+L2zTNUU2krpqPjSnX3XbMpzPLXg6NDBrSXB9V3f
kS04TmHLg7Kxnzr7aGwqjhYrQS+5Og7Gs16xnMRFc8DSEpl+vJt0jzLg7QEizMpm
e7yYOOikuiZ7KrCQMqzjR5qaXpF/rZUQX9I6mEH3uT/oSQe/h8vUn30o3xRTyhFq
X2TtIVghUp3fmDQnrwkVn3fnU+msueBW/62C1NQzEjC5sSFXEqlKCcQAZEjaNjTT
gTntaFs+wHTg9iZCI+aUHtt9dO9wwHfo5enpMqclPSbOyMUGlYRUAEk+1TrV6AQi
bXN82hRohtZOVIwe9GTrPfHlZpid+9DrznMDn0+W1spbR94X8I+MkoEFElMHoGRk
pN6HKiRUGGP0D1Pi5L/xTqrxoYK7TH9xZkuAsJZbuXTTSfl5MSfYMF7z6HoMkRi2
o/umrIABln/cr78sebQdMro004Nw/9f24y8ExzWipctb5sUdQQowvbviifA+iz+r
e7wtSZGFwxGLLGDwhhbr4WvDJo+vlHeYtUI4VrTilAUwELE7htP6bcpyPrgM707+
FNAL+pEIhJ+negYTDhWhHIIAf6V2BIhfIK/vPlvtWgz+rQ+j06PKhs2H1u3YJh50
XglXOW/N7OjW8xOj2DQGdrh+acHVrn+L/9BFXX/IVRbMvpRL7WKHgOcYST9B7fM6
0+lUyakZnLu94zWky1jH3hWnFy1oxTv+0nH1zfx1KXsiHzmiDGQj+xK5ZjvOYlJP
MwqRJdgPlLBedqJwXk0NURzOBmkNXeMifnrEOv7AjAQZx+X9d17yTgndTqgssgZG
QNBwOjZrTgIZ2nbzpqkEIPa3iP9oNvg3NuVypmAsJW+4TybvijIUO9ZtppGkwRKj
pld3shTv6XeWFr+Qm22UADYT5H2BZfOlZvTsnganoWlGKnbRQboWJjYhz+EEsPzI
Nt8LEnDC3+H+YbHo4sSROa+7BeZ436ZEYq8gC/SKs4sV/sOhPAIvfRiLDij65ULb
kM1907XFGoOVAJirCz1oFGcXxt8H2pSX/NLyxDdEpLCHlcUPBeWzSDBxf1ctvCYu
ZSOb8SBwGToOGuTE+8cgmeewRNnk7QK/TsLEQpFknob0WhSxo2Y3RBIljlNOX8Jx
eles943168D3HziCpQ0khOxDuPKxiTO2gsN/DqxaluqmctHxN/o5wgtteLMYBbh9
Br17Jr8ZYThSIFTqPV1ce5k/4hwR6qwx/wFK14Amt/hPZSGHJF3mQZCi4+p2f2ne
X1wx3aDXPqJyMF9gbyFzRQMWNw7rrudQOjiP9OYKXwgobvgeD68FjdgZ8JqUnUnp
FwU+iqk+wBsJCKVN+JsE8MUf/vIw2I5ybsBVSLKFRXQ7O1oPN+G4UA+T2HOqs6WK
dz6SpPZOfy756wAfjlZpg948SUB9Rs7Xe9tZWNDzVtv8sWZdzrh32wbx69fNFoHb
LiSenG+SK5RE2/oozblieIRnmzqZdGQmsrAJE2Wchf3CPLrtSEaznbMKG9X18r6N
SewFIlE1HrPezmB3mq58vtY19XyqDw2H0Nw3Qjp4LGv/nQETvjlguqndecC4g/Ii
mhrd1jzLv/2EENYNnTbZCuyqG0AM3k/C7QuVKtJfvqMrmsK8Gb7+/CcUi64g8/bG
Ugx427kDzSd/u9uVTGd7steFXM6Bt/hJZDeHdnF2oQ67iU3Eq22AxXQJwi7SV9i+
ZR27rH4rPPGVBORtQCwXzg292KSIMM4v+nzEbFKdMDt2OqaqsGY4bLDzbETog5w2
Lkd7wHX2JX6LapRlekaIUYDz/P+8WKJDUPoKSA0jGGWkTbiLIxdtfTeCnLJhJFe4
WLr2/+CFgn7IIjRVQ2lBCw77i6ZCkEB5INeap4uU8i0I2zU7foa/04GaXAZxn8jk
nMFLEbWYW8EEg6RRWniNCWAaUu6jHTXhh124xhvA/OSQ5AroNwiqWipkG+IrDn/W
yLRqQFTLcS9Y86E79+6J7JdCaf4LxPJymnJ06mw202R2fkp81sTdT6iSZwuJOCwA
uCp+Un0AIdRw41OePnFeGaqrixDgTm38SuaGlP+I2JSLYh/L/vIGXul4e4CNmQb3
ZI8cXtd41q5hxtgdqo+j8wK1tUasYoceNx2QpiObbAtViZ6fTJk3tC5xlCJ+aWpi
a986Ouz7qXJGAZP0j55il37VWIPeZuhJw8un/ac98B7GvZZBAZ4ZYgR0QE25ZKUe
xywyq7enni4Ae/fklreRuQvXQK138HQTaYfUCY+EGargZltxUyBWFHGdOx2jtDf2
4Y5hMpoiaCJ7MagS+vUZztUS+L6C6Ia49WYyYLJTqEinVxFsh8xrfbzuk6ClIZEI
Ofp32yjZKF1gFEa6bpUAkTm9xee6rjdD0RkhPqP9Mbr5tnCnyKowaJSEkPYew2my
veu2T77dN+XNSh1USA+LGgTh9B+92MyjPm7rETrGtxY07uOkLmvVYRz8vSghWV49
L+qyIbc2yJgcCMAO1ESUCzHj4r0W8ZsczOFAylDAqYt/pSkWVHjmnRrV4JT+poJG
y2Z2n5CRZ3AnJbs1dBCpk6wkLHP0ZVCClkSdQm6juunYnP47Vm1MpWoVnh06rxfn
tRAwMiNbqvZd+7FupvqSULBg/y2n9NrNye4WCqywr9qv91wf55lp+ymRfoPsvS53
yqU4XQN99v8COEwWxg7BnN82Vbc2fgbKmEnvMHDKcQtt4IzAJRuWL5hPLTgitZCR
TpSheEtEPZGhKFjbrIRrMdgsZ2svVvyVoNxRd2f6CE/PolVvk59lpOW0OBtE8udm
rlNKE7lavG9PmzMLPsWlmdCmFMID/URyuuhs24bcFmTSNrMIBXKysFDFEOcHSrUT
CUh38cK2J4E/VuNF71q00OYrzweb6USya2dEHRCa0+HiTD/IbX/tEgC4TamNt7dI
jAsxfbjrfofu7BZ1GUQh9NbZhVUTF7CTcgZWcwBMSh6xlCiDZp5oKsJP/QyW2ns8
reAZ2jqy0Xs20YQAfr8f93gzj3gx7bc+QavUliC3CtQZt9Df9tpQRca9sa65p27z
GH6crLItSfFGRu2m6LOSLsneTOtCB+V1Aj+LrJc/GuPjp50J+Goh2aOZaz4zSFaA
d+KY/f6suxXLvtOaQkyyUqkC4f9j0n9AMNkQPGqiV6A=
`protect end_protected