`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
ddtXksX2+yylW5zu6QL2Lhnb2d1sD00763mmSITNX595NcHTEkwn0zB1Dry37fOW
FufOhVzEJp80NC5qZ/+F0Vk7Ik02dIR0elf3clrjeJRK85K4e3Hoo4xn7YbFUIms
l/8VZSb14+JVGURjfswrIyCUotIzlzVYZ6gzoZwDXIi5gQIBf/gI+KxNXPaKV+PQ
Ufys/12rjO6aI/pPlqSm0hCvftmBcnezN2hk1UeXgOIuKZnogjOsf0iJVX2aOOWE
6pD/psybjbnsNB6kH5uFTA5frkzIzkzl5d9+YDm9OyC+k84E83I/7/j+rk4L2dah
QJOvksSIzN867/4Qt8qYTQ==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="MvBXkzurAa5VTw+1JJ70nePUfoQXBvZOku/SMmg4TwQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
oRtzZL4VJ4iwysPsC8SXYCzXS8Fw2gtZTOskLcDV+1B9Nzn1zTyNtlo6lNICRmmK
ZRVu2BmCc2G+fmzynYlNTnSa7C0Cuel6FYpxCBlOuk3OF2tzAmLAuDyOH3Z1Yjzk
a0aHuoCdIRKv7BrZCdALt03JeUmXKPdOmIlkVGFl8yw=
`protect rights_digest_method = "sha256"
`protect end_toolblock="Jn9CQpRhJt4rnzZPRk+dOpzAubz7omckX1MrFd4p81o="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 10800 )
`protect data_block
gD6l00tciPUa6pDNTk/+t0OO0nC/UTtBwLB41d4inuAUA3i/ALrNyoJVcBnAmEQW
ptbcNp5fxEUJjnOxnedyZEuEBxWRieZFQnkRdF269oOGV8D+YZee4u2iFzlgs+vC
kjLsW6unhVIk8WRp+xgHZ1woL2SsOB8nEnoshjZepv42Gtwz4RLXFQ4xvT5xnr/q
OLopzW34SBfmXTXtIMJ1LEGFD8cQDFYKKSSHdg/K9uuKztIhE982lvkShNqvoh1i
+RdVQnrZoJMEk5aiRqrXfzDXhbxnlfhxDvH7vgBU368wWhEOSNzG4+fKXKoqYWKE
gb5saN9M4KBSKIOZMoLqZ+e6/zPdHZFCd0k9lPEP3J8if7xkL8r/pvUmNJLpCG0N
uNWHMoMFRhb3DmCrDK5cw3fv1OxB3cbqYWV+57aO6qwMuZjj5jy67asH2dDOk5B6
YxX91NE6R6Vc8IG0FoDZ8VdGeeQxoaN9YocBUSUwyBkmC0GTQIiX1/HgHlrLuT8U
aKQWInDVChU17L2bmvpTz3f5RpnPAcy+6JgoTShbDmLt5FugxEXYUNwVGPFPrtdB
TjQ2gmW8JpnJ4d18tVMUKvAyYqXCUQKyl6tnwvj/Y8zoPcKuabqclnlM4IE+xFEL
Y0SGNF++M1k49d9wbSOMOaWT68v/KuTjuVw6q4X0EpGfD7D6zmY+Gs4RIhOmG9Dr
PfKZfldyiqYN+VjDxZceojqpyfnvN7B3jz2+Wl717foWtQEBp3SWsphOu0yss4K5
GrFjwel3nQITz5jW02kLrgldGi6ZsxZBbmTLB8UfopNKg59uTJlhZin3HMYhmtp6
r4YJ/HpJK1LDXQcihH/qPIO93MyLTn4yBMkQjMhvjraxyAahobedexvOekuHdk78
/zsLKYKOKG0usKA+HjRNzIz+bAhMk6GWBN+keMl4uEOUyqkfr8S1PA8MIvNE7BKR
24frp8D/xYaZ4nN4X7TCak1qrv5Ilu8HQIIsFDO3ErWV8Xwg8V7OpDChpJmhcvAI
MsYytieTypQOtzSh06fTkWZi93IDACAqqz837MVkCO4Z3CwHcTGJmJNlO+NXfMt7
fIRAxFll4wRUV9ICFaOTg2pdl/OA6RmJhQ+cqT24Zwhy9kRU6XNVv/VEG6MXpyaJ
H4YkWQBGDDSJqX682nBfqZpwWo3Hu2FweCl8YXWpjW6yUzzf4RuHtv9CDltrptrr
c6vbMI/4O1aZGwqGiAG0glGwh0XTNK2FO25HYlWH7kOdNHAmkClzircgOGP7jif4
DwX2mDz22UeyktgdPm8NL1xHuZxuRvg/7xtZopeiYTmeLgxbrLI5XS+quPDgdvL2
D9uMCXiXpvQ5p6C3cZf3pumFf21IWtBQtBsy6z4YkBwbM1DB0EmY6YFv7saZR9At
OfsjyWU9Gp45uWzxJCoVXAt9cCcRiBZkvkPdrv1kxsLe3/Up3xbH86zwg34tyjYQ
P9muQ4b9jpcD3Xh38WctE3p9b7b3DxMlOws0wmhvmu75eF1QEpv8QDyYitQA4VLy
fwqzJJje5ZRS70bsgqyXKvvLfvALY21p+cuf0uV+GRo+z6wQWH7PErwUZ6/4l1pf
ZOi2ut9l1vXs7TXaZZL+KMTWFMf58a5Z+h6ZwH62FBHB4IDKio8HF8GX8HQjYOiQ
sqtcKluBDcwWG6Hk9eF25GgwJhhtlAQxjlYxe3SD4xLH7uoJV9BYWoMBHQwYf3uN
DS/u8eEuOetNxUf9m4rcqWmXGbCwdlPo3d1V973zePruJ0XU0Kj+ae2rDAES6eUf
GDNjjPe/IuzxbYqFCYpTjJ112cVadEb4QAg4I4GZ5HPws5SE2P+24QUS67/cgCgi
BZjcEDIzxBa+9E/eRcg+KnO9I5f39rFuGksoHvXSTiP0XaNGRwVDPeGQSiT/QDDM
ZA7ZNC6tSkn2m+ieOhcU0vlo3StnI/Qhx7TAv1bqa1kB3ifKNfXFh5AuSkCgPpl6
6SlkP5k2tIWWcCqBKFtNEVTJlHaBbbY86K+LwS/Yy3sPc1VnDYTSOXRFCQ5Lb9Sn
N/awa/1axO9YkrF43jWU0ZpshgFLOJltATEcGI3TujT4B0il2JX12duBpeBvxWp3
jOnPbgYejehtda2tDQJ6afrWeL6AMR/E/NcZWApBJC/9qChmHgftNZO8GobjAFEU
zIkQyJoK6Czc8x0Wrz35PWJDlEDyDXCt9vp2asOPy/CK0ogdl4JT6VjNqjnkyYEa
7kTHq+hWlRS0g8qibcpDPxdCWUvhwXfDtkK62nb8PzWJ4t+IPVtau2m4SmzdjYeM
A/G799Jtwcn3jRHRGpBNBCSmI+sV+Wlc0zy/XHyoHB/O1S5hqtLAhV38DjdWGGXQ
E7G/RWxZWelFAfdq7m71Vi8WNbN6kVKke4BSaqg0AWdmO8j8OW0qNS/d5iOIzWDm
3rq18wSOxEHSuYCY/UOyAjhl2f0bNcAoJFetW9CgSFoHIYhBbmhyD8JGbpiMPCDE
8JJNi1E7ZKXwTBNZpOhV5i+1Mj9jQ/CPW1PnlkEASTelP8R/prFZkzltp+D1PLXP
QAM7+8wimAFt+Y91bbN/Qi9byMuitQAqC0SNTzOKl3bDFq1Wm71Zcuz+RXr3iAno
IIivxsJeiAl/TBMAB48w8vNDL7WKIniRQ6xUPxoUjWrNl6JDMMIOLpRGW7x1aI+h
zPm6WT54OlevccTWf+SSD8lVwXIAKXB97OeyA9jwhYOyHFDqRY/dN6MW2WP8Ve7m
3+ife/Srt+2wrCYQSgk7evhWEk01Y5tf/JPGmGy+AnLjshlxhzeHRIiSwZOWMmVr
Uwjai9tR/73Sq4wxuAHzxMN+G9yCxpQf8L9oMHdE8g4eUeraaLmZCJV7uHS3N5iC
JlUnVMQT6mON3PXSL4pjYs4GOrRE5Mtez4gKe8byeqG4PJP8hvs4w9PPoQRB8MIr
TBO9CKrH3lLY/vCW35pwtY1GwiGIkOe6uIXppulIpLSDCUCNpKWhexz13RH6jx+s
pDXLKKSVPCnvzXBvrSoL6MZQ9/OqsbMUMQzW3ZHUktBF7W5wjvDTA/cy9OyiN2ps
0Zucl91MSeRn/I+6RdWllQySIOXKNhoorKzo+u4z3SkW8hhvejbdmdXD6yPwKiUB
SP24EwnyomLWJLi1NfGPZVXNIV+rrufskAnxLQTw65Z+g3nHwapnaolVB6vxX+7Q
bepiM8YsJDh7+No/Zi7Cf4lxw8vyI2XMhHW7fuh52LifOMhguxjHOLMqyP84WDIA
DZYh4rnhhmgmr/7k9Q/R6doAuHva3J9yOwq1R+0oPf6PHxAW8AGVOIbm8ukIf6Ea
zhFLJy9GCpR2uHhP7NrRPbqL+HunUnsGJrCufjqkg6ZFB9tkyMabIxURZanMhYdM
S2xxpAPk2wOiWhPhV93yHKkCfyWc8bKBmSKMCjC/KEjZylQiZk76MhL/yDgzZCAp
nhQYUCNL8n1JH+wqyesiKViISP72DJUQeJTGFRaTUUABq+eIJUPvxT3aCkRD+6Aq
TW/rhH3LOuIi2OHDf/rN9433+9dIMny46j/Y5AD66MW30Mo8Tx3zu0vZtoBV6vWM
WIP4J4GxXxvGNTGbiMdOys0NGUJlXknpgMmjFY1OS45sR5sNIiLLVXfOG0Fvpizo
9nW5+ouAF4Lcb8KPBuap/U04BijLBYdnCuLo876WW6/Ud/NrP7lDaQZdBZ2GFwqB
XnLAbESCQ/22ti9OthGSVXU2Amkaaox71Tn+TRcRjZUeVhefp+9F5tcZeDXN4GNa
TGVNwXv7Iq8clh5Cz9I6YBQUyjj7VgFMBGZRe+Tq9mgmmkMOdc7Y0xQAcs8sdS8a
AW7lo6MaW22wDjDD4ZJ/jhJvGIIT2yshfqnopmeRQDIYRFPvC49xNRQJFbdacaXV
G/NNwSWpnmSDGvuuuXwBklpL1RTgbTcddyKRc+P/kuiJE68EEW7RnKH3/QV7RhLh
+OL5NcUpt/J4XIL/dO5M19GA2ffhjBpOTaHlCUke/LGSJp4S0fT7EGVnIjXQZsfN
WO0xd1/NSvk5shuyO3Bs+dhfOWZduOKuL4IU2q1+Law1t2vlKi2ncx15EH7Ii9Jj
LdaBjuxDDPd7o63MeIYTdroj72CGIezuMvATnaQkkkv6yBRBgjVRY+lR8lWyi1HK
fqDrHyYb+Ssw+AoavvkExm/5lP1RSfGFm4/iwUtDYQqvq3G7BaX0dmEVtcwgumKq
Qqi3bEzHcVsu64XQI2ihZ0iYYF24UkR8q8XtSiqzIi4wKEsuudUkf6VJ/hi9oKPs
8mOJZTNAbQVVyQbVzPEVRiLXce6/Gn0lhOIaocWP9Zava9F/rsjS+1m3DB+aaCSH
7/tFpwufbU2+gRMs4fd1DRWsB3FNxIJyw5pn8BHjIa8PLbTBVWbEZBheDKt/jEOW
TBC4ZDkfZiIYtcXh3oGi4MqEWyoh0O3yO9q+EXmrC1fmOyAFaOf5KsiC3OeQii0S
7q3RSc1mOljNUdyV9xnSF30jnzc7UfJMg3ywjYZAZkjtkYdMj6OkJvy3MvjKynDB
aUa/ECyiWenesB70r+pN/POt1vpGQgC4cJ3CA07/QeYTPImDSGb4qk56A4GogxbT
o5LRuYBASiCdTOkz9yrfiUAGyoKqWnBmS+qaQqJyRqqrQlhaVLZ355L3usQz3EAA
van+1pmsXZIiRVj838mQpKzRxVoNp86nC+U3CiM1l+MlPRVN7o+gpMpes0x7HhKy
4iAqtGgb5G4xS/taFL7fo0Yp8Wj9HsEKuZ9xh7EGZMl9YSbmGphwIBZweH6YYdmw
TsYB+f/8DQ532NN1gg5AfweVRGo0KKs72nF3ne+mGvpSiUDMGjHz4kPsV4s2eFI3
Vwua6rBUiWuPLWa0MOPM4JhcjKGRnB8A/a0bvr5QT1sEJMUNN6CMeNhgTwhz2fCF
GR3uzxMpCJRa5NGlib9HRrePqZdKt4wxBuj+ep/pROGkWmi7Q2wIjAJJKMbdclio
Dli/ULNH3Ab4br4vw2MEJ3ZvL8p5ETACM2APZmAQImrmKVBgk0jPrlspxVFg0hLI
IohliLAA+qY4zAhtlRuruUeIiInMuvHJfRG8kEtRHEGUMxv+tdqY3BVrExhcvu58
6w26F37Bjo2NecpqnzI+4KuVUiw3RGW1ZpsNGT6WHYQgZpC679rDUQY1oBKZDmqv
zgkMgIoylZQAZP5XgrK+nXGzndT2gOZXObrFgdtXWi3gweGHrH8tgRV83kU+5exq
flefAJzwoYlTDzU2Hu9QFQUv8TZcXLrlYBdjVtlk7iP8MuulnVgsl1+kAwrbnJLd
nji6YkiK68isecXX1QWBVTLpGJ8WJAbrsbcRxQleldBzy6Pr6+AFGn47cx2nxnvU
X7IfjtsBb2Jt577m1Z1cTWyp61/Ly7+1naPp8hOZ3u3AqkpZ9AKNFRwdkXJBnKBh
9TSl42wkSt5YzTQRCRaHZ82gKEnn1O6bWlWmmRodpz4hAuX5MFAQGk4wTaWvTbk8
xSXZTYgm0F8kmiM65wa4Dx0LJFPXxdWnCAgKXPX4Vk0IuWvOxhBdzTzcb8vQ0hQJ
AyVt5pgg4M7DlcWpYV45+P0uL+KqCqUKUdFmx6UVWhVRujc5hPpvdkECXdHpkkeo
rRRECWEAPg4VC1KYwSzyhzeek0aEh3Wen5uyb4nVmt6EOMkq3CJcFGv3T/Kc4Lu4
Jo8wX8RCgcHQCfI8xshxvlBAv3p181Xs5UE5JRApPRJnin6v7oTFgnDC4suum3Qz
CTaKJEKLKgpY8EVwN5KcvzlCsTsdkatUuo1QFO2248ca++1v/2/7xCEntTHumTSD
ee4Tbfx7CVwH1kHNlEc+FK2HeOAuwJoxKrTa4UsTDuno4eTsidw2CgPmnhGVIgHb
QKjp9sH51/yHv1h3aEF+bUgNOYH+L8hJtESiAo166xViuQQg+rwNDiB7lWYZWMrf
LuGNK2CQ6oASiTkmQalxCmJDZhmRhNe0aYKLYXBLm3gHh04oQBsmg1fEA4H5EOZZ
5g2vsmu+g+UlbQMgf+saCvzOYvmz8QjhJTe4BclCi4Lz5eL+BHmH997ImiI9KHDf
zgVQxGdIUJsMaVbCPyqI+nyF5UBqEPL3AyMto7zFZQqfLd8HcjnvwHJGNOVjbIvt
ZG//T1JMZ6ZQ0Q40CS/fDJ5A4a4YK3+OGPllW4eTlcFH+C+azENe6jh/w2drdbB5
NxGwAv/bXcVCV57MO3U6xWA4ye++BCIXrdBhmeilcLEgkrHnIbuWI65yYtaaf0uz
Bk+1RdiHgN1M3GYebpF36UOibnWVr1buRYtr+kZDG90//9AXJIIgzzLKgN7ijXgV
gyknmjfO9vVHnY9gJ3YhY+9Z/JPUK6A5BYmdlqs1FJ6ubEW7us6wArC7/N/4HKoW
UPA3ammkjPVdb05zsffyVj9ziWZihP+UmgcrrqDeSnz0oeLpyNI1/2HCywjVQR25
nkdutTBMuPsuI9EVuBFZXxhVgd86Wr36mMsiUDDsj35s2BXgv2uagM2kqFGakSxA
4/j1MOWjDA6FK5E+895uI/0u46b3SeSEyVz1zL55jeDMR5JhoDO9QLhcWZ9jDUXv
okfISgMFK4BLiLZjp3bOKbrCS84ds6/dZqpo984+dP0vSgT2uetq9Oa4Qo+hFvan
ZFg0BsOtJ6uISx4jen4LCgIKcaBpDbpX39htPQc93Jg7gAdxEUG/BnWi53BpvTzg
TSSUJ2zUneqrP2eWdyvaD9u8TM2CUuMNK8+N9Je+ckd/76FnTTUzMLB/3dzpUMaL
wFU7fRIVqHW2Qjqh0rCuofcXY9miL6herNq7JK3KXnJVZLR3mMkWwpifRtlMGdfB
OB0WA8vjrVnFR9mTumbx4Djn5fq2K0sp5BlDZfVtkDYqhSBe+4zyWlh/GDqBlUQR
NlZ4LeRf7KEroLB6eKWd+Pu/gPzCaBy+iGoojQh8de5CE/nRdoZPaYA1eLKE9pKC
vH+RVcPJ/Eu0JxGZxm7Sbw6Y6oGD3Y6OFBxvvDfrDEaf/0YWHTogwOUS4SEXdVpB
Od0pT+TgMvnRyFgS85tFCcsy/8Wk5mGvH5flQfrgDC8ms3jbFznKrMM6Mo82VrDG
VHyObn3WywYKhPxoc5deDQbNFcliSYO+RJD303IG0lmojm08aGfVkv1Hk1GjwSBG
+0AFk8A1CLdoPoR+PYbnff+/BZB+gkeHbAj0j9thiiiH0Jft+YUb+cHxKJjCng2q
3xOnaDQbDganN00IHeV/5wJo8bG7cl/4wRGiC9PbGRvbmuAAbjFYWo7dcPh5ojaG
BtbI4DqsyIvSc8ZlRxmSmR4LXAxvqyGDeBWLWLpvIJc/mlh5iZGB6fgz1JFnymLd
pZhPoo1VmP08BYYaxkJ7fC9NPXik4Rc/FEjbPMA3suKeBqQy3K5IULLXZ1CDUMtO
GYW16IJOR/3kQRoWfkPtwUYnjo8YkWyucRGT2YYuU9xTLbjUBRsHOYr8Ik2e8Enu
70SGYx1YOlDbyBtMOuQ+num5ADN6ZVOcinQk04xdTx1op0plaTDG4NbffguHp5so
/sMZseT6IB2PTAGqSep101eJtAILzybWxIZBAu59ZZsF5GrOX1kZmiNfydG3EfxH
XS6sTdHNQiD1WzKzfKbgpFa3Tx+JEwY/jMRQJycBdui2lsOcixRLbPfLIqspmo6a
HSP+0jZJLpRX5+8kT560lBfreu7CXpL7kO6enkgXKqo+yOJ4iW9yCeiRMHvdjHT4
UK8fzCmBFBI2W9F7E1Q0GSux8z+mDuBleS1dju9vG5OXefbRw48NTuoH1GwL4I6g
w9At0PRn3H3AwbUdUuc3LmNyy4VRIuOGffFfFjiOFGRD6pkSGBEcPHe6oIw3sqOt
aRZV5VwmcR4T3fXCLSPNndX+D2j5RuEM/zSlimtDZmfNXukBr6uMzB2+sa75biT4
OjYsV0eyhHtMcYM73xBf+Oud7grF4GMJPMQhNgFuNnSj5CNoQ6Zx7qqqEKmN0rvf
DdDAmhnlkR/+eyrTed26Gr1knKaifDZrMj4khngU15n0V+z5V2mW5jhfMLXkRLOC
fob92ZQetYemy7SvHMD/WhbxzEdkm6QSerWporiodFxh45YXL81TTPcDv0NMtCRy
NdXkPDPFQwGMdu/rjUrBlLyCOTPOfresMZRyb1b10ZyytW3C3lewzOQICx9HdpH7
SxOXkTAIeOL9Kt+g+a3Vum/4hp/5/rGrPkOQljIec5lLgYCkTYxlaagDeQlSnNfp
drEAV4D9AL39F4o/HIlskgOzGVguV/vnMkjD2p5Nd6luBco/i7VI4c/og3DNzN9u
aS7OiRdVWX+2NHArMOP8a80J44USU5/kMgbMj5ydeXHG+aF0UO8RMIbkFTfe38O8
4A2YHCerO09SjIr4ZSgDJpOTfvuKhyh99zDiZhZZbW9baGz7ogZTDZqGIitLBxAY
VkVY9D1j+4FCzXDvwjHVjrejiuGynKV9B0Ybfx/dn3RSWsEPuR7osisgMfdgCdqx
4+ab9sowo6CMMpSc84YS900B/w/VsOpCSe4OxJJzhUuxXw7vCm1xo4joeWXAGcLP
WKMtar99J3FiC1kri0NhwPHL+rymFuHCWR2P/6pOeLhwHiI5bYGxA5QP83BWaALo
OBuBzxBD0debCGiW2Q192G5/nbp+iw0slriNlJ0x4M9qdhlOzk5cG/Byx0U5RKhu
2SY9eb/K4LWpf3KCGX9E9Ul18VyNX7V/aeG3mAjf37PgRT9j9Ko5bvikQYslF/Zx
wzRb6qyHD90bVk2LpzfLLYBE1GeLWVLszetiD5weX3EE98QT+uEXcNNZZWtpRKpf
IoctownSpsPXdQKZA+Kbw8/lvMrjIA1t3A7YmdmsojLKaKXkHFapm1x0zABnI54u
DN/2v0RiABuuMqfTPHRIDdRQadycEbApkii6kL8FI1Px+b8sPw93ocxuZOVYvWew
f+kyBTGbBGflALA4qtanarPaljhUptIeKntB1CSSPVA8expwB81ajDXqND3yyOP4
b5sOqiMLdsWCs0d7dOzUOBMJM0xKP0JyTQmlLMEvVSocXwcTGfzherScwzaOZagr
WGkJK6FI3Ac6wEjI7GVokXl6F/J25kyPovg2IIQWAgHVZrqvrO8DwctZz4+wHNh+
B1Ld8SN8Loq7yGjTcscNf5PqeKmicpfzkVZo/XJ8+TGKqUvuKqVq44kxFU6mBkSY
32zMmyAni3+A0E4xI1Yg74GjU0b+Yu5I/XYv+PNPQH4wQsALvRAw5AFaFAjyB4Cs
AMFcZVw4tEOaWhsvTk2lM0DDzMbV/Bu7469pKFFL5aORW+IqaGymZ8Xr+i3Q0yvQ
VJX6fHSrf5UFd+UCeLM8/YdV6hE4yXA3xbJsmQiSaqwH+8ez/WaGx/yWKNVfpDKr
YTdKjDeB1jk8r1wbsEkfZjyPI+CXuJ56qfNoF0q62ECNzVy2wNb7Zx+RcKq7yJfI
cxZE8WgZ5L6lyq08vcBTaqRLyXC9WmStFf0fzslyyqLMjE7bPy5TJ/RmUAXjqW3n
DAPlOd8iGVHKyEWUcjqQ+0o/N/bRDxyRV7k9AGeEDW8hfC52Fpkbyv3vf2BB3J3r
Licn/I8WYqedXs/8RTmsGvN1LvYwopUiTf0GKMJVTcozL2s87tkAlSnpWCyuAJwu
HEaIXgvsLCy73KxHpSzGrcGqPuhAMV8W3m1oaswdpauQwgNlWBQcjbwGqBZ8dy27
GAfjCA6safb/gsDh23+yVc7YOix2sWMPDZ/DqolU3GNRNDjnazE3fsWDd866a+jC
Tnseny9OdavYK1Z43DsZwZAIGocea8QN9aKYnxtomS8+3viOol53qs9N4TwI8HPs
UANNEnmPrzsN6hXuo6nvO07Kggi9B5C/FkdkjZjs3mA4cr7rR5qu12bIZfQJUAH6
LneNXi4SgBsdZIpTXUCCSaYXjF2ARP0wWB9HL62oW9xnrT0ql2spOhncqlqUf21L
kUsvsVs2KG3B+sp6v1uMlbBJTcsVwIaXsBTxn3UmepIfhu/F6wrF5fOjMVyvFVis
Bav+7onifpOUuLQRNkTp2uC1di/qi/tmalz+Xo2j5h32kgUsXoL7R6/vcscRYvv4
W3SbOfYW2cbJ0S4CTNmWo0P3wSN2+Ag3nR6KCskQWFqrjLqqUvnFoaTci/1q0btr
EQ1BLhG1CHUWoVoZlK39MHbBYYY04HfppW7/GpJbcQaKaFYOBUmbBNSAP+0wy1kR
MBVhsWs/FrHrwcl30vil3yXu3mjBqqhLGEaxZENPLSZak7+AY3W1JiB48wij+gZf
kORZoSXIJhD6uiKDooSVHm20kr8A2oI93iGSIuoDWN1n3hy1foPLnHWEXyVWifft
1qqdI3jJc6/Wo9PZmiJFjMZ+va+9baFetd3DLtRvDb4obfXnF12vQr6tqsQD5Oga
slug4nf4NodyTZeoZsxGav2qZNpz3KvV7oK4kegDYWCWlp5jEDB8fJlykyuIVp6Y
9UneJgSMJbgQ6CmZS95qOn23BG+0cDMDgfHB7mEfMmDFBo6K0R78aoLH9jPnhlr3
5UHGI4DFn8o3yl4ZFU3HWBB0SgHjkFI7hIV7967NMzSHYuv1f11NJ1eEQRoS0EGV
r/NV6NrId5KDUm5XDGZ9VyRPar5uYNnnOC6yf3P7CGwzcPWTj6ndOCZd1imL7pTG
uh+Xpg8Dwjnd+wqphN+YZIUXF+WXK229ig3OvD3qiJusknokKF4PA6WCzs9molR9
bEpxTtZMxctlCMk4N4rFKwVpGil9e59dxAYNpqm8ZWxK9xdeFvhRXARKd8r25Ryd
GXGjRwxHdPJoNkOP3peXJs940BfsYyKKYmmO2eBkzaDUqtxoZz0ZjjLNfOc1whMs
ARoTjIImiGkPVwyhqoMPy84t6b3hxOuDrBYTW6JFwZ8xI3N5yvCJ766aTNHIbR9i
aiZoiZdy/EXWNGgdnfinVR3Cf15r+qh17Vghn5nWma2FjoNWdyDSybDS5Ap4CCSL
jUjAZqd+ZNkiVHLjyoxZKiV4ljCXtt/MfIKVeEFyQ0Bm1nyQddKe7yHPJ0YDRz6t
WmKPjrHJL3FQ7g4vLvFMKvAZJassDQAIVLOZBlybu/X8LiUKwPaw6uPW1gHW5jcs
zUAfhSpFhx+tzwg96je1la68bpHhoxXzinKUUGz/Zs+odAR0i4z4i8r/WcprPLOb
OcLg4h2n0fydR8ZHzhe1ZHI7yV6Q368U/XoB3uvM+mbCpReJxWz6bcrMvKP5B1Wz
CYVcqNUAtx9Byxn1QJCYWqevFXMgmzLyEbELOqHDpA3aho9tVCP2iK8rB7498LZ6
mvaGFPjrs7HpZ/K/sYXjSfZ2QZ6yjbfFWJO4UWqWQTTfWk1uIHtUtqQr581bE/W3
ZJIqAFF4cMkU3nwZ/sdP3gQanON/R+LHaGd25qLmuqpH/FcwcR1O0PSXk7MGfSfs
9VQtR3ITlVw6palYe+hTvQfhY+7ejzZ7XAO8+b6KAHaIKIynqTUV287DVwo12WVf
Pcoc3IIePiUUKHlrIVVVq1Q61sDbQvT0re4NYlj+KNzJ+NsDIffJRAJ87CFi4sYa
uIKtBEczx2zbc+Bvr9vqtZFfdess6SE1YyKUIOUqgMCc1mPo9yL4NVasJp7K55zs
6g2YKhHY0Dj763f4bgHr+ARQEAa4aB2NvT2KJ0PrnfsP3PIyuWMVJlWsasy8l7UZ
4QHC2QXbbTy48yil+r/HwWoov5/xGhfe1lWwAb9pa1JoBU+zzINunouUky8B8dy8
UHniBZod4XfUNZ2urCZ9IStNkTboTRjSy5iPPPXR8tq5g1M/kyU3N4lqcaPVrneh
uUTKdo7UR7Upr5vt5Lq+vfgI6XKfpDyH4dK9SlaSD6G2PtqKuRQcCOek04C1sSl3
3DuiS4Izf4njTVF4JuVuoOuHhO2t0PP/BYWvA/j3SxfxNfMlZM2af3aP7/gaPXao
CwFkCZp6+QCiYzpENRSSsXhR9q0RsMCu4XhBsveAWzdGcl2EGhpw8srTULfSlgAV
EeRoLFVpy+AhyCAL93YC3Ys4jtEPHap7HrMNqOIOnUoyeC5fy36jodqjnYakH48I
JbXnwjiGAhpTT+2xJl3QGh/28B4eXrDTltBv5I0LjfPNFSShfMW5rJB2nZCc3Ugg
SWKsg7WnmZvWdWbjdmIdCHyt/xwKhz6TAKxeIBnUp+mmR3ne4HQAEnKM3ZqY28h2
gcwnnXGeFMoXkWYbEMn/0I0DC2QyzoVWLfJOayJ9p5oWpTyc8f+O4uHurYFURRGl
pyFEB6/23lqJrc2EW6ir7oUj4kP9ubp8dcVcO2LbFD8osSySmZhjQuAKvcPYL9c5
tA4dB4g6ZjVUkYSV/2vqRNQ0YbUW1g+JhoJKyU+AiuV8H34/KlD53tsbotpnNeVm
enSCWeUlntFYfq39MoJpRt9JGXdweCUEFJxD6XdY/+pZhhrxHZAN61cjj5pmOAgg
wjtgjIbzVD1qVlPtgn8y41N1pxqLxdktihzGtuB+W950BnjxOnUoDjju5UWN9x9S
voOIIzUhfDPnHSRYslDodDiD2BZ99STl+kuFHUHUUNM2T9YD1nq3GRTJ5t5CAGzO
Hc63QYFDfb1oUF9haVdgrcj0kRtzbEk9jT2KG+6xGWspdPCzGvkMVpdcEVcahAyE
7OnKJGz/Z1ga+5MHcrnDqisHUxi/8wVeCrwy7saaK7on9iNHx4hozlRJJjbNd0xH
Yl65NplLVt2gNy4/Zp38dfqVonazOuLaZFAoiwbRmnzeinslhgFuqCxjMg3qzGJ1
LjUKFNg9g6jiykn7vhSC85ssW2kgh8FQPD9c86vj+5H+1Hh6XUHRXIuGhdQcEr5Z
5/lEa/zqVo5CBZN86tTGNpAYYxcZHLu0KdIUalKdaoFCCQVZDJUaKssOVhdEG2Yv
BsNuoz+2mnDabYEiyEktSSoPpegAiU/eAxx6wz5rWhpNKRLdqFot41/S+sPsKpOo
7DCmw4l9vSVbiMwhEwmgb6qnKTsAdsdduXOogA1BW1PzFYZ6CUSrSklfVlrDJkMN
edi2L4mViybPrCb/I839HzMtZMiMUwEieFW2VuLVlqRX/7gsCJlpvIAymDC0W8aY
6A3BJVX10m9Wc207yr+NBYoWRYxUSQGFvp9lAWrVARr44J8vGDqccOK/98E7r+BZ
c65BoUpBV1caiIQ0JPKnHrD2h2LgZ0u9/zzs+5si3a4JXsW7tCXgpy6TTgfbZkjC
9JMloEZFqWWyw9d7g3XtfLHwlNpoknHSpOLi7pZKmgdrhpEc8Z9CCD2KyHILazNI
KlS66bonI7LbZCGvG7enVIZKwdzFLLsLLA07eolMZS5S3PYSvs8W0CUNqsKDAMmk
AG7/Bqah15VUKL9rfBLpoR8aM/Rt2wZi2rUJ0BvBtwuxXAM3SiqCn61HRRiRmJtp
pUqj1foTz7LSJLXYsAJNoFpfhlEkX9iN3c+Z9x0PjSWcElRgHN7tcwJmk+LbCOc0
Q9H1rwZHpgu41Ohd6bQUfffSg7cp6BOfec1LtBM9azjnNGrRcXsIFMFzKjiQ7/RF
B+8lBT4oSTa8GGNqcaTRDRTFNr/Xf4xM/eA5PcLBtjW+wDl2RxwY2riVtbyReBaZ
bUIkfiYbZ59qA4LS5q38SfK0StZng0CykR1rHaOe1ipNoo73zHjRhe1cbEvEs6YR
8rfgkOvwA6Xj0Bk8enDuPu2KJcb6ciNw/+zrfqyl4bhWFEAFs6l4jg5hzbERmLCv
GzJ+Y+fc2TkTAcsuNZ9zffO6xo0jF2WnJ72TIuRcYUVs66iIbbRk67ToJ9AGuftL
qip6Sj01awo3M1Fxdbt19nRKM1Z8Av9WYtXYdZ47PQrY4OvQyIvMgl7F00U7djdM
ma7VgedCTi+vafEeY8SMBh7H2SCqBz7PFwYqSvQs9muDbEJdFXnfwj2Ztxh5K54y
J4CTvG23lrWToVpNyJmTMB4YLPfM1jNMobF9dysIADkJt1RK/4oQsm2ZI6yABOst
aSD6YQNuCFakCkTHtuVZ9JvU3Mz77DaoQH1r/qB87JIlvxJ1fdLv/rTzmCW0LDQr
EgO77N/FBkovN862QDZY5J63DHhbIUOJVadUqOhr5NQiulUZIixXPP5+0SYpDc83
CTxcGTTvzJqrYjzkA9R0VKmOY0a7MJ3RvlsreccBq2VmPufaKc4rPKkVLMHlMtCg
fR7XibOtbGWK6+mlXWQ1+Zza6bYLeTclAs4uyw22cghe2Y8MQjTdwphhnHoZAkIN
rupKtV3iFduacJELRluf5PEooOQ1XdlfhtUFVtfGJJQOi1WXgi1Df6ELFP8kb1XF
6xGCxoY+g+DB4lxKJuRCNewFAG6GLd7+4lDVFQI1xQZCrGfWnzPn/8dkXnXGzKRS
`protect end_protected