`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
ddtXksX2+yylW5zu6QL2Lhnb2d1sD00763mmSITNX595NcHTEkwn0zB1Dry37fOW
FufOhVzEJp80NC5qZ/+F0Vk7Ik02dIR0elf3clrjeJRK85K4e3Hoo4xn7YbFUIms
l/8VZSb14+JVGURjfswrIyCUotIzlzVYZ6gzoZwDXIi5gQIBf/gI+KxNXPaKV+PQ
Ufys/12rjO6aI/pPlqSm0hCvftmBcnezN2hk1UeXgOIuKZnogjOsf0iJVX2aOOWE
6pD/psybjbnsNB6kH5uFTA5frkzIzkzl5d9+YDm9OyC+k84E83I/7/j+rk4L2dah
QJOvksSIzN867/4Qt8qYTQ==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="MvBXkzurAa5VTw+1JJ70nePUfoQXBvZOku/SMmg4TwQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
oRtzZL4VJ4iwysPsC8SXYCzXS8Fw2gtZTOskLcDV+1B9Nzn1zTyNtlo6lNICRmmK
ZRVu2BmCc2G+fmzynYlNTnSa7C0Cuel6FYpxCBlOuk3OF2tzAmLAuDyOH3Z1Yjzk
a0aHuoCdIRKv7BrZCdALt03JeUmXKPdOmIlkVGFl8yw=
`protect rights_digest_method = "sha256"
`protect end_toolblock="Jn9CQpRhJt4rnzZPRk+dOpzAubz7omckX1MrFd4p81o="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 22816 )
`protect data_block
gD6l00tciPUa6pDNTk/+t0OO0nC/UTtBwLB41d4inuAUA3i/ALrNyoJVcBnAmEQW
ptbcNp5fxEUJjnOxnedyZEuEBxWRieZFQnkRdF269oOlnXylFJBHZJKrFbrFDZD9
HRW1mbitlPJVweQHOcsBJQSj9YFpzalMp9f8zeETkRu2DKTJyCOtKNdwUPnsp+p5
7HaaNZ1mGJAZOhaEStlSMZj+K8yE7BwdEvrqd2x6Zm9vBWxv1ffPCoua5Nwl07XK
su49P6WsPZoYqq0MgC9maLjIQ5bLvt5BresfEPUuGhBiJgDjsdhXd3+PTdQ6uBks
7uYptsvDpCIrkpPaJxjJ5N+3OSXynzQ84Po8Q4pMSAckFz+nGP1+ntaQEaRKovK5
kKSAOwb5RNAMOSv/tJrGg5GwlEEyfNEU5RBAKgGFHy4AjHSqP4G8hbWkUhnmk00X
56+tymQO/z+M7zuKxxJMT8xsz5IbAu0RoXEQthNAr8RpdAJlX4flsfMrJKG0RQux
sGthdLjTnmD75fMwse3jDTuZdAF5gkcxgGS06wAklaX/lw6WqylSfCHQggjcF/XG
WI/sO/YPCFMWmwmGPC4ydBp1seeqJZGcxGBzSJ1szRuIhqg4dqF50BXrRHyst51u
TeO1fqZmryNKhTE3L3PuT5sY+TxE5xz3AZVXTrYzcY/LXipupaqcg9MIdxWJ5Pil
g5UW1WuEJH77bAalnB8Kvx9CEa5t8YSN/raB9js4nVGTaOf6YcbWouL/+u/TPbk7
LarRVLaQvsxcteJPn4tTUr3sZ+ucFLswN4pfhSmdbuWWjKG3O5+wdOJiPUbenaLV
DA8RRZXKqmx5QSZegsj9lYZ0Cvv/wr/LR7xGjYK4fqlb9C8YaRX4jWexvRGvxiCk
uxspHbMj8xc/WK1C7RIMpTH2Z3RYL63fMsGNCz3tirr6chOr81ia1XLqCP7MwSuc
mBhtiy5rLqBxIS1++IHqtIkx+5s3QZGAERkXqfKvw58wARU+j+0IGwr9ehKMQCov
XLn+wN2B3P04TFZlzm9eAqY5IsoSCfHDMdEfYKYsO636oUj/OA2OnIb44Vac03oy
coX/kIpU7nPNrt2947krHAZf40punlPOIEMt/7feoXb2xyCVZ4Lok8ZhwoD1+Au0
FNwDQltMWFHrc4m9Q3+ZXvtgWct598oO6ORqoC6E42lIlK+ClDnXAGLB6TRZlh0d
HLBZm/tZHdrb9/O8HvbRPm74UFAmv4+N6mph3LPhWziVSUu2Q7DePtte0T69/JRq
bUmsjz8Q9+zLKP2CZt+811AFzItORKphbkRrsr2vkQ8xOJqX3nh3hF5FxRkmPyCU
msVGLTZd5O4GwKDtuPiar0Ns2kAEeavyU9xQlDnEygeSXiLOCJb/P2pQPTdY4p32
DQIV+8BSDcLWHR9BQImOBm8Y4IiiT+n/uSduL3PwvGQfPdZIKWqBS5lC0mecrJcy
Eo3wxhYD3AQL6bUkcP8LNMANSGnODwaMDDEfibPnyPE5ewojaF2BwW7w5K1Rtd7J
ZobosLhiB4zi2IF8G0wnqR8SXjHlLBI9ZujxH7RZ/7GsNJ2H7oavmHknBLd24yC1
VrWYJ8350LpdVXBYAHCusJJnpMpjR0gFH49cTX5LJTUIk1Oau+Ls8McZwElsPHPY
6sFzxayLbf7SvHqndR3hHIoLbrHCjXQq0jgJ+LuWmwb7E1BMWkMAtU8XCgRFtwyk
v8JP6BTjjlse0E7Hfsnp1R2kOQ5Cs5n5JZJ2IdOaxalpHHdF/yOigdnbftp3JXrs
S+MBt1Arv1emEC4DmFR2GxqxyzxAeT0EhhdNCajf5TTkFkAs7DMuz3hyN+qtJc6g
TC1Wu4QNcA1KqAlpKFj8OODAQ7mSZZ0hVIclBnE0NCPDhhLRdkXEZ0oQAKT4ez3v
ZfuNQSp+i5Kul+HNMVaPnXKfjsJQSByGLMVzfDtfXVQgTrWDmvJh0PRQlV4Ezz9f
4CrgqakgMTdX6V+VluoPs2ShFVKNN3Tcc05s6ksIyvXG/TJLKSGnqDlABllOUl0o
4eYgxlm5S6idRIrUEO8HYIt5Np+E1kfWL5N98CewUC/Hl5Yt2vO60E0XTX9I+nxb
L/KVkGyjpHuG7CYTUXb6lNsY8epDd9YZ+p4W3a21QyMOk8dJw6rEQDvB0lU9Sxp5
KDZ8xLD2doZDxhQbzJP/OiAdZR6V/wGBaEsYaLAG8ZC3+dw8A4W1nMZPHxDfuaQF
kzpjVdjyB2ljkMmQOflVkoJawOpmppFU0AXcukPyVYdV9OMW0gSysvB83tlB9pjj
S17C8lM+zTIXQG3Mt25S8oEa2mmDiCxirwxMyR3kDMxcDasE0DQYt9i/bAX5MzBw
v9WoLKdVTJI1wDbhgvMia64Kir2qLCqNRAczJEVy3JCCoMGGECzlnqy5ocfP8z6K
vBl5qT1ICUDanmzfF8t9JyrrQd6nWm1yin3A/HKcH6HCV0yAdSlbrkGePjqN88H+
cCO6Rhtr49iCKxLBpkcfwdt6Cy8syUF8M7l6TBbUSSy07dqmmL8z8Gqj+WBipNwz
GgH2uQbraepjziTPEXx0CNge+eDuOjKmQp5olYDHiC2d5lloQScXszfm9t1dTiFO
YEuhMoLVGHOoDiNV+C7tVOWDys2rmy4/+QBEMmqSIGx717twrqe+ezXpvPXl4ne+
ENZ/kp/FquqPQBKEECmoJ43QV1aA2jx8NSo2usjwdmFCtNs+8yI3ceQiWBwsdxGl
yBW7phAhOEKTCe9/g1gfHiYUktRFToR2rriuN9S9Shjjju5kBzf6OOMnimJ+k1vf
rghOyX2m7JF7y5d07oP8wSXZeiSX5VJ63P/e2Y3w3bb4Sg454AkIbflZi3uOIdc9
mecbUerRYvGZWjIHGEqBNaEquIvmhEZ9VkGkanMfR+mWxUgnadFKEelRAGRz7qSv
fBW0colGdNG+66hR2JRCaVSgbMFYySKBDBE7j4Z27MqUl1aknMjccXoCLYF84o7m
t6F4M54+aeo+Od0RDnEbnM3fnVZhOqgLQbuF6k97akWuYTzyMzs+bwYDHDAP7Ojb
EJo2PMp2tebb361I7+K4WdsM2RI+xeP9R+482lUHjWgbVDkDk9nKS+d4ggXADlbn
nJDYENxM5lEO0BBdH+XZ8KuAfCdFLypgp3yQ7dt6W9Ahj63JdmVWfWxhVAI0YP24
N60XHZQgTWHrFs3S93JAv+X91uhKn8mPEbUl41otgHImf5GaNJDDsBpMY9woAKfL
aVNSCQAleumuDjj//zFa1sx7Z4RSLxdUC1r9YHzq4viIs1BD4rX1qbKuxvgR6Idp
MoZybwFRhVjF06rVDiH1RkjfNkN1UALuXttg+rIsZ0lgfo+IfEYNv0GvwQN4iuBh
AB4AoGLKnHLB1kXYXERqrEvXtFxAJy30SKwc4wG79v+0gAKqOtDC46nqAKRAbQXT
m2cAfZAK+bilAVswZ+nDHYHG6NPps9PErLJUc0FY3g0PcnMJdnKyOBJ4X4doz7kt
3opK1rkQ/IS5oE4i7SyZvPjASRIRxAM+vWcwv9cXCQi8jdj6EcrJEdGSze3Bav7T
osgA21e2SFHZ+W77eTZBOqUqO53KyNBIdomo1Kcl0TYfp7yJGfHLpHyaku0ylLw2
LgF4wxwfgSRzaqTR6evYi3xnBNUilcFd1vE/pZ7Dhp4bOrfwl9s9WVusKK5EsP7H
fidm6pwJj7BCl+IK1T/yJSCigunGpoq5BXGV0ii/EljGl0ACJYmgpyqLtdNDTSmf
IGp+ZLwjYyzt2cekWly+zQVu6UFmywO21NseBNBcV8/eZ+0opFJf40sM8bc9eyCP
0Cy0mT0p/bQO6GNCE7ACt0ZG51iwyjXuCRi3//xSuB1YaQRkKpY2xPTBS1pa5paQ
lP97kmOmo2cUK6+O+N6HTAJlyVNLxpKnJhwXwDv0I0GiOXqWBIlF7kUKMhtmIyj0
imvBZTI5BRI63kRBpMiirC7ANevo1MRVuGWadCtGmaQ9sVoMPRYHsCwJArCBGjb7
MUk/+po18T2ByaVOYHuDKPtnvaGofmttvvjfq762XtrFNGrsbEMZpj0iKibGskLS
oAgWGNzsHbCcqnKjNZSMG56l2s4mW80FrkkEQfQA/tb5Ea/9KCiT3P02vxmWRGQz
AWrtzXlZ2d0yasquJCu0P1RaFbPodq5FkDmid8tLWXvpL+xE33itOdtnBZUaLc2/
0rmzPk6E9luVIBQhC6uR7qNRgWJ10IZAd54H8U9iQIXyGBnZDWSpQ7T9MY1i/8xl
aQt10znMOAaH6LycL+fGOm6DdTXsBQ6PK5LD3OZoKpFG+nXRXCVGy+xf1hB0QnF+
AK/y6cq3uChITDKxmB+djwBPgn6n2tvBzaygj8p/uDwo/SxQ7D2KmJZJe1epVvOf
l/IHi/W+8QSjg5oajjYcIkxflpUvYCmh5jhjpbDqljPWfSC2/B80yA+SlXHE5ARo
TmXjTXH+JN/nOZC4qKIHQxm52qE4xzBC/RuVGnnxjn8nE4QaHvPQ6+42qZ6M9uBX
2iBZVkHo2bFy7EKCfaoLD3o62dGekdJeywQCSNTDSnRjIC9f7hwkRB5ewItJYBWD
J2yQAQNEW5zse3OwOKmKYanFE6qrRvHUBxvy/Uv30nlyy2jJWvUGWcwsUC19wrlt
JMUNKmSqHXNIT+f10KYhTVaxrED/nzd0k2xW5goZ//SY7W6wgFSMWPyJmhzNpCzB
TO6b/Fh1Alk8IrnjxmtIZzZr8uHYQpAYIlEJu7zWzZY2ibFLyoBO/fMNgMlUeDyp
gpK8vEWrnSmDBq6c4u/emdVeYlN8r8ldxJr5qdz1vIKlFaw+EKzpd6/Su+w9o49T
40/EOtbLztTp0vPGZ1CL29o2tCExDmrhu3zipp35mpVYe1tarL43fxshpVUvue81
Z8cupIVTkFQO6MtuVJPecTI3+fF3gMKz31kE7NVjOczIwhOCvdLSoJaXEUSPILk7
IJSiRK0vOCwwDJaKOcVdOoEOd/UNciShmjsEr3iDBciy18hdA+xVXl3dXAw2DFpL
FCLFiQNVa57eYXVpK1klVqXFfW5PGeYdCfsVv47iVrJqUM3WgNo1dtls7w+Vgbwp
gs0HeyoNfZRwa2+hU3Gn9BiI7aiz1/dF1bOzSVnVIEMUA5qHMmARUtO0B4ORiaIu
x3JjrthgSVTaqla3Y0UoG62wZAlz3JnqkPEoYl9m4L+nUK/nRVCJx48vKVfshb7O
Qw1qzqkiPdKb9LjrOOrR48FnbVdPd6CwQvtkKAgSiIPjjl9K144T4FWvzCLJUKPw
QTZjK2sVexz+MQrjuaDPGH5ogd/ij42r6z98fr25feRjO3XDQKVGx7MxOoEP4+17
9L/3qdqcXJNlWMaQt7ORxdefeMBoO7oM3GE5F4Do+tKNJxhZLPAlhxQErYFd1h87
7UQivPiIPpXkixoey3ySgnPb9qDI94W6nIfLuTsVP4E0P8mo8qwO2cbNzJjH6vKM
2bR8VH3o+sYC1EGeu3MdVcUCggXELUOQjM7rigkf1aWigS/PSKyfUt/Lkau3fOA6
7QIhmgYm+vfvJeQOa/LNu96gw+U/Ia8W68VhlFsFVVrtTJUGjEyLh89pAOe1NXiJ
hRbRjyUjvdSYsjeMg1fPx7S1+sgJRIwrXtB17cTGHAX9iYTn0FcCIG0daUTHy7Df
bpWAONN1nV+SD7tA0fy72sqIW1EJ6T0bxffmDWGiLb6k1h7ycYWpcZ9wzdDVyDX5
geq5Wl/OLZSyWzbrl0NMCwLFwKReCvhySyzLWaqIJOGIE1VFN4qi4RaQe693z7ks
gfYzoMee6Jc8u/jsiSONsXJFeSJndp7d0jzILnt0XoRAfwkRn3Oet3kDlvQoDiUx
1ElIM67K3zZkdXRmunCO4BFDGLRsmudKTWy7FfdF5y3v4vEQeNnt8KKINZOQ6Bby
OlmgT3LK+R5BIcyQV+0/Yn/fU1MJRTftnVq0qsoUiTR+KyctrkIA637/iBKo8q5Q
ojq7cQyqFc2op2s+3gAbMp/O9/WzewHKYB6ykvMR2bKMmwJTwj1R5l59YU6ZKR3k
ThaidL4zDUY10L2MZTC9TSoNjw+oBzVG7xTUj/ARBxbicDeHv8OyK48I3GvzuW+0
c2a2lKiYxUfN6VRlpCAVAntqDt2Xw/nmgArsrKYen19I2wZwXZuJZ/VqElN48lE0
2urBcEH+rfALtjfYDRGgYM/Z3KW0/UZ8tYWeRE4KrgTupRnjR/0gfQjlqwQprFBN
4OcpoMPSMRzkIVfafKOHyaA5VNiIi60GEmaPz6jYcd9iTfLtysJjHQ6FROZuoCfS
hwlFqxgGxKpYJjRenqEkQoZgSOL9f+okeyooyEH8agagVkahjqhX5ujeKlG0eb5Q
kbfK358lvnq1baK0iujq5/TtcKuhQljrSjaRQtqCj3B9dshVm+tLDUxjhWxw840Z
DPFttLdwXwxeda+AW/WDdD6X7sPJli88IGGgb2cDhEJZD09yfLMxdt5ZgLLBdgmY
HYnLxBDNxqEfCSG1ZdGLfE0ALMo2O1KoSK4FQUdRL+KZH194TRNxDZrvawEifpzG
42xc3RcQ7v9yCDzFTM3ETfii3MPabs7Um3o0ZDQuCJA0a98OqDSs6szVSneR2RI1
zZhcFdt+P1QMpLkkOTjYzFF2mzcg0kMKeQCgzynBiN/VXyBX2RzwHIx6LCHRrPjJ
rBuCKTpRPBvE0RB54FAc9H1Uvnaenvo2fivq/Tyo0opHtaJnYFGvy2yV+Bc2MM6g
j8F4/w8V2qjukOtoQr7adNvckq6A5SQ4I1pG/dhxC4P7zIrBVoxavgA0BO95QXLp
EiYP3tPMgay0p+h6wcM1MAoDymgLAv7YVr7hTlPdiaNpayh/A3rrtpK6I9BaxsEs
2D1moiFSAs2fWrbqJMQRiR4Jz3u0hv5PkYI01PJAtssTlc/WQHwOwYBYM1q8PwQ4
EwBZMf1szOGeyBRUKDj93ojNUpowqNNEej7rF5UmbRcpFYnZp28A8srNZ+BPBbWY
YV2+tjSRvtc1FWyIzLVJsEt4EPcjWWhSMGz5x3HCI6tsIeYpYwBZ6fi742dcW2wA
mN1ID6DLAZEsnSQwKrV1/UlVlHA1qRzl64HlSyjdvGhSpSLfirrds6Y2XLyzZ6W6
+UZk7WDZdEYCefEAAjqEeB7ZKJM/GujN/g3HlX3KEhEiq8i09IZZkAWjiPngBGrH
mOXprc/jA2xNj72hu8nZ/Secv3RuqGicAsgrCtofKHkbJbnjCKElOcZ8cEOCmj0D
lCNd8YKkAR573ycHatrMRDIxSVVmw0zdDZOTv91d4eo/6Ul/5YJQm3jJ+0hzTec6
TWXIT9+jrsCRi4jJ7Gn1bZGsuc1AdWgAen7IfTY/b6DzVriLRYT6VDgfh5xtGGUf
budQ1DZIphmVgQL1rO5YQrggqNQKZgDd1yjgShN8XXKSG6eCjoHPJa6UNXKYDws5
yuTxudaoF193YJ0UjBcLOaFbzrQe97UNOHm/n17UA3QmSCughIwYsszlgQMma7m/
Q1bD5YAaKzJDDFKoxiF3d8lqnX+N7CSTPcMNGss7MOiA/gRWvU3Q6secJPiyZITB
ONRF9cpDoXEk2CEjXvAh/wYZj735bhIPW1lxsctxDk5ZUwJ7t6WTNjyOgNzQCH6a
JGIrWiPFawU+8HaUhob2DjQY3qWKfbmjjBX9Vwv8aU1lN8Q3Q9FibzZlFW2490OQ
HnzQ/0eB7coWUei5iMWrdDkc1j1X3zC/HG5D+4i+MnK7080zsFwYIn2MgOX21qDD
ylzQupY67itqttu+KNZwYKUYxJgpQM1d8YWx9bpeQP+jLqnaVJxIkGFUYlJMLzoO
YjvnLzmuuDryo2+g1KNCkIfXC31HVGWR+s9/cxRVU6tzN2rN8HUJUhWA/zYHGvfF
5eFHs/uEprOiyfqSKU8sMGP9bntOGWaYdX+KlN3/u4+BMYkK7veOq5h+6804CiqO
tUcOqcCYWy0zbWGDNlmam97ij36s5kb2QWkweJiF/F6/eKiHu3yHoCoD4TIsX7rk
7+B/f2y1AVv26chND5lGX0iRQwFAF2MFtVllC3cEKW4dHpVZ3a/LnokVog8pVeZJ
kIEXrnxvyQ6L9KaJEPuCibNaMlkCY2ExI5cTqptn2FYcwwXtq0dvG5thRTFG7K7y
rcZSehstODIJ8x6l6EN6avZQ0BNGNRPW0Vl+gS/FHXGwpO8CaguNc6PxinNYZUzk
aa7O+y6zS0cgIwSHNV4DApA7YGYonDqTrMVDi6xrNfYL4mzYzp0O1+ex3hYWMNs/
3za55jzTdgL3mphZPOQ9kUPcHq5Z2G3ML4K8GYJkSU0G1sSizjJoN+lmlM0VfZig
gvP1j+6S3cM14PzfpvEjW9ywdzIToeqiGtZb9euZ7qRFETDAtG5C0p0LZlW3QbQj
CF4IA4ZBLIOZzoRyVGHXdSmPq19MtHyPriX+cme/YDVCanlAPzu5O3ZVam2+vq7W
aUJl9oyfYmcfUYpI33kO+hMnKigUDLy2fRAAfg2AVrUnZ4sstPywcPdef+B/R0k/
QB6q7azAe98z6K3UABK2O4HAAlu4l8vSWwnanUwaZ5TBbNT9Gu1LTqK7gbgCgaxi
Y2QQoI3Gk+QY/6BECtFRKLWR/qDn6EQdXmURkO+lmrAcDzYvnPsPUGoSqBxJ0D/Q
md5IzWkZe7WS0D+Ml6ch6ItRXwUFH7I3PT4v2YnTB9WmLwnm5nPrtFY6GNGKtdzs
1yGnv7a2WC1Z4mrc0DJIP5YnKcbHwIt3qwX0HU+ZcJQthMXc3yCisznr9FWKkm9M
rqeMOvu9EHlpxm6BTryDMjOJSL7TnRAfcEN9+hqWJ3XAoc7Omp+Pg2QtN0AnpYEk
XzpTbzwnYOXOjbdhnbDDNCaVuoVjoNueBdYfOn8mUo0Y6RZgbvcb7G3VSgHRcNET
t9ND5aeIKv4b4vIvl9GivL80WwNxo4t9sT2ZWifcQU/zC0cv0d7azi/0nkZqxI1x
tHm9EZ3WiW9f+1ytmL+Br6AbS5egoki6ItSJo+Vuz9+/yGwe7uLXni1rbu486Bt7
k6/Ybsg4f5ITfK+FRqss0Lb6sWm3m+0pSdB1SL4Cf1yKMY2hANOo4FYikTzn6LmL
hOMpwi2cuUUGO5RQVSh9QtPz7YbodGJ9c7louKviwDyi3xkO0BiCmBrJhKp6G8B0
f7UuJeiZwwzAdOselBNaT7p8p8zhh7RWFBwicp8hqTsVeQR04O/6dWM1QAJCEfiP
Kuj8FcyX1hXDZ4eAfm+1979yNsJEhQcXPeTGP6CfuWZxXB7IEz3IaWbRVJAJ7QRz
dGAyRNuBGPbQOZ8vbVd71RLsweCrHxCESylptSjefGmh9sL3zGp+8FD9wvg9JNz2
YrE6otOXx9uCOWWPrcaSrvKs6EIKibT5Ku5Y23VzYv6hR9RavUa+hVNqmfc2P1Al
qcJAZ3OqAJrdtN4AfpIx1vxFP0qbweX0ONnKiW04AnoalyItfM1c7E54UIyyKS2J
xg9EI2ZVqBPlC+ll8znHBdZIw56QSoviEsawf7cY51ndIbd7hlgGCzGFoPMBEooU
1UwS02TdUvit7qZfnxCZtWwYCiNLXCGayq+6tbub/nFHfblpq96ZdRqriH6a+k2E
f8wtV/BdO7Mz0Dov18aSRriGisNof1l0bcGOyvLtjW4XfMtO+yXgLQWR8BXDNB+j
QbIKRt/irc0rlE9tLW/xvMa+wSRCrroibNs0yhscfnFPFz8FaNJy3Y/iKlbmLODh
wxNlXhOV+WF70fZZKNKq/dbKOWYAn0Ew4Av4NP+J7Yatdb/kd730JzF6gF7YM6f8
dm+fUeo4Kw/pUPIX0XLEc8q4zoOO0qtYtR3cq6tfbhkLQvHwFCcMAbbv0uNvGNI2
ZFXczYsJ1A7xwr5Dcl0kfGkRG1kYtV19eqVt1shLWa+i9bBz1nEHDUueu5NrkDq5
zqTLJHwN9n9ZRs00DbEysVEX3oICSlyjeaO3zVjS2bQ+YlI2J+rDAFqGuRi57qV3
hct/v+jAM6tTsHU1TCzJoGsyt1BotNrQMSNiDDAsa5vxc7UV/cgXceIIbNl2ioa4
ClXpAC30eU57j9GzMDyBb+qkARC1Pso0ei3fbpLc7hmiYADJv6ce58FFWskzMq8K
vYFyXWrTJLTvmzL71wBlXHGKmZoI82pt58ZjN0288xGQSxt7ip+S2poMqIdgsdkc
xNH0bahphKbk4GUi/dDCxbZc1uRBU7HB6Oqini4oVZDAvwz0UcWPtMgqZEdLvcVO
4IHPhOgyMm60yxvP1zdnT677rosV1uE/kYUSJ5S/ff3d3uH2Sm78Ca2mowOrvI9M
N7gjIkoeD+eAl/zEVKURN/7DIkhw/i+vTVRpIse7/qZE5N32FuNWMSxlxR05PULH
WkKJuQzIIj5G3nhsmkITZdtz85oBlDsecOc2wpUGXdkjx1VceJj08fdKZUNWMY0d
biSaFXvolBYVqBkxwzX16LZL1Uy5I71CC1+0D6lH5KDfvSaxOaFrtma92KvKwrs3
cIjx6ReG7VT1vwkWt0OQL7vLbt1N1CMWNtTszf4JmVX6MUjsOmPqftStK/Q0ugPj
RpkxK82FTikISS9S7c91MtCVQNNs2Mr1KfUXcrvwWN7GnDieOTLdm9xiU4nrmdSB
O29fXxs/IzPf8MwBzhlemDjchXK4/kc36uQ8A+crgaA4oWUzwlVlpXIyaK/UTL9N
Two0xYeaIlHuiXSw6CUXSarQvPpI4f8OHfD5Bckuc7kwEVtPIGP5frKZ70AtJ0Fp
MHt9Q+RJWRrtqwSXWwsB7kNgQpvz2SqtoHIfap5jvKngI9GRHRrIxrCI21IT6Uha
FdCVXLKgf0pQ07qhrwF/hkE/ZPgt4QN2x3cUg+6i+/lx10caRUNUaxEfvfSfnXID
VxOuZ38G5yT3eq07XkXGnoxiIIPrHB06k5e4M56biXXgQVRiqdTGMmV+vfay12sE
nE1Jm2O27gA8JEDXDlKBewSYtEz36b4+R5a6Kh/grZNOOWHRHX321FSbKW3ExuOZ
Ov5kb+yiR12GjqcI3WDGQYGH8WVkZl7lpi5kvXoZkEfDfaFf0qmVc8mjklmeDdl3
40bhCqhaZt0cmimbHrMvC0Q2jZTvwF7knoGhSQyGKbWAV3gyvYLr2le4+yRtrF85
5H2mIQXvmvbY+ZA7NYv1B61JinPkrPQOlizzCY6Kg/0JdSffnFAhysa0jT7rSnHT
SXYae675S7PFJa6HCcTEVarV0A/UFpJNe7WvvzVT/HAtwizYtTqcxqw1s/KKfnmn
eEdQSoSkmzFGneEQeV1jKZwHSpz86PKKYAaEc0uWhuhzbHVtwmrM64zxVOjCBYZy
NSlls4PXV9fEw3rDXRpAngxRHYxNNEwpKSIKG+bsMvqADbf0BwBKB+TsjZHyMZUQ
6Mw9lp8AmjD294e61SS5j5/qynZjGQPula1nhVwmeJ+0NTWBH4ICPy+4pzWQl/5a
Hw+ZtXxxibhGVBgd6ceywJwF3YuLc4c1E2tTiVs2pngbTCZ/SK/VGtN0THQI3dKe
s1bY1Raj47NBO55kUuyImDEs8QHuNtJPT5tZEIUB8NN06tZRIqwUpw7hCQpIv/xm
JqDz4nbsPwou7x3+9G/J3tMgYMIIAZ+wFELz/F1nDPr3k2GA0hojo6fiayXh82Hu
JDWfn2EXIG4jrn43yAycVwVpeN+2/cLW0y9OEpyGToAYVoYlOuYADAhobZsqAI43
9o9NOA6gvkux8IRzU0ghbh4c4AuzwWyrn+fQuEtYw9hlqUj6in8xhsDXnkarfYLS
q1PjDbP1jgz4rXFICDXr0pULyslH7z+6s34UO2LN836oJKr5iWhxhwJ10No0Yr0A
Iv+RB6vlysCfbZBHxDam82Ldyx/puR33EQ+6WMj+Fm8GRSQAkMrsNNiEuLHYFHNm
hpULw4lzESm1Fq+n5o89Pd+z5MSLyLk7ICUY+519pAwyCfHg0z/10et3GDSzirGB
TFNPtrfbYFiqBhYKN9bCp6EcQUjk2mC0gEK5qe8R9YCClqFtOK3Wy+SFDZdcOZ1s
AcDT/AXmGdp8ZppvM3Vtrbjri4HAaX4uLxWq323nXgkozIjzHkJKLsNdi8yahJqq
sU7RSde30Ro7SibRWB0Kf8I74JA6/P3ihkYp+HgP1eROG6NiS8ruTUsosliSWAY5
F0EPcLaXlUH2PAxlIF2vx+m6Wb0tL3ilNEL/+KyeEht8omBT+A06iyivsGhEAwfE
BXfl91SbMmXTFeMmIUD+5s3NwWI+APS10SFYj4kYHg+RtVuJtYCJqrPUIeipDpF3
zvFdVGmugy2ydUdveYaEvwWEO5knbQdILRy+WyKiqdO7lHaZLw4WngohYsK3/JHV
Ru/af5Qe+N3nudVKVkoxABsItjqzr0Tz9wjdFXgqFuN+rlvN+ny34qvv0sdpbS3f
P750KOI7OEeEDGcEs6nVurB46tbOrwMK16WZsOZ4e+fGukgmFEHX2t5/dWpFpH6X
njS0GPrvwXXt48nIr2U9traC4+VWtzfPG8YSr/nLIWdV0l+ByvHutTQhyXaVQ9zX
ih6SLc5IuMqJcp5e5XdSBxd6PzzSIg/9F98crM+lM88cSHn9/GxcUfIzzV8mILtI
EEDJkAqjfxA/8YNmEp5TjFALxElMNXcny32wUOHJq6HgsR+qQwYB6UP+jtjsGYmn
XMLw0b67M+QfI2/qFtCqvgKIMSE6QEfogHVW0FegjKnUJHLmLR94FXk15lbIYOvA
tRjAitJu+7LDDlstTAoP27znU9BO+OLs3FGdS1STdwjMGEtmJU7abSPmHo23x179
spwiqQ2ISdWqCQ0a0cJlkawdVbx1ZO19o+wVhseIyv4HW5UhRb2Mg83ail46SHVg
YlL79p1ZyS12j/dPE6YsnaEUaN8DfbitkKEoiH9SEGeble0Xov8ltEYvL7bPpaXM
LaGNlw8KRGkf5EgdXzEAzl7Ev46PIpSbhmvn3k48LEhLBrRoGyneQ2xpvPPjhhFT
4qMBJ8OPiFcRknzO8NFSyNjfZWyX4GpzlWxNTzjryPzSVSwhZux91QsdtniJ4nbN
XErPcFSDFgzIwvTFUP0Lb8X1Bf+oHV+xwNX2MAULs0xUKtqdls9fBQUXIjXptjV5
6ALZiGyto/R2VoRSqqBhxNRShmZYRfxvO2z7TqqLQ355jGQN8md91cLYK1Bg1PgO
pI5i7P44uVjdfodxkjrDmwAtsTw4t1rlfyk4f/JtDWYN4b/mhYZ09ZrALEkTqaTx
125Q5Ubz1aGcls4+EstbaFFd0qtY/tirAllkUuv/ef3dhpd/yO5Qi99idQRoNp00
pZhV8esreODXIStqK1TcEdx4lmUtU4KOerGqjCX6CKXlY1kuXeyT4agsqYXn948a
6wagTFqG03T4N84mITOzBLprTyo/FvWMN57OkeHRSgFNO+GgELfX6gyAzCdVlM3j
sRtw1yoE8LF53tojFf5ExIbDnERMGtm/UqmX8/xxRDvmVcbZSGqeOnQ2KnqZxzTy
OGOQWA77qRE4sOynYEIMv+y7nxxjdJuL/mWIZEB7Ivuj/3gBPyryG+Ood2KIhLAx
mAEhKtkSyj4PGjHk8Zh5dKdimv2fiZFqe3xyeZ5lvemaRdJ0c8d2rYYMC0KRQBof
7zwDGf1jmUJCl020nT8naes39iI02tYRDfxiC/taBifPaEV6BgoTAw7bsfpEu56/
Q1BKoWsSX8x1z6Y7QVcNwQ2eCgrjZfTG36ugP4suXr+yqNGsphh3n2pa+G3T7VEo
+hEaDNVN2v2Lr/s7LEOUvMpB4NnPOk5KlyoOxVMedLsotrk/AkSo83gBPhyUSQVF
PydWVQ4FAuQAj2AJvAMujGVH1SaYO+uOESA0Y+nd5ziNGGLeLju77Ne/DDL4iTWb
wMCijllNfLnNkrsz0LRPKyEELn9bGrY7KBoc4WNxddbOkpi9BjA/fDkTahiKPda1
c+0zNtNhs32CMs7GX2bauIei+4UPqzfu8b1/55kB8uQyXxvrq57dI8nthH6H4QK6
N5K5rYJeCGYfg+uWcNPGyUQLLWhxhukswE/LBqr50nEVpb6woETVNsyq4V3lziFm
PdeBmMyWN05vgm+97zWaA8pAUHq2gzPERwSSVQoGTgqOMAtywaC6iFlaUKfTMmqk
VudPr1pbFdoZqgplxAv5NNl+0cU5RlnC0P6fSKiWEl6m1hvYAUkWRLIYyLSCCx+6
vV3X9JOKz9UC8KAs6ZRrFQzoZaX6GcmIk3fMC7zcGoRUbsRK7/PxbSXmt3Q5WO5E
YaJnr9ZGBBefHBdqSM+9xXPNCOPSj9uYsuUU3aBL0Gmouu6ryO5QF8j7deI8LMR/
EGPM+wfWBIhwGcRpe204Hn2mnD5GvPF3JAui3qQbA9P5jeqLAtxzLb8J5Dp1leKT
U2lneyKBoq43kFirNR75R2JtG5wPpU/9PVm8f78ZhNSjZdlEjnR3MSa+sfIPZPEp
nPQmFn7GTQ16Z2TZdkR5juTwGSuLeY1zv5bIKiB/OsOg4EB+/ikX9rK6LQoTy8qf
gPtBxUXmbogXw2jPhI265Qo+exYqVNaTDvhrPlUtU20zfBGjOPBIOK5vbtDKIvhD
8PcRAJDS5IxK4+XtQmeLOwG0RkjoQqHIjBNGZwMtfqsRRAFeRbr6h6cXx2lojdCk
AO7rjPVtvIXZDo4pdVi8bUGL0CsM83EqOAm1DXVsEVKyMcgcRIV9XeC8zbRLKfZ0
j8H5J3/5PNHAQ5E3rK2bsLyTTfA96j99VmFAz1AUcbCC0qkIt3hTv51KVDezKx7l
gTBTCKIdhj0m2yNR/Oid6kHQtxm+4MnGVMj/4BhGy4LH9Wz00YQgmgZT+HYNj+Fl
GVVKiIjKYFc6AaU84GVmd/Pf/xaFTl+D1MN6X0UcF5uo4Q7wi3601mAG8heoVha2
UkcsnEj6hWocsM5I4f6bwC7FPcrZfaVZ4AXxVn9VpR5IiXeIsVuDarqzKUTkGMgM
CJlqwCtYClq7uacrcxnVploLdnN3vUiKXIlixZK6ceF2oG8YsGou9WC0lFZEo5Oe
43tw0AoGTtYKgZerZYcanFaCiOjoYKSc1xhIip/RZS053QF1sdzpishGKzclUSnO
+v6LBjrXESeJAqXA4ZXbemUat1OQ/zfea1R8HZnn0kgg7YI/M7NgQL+WgR1y9ol1
Y4UAmqNJHB1mc3mQo2ScgViBnEZtYGtw4m1ADYxoeXSOqKvG2US8ucy00u/Ev1t4
PQLjY8qW96g6EpqZdvBvK/qf3VVgQLiK0SVrSGfdvzVJAVXKkK9lpbpSm3WLfYHw
vvg/1r/3K08g7g1ZfCUaSUmARk2Ql+G5WRkgqwkx8buIoOwnU2aAL0b6iY3tEw4A
iLxLLbo8x9sjXtoNX5B5mgvAITtDPUn3WgH2B7RdAMg01qmNxbQleN/9ZlkSC/JK
CSqU+2ZAwxotsMv9Wv/XwyA9tPXS7g9g9Gn4Kpj9TIXIQ1Q1eGgqyUG111/v0DFE
xbzLLhHoStelOunkzA+2xyYKbqcocUamnFtxBGF9YkMsFjuAfbDSns8vQ2MZ9PYk
IuLpTMHJv8Z3fvbAC7CWadCFMSxqhsKTLLK1QqheIiRyly9f7Y4oXY6wf5Hw+wOW
m7mU7E9sfqfi2jBoGCV7npJ0MmC90FkX4MbcIY5dn5TYhEwkP3FRcN6tsolLj1/Z
enn7lmT6HrdQcPn4w2f05a8E4TuUG4ZOh79O0Kl6T8FkqBf8UnhHlEjD5KFpyBsI
qM0bZhm4kmTKfr6G+1FgIA94mIgIqyUnyN7aQh7uE7ASen60A/dUEPFGAxI203Ki
wdaO27ht1sD/4slyYw2mYSuOnNvHZ5ZTrW9Fvw7vhkRGpUXQqBOYn1WaCA94a/5n
RQKYMeHQnO+PvkrOghL8Tgjw1N7EIxhdLy8bRdmYA19Brc/FCAOPHJTzAsOa5EXK
idPPsVdmO8Be+gwTdW4vjg55mPpwSFQ2Njx2sDFg+rY0Dwe01RJn/iAcxGXKegIl
u5t/rcNz4hZyQFHDqPbWi6+ShzH6C6nNTRL2GFXNOd2l6Fn1hdF+ezIt7pLSI9QC
ewuSPr8IYvzueQAo9gIyMlHrydJc6+LMbMcGaGnERU3QhHNfLKC9EQOgKw1zPKfF
d8S09wVki/f2oWFHnYkpVitPDrGQRyPffQ5mcfUYZCLsXtU61wKWB/5Yk4/rnAM2
SvmhiklqCOKQLPD8zxCxjGiCS4GxWIJx16J5n63cXhdkIGb+1zyWhoaixC9k35N1
+1JUeKMfP3zHTTLXgyxJJf+xrqpaKoqwrTaFL1yj14NOSAlq3Am9HJsdNx+KFDIg
Lh87LlaWeMzTZ6WbtXg0WTjkhfzDRODOK3j4ek9yswgMxoytaZLECAxzEb0O+Jv2
fwQ1YJs4zUxtUldMKy7YlIpZNrVak2TbZnWBIkfoFA9kFFhqsW95c13EVpwJcseH
wjHfa8d1W1kQNthPjeknLVYZ2EBq0BWUNUnyxEBNaezsdjg4awCBFxfX1qqZ01ob
w0Pt6q/EXyDMg4fYZxfIAj0GVZG1mhMupRQEfVRffONvwp4QnoouLwMhoTT7U0Nz
VOAXlMk/wa5Gs2WVxxZFEkHxmcfoUVvewVtf/wxwl093v7Vh7pviCswh2lX37PP+
aY3Yhp91V6R9wQGTvPa9S+VyYHmof0B8tGpwDofkuz/Be/r+hGF4Pj5NpH3uzpku
qx5dBgFLSs2Jnqvv3HOvDUf/A3hCKdgoi7qyN6MMcytjlaVxeJ1BEOOmYOa/HUd3
+DHr0YjiTxmZG8CJWXF6zu5JM2mhFJMOcwrIb7zOymMLRk4ui9w0ia63fLcLJtrK
dBuGtIbjb/l4VtiS3yadTaWEKKvZ6BDsmyLkyVfF+ywQ8WlnrQ5NdA5T3mvTAMtP
40FXXXznyCU/o94Em2ctIFi241y0fV0pWg88ogCi5Fwi53/ES9cIN+6zwbI7GyhA
KlhUmxhsLHjd1d+jWrSAGYP8XQE7qUpJFMBUYnZXFu2A8I35h3V+CuUlBnj0LkOk
5RzMeAWGIe0q8ukSdw3l6F31xBMUQySB9IcC973duPmwgymcttJ5RxOznEEwzAwD
gfek9i399eiTVzTqfSqT6hTISLCPSJYx1hnR/22xQ1gT9wsItINHRruUoXKZmzjx
KtdPZVogsbIPqxsqeXUd2SgF637BFx+8NFgQACovCdeYU5hNhyFqD6TTlM5dI8Sa
2NkRRxqfS4tM5q0mH7XhablGHJggtO08qxewCXIUMBDTsRiZdHR2fCGjpLjdXsqI
ggEdZcNyRd1IB1VkIZ+c3p1hnp9m+DjniBgEsQ4TqGCThCzfItwDfxwyIPOLaZCj
zkuJEvM5Ml80BhL6wWt6Yym/3nFMUO20EV0DGJNBxbp/MKoKllHHrvGzxEgEv9SH
lhcovEM+p5kzYnboj/wx62prPXKzA2gdE1a1SuJTY1Borfby6yJAvzWEGcnegN9L
+rOD89V4LE31TgEuX2YCAvaZSYOnWK5ILfFprrkqTTpaqyO3L1+Xo98c0DcOfLH+
TZjb5TK5/1tdgtzSozNh5iaPvFxfjLn2nyt3gKs9w73UqJGne0aaGYvwa63N0Ns8
KzYqWlOOu14DdCxvbtQu5rZL12zhLVR2RLxpvYdg3uyfuMjP2Bd8byjGvnOm+nV8
sDsV30ICWClrqONzCXsNx7bmQ7N82EF8qB7njK52Zqfvn4tCxLL6BfxIiP5XVUOX
YpwMkbJQAXE+ekOdbh6gYNfNqMjj+ctECyHT+SMb3Y92+r7ydrx8xoDtEOv9eXC/
T0n4mO7gfbfzDaPgS0gPinjLLy/kvp4DXkpa38jkoAf4RAc7Li+6aZ8BxN9FxuvI
r3UrGE0BflQ/frSDMqP1bCmjj1GGyY3qR1PRf8WXtncbgeTjpotkUbdB/g5kIVbF
cuNRnvSkw118Ivp73at3abfPYdaklXbczT4KZr0XM8Zlg/T3DY9U4j4DgjKdj/bc
TR6uZrpDb7GI6QP9ezXyAou49RQY/XGltx+03Tzelpgy7SO0kziRWB4wZS+Hpqb/
8Mba+YDGYWm2m8gZ8hmQF+pn1IJwyKcx+cQEigJwGCIrYUsPGdqJpEmhoF6O2uUX
ubSHpmADRxf8hSEeCeFj4o53u4p6otnC10X9r9LX60Ad1VS8r9kxBK6p/7Qjc3Q/
/1QBWBwjZzC8MYnjEh2HhQ//uhYv/FynNCbCFPm2ocZtsMfQbbqyMhmDQL39FLTB
XTFY84qxuuV9diehrlMR8dKAmv7kG3Sji+T9KNiQ9sVGp2GNR5DO7ut3Wucc9NzF
VWrkoZuLMP/TS79gQ7bhFUa6mrk+xqa60noXL3z/zzHb3EB1FWSNBVabuenz82Ix
DaU2Qjc2GCgJ7TJUlWy2c67J7BwkLkfJ1c8tjVJWOwUtPg6XNm2MbWj9Kv/VCJsV
QcBmSkeqvadhRdlo6HojVoyyMxxxw2c6hwDwapeFFGToX0BX7Lx//r8sZ+70DLcs
1MHTOtyxTz7ZPRaQVEuj5TddUBR1xM6NwX4ivpvbQaMRdo4Sl5Xmk87ssm6rVcEP
XUkCLnb853ju++dVHHzOvyJf/OuyWQgt4tjiq+xiNLjQrmQz+SqMMrmvVs7NaQtD
Y5WMC/tWF6NQjRhZmg0mU+zaqQecpEyb6hxUqBBTxm0prblvUzhoUg5zsXD836+s
L7JQ8JqEbRnKIrTjj6PgS+THXTb0c16S1OTkY8l6ZKZ48hQ+1MCicHbxLyrYpbXx
c1qMYQETimTaqgc6erbB3u6kQeM2FQgQvOMYQlxUEeHKSVAxh5Te4Lj+YCiSmLjz
ojgyLh13152Zjnr8duayl/pSIgFtq3IVBUvdvuAHzypB0AmmkSZ/42lFsV8Ty/Ab
XKR/tfJorpcp7KGqbpNlXHJUGO733yYLZMffHbwuDGT8DuP5gb5w9XwAqvYGuDaR
SX7dTY5jXTZLR/p6fz6VB9ZqThD79g6f9EDZ0cuTaQxu2dQwCyPlbZjfjXTvHDYh
BnZpk/8JKT/SmwcpREGnFD41cIm0Ws3fPatR0IyTjZ0xUSNVT5KYVfL0/Ed1aCFI
6cy1HzqJFLJp/jtLyVImS8s2SFBXMYojnou7Mbmm8cg06WcIMGdDZrsNofIO+GGh
0wmIttotBGP5NJ8j4vYVyDf3aXc6YWQGPMSPs62mlhHUP7FLuDfHzW1hsL9HObBk
idLauAdiTc2MH48OcDVr4rTqRBAqQHKoIabZu8mRnh9jG/7zvpHpV3oypp1zOo8L
K7AxeHaQY3s1I9c+lLI+Tr0GHL16cRhb/lKBcEZ1TBjJtSMDfLOZw4UjtK5DXtUW
H+GnVeSx6dePVC71zXiogkOx5bh5L1V++vhveUO0ZRg9sans1EI2p56QTt7YBJa9
K//MvaE58ivz8BeArUdFRciFXk7OA25udn9Ur1GlgINYZaXBSHGejvJmOPjv6UKd
zMWTsFtnPUNr6Xzg4OQ8hLNDiV3dAxxiAjl5mSw8R3tNyaKUFNAMIWNHE/MWnIXp
KxfkuaNpY267mBTchHBLuLcRZ4VPDMoo6Mwx8tXupUZrd6qq3fxU9GqjahoypsTb
C7i9eKuJnhb8GBzMilJHqaI6HtIXkR6ZCnC5xxgFW06jGTrq3g87uRRoOo71TG3n
rISDoykdVlcrJTIWbi5EzTP/s/pwtdLf56LNYh6hG7N5Veib/9w6NzooqVIjyorP
DzuGcak7kGodnPSDtiZ1QtytTVaOUQyKlps+DUGKQCbvQV7MmiRqOOhK9cFkrEs0
KqSb/2DX+HRpG/mOMwbMFdBEKQZaQMXStZroc1KDqN7dOyK3R49sfMgv5asYiHhO
phuRNP/Qcq0CNQMujPkMrKnEa/0JGqzo8UmcAhWZ5nwH7GZ2MNe5XpKOBwOIjPPx
m3NHIhfY2upBKYxuES4LLLwxYl/dWGB11/vnzEq+Rjn3t6mUs5MtjPg1I1snjFOK
4gXBT8RGQdwZ/AjWY5V5lcAY7y6WbUc1w47qa2EDPNqrADfxFnFKopXGmMcEGGOI
0Wvpujlgh2XnTS4fxepp31qG5WrRjhj+3pE3NyN8d7nUmlAYX6VMIJnoET9mIMxT
N1HgDawdMwjqKodxjM4pSYvUryVzv6bcXS4+UZXowG2gtVNQLnkwZkoYmMf/e1xd
f4kBxyb9i132NeDVHRSpomfrW3nsPXibUEuQGM0rpb5SGv1aKwsLE8FUISjtrajh
su/+gaUU89bZqeJuLo9kMYbA7Ls8N9rABjvnn8vV1YJdX+EEQ1uQmbRGc7V2W2gm
6WXqKkl8Bo0JRRFd4HTxvKrQ0oSkryZ84OX5FjqO/Ex/WEVrpdiF3JrgEmPnMFcB
LdylVmu/tpMoztxutl7GtHQDzby0RBqfcSUFVXkvO8CcdJ5xKLbFGHhQvtG/WVe6
ZTcoTExIPZlfXVtPr84oKozMOHvIJQBnFH/9eI4t7kP5LBhfNF+jO/c4N06CPG8n
1VadOiaTHdcOoUqWZkwmxI2oftpf+tKv433eueXBktKpzdwF7sWHDMqfG/Suz5Op
0MM1A2HO8He9XJlfsQDtGg7tnFAXo3GfbHmKaGu2tXOFCjBwrX0vvy2GR/bIjaiB
ZF5MXoZAXJxvl/dzx8C14Hxz3k7NvGq5qGFH5yyNsEbZNVLxSgiSITGbT04S23Mt
D+GIrQwrwhTdgBl9Z0fQ/g/D3pK9HEhbL/gD99FuqAN8ucwvZDd4HqnoUTqO9J2G
kY8uqdZpfHkp86zkB6YBsdmTmhp+SLeZCs5HUzLs9iscLav+J7w0N4fJhUr2v9lr
kwHw4YDfyrGpcGtWkhpEcRcqal7Ksdp8kyaHcdgXMvfsz6m8+Y8JY19RNA6awvqI
Dg3zvesHQD2bcL2JoMjWKUK+LGiNGzCOcC6yjo/X8bcAogIrAs/rbAt/u4TgtxO8
oZ55YlRuPv3wJYDMALrbRLC/cIoC21/unzTwMFegrRnodB9w774+SXfm0rS4iS4B
wk5POfUtKo0jpIGHIR9DYVi/UFPKUr9d8Ilq8D0TLWXAbAovdByjQQ/T/FA/GSSc
r8enMb4Q3d3RYiO61jiKY/0QZD4qDqh2a6dWR6xagl/BcrmniBx3UbPZ7l8YhGhp
uhOW7tgAjsy+uAqhFzmfxzlLWChiWjxy+oBdOpnZoHbgQYak/hVk3BhRFKtiWOOg
pQA6cwLyw8gNjDZdyAUN9I2qu9aGEkTn3ArOHI83HzxcQgLf7Nmc/jqxTetxvW23
DF9/2vgyWbiXPeYBe2ZSZUkaNEEY1tpgbEa966M4ouJjsXtSOBqUYxRYtbittyje
WiEEAOgOr/CvdNJYBdno1oi2av101TUgGon6Azl4otaEB2bFzg2rJxu/+zq5df3i
+fMx6k+A4LTBRBlWaVt83c1v98p83MyJVIlkfAkBIupJsMPodXpZzpkuAoRcYFGm
P4Uzu6dRV5pBbj5iEw74Q6i/c9//CkcA0hpS3FsWJC+dccjKx6OO84cgzX7TllRV
RlZy1Rz5syHVImUYM20xopqbyAyc6pgItBo28+o0xGranV/ngJ4iFa224HwauezO
Nla1byQbnAfWQlhAuDTAMBHwxUBXeycp61ZuNyxu7aRVUzQsxNDCY8hQXwgAI3GH
jsWEvePPX9P4Y4LqNL7wAnpziFu7INPmkUoBYZc8h6BvvAP4y9pK31YtOtR2ja28
5cf9tqs1C61ejSFWGYlDS0MdUABwH/P+udjXgScX/zpVlUV4JYBU8LH0+ptoCNIr
eSobUt0VEs7p2eSo0qI+pkWauazh76zbfIAHwrc2oAdajDnbDnQApbEVItbsXcNI
QekjuNTaNR1uLR9h+fYFisrqYwlAEcVR3mn+9EFlSF6NyT/kS/zqgUDyFP+aqPwk
Ll7lRdHbYdFXMelswwT1NZlvRIxCM6cmcqkUfgfT6l3RKQl6QIzPCBrTO9ChULR2
pr8qDE778cbynzLvGe/qKQY1IaFjbKMElmBZDoDTtuiFBfvkRLNO7wlGFpGQRzJ5
tdjZ53+rWcF7tY/wEl3WYjNaDq0q40sASmKr34fDY6+EzSDXJE4Ts69V0NRb0LYW
E/Q+NUtJRKLcvl/Yt9cUxTtdZLvzvHquEtDv1a2SpwRByVam+x2Y1G8BZpHNVc4k
Zuqlf/1106fkDwRhy2g5Xdop7hPZ54YeHfDNbTuTgKnBqPgt1huC6bz3SXKi0zSd
dg7O3f4AFMAgZQwX4qTDDlbaCmFbvrdZx2YimvET4k+BrW3FANOQw+3xro5uCA8t
gDl57f/rD5j6Zl2IFkGMAuGAptJdRIBDz+rqrbN+GcN/Mx5F31j8iajmdXILLdGV
AnRrHhYtH2juVXC2y6yR5lSrFCeDIP+QtNWoe8u69m15qG2oIKpp/ON4NSutXW18
uEe5/ididTQx9StBHOeBx4/85aE/vinRAWO8rqv3V3Vji1JaB81BwSXWJ//eRfd7
SLxq+ifFUfqfoBBz17amFpNW9xZ1YeEDqocTZYl/6zdt5gqLDOWv5Yw+O63Ut3l9
FbsnB+mDDDgjvwitg0aNMh7hGFf7ZgUyN5pIW57LS3QsXnXCMUEnxawB8xdlgic3
1B+OVol/1/RO6FiPSlJ4/jEHbLWGL0COYaAk2iJqoP/zE5q6CQdMtAFp7ocxQbCw
yjDU4qwyemt9lp1s/FKNygU8JV5y8v/VT9EGWfQHBz8ZMl5MZRzCcXRqYTKUjm7d
J+MGZ54cgVxYIM9mvBmMiIzTYrioXOBLkG7hyb4Sbq7j6u2CRcCv89gAlZgMQUX7
lz92ER8fqvaGxJMaNftMIf7tR82SRhkdBnlplXOq+Q5BEpiA+Q7oqdwYQbLqAKpL
N3CxKRYt7ELw91AiUOLnnMRlW9fjvfy0myZ46rkJyktz5jw0R031qihB8uZ3cDF+
AC4Hyp4A0An0iK5lfsNIv6RSHe/t39uSwJ//lESi5QWh7Z2mVvE+G9GZnlAmOqwW
2NSK3YbsIYu8AlZguefFS7OMeIRB6I2B36i7Kv9acNHRl8lylk6fibvaHVsJ4P91
fl/Me0ddFkuFnCuUpyTarc5K4K10+wi3wp5X3pE9qbkYJTtQtrzdFW7cO2VKnJGg
hS+rAfUnEZ+5j8Spx1DwO5XG2D1pXvbnjhQZ5vV4alnQh5zuFXPH73aG6QaX6q7w
4P0TkyvFJl51vk9zBOUtyrGarOEI7KrH0gf3CPdYaXcOG2ey9hzZ+DnkF3vuUd/K
nVSM5bU9TJdGvttvNvLG9GHXvnFnwTbLRFPW7DMDaSFSFP5GHkZG9WPZdWlRBIqd
rHor7kan8/PMCBJDkqeovZB9A6l/C8lVJbHnAglC/u0ih+WK9x++Bj+KIUc4VwPg
RvLQCOKnpHLxsWLUePfIEV6c6Y58I2YEECJcEwwQoG6Tj3uR4VUNmKgL1cxGEdcJ
8D0SQntU0dlzZ50C6uP40HfDp4pZodaDUOKqHn6QeKjH9qLELBpC0/WXLQ9WhOcG
LBpUz0JAIIT6xw1wY+F3oUGdkFc6dJcsZWTapc9nAzoS2rsqEKzR72fmqJIEQXb2
B8S+ev6QyavsWyc8V06DEQrahdMnjIoSU2jGuUZVMPyM+MZLut9wa+F/A6UsFrlc
BPvURoG5tZIYCSA3o2D4dLty2Ye80rSejENyyIAkICNPCnQsYeMZRWSCglYgRPAm
TjEjoA27bV8Y76CFtdzzVoGbZS8ytBAnD52pcixZsYMcybLf+A/8ocbIYRANEtqT
S1oCS3zKI2rC8QF8zbZf73srEEjV9UzIyFbHDRgKIxRHgvwy5COszHHJ0qZ/o+4l
zalSMukO/lpo1Og0itdMNZ73chF1YK6UltgnQ7pL1EFarRrtSuD/Ku94ytKSrL/J
GofylklmvV0d3GkU5DzHyooHZu5g3eENokMMIAzkZ+cELrjF7HccPVyvAB3Mcmtb
YPyiBQEhiLARnqitWGxo4EbUyMKvoWYGPyLXv3eYNSjziBAOGbJHfpNen3gB5Blo
5qo8ueo2LB5Qb9469ycbczbR5mgCcSuUyMOPU2Tgg+w6kjFZQE+p90oIfNIN6SGV
XdsngyO31HAjoXOfnsat20AFNRz+R1I6qXex+gxzdXy/eFAzFZ+o7Mns6GHheVhn
0833aeV/2elcFgLAlN2hVnXcRriKaQGl+tXcUg8jUEHDD5ntmi4gZhgJh+f5aOrD
041EGTjwgktRWVAhfchQMQ3GPRSAoWgPvIIoXkDWEnpa/BljGFobUyBw9mo5RmDT
aVYSrQ251To/lCxVGikouRMxPpU41nh4V3zW467CrUMIWAQqZEQG0EROeNOFKCMF
yacFYvHrzwoSR13CoNB6JJa+O6DNmfILi1tDdB52KGjXYzkxFUnUYStJn9Zz+NIw
pVYvOb/1M7FwwJtNzK3Sb0OzHYcwZActpvPi51jV3690wKL4cWZrKyetVE2/RVDR
GWaIIicZicLjg/j+lXhvYpgnJNf6BzFdwDMrizA2h2r3bc5OpSYKtgbT9yKfrvVe
gQ6DMuCWmgy+vw2vErAPyy94Rx+/xTooNFXh4s4oXI4Fjdhm0qNduhu7n2i1H2y0
L72tHoQLaf0WKsf864h/sjy/pN2Md+PjlVtIkib4FNd2r6iUK5gnC8wtfZNfNFLe
Xb+GT67AU6YR7u+mnRkbtURbHGpNRGessRCP/ZG6sZ0CtxicoRVkg9BsLrtRM19T
M8cCApBJjz/fFpiB/0Uvg6LdbdDSeLINaQbnYxYSBF+QMCgkflutyAp1Dr/5aFys
dis1zuvxlxcNShY+YgmkcwzF0xVuq3M2YElgcW9/pucN7kmJkWBwxArJxm5gpDAg
v56yieanG+xg/vDAdMbmHqVKFOrxDmYtKFEHBOCAipaGsXAavt8eHHzIMMdgxFbo
H0g4y7uwE+Z94uCARM4Jiw8PtA39blfF85UrWVJzTdpKVer7vY8EgSOxkV8Rl9KI
em7XwbIJy/Q/XCSjN5NQW3daL3c/RjjAOXIM5gaxusVIyQaRUse+fydR8qXUt9L0
SxSR5DU8rLpTYb7A/7NklgumtZa+P5Paq2KHMotbVIrSNNLlkgQi14UNonxh2E8q
cOsu+fQd8U/c0OWvTrQVh9EGZTZW2Fbd1yPgY6+/vdyx9kfv2ClFy//iPFcmMgVw
sYvlmz0/XonRrXBJ0XgjvudwwrYO77DLxwOrfGp+nAhp6us1Rgt+P44mycDMAOCQ
6CSa6u2BT4CRtXEqNgIHPLWwzz54UvnK6y5FTnj64JW/oEKv/2GxVdiTK7wmcZGy
mPEg6nyoCxVX8iGZImKDyQhza0XI82ukfxhErAdFpKEdNgaFLqxjZTb3lE2cSaTa
Syydc07rOGK12O+eZtzzuYjkIJOBPylpHIJe03+ETRiadfNIpbEEsjb9OFUsAFNY
iF8qY5epcIfIWYdm0yjpJvaaT2lmDEGItlwK1ZEM9eEH61rD1rbEKm8qEZ0JnbSY
+wMMNB3TFthyqADBwmeUMgf/xZxtOWimaz01uxmn0G/3rO6fDnbrfUbIsEERknZ4
BmvTr3D9XsYnLrJpGMhusn8oDMavn1xJGMCZ1orJ8iA4/8YK09BtjFo+ed600HnT
/j+qXu99QnwT0XIKDLm9RsVwbIJwr1UkQOQ3I89v9EuSM6HZIUZ+kiNrf+f9XBQj
aJBDfYIdXJdcuN5mk5CgEpcSMj42+HFqvphV014iQSa8XNZoDKEd9Aes/C8oyWsK
2jlpj+N3BPRK9oicShSRH0wXY4wRu9l9kyvdzZIxSz8TI4Cyd7lqWZtZFLLixELj
XZ3FnetQh5d6uK8+qBdxVWi62lzdjFAckUavm076sXtZGR1FUE59FRcRuDuDl9hS
25AHWt+hedYOdvALjcWGVVKQYvNnwyahrInhU8Ry1bu7MIdmyTjtwPjx04FCCnWe
x9hnliQhmJ3XeV5pX/eNDHb1lLIjeqsNsTDNJOn8mLnECANo9k3Bn5BFfRXTq1Vl
69b0BHZ1FtpI7m+AJxinL1afx1AUIHULSQ/MUJWf5pmd3FQWeSnlpMPDz8eK3jub
yvv46f/MwhQiahd6BGSipIbM5CkmPeSSk7DNiG+V7mVjrU4w+GKCOwogv3+ZQ1nN
CPCm2Ixi/QhDPP/zPaOvugU6Q93N7Dlg1n9B9VRbOmgpwPXHGNNMino8uMZzHWYv
/OsBP0rrMobq1S6UJhY8rjUqGzqVI0ZpKRhjM3NCGJrl20VQwTvrXbICHfGJt2F2
/Y+n0bqXeGlCmR6mUl+kiAGXSK2S7pMX2NnZtDdjFqvwB3JXrIDJx2KVqnAsefHd
uhv49eSCAN5MDOqVWw3rJksxtgw01SGbeEL11Waw+RdIzpA+2HVf2+K7Mo8HYsSM
dRYib8wZtX0WtBohsJtiLYTCD8/SrfaXCybAeTgXVGp7s2Kzvu0gvw2my8SxRIuO
7gogtspNXSKLUGXp6zYPaujv/x7w8lJkkMT/MgoV+iR6PiMY9bJaiBWUUGF7urnT
by01NXxxMDkpiOW/tGJ3IctoL0wXedBS6Oe5JC7iRcZKeuuYbNORhW7r39rAtILm
y2d1theGm/aDrg4YrB+JcUVWN7A8HKUb46FQa7DNBMPublwrQoWpWpr8UMBDyHlo
T5my66p0wnGMXiH0n/Qr+U6HjUKBKcwIctzgHbaazWhmxKrkVgBEEGC1PQ/U8oqo
CyoWE+HWLUIWUrrfdeAWodBSzD91nfRhe6I8vEWLGZ2nr7iB5+JzuzQJyUMdEoZ+
JJhZvkobECJosm0hx/u6A2Qy3ls8wTLWaowwiF4mk1pm8db6oBBM4FLxRxxy7Shp
08MkiTTXx0J43K/yJoQTV1S8gi40Ivs5QWJNnc443Jpi2hP9h/YDANdB/+aRW44O
QfhSPpssfEcgkgcMvQcF98pNnKumad0OAmpYDVGyrgl7+Yqm/iEWKzC0HwgOXA4y
A86I+7dLEkExO4pegDWJc4rxxhSg3+bjhM8AeF3iBme5iJy0bFVldxMWS3f8RsmK
xX5vnfkBYV2Hh27LVRWgHKR/0gijdk9U8xrPt9hdlZfgcQrgxC0M4zV86DRQ5pAO
f71KCLpXbG46llGdfNIcgNuqM56D1rG19GsXpMQn5s0E0XTIw1DtF9JP6SFtWEiu
zHc2ULrfy4/qo/dCMNyrzNrVm5A3iglhVDcSihoLYUt5BZm/MJYTxuqwt2mTxgmg
fM47RW6JgM/9A101KAnfGsJRjOjDolBQ5QkSnljX6Uv5bFqH11nRhzMXXoONxu4Y
4ZvkM02fvywZjOTAxLDJ/vjg6J9/hmFblf3R87PvMbpgxhYhZKEvJpK5m4xNYJe9
muhM0Gf849EVZX3nMeakx2oUv4ayzUlKJwhczrJ+vOXk2AiMlOzER7NQLhV4gCCK
36tcdZHzZehD6/Oq3bXO1fWlWBEprr68AY9NynxLqzzu3o0e3MZD1yW+pTPSVS2q
QJ1qYBSyQG0H/BLYBi0pnZrtEuw6vaYrnfS1Mh//ImljlEXk0x2HPaTBRbDTeCgh
ZNFdThzmDcRQ3rKWf5vo8vdQ9ZyNzqC2o7XVXxde/yJyqzwiQ4GvqdIOHHbWx3ak
e5lXwNnhqGOZoEWiYcpd3M9dL0yc10+GwENjaQnb9nSFtfd/zD57uaKW+IuZ6/7f
vQ26O6bEzy7SxD33MPKto7yj25aaKdpusf2xdOfv9yIznbFmJRS8f0Qp88PaCqy5
f2YxjT1qqqqDHrUlZgXFrjCMxzR0Bna6MPfN6N6O/Ju2d92ObvBiuizwJwr6tMMO
YS8xT0XZ5GT2sUbFBCK8l+vD6+Ic5CmEEFW7jHh+t5YTFrW+PQbBUAp7f7ciR6kW
EqHBclRxDCWDS8sWXPnyMCTp47tcLPB5trfhWewEGHj67wtLdGKQ8hdAot+9oOfS
EnqEYLrrEnlOepuJre0pjzjl9MbpFxLFBAKIxNtG9pOrlvKxO4MF8WAxytJgamzZ
G1Qw36eSj2+jFQd5e9RRKwBLAwgcpOSmWXzrejHkfflzcVc0gMX0scwspONYLdR7
C7YZwjQKLYsqBXQ55mfI8UI00tPs+CL4nfdSe5M6MIztDFamdtFBIL8knbbaQgrT
GDwWxJvz1t0fgCu5SVJnKRuHbdOgthcOA0B5elCL7MtFPZBAwiVfUpvhwMS5YpIG
IqaiTe00C4t0ysftI090rhK7Yt3NWJkkAZonHjlBIInUt4sbi/H4Vx459oI9pMfb
DpXpxXvf44vMe0FTnFVvcFH+Cx9W9Kaf+TT+3MhX2R+iampU/xU3rSxnosn4h3C4
Kr6/Sn/iQbVFoo86fKvhmM2r+oKcoiKSaNNmV45jblJoxmHoUnxc9EJGLYkDfW9T
SftlWXe8YbogtzX9UhiHis5R13++rFJ8uU7Fgh2Prot+Lecn/1+snVru1jslsHy3
pDvBm86tbB2bNTDxXtaBHaW9ZGt6Dygbm5t1SjyO0l0AsTp1uO4e5AQ5pG2OF8mr
fvNODo8E66zM+vvoggACP8Ig3GAbVVoWfLEi4ANDrP9CGricM0uIWkbtDjXndqjd
XO/ixc9iMOa6zVjNxjUiwW+HcOnnvmrHwlvuf5sldj9js3Iy8yqqva1RbIGWSDNx
YBvm7L61fdk5JtVAWcksY0qlSPbYpf0NclMJAijtEQAepe1ukGRBok1eqwzfCNHZ
yENtjRfL+RoAwk4FVLGaeBjSxPjZKUezrmkdY27L//zIvi/A/44gvZ5i6w5oQbxo
eSyLV5PMX0MPuGhPq3XSVb5I60fxS8163K7UTnfmam0/B5yEeSAmxgx85k1A2ExN
zVGmLgDazRg3ktmRSxxbrzxWk9bBN1+AksomDX2LAgqNulurzinfIkxJtewNOVSQ
EICvUJG78t5ZpqNi0eLSbUYR3tY+LYNJGFH8hOf4j1cKrDxNKGOFdnakhvSXN5WK
07Jpiw2kmRj6IJyysiudQBHv69U5uP2sGbYNiWs9+OkBH1EivZTewEu23bPns5My
hJ1V5gH4c54pIiRuaIBto6njQiFooaajdBU19S0kZxBEEvKXKBTGdCZCOStoioEN
ODBmjEsjLUD3FRGNdBp9FBq83Xxyx8oM0eMK0iADzMPZcUQ8yBZqYhDeRlNvX1Gy
qbj28kq7TmIuW7jVriUp4MCx6riQ0n09LIljuKc/uTqgKlW8enxC0A6Gub9mOdEt
efKeEyLQeLl9Xc+NlC7Dobjghu9dmI3Ap9SrE3DrWv6Ph5UcizK6qMCpa+gZmkOB
X1Dmsi95FnAq7pOnpsjVw7g3alR59QXTqvl8fyfKdt0jmoT3xAyPFfPwLoLl3dfk
rIr1Lo8h1M2vFYgFTg+2oSrGjmAoBWgZEur4vYSqRqqi1wEE2YuxQpvJSC3PtPaE
Tvh+p+E8kjBXoS5BfJpTpIWtsrDPAq+S9F0rqKDXK00GwtalzadxJPiMLITprrZ2
yOu/zsJ6P57jdbmZUL0u4Otiwn8YUJtFUgmMCnIobVBY4A0yDxexSmvFpFmXYQR6
HLXMVozz4rOV0iaCY53er53W9QTgNC0+xAmeYX4rk9FRLJhq3RfJKZAR3AvQUo6y
zKcMrpLjP7P1xA0HZhDGM9NxZONVz95YY8Gvds4HfEpi0AzvOcAXdJFI7N5lbd6X
LVRWJcU8f8uzGgu/AZ5qEfJxn4lIRoiROCq9Uxmsitijy6s6qOm9ZcW8j1vTuTMO
q21ppb8ZZOCe3IGH7nrJqytCNyEHu3Lv7z3M66WTV+33uSWnrEcQDguvG8kwtx/s
HhWRP12Z7xSH5uf9aHr2w42ZeYfv8j+spGVQVrUD+Om/t/MfW4AXDFK3n2VNM82M
jRI1FvHJCfynX1OdEGbgZFQgYh0U4wRkfPllTkgdteyRyKDntJZtv9CWGyg+pwf6
12MYmSAgWME6OM9o7rKgFZFezI78AkW8ZT6LyDlxILHKh7E3Z7cVX2OEIhhKR8mE
tYZO/+BAMHmSWah/OfOp23PNpep+COC1XERErJAYE+ssvmfGfCGeEj8CbOaYdAMS
pVz5Z3IQoK41rbf1rxfywO0E88bmuu/y6BL0UeQ2Wl0cd7rnGDn+nzYon10urQo0
vDgdSLxhqQ6QSgwdfYEz3DaKGE68q0tiQyPM7xKEKpNrtlO3alZQQScXG6Ou45uF
ZfsE34hPp5X/Me4Qp9zwuZTbe52QlzBwPQqtpAH8IwaP2JwRJR9R7M26xbusSGlr
F3i4xOfXD+RZt/JFWK1Ss0mApAcxb9Yt1xkXmUNN6hc10lZjke+jZtYlRqAhnpte
jzB3rbHI1AOB3mUufWPUiqFUDAd5SyhEhCOLs1WWRTazdleYRd8Lnxmr6aFE+uqP
3WBEBzNDvUCQnRwYluTWOg==
`protect end_protected