`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
ddtXksX2+yylW5zu6QL2Lhnb2d1sD00763mmSITNX595NcHTEkwn0zB1Dry37fOW
FufOhVzEJp80NC5qZ/+F0Vk7Ik02dIR0elf3clrjeJRK85K4e3Hoo4xn7YbFUIms
l/8VZSb14+JVGURjfswrIyCUotIzlzVYZ6gzoZwDXIi5gQIBf/gI+KxNXPaKV+PQ
Ufys/12rjO6aI/pPlqSm0hCvftmBcnezN2hk1UeXgOIuKZnogjOsf0iJVX2aOOWE
6pD/psybjbnsNB6kH5uFTA5frkzIzkzl5d9+YDm9OyC+k84E83I/7/j+rk4L2dah
QJOvksSIzN867/4Qt8qYTQ==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="MvBXkzurAa5VTw+1JJ70nePUfoQXBvZOku/SMmg4TwQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
oRtzZL4VJ4iwysPsC8SXYCzXS8Fw2gtZTOskLcDV+1B9Nzn1zTyNtlo6lNICRmmK
ZRVu2BmCc2G+fmzynYlNTnSa7C0Cuel6FYpxCBlOuk3OF2tzAmLAuDyOH3Z1Yjzk
a0aHuoCdIRKv7BrZCdALt03JeUmXKPdOmIlkVGFl8yw=
`protect rights_digest_method = "sha256"
`protect end_toolblock="Jn9CQpRhJt4rnzZPRk+dOpzAubz7omckX1MrFd4p81o="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 13376 )
`protect data_block
gD6l00tciPUa6pDNTk/+t1gcgy1iCdpjTkA/bOvU9JA+cpFEv5u/7dp25hHk7lLT
6tYtR8HgwcLXTcx68BnPlzdPHkVIv0lwXo6yhFVkYlDWBcqD9ubowgKij0UjlXmV
p4anbpVt/gKvAYRDYe8Q5F2CQ8AIsxOuOcJ2vhCPchS4QF3n7+oG0MKU5ZyzxTu6
gSvrqDZddbupflT1tnTpo8I4fb6B4/pUU5FFdNnmiv7nC8DihQbpDNGTLK2qlS+E
C+yLYWiYwPpASNRQvG+8VaxN6s53TRm/R9C589BsYdl2VyLILV1uJp/DH51Cr5M+
5+x/f7yUc2UUs8+Gt3itiLu0I3N/wcrGRjN/hLNqPNWzlJxp+u1yaCtPs5Wi/p0R
D7R5EQDvDh99uLgvG4i4wAuN0rKBvj2Y9SDvPrNvX9qDhM/RIqby1z1eKUCDWl0x
zekdq3TTB9ZwKCs7w48yqrOxgxSI6xpxb9yCqfkaR5Nhu0vq+IJIglw03zBFQwK1
1/JF5VsahP6KBle8C6u3LnH2uXvqikzxt0CrBOkZku6MY6Mt+3CrEwqoDW6bpD9Y
4Kw4ZV7CzexiwCHze5rJ8pEv7vZw5UBbLS4ctVTajDy/bRzpXAEKErsXf7FDCYVA
7a+x6VokGz4CQfpf6CkB2QgCV1bU4jUjCvlMP6kQIQw+TONi9OdPER1iHVqbAtRx
riUr73AQdBICIKOoN6RGibiMnkalfVS9sJuCFOaFb4VyrqdEi8sC8xQ8NF9pLFml
jS4aJPFILlWAn65+7jzzeIWv8D9u3W6nFKtntQirnd7UdcdB73cLZIVNuVVU4ZDy
XLTs4hZpwSwFoteziqWMEGHU8HBOmVOv/oRhQ84bFsEbaoAytmlATgaIjykKz6W0
fiMUSzdmmR8iIbjPzvXhM0nZl4/s5F1TOfu1o59ZZPDoxfdoON93bdVKMmi7phnu
Ok6vf/qXOTOvK2via0gVxxeyEUptFomqsHQL9GRNHPLhHZxoj7H6MnASIJhlenCr
KjEVYirfsmKgfPMG4Id43DUak/eRO7N1IZfe+lJlW/wR7MjJqB6bcwiZ/5XjDBXZ
b1jBmw5KNd1/Zk6oV8RzMKuVCsRqLRcAIgIFitsTZ0huYU5DdWdkFGn68af7KetE
OI7GlR6dEyzRlGPfWoFXgrrWu91Vo+djuOR9XYTd9kziZHB80d1/VDcXoSETR38x
Bn6cpjH/uGfKmH5fugvmIwvsYQ601qUQMVA+exaSdWJKgaESSfezOjkz96oaXix/
bgozR+kblsN5pkNZpQW3+hDw1Dfx95I0JQnZLyFm6U/SZfjJUzsgoyidYrLBz3Fk
mjECRItw+l1PyYQFhptgDLOcwUeyIVhJlKPXaop73F+Ff6ukPqvdRmxZ1GHevoK8
gktoYSrpVOr3vVM2YaGXh6mb/ZVAaNfTfhIL6bijvfhLucKbBl6pVt3sri+sv8OX
2DeyjFynk4tHTEQtdc4RAesFOcmYKJiATfmpT6CERfLf724OkdH5nIzb8C+2jmIR
8CVGhe2OwnoUxSVnDd9lbtZa5upFZLLTZLwXRyb87q8eQXBCmi3/QmBvG0lcGfo9
KjGkzUnE16H8PFzWb4Xl++O85GEJCc0WAmgKL38oLAMeQKtF5ln+WejUd3p0zIop
4c3LLipAljNFv1do9cMVymZr0vE8mMKYOQh5BVMOnivRJ2auzXZk+TCCJt6pCmys
CSzDuMojzI4IYKAr5G+nxthwmoTZCrWY/rTsofdk8JeDxDkqPz1PUZ7r/1cOGX1s
lm2vW00CeGRDPRfyvXVyzhpIBBNpZ4/l5KiiPmdYI8D3ZKBMvwXxMdjTidX3s74e
39NTKk2Ou2CygxdAoQMZ7gDUuSrvjuyby0LPVwrDnvR/Y8g7PCmEP4Od/Rw74JZk
hec1t5G9SgZfB91rtfrTYo/V8CXbeMgciHHvdc7a3gUFI+wOhXTN8HQYiy3+Dfla
gbnfTbpWO4Z5VF4gQVHOdLnNej7HIlnBtm6EqfulkBAVCea8a52nUke94oMLcpkN
8jxnNqq8xjH65YuoSZIFCUdemaGmBuBShvCQoR5VvBgGSR+aGJqfaU/1J975vEXi
d1yNrYVh78ujVpmyKRAWScO4DqX2fwlET5R4TEkBeIsliu/kh2UPMkLIuCMLXHmb
Scv7OWu9FxXgpRYBZ30PpsnBwqtpuUyp9ZBWQ0NQ341KRs8t1N1+yy5hcbe0qJ5Q
Z+BzGs1AMsrX2FpYr3Btl5OgqlmWB+uKgm7cZPnqpz2B+cxLWZ8pkhmH7cNsIc8p
V0d7G1CAls8N66L2rTtz6GXNSnMuL3IddWvKVewEOLbfWNCbLonm8t8O+KbAN9wJ
bfTO2uJuCeDiytIzGEEmjZ5CmNqFIabFVZWtiH63FQw9H2lCdhEkj7ssB1CgJN3p
O+9ZYOu+jyV2AilcT9YQH9eKQWdYPhv8zAQNmuMxR92nt0ii7RfMwRyumx3yhhuE
rDTfMI03U9/ME7LjlL6Zvz8v7Y7h1hWc7j7upWCA+ajMdXK05+tItbXC5qGVua/y
sm6OHIfR4UcBDnUlr6aq9tv/QkE+8UhHTurIJO23gF6ecLnbXd1jsMdmyojSVc81
cFS926ailtR1wBbq7kv7DqeyigMga9ckOWwTnQenRK9Fnw6/5IgcZLBUAVMZAp4U
3PLipspeJ/+g+t/3y3WVczEnH3QdYlcxKRPwC+Y/8OmMJH6+cQ1XtE8Ny7Z5uv8f
XEgydp+SibXE/gbr7HHdHfdZy+R7uos6Sz0UtanjC+lfEy/4ZTWIt/z0EiQdKmm7
h7uvmRiMoIeDe4sNjQV/LlSw646gwt5KJiq4EJwwRRq/VChvjPwp2zb3kgUKjlie
Vj6yGrSbvGPKBp2TdRe7tTChWJ9G9ulDZ6LhVhDNXcyZcIQZb+ly9bB96wlfcC6w
AA5MGZtXNLgm55swntfBn3jXgM8lyOy3JIaiGxNQLs2m2Rh0FJOinLvE+CN186TS
hQOznulEuLIqG5CXgqtDSAhieBoUYRXkaj4asCJi3vCnBMfZaddCPlQuM1UKm6LM
pF/MK4TlMYolSPy1sKj9kCEj5W2/4o9fFKj+/0Id8YYufuaYQxGCU9Mh29U117c4
wPp3zxTRf074L7zurA3a6U8JqsfyQFIVC7kXRT94fFluBu+kGprm2Tjyd4X+V94v
L2uOlPC01c2QaDRF4L/OIt0B3OjECqllJqCRpjQN9s8pXBc1UZHuFidb1ojBSLBR
mEbM7BNyR+pGqRHMnhw2gGc1y9X1N+a/hUVq5MkE97EvHRwi7QcP1sPj1tTOezK5
DYdIpwMqmMq1maT+VHZomiBauxvhD2yQy1/N1d6lQAoZ/KXYFTEddi8lrJmW7tqL
NWIg5i7B2G9ztFrrS79TI/5ZXDQiZzcJH02AmWUg+Ed5GlWiSmtpTh85zbSpwIU6
Nsj/KOOG2hh4KQR3CMFMl2WGJiTMrjZLjcjrh0K2yI3xQYnw/pSBbYtSkGdwfsnb
NKxemvsWrBj8DpSHp1AxaFcFjeXmm6FEft8FBcb7DE9MOallPzYepGN7AAzLNUCp
Oug5Px2DQG076GEbwP1hcT+Kzvrt0OzzN3Lc4QCb4dpduvK+sWeSaKwVoq6KVAVk
tURMaprdqPX2Z8+xF6+w3uI9uPGhrdqIBQowmjxts70oaz4koPw+cy1HPqoTeL34
nwRaVjSsTPR2XZabz8Sb6ickuASciDHcZHkpUGuioD6mbJwJ2khhWCsscdINlo+n
S6aHRf6Q1Og3WPkPbcv4ZX7J5B6EfNmT4qXT0NN618dNH9SufzPeZw4UfX07D1Qv
F2DA8Qv/6SYizpPOnM9bDYa95IJ3FuKxedBAqQLM7gVCTrODacDpY2MyQlmKbgX+
JnbWSjrosoAq6s/tX75ps3JVaLpfg5YuUnFSRMCuYsjaa6jV/Flb1JUl7Vno1eBy
DqLqHngyxKic5tuaAOXNMP0dVuvd0N5dB7bfzS3xteFDabSiD/e0nAE8/XBAdaPQ
cmPxZMzeI/JKxz5GIGX4EMLnSkoHtyPP9/LsmKW72TeJ8B5FGNpAREnCnFiwiEp/
/cLEFYUnaiEhTv/l1jXIX7OWGQJv+jzu37DPxn8sXoYmHxG3rFLZzH9scXfwm4UQ
QCR3Uxu2sgUGmkAIkwKju3/0IVuDlu74hcr/tQS7KOQUmmZHTRqRVztySpUZNfDW
jULze6fBZpzEfIFLTG2INsKQkFjKUpcLX2iX5QNZqf05mZtvgiSLG3HkB59bmGV9
2uhvkRpS5GJj4QniYP+htVAXJNJZZYmLcaxLVhaivLqoyZm/svMw5lmbpIo/FUeH
XXW0ylO+RpEH67EoiOvl9ViLHCNftBg5IhZNybNZDXMhgqhhTNUmu9Bp/hGjge8w
iF+O3ydfIdUyOje/KadLwEY7lttLda2TDT73Gkl8CZo0FnaBJPcqlzmzv9kiZEHK
MmHg1JaXGizMAaQSWubWkbFQKbsRDwMp6CV5TfbLyvHu/qeeSfGwz95fFvYW7LNG
alNIGv09vc4Ec0MRsOtONIZMHa8pWAOVu5J5WrYYD1PIz26TIQWieH8MaCmg7t9D
gL9CBmmEf9/KVHv7kQJ2K8QpER39ZkDcK8lRzNBWOXRpsCLhM5SUJkc0eXhVnlCf
M85sgGltXMdGiAcqEELZ4TpnlKocR5Ppjc1hJ/5npKESeEf+sSnXWReOMZcQI8yx
4oSUBXNvDBlvQ+9N/uWZOVHhrijOdOBViMu1aYRP1v2c6ujLeFKtdDzFrHTjQXDL
09wEQVpuNOuRXloLVK6V3+Ins+9pe5rap+jS05Ecgbxf3icZNb0xxP24vQNGzeOG
/LbUMYKDVF8/dsA//GPl8Yu4KstPrJLTxh9Hygu7GLhGulMZGBVsSMV7DUV+9GPU
rIQlylVDfVex7peRoDNNhJBPxFvL3WCJXk2/4nrvx4ZguuHUd5VD+nESnjcnn3/m
0ZCw/PisRCQYfbiujUJMw2Tdn+AAeEM9/V/iwxx6SQy5LgUFwzGcojSGUxfWrztB
vzf5GwOQxn2i2ZfSdSFK4lTNikBa01TYu6KQfBaIDiEkCdHifSx87xuJLhO9GLE3
Fnr3qw/dDWo3u68zRlr2pTPn3Mtk8kFwtBFNaeJu88KDcs3Uq9VZw2UT0gX2nr5R
LhehSO0OsGtnwnr4Ubf/TYYu7iKz320gAaNdhB3apd0VUF7xD/5Ym0jFaUd8aCS4
HWGHCP57agyJId91MtKGBFFOMxFdgjzcMFT6ns4RmcCglpLqhN1vbfcZQu1hla+v
DW25w+QBzZUfdcmnPOQHv7Z4SHac3xRtHDqYnXP3ioWGBzJZUh6mlsSenjGaL+oJ
7JD3MVPqlzYnWaDDcoSqBAR14ihiR3sWFgOlrlpRy8rJjHtdttscSXdmR//uAMFF
q877m6DN9Mj1gT5TJ7/yeKxeWWlTuDiwxTVGpaNYMPiWpTHvVORsZqPA1KCRD8OM
18SDaQ8biJ6sC9R9p2lrI9sKfSQYujFBF6o+vXZ+0ytpZxqgV54nG3XllM8GUe30
iRqXMH6q5bogpe4jWYgxM3H04hTFMlamG3nG+UXXXbh9VtA1krEAoemA8OoSAdoR
f5JE5SfC+wOUBYAke8mcYriGU2UOcmxu30L1XMyWRiucQ66jeimSOKAHnx0SEP3q
K8sd0AmCKDSZDPQvzUCIlER2tpJPnd4Wj6ZEKbalu50+juqMwMB1CNMfgoZ/9vkK
+tNGvRmTIrZhRFsSPMufJptR9yBBmRuJRJCtUPzjIpzT9AN83RxJeCNYFPNEnb/t
dcGsgWpIhWRucEWl2rnUgxfIeWcbWhKBbJQkHWH1LNVyagc2brkQiw+bb0UObCD/
l6xRS2QAfWbjOYDtQ0PnRdBvTSGZpAP8TAxFieV89e0SmhmHU7kYqIr/6NI6pD3n
Iov03m5OtlmsjfElSqzgynogPl8pQhZeOTcY4AoegwhKSxJO1GD2oGo2Py5We+PJ
sA8vAfdzg/2YjqHJoMG7nrfODsRkKeVRLdq9dXvsrL0rLuV7MkYHJ0MOynzho3wH
aeg2oXpaUxVXuIcmeq/HEgZnmmLuVMDxJ5WfGk1wR5MiiVPsGNVT4O19Dnr3TM2G
S+vI9Rwla5YR5NGRU1nJCWXZ7vkkcCximFGlyx+65AmLSPMMuB59uA8wYH+ud1z2
/SbIZf6al/1/uomxmB4EQYHJ7+5e9VvY1fOGVZhc3VFRofQhjPY7DA585y8q6l/M
5iYuEJltZK6wJUqUZbgdtjx6kAVfKgjscnx2cPk6LH8BFBG/lPiCTsj50rgNjZb0
UJ5RBP8H/yCHkyJ167o6tSJPlffZ2GnzGDl8lJrQmmVpnkCxkvIEZsh9RzBzd8l7
MFvHHprSei23dHo92PakNWG/xQNPlT+JhucJUrYSL0PTM/aQyb2ofbmjPnvTGQbe
jpW6nGS1PIE/wykAVW8o6dknn3WjYJ02iUqhswPSaTGH2/UZWf3IN/QeQb3txgqF
r/QvRsbivBcqtV4sCKTlXnwYwrKVWUFTKtEbp4ehaEhssX4fTQLSck2YRMt7ft4B
usNhyZrxG8UFGBj0OAJtoBP+yFXBKaG7KgLIN3Dv/2tH12zLGAiM9kiDAgDH0Dob
3VOC8l0ynbz7XChej9m0mnPN/MzYINqUqqI3Q11epyVOIJS7ySSYZfiaAyTCHyIl
5UMKI3m1nIpJmkPYRKlsZ2OGEVmmxx97e5FaNz2yD96DcHKPuvapBq4wWoeE1FwB
3CZYrPf0YnBfI1l08xUO9El8afM+8oKHAP+VE4Tgv01W1M9MjpF1KFqqbOOPfErP
0kPNTbaIDxrv6Iw843nlgTeE4vnGPMasdIXmmaLHTwINcp8R3UDKEH4ohIvcIxF9
cyGB2bZVOsX+6OWscW4083EB4uto6oNJtQLPnV9ZOUCmAubZ85Q9cPa4htJPWdUO
iO+lRH+LQnqncFY3o6ISCGDJrfzBOnvaOBXEbg1AdADJ0dWR00cBKtgF+m7/Zbr2
ocmv6dQICHSyOc6YXZ4YUJafVQpQheQX3ZHubbwUVZD/T5gYkIBAxjcNi9vTgnC4
xW58KQDQBiXHJC+7/Rc5BdtKKtdE0bplR9QcN9xPpYBGbWfhVofbwhFHUFyAf4zv
IsM/Xuqew30mpQSA1kqCTEAKGDSmy/YNG+OptG0DPgT2JN7xteJDw7G0lCTbD6Vn
Ef2mO01VJDgmjcIoMwx5KfCTtpg/BYFajg7LbK087dXjoemd7pDi3+e9O5332bLc
3gwk89CIKQcZgm7zKgH5g0rU0YNNwEjglqrCPeHZ8reEP0rEomCBijxPb1dE9FWQ
xU+TNxrDrT74qdvIj8FTtm1EjV6wbLYIz2pYn0LQn+yH4eEIKFM1g9yXADGHGFnm
FFXgDU3HiYbjHLLDb8+KMh/lIKGTeljcTPB4FeU7oSOkiEbL59dANjFRKyqCY+yy
D7rZ9Q7p1E7UK7GUJGCNxP+vA3m77ffDYagRq2lzJkE2n6D4JX4aK/6iN7NnMu9t
Ksp2lP+4/SIN4pFlbmdrmOzIadXfCffLEHJ9Fe24g3g0hIsY4K3ZBAabsfxMQep0
ER8ToeBLAe1x1GQtlpZJ7nDHWORCiRQLE0xNx+76HVr1BwQ9AD7ceg75xWEKZfNB
sl6KC0UTnf7ge/sRC7mX9cAPnwIiBzcZ23UToniuzHhwckPPGMyeZlaqiBGZ1734
Z71XVFGwtIZ44QwB5Xev0j9GSjNMaefmuSAszAZjn7AMfpvLtp+GY6iLPsnB1Hb3
7Y5aInKJ1l3NwUO6gvjF2iOSIaAH6EdaPRlfFAd9u8hC+kT+mY3owLdyoK8YtGc2
HHxxap9QBFE6/o0HWtFKImSoSkefMw6dCbR4MMQjC/PiQXhBUyMv+GIRgk1XD/D9
UjzGMsJoOeDCsL5SjQlEPMVrSsLYkNrqFaFXndp2AtBjQShLtlzpzbOK+MxvY1F9
HFAmSF0mQhhRBJR55C+I+EHm5/Xm7WEHvuMZNsbcvZDv5qpiB5z/sdQFbvNGQntu
7Az011Jppf6IoasC9DYmnM/QjbBHoHuldmK5MWkLxJ41fioCD/SR7irjcN0vkuw1
PDAOWbk2ZbsU7GUpTWjTEZXjpIDykrlRPx7Mlk8+8frGdk46q1RadHun2h1z+Hvn
hw1lA//hgYy3r8WXIhOYX0RdKzCqrYwE9nlosngipJ5BpfEMLROWffZJ191IbKOV
LtYypNmYQk1Tm5P5REjURmlICOJWxGiXnqpwC7IyaocvnzqqpwPUXgOhVk+lhFWR
TNBfJkxT3cjBhhTzZ1rkHsdCpcRjneoWKHXvNiYG3W5Fx17bKGlyCQ3M/aODF9Mv
RGYO/9iAbEcPist++l8j0gzvFGrri32W5MyoO16QVmmPMIFVY/w3qJ8nYBHPyITN
l8gez0HI/6IYJ+2UdmKDH9hnb8hl4DuIJThJuYRofVPO1478d+8qoCQ+JIrxBJsY
r5nCdkBR9ug66FO4Nl/bWoSpmnxvOPqXAF+hjdiKUp2MXheyJKdMGzXglcTnRT5T
KRIMwMWgQnbYJF5t5xun3Ue6/++TV//K2fmbiHmzNO5K3sW5XQvn1ywnf15xtF7t
ZUYTjx6e528IhxfRhdPH2N7aimdGEolRSJvTe4saSU5KZhXA8D1ZdwjiiwW+ILO0
a/W2hZWEHUvfNGTbXYSBmhcxAdRliXn5RaYEhBND8/1FaCrnIqdotPkXtEZ2IwXi
bPNHDTemcdaf54oMObCRlitios1FD0nlm7mUmajMaobfv0jwxosjwuhK81dp1wY0
l6wZ+PeYAUgWsVu682lHhiVYg1ifW2R6pKgk/l/K2EnwdiFqPSmuO9VNt/Z+/GAV
k/PTlp42KcuF5BIK1BNQ8ef97ODV5eqbzYHbv8V/8/IzskNydlUaQj149weu2S8T
CNo2d5cWeGBiQE2jUNdauqB8V/jN19bCWUW6Oq1mlTK25/I0wSgZyCtCa3myKTfR
TijDoXaITtX44tq+zFiah6bI3UBcpC/svk/o4LBVtlCbjndrCDU84DwxbXYXKgmN
8SmcYKeqV9PNBoVfj0xQjW/G7PtqnHMCsw6oRENoCRB8+AEj+eNselojaKq0JIN4
62bF65ioMC/Bub96qL8pip/CmlVYjvn/CRBcZ1PCEDGsMQntZ5Mg7RJGAs6G44m8
ak81e+g0QCRgf5MtWulkEd6oidkudNru5Yv0AWzyGdrEzVIqWpR0OW0e5VRd4Sd9
T9VxvugbZ89Ww/I6AiIWiXPMQtzlmC7ZHkArqI3yJbOV5RJiRPGxZV4UGzY0VuyC
F0IoYAe5eC1SNOsyLl3IbJE5AlckK5qAEtClCQdf+K44f5JCaYwRT0PJXFKR7o6M
TCYVYz+4jR9MkWtxgjYSf/MBh1d50rDFAqwvu+7NjayzeWR2FTcgD+DA8qx7LkZs
N3QWcWo4uEvQsmOqF2PBA4O6eLOh4KJQhXmdXStJ5jkfiJ9u02Ne3j1RUlqKj704
Ll5tVdS19ZtmjxFbYC2VNr646ZEu+xXyo5q08yPzyadhQ72geYGqIn+wWK8qHenD
9z5cFUcqlukJJJMD0TXHQ9AyMsXMx1Tah7w8R1yRpOr//J8YZSJpO1fzf0ntu2uH
wVuDo2lvokXXkzJbjNnrQaZI1XLIlwPourAbb0BTN7iUGLnNbTgoH9USkjjREWsD
BSQiuLz5bg2E1ezGJFPdQVWeplGDFq2vOQrOfCgVPCSZubdSDzHkNHHjZbw9Hyq3
mDVdzYxSv+heBmGPMJtl50yKq0fsAg7sO3vkrZtkz3fvRYBR3m8uQg9s2nMDjVZ1
GFGSMxCN6pbK1+QiuqRAWzp2e1X7R7Fep+Py5z4LPbq4UojMjuCMDihUlX14BQ4m
1FHZsj7yVvdQFeTJeG3LVfCiap45JJ/tpcCja02grbnx3os3l5w3ANEpAu2G0m+0
RW/aw2pK0K6//m6JXJerw4XzgJvyGkVJgEtWI8rGw5bxYTk6HuTXHqRkcmHUanI3
F6Iy/gxfw0XnAmBfF162fsU3bwxPoFi44Df6v3Bn4pFDCjIiBoYsM5jZ1T77ZXZR
IthdgZ0mf+6lzjABBVDlAhysJyw3STiDTwxmc/VD5/tLj/0peX0Hjb6I9TJjGzZL
BKtRXKfD8OhjXBzY6E9wD7mq5KJ5cggebLT25drl13d3BEyWyrnFKqPk1YqYj6pP
IH3cmPOFoOFUBAltelkTlL8OwPPLLhdnB8N4ShcI1R3YCpvz4O+3tDcigXoHcqVY
Mmzdt+aBr/3hLl321NZqpkrvPpEtc0LB1HYAzENRyvvsmFczD3c82wVIgokuP5m7
yRg0viMmbXJuzZohEICye1e24PtSx/UqZJ2YiJroCbMXsnZzh5Kxj2OfPnaxUo+x
0g6Qb/jsKiebIczvE+GOePhEC/2RF4qMm0FRdUdMmYsMew2ht/aVJo4y423Y0kcz
896/lk2m2amhSEsL8EdrFOUptOWh6pvbfguSeXyYrj6UeakkTtvhn3iXzhOf741s
VErhy/tlL2rx8LeTCe+mxF31Hwf8IWx7HxR5JfKiHkqeEwoP1ggReFLMtRHarrqX
N3YPYarZUe1ohwg4uvLjT1qOyha1vs1PkhXb4zYQBvPT/6jYY4smA5wKWulBi0J2
fEKrbvshw+B5dphvQv2dZOGGsA94twl9r73ANap4WOdE6q5Q1q/KOymjPhkDOhpv
9m/eymAzlbG4j6Qg6+XHp66yWnzABFAYrwkFXLZfHfc+dDAZqZizhuc8zmbTLY4e
hxJaGvmgGo79LsztK9jlPRVQZ/xy6YS1u+kCF4xjh+0liqgkUIvJzNSsWCgcJuvS
97XsSGrMWZHKytl/HgK9/4RLAbbBOFylvBCgWPx1hL1sGNK4lZO8SXvNPzWJ/1LB
TLYzBov0JmNLYk6Xivg3fkiiGqDTcBhWoS56UAeg3PXMpgMeq5m4GgD9bMtjSmQv
3ekF5FQ8kQOrhBoNf6FnQdBCZW5MT4ryysO9Beg21h39v477VGGRU8dbhVWpWnc4
uV+popZYQYS3O3j6EVn3BYRAry353xj5zo2H8AisFAb72mUbKKSz4M5bv5PxRg7G
2AHcsSyUBPrupzX0Dc/qdVb6i7pLb1jVSSyiGRW2nk0LtCowy/oHoE/vhsfXZCAs
hOhsuVSz7keFYyqX2jskN1d8iUXODHazG+1bBpgZcyuiL+NzuFE376/GqGw6vfwP
UFVQL46a/6O6mWdyaH5uh/jBEB7iS/MCWgbs2YR1QQ/D0bkYtTBA6EEnnR+jkvm9
7c3Y4i7ReuzuGptMt41zVxmAbDBcfZdz7SYa40OzGeBtCsbs8Ql7kLMseGabnCMV
tvSQelp7u9zQTgR950y5ORkCJ9JeO1yKO52gHLIYLr0J+oh97fk5MEj0HWO5oHE8
LEVs1TKvymDsowveaVTnf+nROj+tS1gj70Ttiu3aUD9yjAV7yQkjhBzFyshAWZJ/
o2fDf9ELGdTkPUE2OaA/YPP+ffO+a4Io8fbwPUr7OMZCGXnGx/mrtV0gKeAFITWZ
yvmSd7o+Roq3MEKL27APzdA0wQ6LDFKJDxouEAOaZb/wj370967Q92aTZj8JcuEN
c4bcmMshYQnhX/wr4/2q6h+ZGFBqKSMnCfxGCaPyivIUGPdApBtJRvrtjgDixvOV
fQc/+ngFkc7tuH2UIaO663x16xhMJU6C6Ru8+oCzhET4wCsV7JUGFmlT/apu1XdQ
833aAPjFVrhLTFmzP9SWiZXkeJakJif9+NAw7WGU0+rW/2/qIrF6bohuJ8dzlSvd
B/gZxe3nHH+39MR5v293Y0xketitgod6LPb8t1FZhvTjGUEMSyVKbzm4ujmj/n9i
RKw+CZBMmcJ5A01BPoreYwK95T89fqf47h01C29AmdyyadcBqdKbxnJnAuGR1zCz
ZA3mdq4ikjjJlLYh5aqQTW55aNqUWYgoFIa8EvF/aTI6431+w2S6Wpnq8gNwVq38
8tUSyVJ2+4OB5s+foAwEbZeQObW1n5ipqpHadratCNxg+pxdXe/yN+ZrPa6TAt8f
jWb9Dv3SCgHlCU+RCbusBIopVs4hN0BKVHJMNhrmzbYiE0j21I2qPqtI1jpJL7vO
mit+mZ8p7FGTbS7FyAL8NZY4nEGi2ok1BbtTgis1MHDdxqinL3np/nSW687PPFsa
xgFOZOj5HTp8Tx8rD59YMKF4C0gOpdG6uU/DXPl6sAkjburCJxY7VV1RAosHkXku
5mSvMscwsiK0wkviFnbv0ZO6OG9HMjedbZY2MsNxueBcp75yYWhA6aqf5UBnG9QF
HcR8uJ/Ri4YhKwOf2wv2R1trEYTVpn6pljPHBDV+5RvJ2a9gh3BAt4F3QFf5XMQx
SeVekVDr38yDUvWUfsYGYzdKAzTTGikHA5O3VX2Eds1Xfvz83ju6k3QbaKFJSqZo
CspJdneX/4+WujenC4rQN32crCjCW9C2eQSj5DuaQ+IAQWJIIH0TaAgzGCuxzcUY
SwKxEggCXyQLNmTIYfQc1Er5F+ZLSJmbvw9fy2DnOdJMJPJSmTo0vWHk+VXE5h4b
eAlIGpy3sPRoegVDmNyId6SPg6bPeiM68p9ZhswLckbX03eS1vIB581/lVt/S/J0
rifvKbROvA9yUBIBTUk78Fbx8xEtaie5yuNM3wYjUInbFYIumCv0U+rXa9V1GbVz
vJ1O/PEAMJC5j7VayEk0aQ6DopqQcCPi/GBHEADtqwBzCurrtuJ2Oadydlf9/VdL
AlavbCDIggwMNyExsDs4H2sXaWvnQFhAdpg0i1aK6AlGoCse6HLBMzYjE6KSwXHf
lJQTeKSfXwfATfkDXwbaEChJm38uUyCHB0ZsXbiPuCr/6tr8uIZ43/RVPKrIy0Fl
q+pb3tClqpkm3pbdiUszoBce+O1vq969mmptZ485WP/S9SWUOAREs3F5RGLWeiSQ
FA1NYqokaLN4nWRC5VjNSUYbSYOQTwiiXwStAB4MYfufnbwGnd0BtUY17wWZ+ZFd
UgHo3cRF2Swl7oTths4YknN44xz+WrZBjpTVye3TMDNq3b8fJzufX27+xji68tkT
jb49OdRqV/jMC3PaATiaPbUcqHwIuymJmWZd46zr7UJOnleCd98w/dasE0BRKsVv
isF1lZ+kwwfHLC2zrehOpMVLLss5TJ6xWi46x4mphQHCEty8SHy0NYw/4hoLtSgz
YAP/wq9Bw+EYviu54eiuLfc8hqa9jsIIiQ9Q4+Oi56tBm8MOLzbiWLqv0LOpkFLq
Ugg0nIKNZIiSOyhrikV7w0F1AVgvJvfGwzWYwScj21SqnUWBiQxe82uVnAUY2q0b
Kn6Si1MG0Fk4ba7plzdiRpnBxwMIDdj1vN95u34y9cW5YOdYsbQv9ur7d4mfLaP3
7eRkQ0Feo4T2hN+QP7mOV7B/0dzVoQznhCcmj+Oce2TGlFzBnArWmddXrvheG5x8
brQXYPkb1TA/8/s4LqprmZBowAXvrRgo1XUbAlzMXSCE3DZBeZvRttV78vtYnJ2s
ZpMrJTe46TMELHh/N22+Amed6oQRSj8Y0OaGB0xdXIfnA7u1PWhM71FyMcfxwmfo
VBlzUa5rfSfP/R3BUgWfBBce1aJhBqQ2JUBEgHIah/ZT1dRhIpfVnWWHUJ8YpE6k
BN5XEssuQtUEzu0SuCbZKNAbh3S0UHc10ZWZuItKxShYClKewQJiA6E5Opfq758r
O8rdt7i6bFGKdVJXR1ZydLx9Eb0yb06UMcqreVdbb2J7rRZCxDt1b+SfLT9ehb6c
4xtIcnN+dmeNsfn8TFYSFmoggXdyB92j1EMc7u3tGS8PP6vnzjjh0DuTy45XTPc2
2Vve2irMvAaGr4/ww+hF1NMHo0aW+5wB16NLMYI1g1S0dxZ+64QPT+xSwV4N/rxF
bmj/4zg8eG1QOXiA81AdJyUBSmezqVN2xlBmMC/9TVvxlK4ZCzArxeQ7yrEJdKQB
fkabcByFU2v0HbTNmPC9qDsFFbUn1kcYQ6KKLD7rf5AnfMZs0o5cuIUfHkOJioYA
o69p4yB+E2MImqRCBPWmVf9aV1lfJWF5x0Jvbn+g0uEHncco49nIbcUf84EsJYbD
zGpqdpVdpk97f9BxjkGdqseY7vLJNhn02CwQoZQY4KBbDDoLR6uxfaN7dgdfHSzk
Ec17Gk77wSs0iUFwfGu82nz1bKAd+VCierHp6jCvgRaVR10W4em7m8oPhkcp6A4t
bUQpcPwAvlWXXVTz7Yvn3gkfevyoRRbt2UXV7IL9+t91NK7ROouml+ZUIEbbdudm
YsdUEtfHj4sJSMBvmbNeJ2ob6DOrven5nGvOqJIBr4DptMt1vzM2wO/+lwclMJd8
9b7+kVlUCeMX3hBbkqXhkXtTncBarVI/CUw23+wycOXBUFZ++C2eKkGwJDFV/uQS
aKP90vEWr1CJacyoc1X1ieVDRE3n9GbVzce/rfRDa50DnmxPtMaFiyK5RW8FRRI3
GyaXIJoqopeJuEyivTcE6voMJT4TyBVbMQaxpV3gfQkef+8xramGiHbGf19sSSs8
DzzUv2L144v9lZuTFpv30HvB0R4k9UmyFSsZ3+CRCx84zaT/tHNpqlSdXS01/oPB
T2kr9xPr9bvyTTxNek/hL9X1JlxyShc24PYplqs/hh5LBs/MN4p1tQgUDeQQqWoh
xLs89lmx0VxthP7I23wdwjgsqIUmh1tQhWooAHMtTCoT/I0Y8/9ur2PtZ5p7DBs/
+e6ommH1OV160f4XAWd/or/05WGM134GpH3k3DvSMLp51h0fvn/dkEbdgfSrys0T
TNARP1LtPCa1Omw9JWkwREAbZ9fwXH0fWbBpm0IANvmFjD+ODNoKRaVCgE4CVeSL
ayMp8ZKuFDVVNFWgZx0ecBHWLvjuqzfPIaHzfnAO4p6Mp2WZm/mkdPWsoroJNF73
dnN888iMjSkP9rJdkz5R4toHLHtQt5QZ4/QijbCUyXGiNA8d8w+7Qr8y8j7Is/16
9b6Da1rBSvm6AKocdzukm/5eWV+dLWTVcSujLJEDglS5PKmx/oYRrRLKtubB5Y6K
gSKeM0JetiPPID6dYwckZG07D164mq+cPiRcu1URrspn9WpdlGGkk6jPvYflHKZN
S7WarrKSaYncV07yBg1r5tDDNwzq4V/EbZ7yG2tNn05YPuMz10GfR+3KjRBQEgkT
4n6ZKLibVwYmdY4vgmUOu+pNBIq+eSWUlVaDbKrXzlHSY9rVBKwpeHrlPOwh3A9b
4K+spyXYUL2U6SlTGENBexEHS5L/tv9ZvVT5PoZ5WvMeteYypiQdRknmtM6pj3P1
kQD8Xubw0drrrjnqNIm6Kos158UxbTTUbeVRh/Jl7obbGtRdeXU4U7ODydHHOxNi
kxzBpdDEidzlUx1fTg6oqlWYHOLcQ3lOHFcYZjIfBGMxuKJ/jObLiY0jNSTOtZO7
o2QZXZq/EdBjdGSoiRq9ZBAEHYgxeLKqkpVXQx6FiorPzXrk/RgvUrkR6uYW47MA
+OX4LB1oKgwPXolK0muXPcrsf0rMGVRISpXFFyWNO9qPqkHOXGpmyGYG1n8vOgvg
Dl6ermqlgFPJPHgKLrC/q0kIh42J4RC+H8UzbdiJydjIJ83qrClRUeBFcrT8k/qX
KxTe5g8jONOy854BAIuM8LaCkDVTRm6zFliOuVA4DqwsvOVOOdDZABQXWkbyl7ow
J0EhI07/wfbk+uDuXY60ABO8UpL9Dg8yjrLUe6wlFcKGka/3reUmyOMhBMBeRxU0
eSIFpAaDdPJQrcBxfV7ouJ2REXBzopnKAoXeMEbm4Vrx83/ZNoub9VtnxVr6gDfL
T37FGndaXR08e4apuHG74+1Nj5t5jnULPAy3h1SOAqB0k5lV5zZSGM0lfiuTnT2B
H4teZeQiHanweffBijqDSeqjZ7JZ/rnhAimm5eke6fNWfEYuLgZXgnGSj4hv5MrR
9ringNuJNQi10K/ZrIs82mg4SF94uTjTVgQM4LZP6Ye0XADBAyjOu7nUNd+6YKpO
TDIK1JeVlSsIuxAixhUaaXaVDiElqUttu5Pu9xj8MJzYtiuiHLD2pJU1FHfANyXD
jbbTGnOJmZWmmnHnSoRvPPrNN3ODrY9bK2N72as0EHWb9+UkmOdRf7bxxUSlPbnI
Diawcy7bXj2zUEGRTbam5sK4+CzSeQfQ4fZOMFW/HX6fih4b3zg0F8Q891B53eCm
z5C7nxWoi6RUVJH5PT/Vc3S5kd2PQ3S2HzHChzR/EUMTR3KDbzH4W3LtClxeiCXL
hSVAPRtuWHGgX9eODWlcLykpNKQTRuxBpmPjDdvO25rQa/jzrdDo5lsZPumbTKPC
YCXYYIjDIRFNjBCvAS6uAcpqz3FVICLnYXHWoNBGx1EfY92bVksO9srWnM+JzwIE
LVb41hns0OBJ+E8psuz0oaAQ/EpUlGwhWeJoCo8izyEAP+3xYsURr6OolzpV+P7g
ipVXIgEu0oHcHoy5in/biyXgbAaO5xmUB2IMOnOEeb41N52tH5NvN17WRVvELlPq
ilMan9s8eKbKwJykcPPr48Yf4VOY/OTSkFwa4Fa0YG0KacvZmmJ2rmsWMyKmyT3D
u5+5EGbIMnpYeTJ99YuzZ11phlPHBkzROPQyYz3Lfe0i0Jvl5VFGjw7ZNwmRjnSM
2d9ba4IO82A5KFWes8kHn+Xsk6TMCdAn4nhUNMgV2PGX0WWG+UvQf4B/lDT/9m3F
7ZWe3EvVJKEf+71Vv1ieM5kL98uEmCjnlhXWyZZzyxXePs1DaOmyUX3UxCdxvOGj
ST34QSaGGXQ71Bse0aEsQl/Tf8BENxDTzewvhIOXMTOFZh/G+kcvn84cq7WSmqey
fVndCq8NGxOqNzOIyHLFzbP3cTyIzhpVChui03h38Gr0g9GPI1cG9wDpu/YPrWH4
+iBtouTQ77jjuHeZ+c7IjyN0J5za6q+Z/RchdC1ZOU2LuSX0i1UiLtrs7yqsB+rp
k5h4ejXbLb8lAFXscFBtWOj3prOuvHQDMJ7YJQj49NWBYYucAVTqFJlFgZCsihUO
WObkyWRJBSF6W6fwpUMCxNV8wYcX1HKK8yCnOgC5v5o81AjsEjC2jzPzRgYLTEv1
FRSE4DspZex1mFmSaIMotSnj+qurZ7+k7yNF3psbGVaN/s4T9np69ECWtV9ps7YD
v9vi2w/0jpJrtolGHrzFMo4JwnlZ5j2Eyr3mrLf9QV7fT4VP3L5ZIr71TzGeNvGM
BO1uAL06AarMpUzfvjHbhpGNofOQltX0A2IrpxtTc0ac8V3Rmol4tmAWK1KlYWi6
qx+WUasFwbV5ENsbBDl2e51XtK0b1gbZJSnf5g10JM4Q2Ojj3kolgJV0NvmahKmO
YNc3bm+Gxh/fX7mek1e5IWM10Byc00BTc8CGuBxFHDAhz+lPQ9NWoNMSY8dUIUje
eLSlZ9L8xLcxNYXuiGEZsNmXVdp3afNOJ+RI0924v08zG0QYAyvrvAZk+jsUoicI
llCnQyLJa98LH8fGrLNqqoOjOlv8UOUGRJ/x8THzUm8iWqLYByx7o9roRcAZXpkt
XC8FMkgEzijlm1K3lIe3PLqIFeaq8zHRcASuk2rOUpa1l340VZIecG8ZKkBAJAfW
ImKBsDLfmK9w7u/or65jnmNeckppVEW/mvKeg52GClA7PcLeX5f5c/6A4ikM0PGy
8nIuy/3Auooz+s+uYfNDIXPGFUyzdttoA3cdKwvmRJ3ouvARodAftX3babFSQi0d
MAg6J8eyS3uHM7FwHcNjAM08sdHR2T9Vl4sWBMJfWsw=
`protect end_protected