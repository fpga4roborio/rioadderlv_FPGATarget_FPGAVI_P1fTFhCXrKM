`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
ddtXksX2+yylW5zu6QL2Lhnb2d1sD00763mmSITNX595NcHTEkwn0zB1Dry37fOW
FufOhVzEJp80NC5qZ/+F0Vk7Ik02dIR0elf3clrjeJRK85K4e3Hoo4xn7YbFUIms
l/8VZSb14+JVGURjfswrIyCUotIzlzVYZ6gzoZwDXIi5gQIBf/gI+KxNXPaKV+PQ
Ufys/12rjO6aI/pPlqSm0hCvftmBcnezN2hk1UeXgOIuKZnogjOsf0iJVX2aOOWE
6pD/psybjbnsNB6kH5uFTA5frkzIzkzl5d9+YDm9OyC+k84E83I/7/j+rk4L2dah
QJOvksSIzN867/4Qt8qYTQ==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="MvBXkzurAa5VTw+1JJ70nePUfoQXBvZOku/SMmg4TwQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
oRtzZL4VJ4iwysPsC8SXYCzXS8Fw2gtZTOskLcDV+1B9Nzn1zTyNtlo6lNICRmmK
ZRVu2BmCc2G+fmzynYlNTnSa7C0Cuel6FYpxCBlOuk3OF2tzAmLAuDyOH3Z1Yjzk
a0aHuoCdIRKv7BrZCdALt03JeUmXKPdOmIlkVGFl8yw=
`protect rights_digest_method = "sha256"
`protect end_toolblock="Jn9CQpRhJt4rnzZPRk+dOpzAubz7omckX1MrFd4p81o="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 3872 )
`protect data_block
gD6l00tciPUa6pDNTk/+tzLxvdHE2s3DQL3/JqqujQBC/Ei+vcAB8wM3doqg5vTg
mdfn9XB1bLOis2CVSfu295W2DNwHfMSTc/8BhCDRnTlLIX0UCJs9Za0+LoM0rMrV
T7EjVWppbP+Em6PkVKCwlmIQ7JKaifJ+Y+kjw9HCGboYo5074hY+K/CBbfsBQY86
AyoN0MKhsIx+eViNgnWjA/InyoSYoaQnvM/tIPtai2rOw/U+wWHG3gc6+NXRiBTK
9qXQOmlKl6Wu7yNyL0n73ONyFW+qrE9iYh/98o84rTdk+oNUzBqcysvi6Yx1m5wD
gm59ma20j3v+QkIwitPzVeJ1AGFekBBu3lMCVLyoaoMI9nRrvjZ7BN0rizTzH43E
hO3DwU+oTHECBwE5f3kNr81e8LZ6EWNZ/hblJbSBBVdHhnpjnJE2hkiG1e2kQlU+
soTBSWxYr9vpcBESxJlVpwhIatqk41dhQpysM+LAmTtsZ5h9ZnUYmmEWQtJtkDej
6OB55c+1MaI3TAmSCK/z9O/eYv4dDWADYdnL+pih1smPF31n0JjP4CWOL5flxvcZ
pLYei6OsCMKZqqVMn1H5uhuYDMHmFEvGau4riR8AZhCkV++nMBzHvnoxuvgd9ecI
MlMyX8xsG2jCopNeuCrNxOxcFhn0jJw31ewW7u139foLZxASpMW7kOboUC6kESZU
/Zok70ZUq7URKL2Th62cmTdQKs7VeW9jdFRRaKMcXpIOGdaQMFEBjogOQtF5EuZK
FmB2AfbQ5gG+eTOO9tjVVtrOpvjn8FQwbeKZLmoFj7d5T3ezOTHgsDtLil+kpX/7
0EeEhNiPBPNQ6cK3aKzYCmweXltNDKQaRtnHB1ixmcXmp3gPpBJBKpyfipHxmI/p
20SeRgl5Scyrw4bKz6t0c0GvDx90IRuDMqfoveJkGHPVutfpUIGXFe7s14M9AZPl
QVXKXXtJMWgye4SWi5Rppp3RIipRhkXjKJoMarRamhX355HBdamRWB+3wTTf2n8r
8eXZ7dFFKLJy0Tyh4Dk/euQ7JYamWmDeyV/TrXafIg6Eu/jobwjNzUn6qlE8fWaS
CcsAPe9J+p/pX4Y/FECyfzWH8k/cmt6jU/MQyWSwGKeXLG3t4aEUQGRowII3p9Rp
sYrdxKgrkKyyyWEoeLZKmeMh/e3c5naY2O/VL3Z/45aLANzBT4E6K7BqIwyeHaBx
rJwoORZLwGg3J5p4Aa9jXOtltBv1zXwZgTuj+Q8k4rF6qXyvAC0kq7Ql94ReDBce
ndrHRu/6MaSL2SbK0AzBz3iMdwMUqs2yVK5Slek2G+LieFtbY87wJeuLMA/gt/xS
h8gZ7h2PqNwEnLqy8Q3KgjC0BZ7bMNqIH9+1w8m26A7BmS0HVxqOOHDKCJ+yoFJ9
bzXG4gm4z30Wpkbcn9x+fk1EW2DsSb0s+QUdRDR0joo5XhhP7u11ug/L71EFNxNh
geqd3IGNZB8Pdxe4DbrmvOosmMoifrsILb4r5V+z8dCd3Dz7kOoP9dLXlsq4a1k0
p96e/kwQKwM50hoOJ1fzJy+zazyPz/7laZv8F+FihKNIcdM9NrJLxSQV8RbUz7u7
Y7iB4OGjyystXYZuhEE2Hv4A848QXcqBs/jPR1IqamkTWgZYor2x89uLTqJ6xI7b
WnTL3T1+JRc55bzLN2dKrY5yX5NpY96Yy0BqcukTmZ3XbCbgmlhqicyh8vDzRYIR
3htsOH5nFqvpeT39NtSIv4pC4Rbz4fu3qVQqD6v0CLpPsaTSFKqqb65A9IGhqB/Q
bQ+Qn4XKXQj71kkX6d3A38fdYO3G6gAhEGiAa0m+gHbRq9e/rdel2B0Jqmw/f1m6
kkNA7aAp3wjNmkWCiGRivxEfcPjpzOVJl0UOVkSi0hGmI2QAadjQGDEKMjg7JgqF
cgdrGn/wf8RfKGVwi738CnXPuKhM99Xxt0O+B0uRASvU81fy/Ry8PR2hna3mna0j
e/cJgAb+m+c6OjtEGCq0IRavTVxAZH00ohFvSAqvH9n9fb3YpVfy/R8VRVFVZo8m
Tl+d4fWJXdcrcORtSJ7Agg709Q3/pnL7mQTXff6x+mozncC3rUmrmMuUh2vUbSb+
y1XU3Zf5A9BPQP72+x6s43Ok100DbVbfVsLDu2wtclRnF2C1zij0kPUu1IWMOFkQ
kX+y3K0W6UZ513Nb11RgrvdnIapsI0/azhkwsxmQsa3ctpllPEbqdRQ6rYKsPA4V
QR7Ag8V3UMWwlMkhltb8cwzN6ehgOQkScSQOuG1JyHBsR2zZPJBavJ37j2mx1ohb
7piywtc3T1F8tWg/xVg8OdqUDHemCZ7nmEZyljcVTjHx+3HOu4toJ1qqVPaDrljq
xjtjlJOnwG42Z/s5RRL2yf1ojWHtPdMb68zJlhQsa3PhK2d8z+Z9gW7m+OSV4MOu
mHvdKONxpNr4ZsoO1YDs1+zgEYm8IhFa7NBuuC7xtMvqaDE2lmTs+DP9rnJtEJes
1VEqIwoEUHvPaA7uAFXPJEsh3hz9Pcyk8LJP1oAd1dsUgNg0wEcMr5/Qt8OdK8qW
PQBNg0D1mQRssmoH5Tj4GrdjW1I43hHQvK5eePq5PBx4/jN41Yo1WTy501V6/sRJ
x+bSCBzvXyHsBa36hxpMFw4cizqiyeKp10g7hOnBZr9hkuIrs7pfiC+gmPzIdCXh
7jApHeBPiTPTpLliJ6nAPrYJWfB/S0dlYsE8Wx/rV2wpAdeaJDOYKDB/gol3P35o
VBs2d1sK/XRMdV73waOwqSWStks49zmlkeyfC08/UO0UatDStf1s1aLwdWKxUy8/
Jx4RRw2neFOH1Jz7UrTeyaOqp46jEfME16oMd3F2G6S6uU0hs6Ckiwz25xoq3mFG
5VlEYeBYnKLTEC4MzaerIqMILPgbhtLB+jtYUuXXkn/qC+//oJwc//8cFXbHJ+9u
+cdkMWdH7SQeHYaYITkJovRToIvh50/ySJylOX9CNwuLSrkH1e0g82DAtmx8e8kp
qWd9YHvJ/lEQ/JO+BD8zl+mCEzhC3Vc2wMOBYKsy5sIlynzDexGUSVmz0rTFG9TA
kz+oC9Jhy1I66Hg3HiL1uF56J3EP5KzMN5RYYOJg7kFKjK0fknVLkRoF3C3vfdpz
Cw7K6VU57pNzutcpxeKwTxXw5jCUpGJjSMJ33Jm19bK8nMJYOxrSZE5Yq/0lBFM5
l42ottX9CPzuSM01pGWNXywMVovd3Qox3GZW2SF+BPWkhHw8gzYfe3fIJu3fX6k+
N0++ROAFguAtxtB9L74qTVp2qg3JDaZoAcawxPCs08Nlr1ss2R2zu961HzlTAWkZ
LvmFz8U3/AqXGF0KojQ7qWS7SopVPzmYZhFh+VH6fdvnBSCl0Ye56cVBpYRXp5NU
be5a2MC2vHAw3xwOYwybVrjdCdnLF7tJNQCCVF7uL6L9GjBo3N1eMz8NW2dFcrA+
jcb9xOUUEypINEbJLkAL2Br3ARboSK500JFkR48LFA9UuzN4P5z/BJDkYbocTKoD
j6ODaHOHr4ALZ9jSOojedtw8poR44NvNsvUhXpoKMPzQdOPPnojM1c9TBaguEGKx
DXjDtgdnxLShEDN69Iv1KtUYPpIV3LnJ5Rzwfz+tsqxU+4aP7KPIsTDvh2VZkjHz
7XSoBNFalFSzaPQ8I44EUzFfbB3SBVFI19oIc38+CzPPknBiB3n7FI6f/aL70cYd
+d2huPpmSJPBjSjT8jIX3vkzf6ptBtlBfQTXd5DJ1iF1/+0wFueB8GEVrs78B9k0
wpqk5AWG7s5zwSoIh/vbbbM1Hk/7LfgCSPP3SHJb0KAHDcLb7+kjmOa79f+RAdSJ
34hg0IUqbphaANuk4tmYTXoV0tJgWs7i6+rzHnqtARXA0+8A+dIDyZAL02VowOSc
ZtM9VlNHdmq6dwzZ3ZamoE6XQF0JJgaOIFP/3Q46UVBmQT7OcFfcMvUiZr/0FMEG
3xD2yMUQO/zfA+8vhh+WObzCS09kpOekaH7B/05fdccQ6UDLMhaMujUi8GqmIiuf
RHRinlnvWjJp/E/fZSnqXj+aDyO2TjlbZjmHMuWkr9PYjXTAznW89WNCEWdAfJ4c
9BIKAyaPc9EuoBA0+gHnkCdDebgghFpcS0Hxl6pgnH0D9Em4W6d4x4zxZOXYdJE2
al+T752BdJOZkm+RQnhaALesM5VY0zI3bwfCPvDJICBQWDKqUlbH7xPbRRpPfmn/
Gs4m1d1dseHJ/Hdsn6UxO77kLsRImZLktwWHmLFeHGCsN2nTZmQgO8C+bY4aGAfx
IxM1ug2MdcMvaiHfvFXhw/dRXQZSQ4n9J7n87/kqbG1rx3teUsM0VX5GPrMzvfEM
h4y3MSgkue/XkkW2qXFhERerBWGfZQVlJu8j0Zg2EM2au4MU1BGkKga4sXLEgMy/
ryz2nKBCztXkZ9h30jQ9Za4j/tT6w0IE/y1pZ1vLLibgrWIkCsqOurH0OdmmagKN
bno/C6eDqU+1u3b5xKtB38l9XsTAvmmoLyt/E33a5SF5WZlRMSumYxETfbZxXGeA
TvkO+DN0Lh4Bx1UEF3WPJNHaLwitfvb5EWwvobFmS0SeSmxaqgeJwQrote9jZpus
KYfkjxvdlIIlw2CnNfuEIpVCuXuNjI3b/KSR5qcUObTDa+sHZPCIHgAOFzcCnG7A
P/pZAmxI0tu34nCBFH7H8AtMgsgTdhNtS04ZyVcJ+12Os+90G9pUy0eMIHccyz0W
ZyJ/u5qFzR5iXLwRjAwF/nOGvlzgAmewwnhscx8QXdwQfTfjCbA2FJ0LezGjQCSk
y9w4qCBhfhSY1dbT+45vyjNLu8/oZY7eAS2yMarAJTnG3/IBYIPdp/bNgr61ojNa
mAU1XMVNSO/QLaTYFcu8yHmouAgU11Tg1x/A6wyJjUmw1yAzzujCOIIqeHPHJrwD
Pq3sLvHjCJ/JPnogfsTjJl5rtPAAlFfTgp0VItNHUlbXwCKYbg7EsR3wq40snToS
M74Laotctcm8SqJpfGTUr7fD+I8tNd9kr0HliaUONHwQmRbvbfUk0RM5H/Z0XdnM
zX9VnfeCSRD2N6JRIUASs3qLyaRQKU9Hc223JcDDUEjDvgl14O1ZsBzuhVZXqXPP
0PUeteqMPHxkejIVVusukJ8H6Bmz+OXf7hZeD8fO17E=
`protect end_protected