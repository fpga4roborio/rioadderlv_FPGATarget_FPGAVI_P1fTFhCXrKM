`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
ddtXksX2+yylW5zu6QL2Lhnb2d1sD00763mmSITNX595NcHTEkwn0zB1Dry37fOW
FufOhVzEJp80NC5qZ/+F0Vk7Ik02dIR0elf3clrjeJRK85K4e3Hoo4xn7YbFUIms
l/8VZSb14+JVGURjfswrIyCUotIzlzVYZ6gzoZwDXIi5gQIBf/gI+KxNXPaKV+PQ
Ufys/12rjO6aI/pPlqSm0hCvftmBcnezN2hk1UeXgOIuKZnogjOsf0iJVX2aOOWE
6pD/psybjbnsNB6kH5uFTA5frkzIzkzl5d9+YDm9OyC+k84E83I/7/j+rk4L2dah
QJOvksSIzN867/4Qt8qYTQ==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="MvBXkzurAa5VTw+1JJ70nePUfoQXBvZOku/SMmg4TwQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
oRtzZL4VJ4iwysPsC8SXYCzXS8Fw2gtZTOskLcDV+1B9Nzn1zTyNtlo6lNICRmmK
ZRVu2BmCc2G+fmzynYlNTnSa7C0Cuel6FYpxCBlOuk3OF2tzAmLAuDyOH3Z1Yjzk
a0aHuoCdIRKv7BrZCdALt03JeUmXKPdOmIlkVGFl8yw=
`protect rights_digest_method = "sha256"
`protect end_toolblock="Jn9CQpRhJt4rnzZPRk+dOpzAubz7omckX1MrFd4p81o="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 9072 )
`protect data_block
gD6l00tciPUa6pDNTk/+t1gcgy1iCdpjTkA/bOvU9JA+cpFEv5u/7dp25hHk7lLT
6tYtR8HgwcLXTcx68BnPlzdPHkVIv0lwXo6yhFVkYlDWBcqD9ubowgKij0UjlXmV
p4anbpVt/gKvAYRDYe8Q5F2CQ8AIsxOuOcJ2vhCPchS4QF3n7+oG0MKU5ZyzxTu6
UFh2tOZ1UkjsCcDisYgJ0gTt9OZ6ss+TZh0Qz7aGPb7pLPY4i3hNjZlQjDZdjmNz
NrTcQam58xUqbtxkACL0H0tWrMqljIYj3f5m0V9vyRgjouWRPULNPwwLzzK+FD0H
mZOrrmrNzpLjnYU0QtGwD+l5rdK/dRwxPvluSrIMlviixBfCLHgBHoK66Aejdvxh
h57gxaT2UTcho02jUgQB8u5bIpkbnHwQwfW6LbKVdxTZ7V0Ek9J6ixmknXBRXanq
xXI5WFYkdoOzS7R4PcFUU5R15l0aOEKbe0Bf7kQEDxyd30DP+iA858wc3ljFiaxl
Cx5CivqbKgt7zgLxC8nqHJYqyjPQHfm24V0ZsUG0r0R4TdAzXPxAmX5KMInJdYHk
do31FDjcDLWGFRoOcsEhljUewyNW/shK5suJP+D9an0BTyAZmXJyPKScuC/4hEBC
r146dEiZwgO0xr2xEQLq9/IpZPnmFsBcUjq7L1zu+LE0eHDzF7TxEVuIoy31VA3A
aqpq7/Da/pvFUhfnVVVyARdevgLLI7ykuh97Vc2z3alJFnZPGdzJguF9unj7cpaj
z+LnSsoBPAiQUMooiMP7SJmTuw7ZcSDvArPmAFN3bkQ2pRScde8V5DljJoa+Sm69
mIYnyVYiUYTp0cvQPKCttwkYQ0kMEe+32cVWIqWkFTzCcSeMHyzsCe/tX3IQSXts
id+Qg0HfCTsyId+V2e7i8VooJSO0G8TlvXebc6x7mpl4CFm7qugXBGhWj4xZJBax
jRakJc/0/4L9XYYjIsPcD6VdEGC281XSF8befY12HLbeihrNx/CEt3NK1myqgPwx
VvoBSy7TapAIjZOguYnhzOFUoH30S4SOSS4xQcb5trtsaHnfapz8/aszuIrcIc7N
+lf1aHUIvMMIv64uzOqOwdfdANouD6cGtEAhAmARgEj9i/0HEUWXFg3LqA9triSy
b1MxVT/DKmKJVsKtT895pvUK5BTfkH0z/jrezgBM73BjNMIAV/FPlgJxpQdUmPZP
oXzfQDt3LrcgnYEwSZxcduNZxsLRe7U6oIPx9gUYJPxUNzhGwndu1eKvButj80aF
1uh09xO+mRQxGwBfir+UtZL0/JJMZ/tC1XlKzZ4OR3QtC2AWym4PVe154IHeHzJw
HF1r6DD7IrQYVB33pO4rd68aqc5Fui9cSPP+CQSTukt/8W1fx8zRgmAEMT2VHn1n
EFh8+ypPs8KyLpWysXTg5MfvXgD3H2bItNFQlbLhTL47gwwknPFUcxUTydWDIewP
Yt/fjsTXRRB6huzW5/CSYUDcJtKZAwSpvlEXhrQfz8C6deyTj9O21cwz0nXVToYN
Bn+GDZO0xL1TMl+rKbB9II8S2Kll5beS1o7hNh2QfEtA2Dw6v5Bz3hyaQ/xu6dHH
dKSUpx46TFOri8akKYVtTsMPn8gKWu7ZHt3McVppbkGUkPnd/bXsVcFc+WmyJzVD
Uqq3M0uLiLkUroR0QCQ5hAB5mRJskt4YIVVytlu4D8aUbP+3tdd88H0suCVBuGNA
chgruJUMITBqx6T8174OpdHZUceOXk5WuDcgIcZzU6S3dj/b0Uya0xH6cbQ0XZOB
ILUCDPzmHt+70xmctil7xvZA7no6gTNSEjOZ1JTuTA3itWv5luaSOyw6BOGJPxPo
4yEmbzjPDNAGIE7FZYitokEsZTtBZZIhaICdZeo55wA+2ioYP90GhR9W5j6colSy
VhCDIjz8CNSKXAt/zwwsAMVeqC1/9bmgZDNF9goyJxqzZGaNfEUhC42SbEjizqSo
4eyASD8lkFqy8I9S+a86UeFToLGVuzIAkHpDBBGFI5Go+L1jm+1Y2JoyYXNBguv8
pxpPZQEcKquQ3b5oUE0NcktAmKVFaiMc8fDVTZAW6WICM9pFt2iAMaAfLEk4uD+l
Ege1XvDB1HEbREklQyqd+vXfgyRmrbU7T0+BB7ofzzxUq9maTv0S2aUKDf97bJZB
A5SiKIF6DML1CYSLJ8PgDqEapizrKiDdovqqihlg+lH2n/NV8mkvEGb/OsJ9GGDx
CWK2pt8l/aaFwVwHudnmx6XCezbpWEjtKhCHS/FTlODirIjMWDAgWC79IQIkKHj2
T8xi5NQbzu72UxWf5PqD4yNW4m2GIAvOxZXIFEHOI5KjOhS0l5/MumHyUkstpnUa
xhUg2jgSpd5JLWuqridaFPEiFHDm2iTwM7Y0u01NbjgOPYMRCpXNXXlxGwfhuPVX
jXrIiT4dmP4s5DBWM80VA1E1Sbxjn5rnrER7rZO5lTTxOgod/MfMCEbj94KcAieA
iD3JrAWH40GqDGNwN3TMq91GBiQtwysohV7vxr+fWFPqg1ldyhUSIAyWFL1rY5G5
/9lhx3zLZMyEFy7EUudk3pqan2CGuBK6Cm6MbOaXNeRSlA94G+Nu+cvhY2rOXIjq
9/vQOIuDQFzfw0cpCuNIhIvX6XPFSrV3u0CtdcjuXZEXUg/mz2H9hueltNTFfWyl
qJQ3emrFbfk6XLLjUIUayEYpwfwacJh0GPhKu67DtUwouLm9CB4uTV7LUdNw13DV
7J+0AHSjwGYWuNrv+stzPPKTQv7AnBfRyNDejsWggx2GgfyMs4696JD+uBluoHkH
21O8X6KTUYDrAWxJGXplDOU5zWWyrUb3q0t6jMWXiXusJUvOFBN6qzSHu5Il9zAU
QAcuE5Vh02NAIPOlbdn2iugbVkiouYvcHLPcVglZuskhBCnqOvRgTYdIZNuirkYI
N+qtCE9njZazogJXEyuQPoiwCA1PTdqFroaI/G9ilYrTdvfUIt5vAoSSsG4tWEAA
XryPCGmb2TS2azeEdqCsd1/DcG3FoaGMRzdtx/++nlxKl7GN7l+1KPeFIBg3qdJr
h/6vNRrZ6rAfIEhr08+6gd0aooNVCYndjJBZSPffu7rHc8rVMaFdpPi4jcLgoYe8
vx4BOPx9R+HtNLfi93WFpPYdmB6Txdn3OE+1RTu0+qmmP+XZceO+zPEyBVeBbrL3
bUzA1pDO4Fr7C64PQlHSiTtNkW5lF8wDbRjegJrExjBroBO2HS+PUHSM0dB7i1wU
UPDNCccCkOHlFT+yBO4YozN5VNMjRBoxaMXigM8peYNC08jAI5wOxQI3kmq8cWEi
qlLy7uSDgxUoH5dmj4nhkSHOfn9wT+i09Ud/VI1H35/5RzCD/EH49c7V2lkF99G+
EsWlNGv3A50qp0nxdZMe2u3FVBDD2mDCZV2exHCFs6JFM9QXzfX9SLtJR/u25rjC
OAvTHgvr6oeGD9BjBdlNZ/cYkCyGgA7wnRgU5OJ55gyjdMoWg4gjArltWcE/NGP4
Dpo5s+uVhjwePKFG3vsRQVSf5h8z1daTAZOkBWg2HrTSia/XWH5xb5T3TaMBnAlX
m/LHfm62E2YegRQVV2KVmxlxmUEQUrWk1HTFbvJOOMmrvZu246z2q7EXbePVUmLC
PuMzMhs1AOhhAi8ehnTFJNNgaQcRgemPtzE6VrGl0YODizHUOkwhX/pxxaWxRPzB
BXqjd29mYwGx/kCCSCErrrJlVigyRg7eEHunGOiHd79w4k3qx6b43GRrrBSs+sWL
p5f1+PNSJkTFx2XJjvC/fdXYL57HeZTdb/n1Dx8RGliA4iGgtgXA0x525g2dPRh2
xMLUqwrPt8wWcR5VgVW9w3IlqQx2CqfSzbFuaCZYJpa2r5fSIgV24+jXhGP76Owr
nUuyA+VML+/kHJc5CMKNSwK1p/8jmvVPKSy6T9qQT8GkJS4Es/XE1NcLaHMO+8UM
cNpQa8b3+MIIkEN/kMsTqsh6xz+ojpkwZW2HAb2l111x7V3e24CyHMzU0F2XiHoe
XpL/bPSbB7vgLKaPam6D5jp1dj0Qoi3VqeygJKZUoGVOEhVLvCca6oIp7AtilmA2
9XmSICrV4wIYGjAD4tgPUr5QfrEsDJO4uH26voj2SA2hYG70xq+Y/V1tp+WnQ3ok
VGQo1BtjFZh5nLtjywi3V+jNhabqUT9td/Lwp/cMhOPGWxT4M9uGkTQPO1JZLKym
CRgmWNt+XjbLC1rbXCly/HI02OtKX351hNCwVuXbSbIIHBJlUcaZZHhr6WKMib6g
RivqfDk/j7FeunmCVv6C+kvciZ1Glel1tDBZPa2f4KFNkXDj2FRKgiqwO093m9qp
KQ+0i4cVsAfE2Au1rqvwiu0d9T3ZxQ03MaV/COTrITB8GRw8rTQ5DGty507pK1lb
hIYx4vnFOZJl3qGyzVi7JUTkN/gFm9kVfP4CgyGzNffw/vBkdKdP/yJTr4TtsPBm
3RAdzcwUP3cKEyDohrsl6yVx6W/rEUvqHfje6lW/XRmbj5GOC9e1JDiXlNJs8IDD
K8s3gy5kUT4P/tRAPa+nJqhPlaXM5PIeicuoY+zHmYRvesobQBsm+FSslhctJbEp
bo1lSUOL4aQjoy/gKph8wOCg8rgtQanY7WmZVBXLBJAfxGmnpxDA3IeWys/Kd7nZ
qF2KcZ1VGA40ud5/c3XFMiVbdvYZ4knzxXmon6wB73SQK9VgB0wTjFTb+9GrsmRy
0nsOlJ1Rt1QDZkJpmHoeabNIV/rSzkRVon7e9aaFBUjkdWXQtmIC/a8XiEx7a7lw
nQAPavfY/iXkXzW4HuunPeXjiAyTlmjgrLywZ0RiO17n+41Zp/R5lbhqJFdDJo3o
WoMhjOnUiTrKFtlBSCC8vm5aR7Pi1P2uWRzZ9t5o+FQ1+uIYWigp2TggG1qIJ67v
Z5YAfSop9Rv8UziO1p7VDKQHVQmlbeEdE9Uin8FOD+4HDpkUXt0WPzyj3kmz7hf5
kuJq/gECjyhcwuQk1iS/TswA9bEiFNX/wJE5jWpGJPBC5DwE3k276bpug23UWXAW
iJW63GwT2yPmEdDXtFoQa0Hw9TmIbsvDgZCtNgZw2IxQfmFwWGt/LryBjxkDRPLb
hmobU2h0oaD24+P8S9FxQ8NzrGOdlq/6SPprnWUMjDPGLmoVwKYLOSh3LWZYhoow
GtOTupCnqZr+x5VvlLmNFp9PvtwC55z2Afxjo+ZsKkMga5E3h8d0s1Lj041LcHPL
uAbiHWbbcx5cn4ud6Le+fk5NoUCPMLQGFYZA16bFoi8BBUAtIgQQYPa7ZaV7jQZO
U8MkfDCp7JliibvImUAAgZv4lynjV5jRtM3KXQ6Dt+i4OE1os/5S5vuVkbJaBhnj
yKxXGezVeUeAHXRtp5+2ch21lBBLtjhCuBOJqrERv5+sRLbv+hkbnWt3tQ0zsXC3
XAGxItxIlAONEe0OTzfCceMfsb09Qy2svnnp9jk/MLltBkNOgfCj05zZBFm0UPlJ
SOcl5PdG5MQ8EWLKnf3s9ynuANEJlP76uVhH+NpgUhUG6lUth9pgbSaQ0k8sHMi2
nAvykkpe4xK6kQFpLUNr5yss64i/AdYhW5+V+FoXmLxVPRm1vpAIlK26W0T3q2mP
fXPBD+ONJbJ7WYBb+OQAV6ZJhkAjLR4Y7MmR2sXcOFAnTOfjkfSVY6kC29MkXoiO
yxtNDf6FdjIRAkXP3+pUOsS3hgPhysP+rTrHaWUMg+K5UngtUUc0wQ+Qf21560sA
ENhqYm2ld1BZSfJ7eTCHERcFxPFEUHCIEFcXG0i4XpE1dwGx51MS/5GrVvhic390
bAebgKNtZ0T4/2MrFcwbbbH5yJ9OGNywuOVixdY7LaH/O9rIVlXd6ztUwmJWYCDd
WVp+qJOzrVnGzfsbejaSJ6ypS7NaH3ruEd3lFJb5SegY/U6AyyWUpVvSLs7d9zyw
zFMWkWVnzrspreqFyX5T69FlZszS9ln2RbZKOvvTwOo1bdZt2CPVggmLeK4JDwAu
lj2xQiMDgrpWNaw350nGPudjdwZR/LY8xYoPT48YLPH80REKh/UnsSSh64ork+g7
Vk0TY1/Tr8ZLhwMr+C1o563vVdCXPuepcy/VzFN0fTOYACyd+S0UE9U2F+nTtwAB
TSScLoS0Z+Qaq222QUYd6sd0vW/JF1DWHyZn92YSntsTFh0Y8mdyYMe5w5qkuy3m
Lz0x/lVDmLSE5Giglg6UaH8rgya9N4oCgPrLX7BQdF0WPFD750oFHmZk13CJEBxb
rZjxMOnYHhG2wRdsxHnbFF9aUEuAsKJOTD7E1hjZ/edOjT19SVlrDiDPZUuNAdj8
xLFSQlAo+Yl3r6YQiUEaLhP2EBYsLgiSlcpk5+SSloskOSAcnHY+0SDCvPfmrxi3
kmlluFqJ2WAtMiSWUdMalgDEFbC7Lh4u+3fyx9R4lPNIYlaL0mfT9Y0ARcp3QxgA
MSu/DFhKGkUqS5RhhW4RNSt63K1HYZWon/OCe3eELST+lVb5c0wvARnG4zz2Szl6
iQ9bvIK1QGO6y3yCZT7DWqyPmvx7z9QnBo2bV6H5Gjn95ggJZFihRHcnKkjnEEkw
P9JcOoJUEN9YvKpZe8Qnmz3UWQ4fZVt8kvn/cgu/lAj9cTL7vxU/yO8SGrsqsmoo
PIADpc7F9wGKM9bdcl7lWyvAkw1MHCm4B0GFogzVMlT5n9xA4G2t7CiVVoW1Er7i
1/BvJBekcKv7ZFaOGX9xHFgqBxjaWhA2j7b+FsYYWMe6Pu9+MjTS1ZODrU1/Qq6M
woxMhDu3sdCmOykqQWZ9RKXhE8mpHEz82qyEoTDWV9mIVaGolApISApWZHvqdl/A
Fz38ktnlRHlO5N92xX193vwcAD3F3UIBstiEecUMC7cBtYsN4wMnZv0I/YAscytM
C0z8XueDbsgxYPmxQ/RMOSKXos79j6I7tJjgkY7LTihXFAil8W5T5jKuUcCg1md/
K3O0oBrJlKABaSaxhGXyvdusS9wNZ/F7cNHpOAhbwa9tg0D5uqdImF2n8vGVldtL
mrb8xWFspzD0kxgNa5y8f2dQ9LPX2ZNLkwQuzZ4MdxPPQ2/PYNP2ZDEaGqOy+td8
YlhL81gTFjiSCJhXlBvjUFOBreqFzS7+a198l0nDow9OIWTGArteLU37sT9a2UKZ
ftkWHnrOCDH89gT20uwPc1zio8fFaXOfMPA31Qxjyq8llj8X57NU7N8tIPhHNxqT
oBQMqoqfXOTgfD2RMGNGgjpBol1HxL0J607ScqKdvhjUyds4xS/0d599XYQvfFLs
ei0u6oDRE+Iz5tfq0zPd6YYu4uYJdPC85mFOR4w9EqINc3Vqzgu9osOUxS+NmAKl
bPz96CEjYgQuboyRgAG182QgTEIjI+7UUVM7HxbotUYVY7jM2SL4lOvXhQnJUyRw
qFkQZL2VMIwUgVvMEs8mEBCWlnCVUAnkDAadsIrDK4hNJzlpb47ajpDGzceMjN0/
/vzGY0W2GAI2dJMDmsMo0tbxve761x7VcuhdJbx62F2FApv1pom/fS/ROj6q3znR
kbbK+wJX4Xd0HbwF/V51iBY8NaOk1habnCm/0x9ub+QbZ9jgIgPVleBA6884+AnL
jfUZJwfnZ7GnfIZTdwbnmdGr+OjlTgBvBRfvxX4vrHTW3WZf1t0IuPvd7U7o2nVn
IrsxzfXeObUMo6k7s3b5FKhNG5opH+k+LPSQB2HF/m9nPlhZFblL5My2/IfnWH/w
kr9VhOK76M8fsgmmDKxnOWG9zGoYO1wNFeOHfGowARx+RZDCXL8idjpOPFXRgEaY
KfUUyWgkOKqvvnjtB9AB0mC06/lULIOQzQVhUrbydhDn3wr0+uHbZ15sHnl6LDqq
y5EYJ8vUF6mhZ6YNZdW1eqpeWnXtBgE3WSIT6YG9wZFDG/faYoVF8JGSuVjn5T6b
K9d+8f8D07+9MdDgpdbvDDTyx2tnW7AUviIn/UL9TFsxdZEhsYNVoxDJXGNP1wTx
GtHofD3arIPqbDaTGTJmMWTUt0Jt8PBAuJ1bUGEw9D8BjUj1y2nTSVvtfu3m/KCC
4u/cTNu4s4Yageei+4zFLzma9m1Nlap+CUkEzH6zpeorfk29g8f4/PSjfnRWr9la
4V1PUZpISU/I82wH07YAG4Yk4dOZ8y4g4sHJW1FmWK4x1KZKPq0fkK4huDNlH8b8
9phMb/ODvZZXdkAeJGvXhTHALKIM9CvtyRQSrNFbdPtF20efr0W/GIwzwO7PU5Hb
S/sCQZNQA0VvREpSh5HcIzBoVrARfJorxGAxxiuGIkNcDqSTIO6OHVye2K/WoXEM
PWuxkKKhRyJuSe4/eFV9l7qizmnGsTncdXRzjA92nAk1gMWkL8NlYkIXila8M7TW
KaVZdHFENd0+9PsnCGTxXn8EuVOSIyxUDzku9qMC2OEzduVOdUAvPdj6i8Yy6yDb
G4EcYLd3AwFKDVrvvbiQ+HbMYOpTt2O8RnOUWUTxAGWTw1SdqUUsNhV/i2O+RAio
l8ZKgZUR167A0mq51LWfcocRtxN+Pc6V5i/iBrq7snONxC/NVkiCXvwWI3xs2ThM
B065QqmzsLRFD5N6t3xru+Rwm8Bo/hfHs4vA4WWCTLzySsJs64ph9h9xP8Y3JJ/j
VsKFPFfNSEKM86VbLQ+DmNslSnkigq8VcZdbwq5KNpidf/0pbd0PkPHoYWSmkYz7
uuURe2eVSf8GVUyO6CS5pXxzTuHu7bgB0XaPcQUQq5DStS5LJRIQvvtksH7o7QW1
DyYfRh3ZPylZ/m9pfCADCNgyj8VMrwuy5ICr+EHV77nHZhrqVf2ZVgkmPWCOh+IM
6325fxD7M4NFyF9xzekCPvLMAY+/GKES7OrzCklCisYxDUiGeIOT6yZrE7lTRrzn
JpshS/N9BwbnI6PDjwh1nsM51cCbyUCU69Y74rut9LU5b420p3tq8q0jFh+L7n01
zavtvSrRBbE6qrlB7E2Fvyi6yEvu3hNM0ngkyeVfBOh9MeWXVW+cB656ozuBzYTC
8dpkrkmQUvj6FSSPD9/P6o68lnhqWGaYErLkygoX/t2ehebALWEK6yoadaNDNpTt
YNS9jYJR4eIAPLmWh3TYR1s4qTjvvRQ8hjektzFoNbfm2TF5kDOAQRzgke8bkR0/
PXMluRBpFw2B2qf/VhEXR4zn5w2K1FzACK6hhqb/NACObjwor6Oif8c0RVQOwxLP
EBGu1UVxn22KF7pVoLztwauqBu0N7oQ8oiu5pUuApF09m9aRcL0gWKbriM+wd/yM
Q+6okgXqu8TLFDVGksS+Qps+LYHcf1joUVvtQIcCPmSLCU5BIGfuQReZTBYpB+NG
PjKBovN93vqgxOw+rpnRFOadalmEDDoDeZy3jjJCByYVPbJ54+c+7t3FH9PFpR20
jDwqPD5Bol82CehAsrsITZLu4i+X92p9NclidkAUys7+P6mbk13h9iAEJNMUirLo
KaThFsaU3e18Bg5msl3alDfEfuKMunXN+qjxF8jPT60UcktQCIwWcw1z+QVlE9OY
y3WVQjiCISItMk3K0dPLir8pKn9VOe4clW9/iiHunJVa4ItzH508T5h9TM8f8Cy5
aXjSIYMJd1UFuGuz75tCR+qNO74i6PRlaCpHdRwcgeBf1JL252GN5syPiOLIS8gy
25UJok+9xaoqdvCEpCkJSI4MzkxG3jp4eBBA09X8YCbSZm8LQBGaPd8NhW+X1F7l
XRU81MUp7Zxmc9g3q3QiFjvt/jNd1g7zCEMLHTT3zvqYoI2hCF2G/4ME1hZTwOy4
7zcgsya6JfMVZI4eGGvqhSgWpIUBrhVn2Kx6P9wTLzDHDtMHEX+TQtRIQSkGkgrg
HdYTD/EJ+60brOZQwmpuxxvnxk1Cwldv3rFzjyQaMsVAGN5JaKcKUOeLWgKxVvIf
xrzBi1twK+Ua3w2cb4X9HAlKkrFYoPYBEJV6NlnrV6uUfe5xYoDo1+4BhwzNtqX5
CyWDghGIhOu7dv2mPMpigvjSiAYLwFtmHfwpZPiMC1V4I+xfzcWgKwekxuJnBTQ6
4HGzGed/aR/Ryay6qr6tjUvP/TWXWSNY1gU/LSQCMNn7ZaFijFtpfLxAj4gznOMc
ztqBgRWjwh2SGAuNW6V9ta3FsghaQj8KNvIDVDfQnto3UsIbCP/PFZY0VOc8+gSx
p83RGxF2Vt+N7vlC8IBpX/axMZJgCO7uFcphpcObkBeyoFT6NXNsjLr37AYmTyLg
kRwycQU6IKBYItrltnromwUhC19W3b91O+iZSpWL3vGHL9Gz3QYCL54FFmzeq6Xn
D3gQQDF+rsBNU0Mvx3D3j/ZyI/bLa2bxPzIFLiWHuyn8Tz19QqmrOyT9OXyQp2jI
8WTJ8git1BkTCUa9HJRb7H8OlvTWvsl9GNWmhHQ/YD8pq0kUfEkTU0PiXvUhjQ8C
CUI3L26E5oE/2kS0UCgkeYnY+Yqy+yArFameG0Tcmpe3gS+xHlUhavOyq0aVlRfv
y/j/M01o8ABp+wNXLlJEPNBHXBzzuUBUo1B73kQXu76SK+9anWwGGiCScmV0kqoU
ougL4FG2d49bTX+nRzKbPw6RkVnA2SrAU2ep+8NoQt3ByzWRgbcPvhQlM1FYRSFi
U/C0qycQ9gIZKKTBBm0h++rNZadITsGsmMWE2vlChw8fz6ZPP45PggLXR4abtS4s
uTlNlG6/H83gc6Ho59bbiVc1KTKXYKfrITl2nBKyBQEgnTFU2AU+G0MiJ3vKT2/0
FxNVsV3YqrPI7ZezEPf3M96c2i2jIckDzIO5mo7mJom91pw03ei6dtSn1YwMWnSF
WuCLphEl2NdJOooSdwnDbRAt/ZKBb0LuRjKysccFvIUMx4mDLTuTmoewvAukyHbC
nO0j3992TbIG7qmKuI2Ik7UDTolEZQv0oWNM3yN0zSVXu8dfWYMEpaWHBL1rDYJO
wC4Li243aY0DssXiRSvhsIAFlIO4HXFEwUlb2fkkfe7UoHWMfjlSPLb+B4AnLwtI
8WeVICUy3nVt02SW37Kc8e23BOE2eFpoa/wbNcobQEqbRRD6E8JwkT4jU8BUqn9c
d8PzVxivNMYAS3dQA09ysuF7bm7EOji2x46rGOQfDGovhejeCRRAxF2A9sJW9ULO
vPlyB4eRyXjAKQwpe7/uXZNkur1bYe1/sdvKdPMBnahBmRx9EluvNms6SH98mGeA
v+vE7GntC2W6hqgtr3XyqP1NurlIQ4OoKFsRBywypFDD99UdIy8ccY2zX4Qr6v0H
KIk2+ymnL6s5RDurGkUY9BCwXrbGcIZNNFid1zv1Gtt2JVjJp25r432d9TgZUqoT
JO5cDGHs249mb0XaFczKIGabY9xCKqzAJf69NscYa8cnI6IFvRIOYYAEap25hbSS
UIT1quGNDZCp9LQqdWZ7m70J4OE5vTRAZENLWBYOPet4z+Twa1qqc+tbF7FRlGiH
cenSAKkZJc3hlwInlY4BcV+fCbQCzkdUfiRRfrFzjrjuvXYtVp3sRaRRWRdpFnYk
mOLVIAYs7y+t5yejJwn0i3ruv4hjEtni6pyTQsm31Dl5WqLUe973m7r2W9wg029u
az7UxUG3tikuk2pcrtkvxFzz4m7JtvoqksRggtVDYZh900ZCD793ozLkENW0WD4e
xwZimWh7jBE1/5TykKBOeJujhi8bLF0MncZ7lrzYcyYz5+2w3tphVi7ZQUoyJuCw
TZZ1iOXzlpmu0TpV5TkBPcANf0qdB32YLQsIhf1xAydr64B5Nq8tFxxWpYWw0pBs
mLSLAgDQ+t0T1A5mYVUviqAkLjHvpdNodB2PLZMb6o/8uq6KFVQe/YBgUgZAUXXF
eVFz/uPJIPWR27X8iGRctgr4L4/LKLx6Yiyszj9dtvJhfyr2NbNKQtiVABJJVlkk
//FxQDxqUOM5rA1SQs9EnYBaraVvNxeeZfwVlQFv1MkAYkJkmDrD7l2j2cHb23yj
2KaXjJn3KAN/3xGH11grWKTPaZS5ttvFrGadVmWyQhSncwW3gmpjgOHlxeNMZ4mG
2Yn9oe3sFnkliB4bpknMQYCIzwmFx0WEJzZmk9AhpqLJlHfndiTenWom1FMbHG8v
`protect end_protected