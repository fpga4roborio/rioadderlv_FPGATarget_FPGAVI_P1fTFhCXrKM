`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
ddtXksX2+yylW5zu6QL2Lhnb2d1sD00763mmSITNX595NcHTEkwn0zB1Dry37fOW
FufOhVzEJp80NC5qZ/+F0Vk7Ik02dIR0elf3clrjeJRK85K4e3Hoo4xn7YbFUIms
l/8VZSb14+JVGURjfswrIyCUotIzlzVYZ6gzoZwDXIi5gQIBf/gI+KxNXPaKV+PQ
Ufys/12rjO6aI/pPlqSm0hCvftmBcnezN2hk1UeXgOIuKZnogjOsf0iJVX2aOOWE
6pD/psybjbnsNB6kH5uFTA5frkzIzkzl5d9+YDm9OyC+k84E83I/7/j+rk4L2dah
QJOvksSIzN867/4Qt8qYTQ==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="MvBXkzurAa5VTw+1JJ70nePUfoQXBvZOku/SMmg4TwQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
oRtzZL4VJ4iwysPsC8SXYCzXS8Fw2gtZTOskLcDV+1B9Nzn1zTyNtlo6lNICRmmK
ZRVu2BmCc2G+fmzynYlNTnSa7C0Cuel6FYpxCBlOuk3OF2tzAmLAuDyOH3Z1Yjzk
a0aHuoCdIRKv7BrZCdALt03JeUmXKPdOmIlkVGFl8yw=
`protect rights_digest_method = "sha256"
`protect end_toolblock="Jn9CQpRhJt4rnzZPRk+dOpzAubz7omckX1MrFd4p81o="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 5168 )
`protect data_block
gD6l00tciPUa6pDNTk/+t0OO0nC/UTtBwLB41d4inuAUA3i/ALrNyoJVcBnAmEQW
ptbcNp5fxEUJjnOxnedyZEuEBxWRieZFQnkRdF269oPGHH3Aq51C2Dw03gymO2U4
nEffB4Jcr1OI2BsoJtoztumlCcLLSssZmJ2otKWDIs92oNZQWDhryN2FqAP6Gp2E
fH5gKAAcsEosTFMSj4Iz+1pBUwxUI/FsREb+e7tfd4nOhP8xiM6XrTZO95SN3Jf+
5xmgNiUcuzvtJp05/yIW6Vd7s53xYAl/Rr/TlmrlFeitcbYnNp7aZ65/QhRFt7g5
RrzTNA944P6BcL/7BIYG+ucw+Kw67YKZqwwtVmnOrRiQncpE8TLcruGTDiETCHrB
2UtETMAEAwcITqtddu048V1hKwcvrqSSuFyeZdaazYg2kQytYNJI/P6y9I6wH1KL
BdNC0t/igU+9aCxIk8aoK11Nnhv4aW5w7Grsh+lh4Kn6eKydc0wuSMhUstkjSnc3
nBlpYWptWWIqMY3yov21Fqdl/uL7XnNsOnOSpUkktlZFwo6Zbs0a+TkOESGI7Xsp
fNFdbYBe1/MUE0Se5GG/Saipp5Am+p4EpHQ9khRFfURyR5zGSjpHhH5HkkZ3NmJv
ZR9As4p/7cAVgW4HWuNdNiSpBLpbe4Qhfggsoa3/PDjS+eqlOEKYu3zEG6Dyki38
aluyZ8USgTCJalrj0VQy0F3n9WJbfpSIkihRYU1yDsVdLydiEZXHDA86lR9Y9/6L
GuXmQ9fXB1z1Xpzg5NZdoIvZmEsjn3MfWP7rJASvFKrAonf+ffXRi1Trs2GY8VTd
XYVn6bIXA4wvmh9xX919KF7AajiqZIJ+vyRyBQlirNZlCcan16LarBXBuqpegMTW
YTR60RQX9xHom5iNI0/GZ37otEMD423R8Fy1DWltY44hcy4PoUoJnOAvtLaO27Pb
YgNYfXgL0nnrOfi2dvsNEhzhEKWYYLNYeKsHeabty8dSgOq8E1G0i0I1DYdVktL5
97MIg8xxX1gMh+EQ90eZiUBGMd96ND1T9iiY2TxVS8YH6ORU89DOOLKqnvbDFR7E
elXQ5uX4z2xVlowWTaiq4J2uBrAsAZSOZeQz34GXO7Ioq5/xkZr5x+CrSH9hUH2A
DnmB0DXoQR8uJCk/SdHJf5k8lhx20b8vsOjCZ4Fz4bx47vumqJyxXTZ8UIWMr9GQ
v/pStTlBvJrxEsYZh5QV5n6IDh0Up8tQ4XClO/+ZUETyJJOiVi3ITWZxaGjsx+cq
UeSnXi1ehx7/buhvy5Oe7D5f9HMXBY0W1Ytm9bineJufsEC2O1inbiK+C2ZlgJFr
5zxErJ2t8VAwk1azBCRGvh9W7BPUrHQfcS3sXxNAhEVLkeEVa2Z6eNSYwwOGcfSx
1Aquh2/tpUiJ5F8NgpxLo9LBCWCTKgKLCFijQWkkvUTs0ehD9oojba8dRRkSpMj9
LndmgMCgblazA3D5kekQ5a9JazhX8sOY51rURjIaUaZoYxPOoZq7+L0UQw4QCRR8
0t/TO7E1/DqFYmQoNIQAg8EfsW3+rAsttRwgKeL/U4HcaBLDJ+0sKe6gSvNbS7Gd
XlK3n5HvYloGQsfZbNhGIhaX1l2/ag6OpJYlqNWazs6joa4bfP7T1ynHafi3Zvgf
oYYjxSQ289uGExdmCZswlh9nUTtEKoGtbr+cr3kbheQcRnG2yYbVRswpcAHQj6Zf
gTPV6RZATdVE9mXI9R7NF4osIyf0X5R0VKmpSg5bYJvtkjdvpt99WPT3zeqom3Sz
YOTYFRfzdZO60oHERM2Nbbn6/ap3pJePdAAllO/b9hZ7bdETlI5jsHKgssppNh55
LI1r+6QEecBT7XVfmMz5V3bgxYFBe2kdMEF/iJsH3MEDsLMfEEz22VzGOlKQzbnD
Ui3qJ/DGPnKE8vsmOBEIwMMhl7sGmad4So5pzzLFS2eDT2hKEdxFWURHE2Qbjs7l
5spKvp0wlcw/7Her5cAt9GYm+0yZUhXdfWBuxxpZVEb1cK4FqiE72IDEhd7ZqoQ3
7aM1Na1cXgfkME1agej+dzb56PeGdfx77jLzoy8wIchSYvI+i/5qYvs9cSUeoaBm
wphYvRdvkipvQAn7mfSXRUqrwBMbxtFWr4iId3FKPDNAW/debOwZtQ6mA9HSZhuC
Tr+GYxap6h4DA/SaJVrBlWq4evi+TSXbM2pmgpM13nIkoweZM4az3lTbRiujfg2e
Bcmf69U7JwV8yMFcSg3+D5Cuys5LYtX4JOt8Z+bkVWSL9uHH7VeSX/4bF9Lf4wLW
CTXbyVFZU3PDhQt/bEsJTk61DhP+70D2gP/6uW8baBgBCC0BiBNEmT3O+ILAVDsQ
GS/I5fxbdomAN4Fl+4RewUwI2CwM6gNuHYvHZbrE8gbKCsDkQgfZVa3gl+kKkJSC
niVUFXp1pSCgCvvnCNKvgpHl1RxGVkoTmSaEwYH2XY36Y4Ow/87RuL67UqMimsPb
AFNP8V77xPFmf16KXsTbCpAdiCHWJbiBwkkNC6VZK4Ez2oM3mmkMZIt12BK5tuxy
+xYn56XMu5d3es4CELUOs6G1OhNt2bKaZgBpvTqpD3oSzseD6T6kg6mxHbVzsSvf
RJ4JZdUNDxFfKhlsGJAMiQ4H2Tdc3h1HRCKvce6gAMcWWIM2I7Sia82WZjJOwkGR
9YVh/ZW7BD9RbwkiyaDyxAxaFkzAa/8d+zaBlPpX7al7hrAd0lDcckABepalhAYw
c7vRvdQgFXyrV49qolXAYNMe04qLNqUBBXsHabiZ1BPfcarQ+QNXmLlyzb+vUFa1
D7io0HfymPV+sJ/SXdTIdLs+rG1wIjdQmZEvgHB6B3YK+2cn3tJtO+cbzFxXF/JR
1Pz00TnK4/7GQ8EaevykQ7TKOnAd65wvN2ukmk0cUxXWXgGvswM4u8h25kV2Cepa
/kk5h3GSXm/co5weo2A8iLod917s+VgeCWaQn5zLdP0ILRSIFinP9nwa5TF+rExb
LkanejTzgsJ1tsUSEEYMSFGYcppDbTOHU8vVccekhBonDbntMdV5DI5VMsBHyiDM
LnZ6VM5iegpvojctUNbtNk2B/Uj0/UzxeC5Q5mZI4389KYJiWFnmfjFjT1d+rgK/
lo08qzHd9GmITkMjVoc7DwZXc48inI1Ak2jljcPOM7YuwJjbCi275Vr+4R5pEXfZ
XN03a5+or4q5NlKr0VzKPcZ8WVDomqyQQUov4pZntgfQ7d4vNLC72ulm20KQw03P
3bU3+5Ps3rlAGcC6X3TcDk5SwzCzdwmgiIHXyPCaQtReXkGfKyNkwC7T2ThwOwGY
Xbqxt5JDOCaHuY/N4M94tOm+F76pOv8Mvxp1Wnl2aTrl+G1Qz+Nj4pC4wCFzGP8H
E+KmyB9ACW14Ng+M04864JvGwJ1SoBL4Q/Yygejci7ijcmWqzlUg6qVuy8EcI+8b
rcoCITGys4h8JXWMedGTHSVvIRInwtos58K9OPBrJUhtObG9xNQXiPXS2HAsRndJ
Zh8TSLw3GdyKekN2RFHac/pxHZQWRVFAwp9PBVWfGakHmxJyKXxPwfBP9nIvxla+
66FFEXlrnvRJxx86QOedQkyLfdD4R3hnmhl7vqh+u5mJrGbCvVsPxc1qgHqZISNi
svlPaymbg42eFEY99KuH42quZ6vpqX9QAZgAHv/cklZOoVcFp6EmhpqqrSxsEZHm
WTJrBtUPmvjjOw5YKkdUelPL/FAnLoF196FIbq2qM9ct7SsXK2EpRCuYSN2Zn+E+
iFWsNVm/glKG+i2G5L26lpHKdnI0jLyAr9IXS9E9mOXea7vxQHJlRTd6HuHWwX8q
HUpe+qmUZE/8BJG5bjtmrXK5dV6KlCNbnGkmoTElI4QmDwt0V8a9eooEorZn+3rc
kV/tQqprBOpDrHgSb/KGNk6tOzX/recullACiAX9HyoBneonyzu7mmoOLe3Vw7wY
ayGoi/wW44WH94UHIp3TImn3Vwh4Op+zgyv22Gqsxe6CDfhGI0NgUPv0d0/WiujB
G6eL5+ymHatW3OZltkmZJkxKxUpO3LvPFHDjOkcRwogO6FNqp0F2vfv0ONp4vP/L
WmPtKR1hZNKxQkLT0HZ8mEiVsosDhRN20fjOWwVUjDi82GD4v6De1Lvov8QpMvIG
b3qkK3AzCy9L08lck5KX8+jGFqQ7bdYhQdkFI+OI9BtRN7E5coUpMZgoJxVYgWfQ
B2b9PLOS1dzz3rg8U5M9JUQPHhcyPIeVlb8JXC5UBTSu8G9yDdPA3NofXkZxoHTH
p8UHH69WFNELSraWbrNG/Yiibqy1GO0a7gC5kOqr0cPtZIu4/lKDd8FIY+UIkQEV
bMek15WTsAopWLQ2CWfJpnzjnfDZRaqoUmZeG6ALUZ9fLjxlReM1ONLUsDKKQLyD
fvE1G0vXAf9USdfiqHwddF0oO3zw1cIUSfA797plT3B13AIj04zgCWRarIAtzGtJ
bHGN+OjOeTxvninZVCvu5v5qCVdatgio73x0sL2U96K8EWfepHW0kV1t2x02tbly
bqNCGyVxvDz8oFIhAsgofQO7Q1EaRZnm1L3F0gX0x+AogesgCe/rq9Zj51tGF0ZU
3GKDXamRvAUzyO9BaE17HCZHZ7DDlKlk6uXo1iTz0hNstdNWw+vVT9/I3SqRv0cU
a/qcu7qSt1477hi105WxQyUY2ZYiiDDswIz2u4dqo4K5HDNHGtGj/vdNAJK9FZAU
U58wDLe6oxvGwh+ED9fL3n5NWA+UamqM/M9lIFBrwgRYzCCKRhNCYE+OboGb+Czg
0/xCRE3hNa2bDPd6r6rbCLkGx4ctadJm7ddVb6zpuLyJrjxdq9wx0UWwOkEYMh2V
PBlV8QgHceDlTVXaf0KfOSY69DqQZyrgk4iUxzmVbCpu1QHJO/5fkv9ORWl/ayIy
v4X7/2C8c3Bv7TQP2xcCCMTbIeJUp06WW+aHSDw0smhH/9gGDPlcb+LF9LBziXWk
2yImXX8zDyfH9R72qfF6nDCzX5ToGEGfBwiNWjULi3IC6hdy8nROqbTNsI9/NlZs
7mTrgijAqVpbHXDq80xZvbU9q+/5OyOoZMlPZcQNtXBsq/nXY/GB9E5LyyO7uhXQ
l1p9E/6PiyXA/FtxikA0zel5k1/Q87TcZkudDC/BT7DJHWTx1eK142kNht1+PMNQ
xXOgpV7r/5MpJvBAAHo/Xauq/i9Obni9hFrTyezft9fFXlyeFMxOG7ceDWeVsphH
5y44sZlSe3tmeNDSvKQpwPvpchisOAo7KWgcZ1qLcFR49o6fEwZmFd8ZEcVY6meU
iP2G6qlEw8eSUtipuXJKbA3U6f8wwWjEwyOSo13/7C+mJHLH5iY0/QCg6d4nRe8q
b/HARnxeDBR5VCWXLWXHhZKEHMRCpyZd48bKdeO74Ax4DGlRZXfOkM01Wvskp0sZ
8ppFZUs1jymeicklHTGVgWwYw1z93YdF9fXkDs4ZU3Htew5gHIFy+G/QuD8AXjOE
h+w9dqLg7h1+te2ij6ffyc8Nb7FnK9fBot5C7b9grdRTtqmYYdyPkuVRFwDOnXG7
/wyQdegUVJJvonzUaclC9EA+2ZWTLMD6A9ptpNN0UK4MfvVgZP8+8FHjzOzRjon7
CTfjSOoY+KDnHiemH2HItAaoAnhye20RnheKukfsKxmu6C7OLFxuSDwOtTzip/5R
pVuXdJhWJcwRMScRRFza13iFyGmj3SkJipvu3/Kef55aN1f2XeNW/SdL8wW1VlsE
QxBWVPzxb+zHu/KRhjQpa0XupNdlGNPbKv2zKgbqu14XC/3LC6igjrGET4UNpTUx
yfY/fKaMkblk4Sly+6ZFeHk3z8/dgzH08Dp2vhLjpR17KvI+0rmvCoKLRds5VO3a
v8MhLBWHG/FG1vlMCOBolkiMG+XmKiDf2kEbfy8nHuZZatKWbo9MuId9ceB/QtVb
TLwoqDS5lth1SmGLg4wBbaOjSGaZqf9YdW84Gf7Pam8kI19qJ8ed+b+Lj72Mkv4c
OZQMfueKBI7Z8clNRtx9N87vuCtQ2KThww9r3d1MqNvoGCv4+S3pKnMKkLNcBaIz
efRhufWUNz26fWm1uhzRexxRJlvEHK3J2J1meLno2Jx2Exj6WqRuXCmB7MQG6BZj
Jm38ju2eb9gqo/FQuNXxnO+nOaQ/76kdWV6CTvSP62p6Wyy3itiR6MYHl2uxXarM
5QtQANn0Q8M6t0pf1BDGOydPmWDILupM0ivFavjX2KDlJUFQPZpMnKIPCL4IxlkH
5gw3GzN6P7IkIsyh+foaq8LipvLxeTsJSq/twjyD3gJ3XtFhzglZ2leeaEAVpgNd
VYXohGXtYqMsCGn38nae1AnaK6PmdHOgKgRiKmSl2inP+LahTKWEx4QgMm++RSV+
DnSCffBjjznT1RsShbN4PBZTgF0bDcnLSJWD1CY1Q8WJY0AzqzF/5I5VnMEBSC7s
t6uetNXfEt7mF5xCeAOx0Twvsp0c3JPMsUjUUve5j6nnMsaKa9Zyb6Qu7eoaYTN+
4xm0TSzEAsbV9fPNAdHAU80/YXLmj/JirnumAeZAcXl/7fU/o0DQ85qJ9547YcuO
ArvsRBKBdIsyXEjj4n4ogI8QgzXufOxWtd9kooxQgw3xyheXDegQJ6BDpysctWxN
kdU5/SeAthnggChbQQ70dWduTroYmRmDiS65XIawo1s4qejgbvJQMthhlXkuN3C3
38BoF3jMK3mWNmX357drzIuElly3eNDIeSpAsjTwvyrfKiO4dWKky2/FTsuh1bdK
pwXPnd43djAKv479mtOqCoYmolwu2xvjE88JwQ1BceNQ+qC6czM+tJD3EG/Sr8fv
9OKP9hizX74ER2i95u2PqpgP/xmolVrLXtmPBeiIA4E=
`protect end_protected