`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
ddtXksX2+yylW5zu6QL2Lhnb2d1sD00763mmSITNX595NcHTEkwn0zB1Dry37fOW
FufOhVzEJp80NC5qZ/+F0Vk7Ik02dIR0elf3clrjeJRK85K4e3Hoo4xn7YbFUIms
l/8VZSb14+JVGURjfswrIyCUotIzlzVYZ6gzoZwDXIi5gQIBf/gI+KxNXPaKV+PQ
Ufys/12rjO6aI/pPlqSm0hCvftmBcnezN2hk1UeXgOIuKZnogjOsf0iJVX2aOOWE
6pD/psybjbnsNB6kH5uFTA5frkzIzkzl5d9+YDm9OyC+k84E83I/7/j+rk4L2dah
QJOvksSIzN867/4Qt8qYTQ==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="MvBXkzurAa5VTw+1JJ70nePUfoQXBvZOku/SMmg4TwQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
oRtzZL4VJ4iwysPsC8SXYCzXS8Fw2gtZTOskLcDV+1B9Nzn1zTyNtlo6lNICRmmK
ZRVu2BmCc2G+fmzynYlNTnSa7C0Cuel6FYpxCBlOuk3OF2tzAmLAuDyOH3Z1Yjzk
a0aHuoCdIRKv7BrZCdALt03JeUmXKPdOmIlkVGFl8yw=
`protect rights_digest_method = "sha256"
`protect end_toolblock="Jn9CQpRhJt4rnzZPRk+dOpzAubz7omckX1MrFd4p81o="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 12048 )
`protect data_block
gD6l00tciPUa6pDNTk/+t0OO0nC/UTtBwLB41d4inuAUA3i/ALrNyoJVcBnAmEQW
ptbcNp5fxEUJjnOxnedyZEuEBxWRieZFQnkRdF269oMjCtaIhWZoCSQ8PybjFUr1
sZPwgX4IFEkpO26LWyVMESEMPKLm5ZJq4ru/HsF8lrUHJDtZKYYN4Kgg/ZFvyFob
Thw1mMqr8gonVEHo7gxvvtkFacoJwfymKZnziP25J4FnnccgV3t7OzUbdvDRI4x3
esCzay3R2mmWX6szTREN6HS95vEILoGMrnUvscZnQKl7d/cSkObuQVYVz3j8UBRT
MHVdrmvAbUGpMmLVPgiPEAKi3wB2U75I//Uuxiv5ciqUML4SdJMh+uUQfq7yln8a
HFsUSENnhMN9qodBqR8xt/eCO9ks0MeFWn5M+3bdzT1F3RaHbXbCjZXDEtoO603D
lA6faqYZD/6Oo+3OE1A0mjRq3m3aBl7D5exaxsrBs1wW9WlUyEvu+3/67FMHj8K4
fxnRgqgBsgh/PJEsFU5invYeqyDvt3LCdAz6/SDRV7oj8RBCi8RVYfzdpjAtsUwE
iGk+HrMlkUzR0beOfu2aneasUaQqac7Ubjn0G7C8cLyHL7mR5UZiImPennYBpOja
8ANF3e8BUrPtu4/eG7F33KGRgn8nrtOFwG6vmYx4cDoBN53uZEiALZpr6q64t3G1
WCbo1bloDXz8JqyMOdvWYUZvpVyh39aolEBjG/3w6qpAeBmJgJ6Ai4V7+Geo5N9A
xA6rzIdYbTXrCbM8W9UmGkYFKus9yuxdIBWhIBupDcJyIM9l1L2+Iz8mVbKUQzga
sOD5hJTZis9FUDAa1/WEW4p4X30c83InFOCahlY45aYuK4hPVmvBTxhSOUkMcnVY
V3V2IIxGPmkr08hO518X20BuaF22RrCTulTDRrN2/Z6igj/lblpTHqPKGBrM9mFI
0rZZYze+8CvEPrjKK09Fw6esBGrgLU6uZWkRTqHUYwXH+lcsRTtS5WL80nRymgV3
zYRjPFh7YFxaDo/89MAb52pWDpHaDpB7JY68jrZLnC7IEFUS1ksAZwnp1vy/iaLa
hqvwdQsPNlHkH82XYjDVQFEQT5iWmqB1FzwgjnmQmuIKthvB+ySThQo5yI65i9Cq
V5HzwN/+DOuW05KRfeH+t8Gjtqe9ov2NB5C091CXvw66kOma9OF3bvbd5lwIdS2o
gyEHDjWUPF8c4z4VgPoaSm/xQvQRyR99rsX3E6eggmfz6UhsYSk3U84rUb4J7bKw
RyBuenie8eNWtkzoMwVq8dh0zP+H2GuANkf+Ft3a4UOVD+rowHVFWeBLiwypRSd1
QY+zcjakCj43HXnZedQlIBGrg4ZTH9bMHUOL6UjWkVxtU6V5dk8wSUqTVSNKD/bM
YoJTNs/8dxgWXFQpZq4xeJY5Zvs6Dw9cqJuFRHi4D3VETbJ7NNULEVKQUzfEM0TO
YD8lOrB8AgD7+m9UfnFjgktVsDOhSeSveIDfJJ/Y0+uhObevKIIlzlKUX0v17NcF
h2wfNLS647ygX67e0ef0cl5NpI0V2j/9Hqol4MvI8cdrrFKH1uA5icrVw/YZL4yh
Ogm25Lq0K8N14j04ZjTs0p48XrHAybtAu1jrkVKHpagpWwGZ1adrDT1xP5mtE7IO
mvJPrnKcXL7F4Hpnnp6gJEjtQYbMpGmx/9uyabcHPeFI/A67PDXdaa5UHzl8jH/t
FXHGxdPObqFoU5flERfNKnzCUSu1x/cJz1/USld91W5+rl+HezXhzKYu6eKAXwFd
688jXr8q88xnnqrL8x3it8SZYO06OgPOx3Rr0jFIDUiqzEo+rPx/210ppxj0vybc
ciX9QIGIbeV9uvqtVc6BjZPBaBJtmqEh4g/nFqYHjHJCPJPekNMoy/nJcbkJ0h0c
5OwwuZLUiTxyi89t4xxk4z7Td9Nc6qJ54iSuPeunuWRKwiSWT6Ae5FiqgaDaAPr0
vrZkEHMb+mjfhgnDVKbYY3dFq7MQqwo/R1W62LHQOQk5vq/LHs+nha00+Bs4g90q
HBdr3hhrSjAhXI7ANP1frtfkVKKPS8wE12sxPgnWrxYA4o0YBvQLx9bd2buaRCpu
HZCwocLZv3LMTAIV+O9a4ueEVvAftQ2QzSnHMHTsQImdWtNpqonxLEi3LnsJjpmH
3yM7B6z1wKXb7O9KUMi4hhTuc+SXJrFCzjRlgEvh7FoRInp2iEPFC+fo0gwbd+wv
1cC9OU2c9rPd8h1KnbYB/xKdNbpUbAs958EHxhBotcSMFQ00y5nnIBUkDKYJi7uL
v0QSjQWY0DFx8LQPJJPBbR4on4c6YypJmGpJ1Z8dxTkhJ9XXjhhEgK/fTFZRuu/w
MWWlRwK3YaBqZ3rohcsDY9fjqtnIUD7UlPUiai9e27VkuAK9UX+KK/wfuN3+K9dS
ap+0Dm5o2CRrJP80qmpa0frE7xr9BaV1vNixw30BvlmWPbZ3j9LxhMQRW81K7rGf
C1ZAjsURztvP2bjWJrjLXKZJG6kJr+NqiC+s3BubDSWJJw50jCeDSrJFfLuStQMp
WL5Cn7cXJafpobdpld21mUKbSHYBj6tjeM9bPQ9wQ52yxhJ3FRmHvjnO7em1P1In
4L0ftVXLi3bWVrthmg+L+kGD1wzAwsFDJDoTWDut5nltTemd9EajWt+3d8uMcs14
l7z04utDC/7TGUCmz49cbouLXd5TWVAt5RzBK9A/2n4Kva/9cgeXC2Ngq2rTnekY
fzhZSib71zh5ZZWELKI6uf5MgjVE/rZPk3g77ByaCmzIG6lthTjjJ1naFkpi+7kQ
oH+odkCKyb9v8yG/QgBQeFjOuJrP0iREH0xspJlmzfSANc1eHK+QNMS/XxjQ/kvG
5gFUK738Vhk+Y9fxZx4jhZ+avvR92Aopp3fAdJQ3fwXllKuvKoorG2VhuZAEPCPn
1KMXHGbSN3Uzz2B0fo3jST3IY0g55o0Lll9/aTZr7KnJU9VyyAGDuIqs840aC3AK
jUFFpZLpbnug5KBmMRySNFtxxEi6UieL7O83iJvSlK2SI9rwTjeLMJfSn6IRVEof
6sJa0RIWChFtpGSlKg/m6JV+WTlPRQPByC02RMdnAox/flgKnmsMKe5UdiqVcrO5
bv6QRRERKdaCdm07Fq6DTGPnOnxG49iF6wNxd+EvB50dqZwEfG83wWNbEHP0XL55
R+EP/AR5Jyf/yoDZ3cmo2nD6l2KHYh8qpfNsVqPCfbT0/SEv6V8Z7FLuqYeNDzob
H8vDXvldEKXeaB7hyNX7H0aRUmjeBtwWsSg4MZW5SR/2h8ToazNf40PS5pa2Vvyb
rP+qvOLQJY17KVHSZLGUzISxxeUcOhR845xrLpv2wALbl32M4eZs0ujamaYW4gGr
jb9mgLMFn4/i18tCEo8JQwWbtI4oncpl4MZXBZctuYLcSy+RFJeek7CC0imPmYOK
lAaYrGrGk+TI74f17ub9nXP8VFNOkLF8L973z8GjxsuBKP8rGdaqfCiMoaQ/JfNT
rX0TjHLv5YwMkelbFQoeVkWbLrXey3tKSonRqd269NpXSAGVvoEPDXb/6PjeQ86L
3n0kvUIl6IOsOI48U/4zbtnGGl4oV0oq+qoJ7MON0K1jDVc463Ffa4GBKvXPeXRC
9btZ7x7bpBRt5HsBrKYCXeCvltTBtQ0Qy7dtwBpl47yMYUqVubRqbnGZaib552Y/
7FJzNohEMLjYkjfNZls+6Vflu1Ja8KbJWbZelGd8UqNWi7NnUflle8Wco7T8cpUZ
hMnbIybh6Wi2bS2U8FzHwyMBGbn5NBjazr6OtFPQO6e0p0ksRvRVnpM6ZcOMuCnG
oICMsx+zswQQ1XGIgw480UWZbCO6DBMnAYfcB22ne9y/0wjU28M7Rh+tlUFGIKX3
sd3Tqkv5V1sWcMOL4j3ByGu5bMgiWWSefO+8PrDc2lEq3tvQgeE741q1T4tekhcj
dnONTNlrLpUr2kJWHg9dhDzJMGchYGBJWkLPjk+l2/mg97KYOxtrmGuuD55qFuw0
u/Nrv7evnzIxxumYDFQYFeg5bQHa3sGv25xxF6pgVwJ9N+Z+pq7XZDYraMdxhK8v
7BRHn4Xwq0W0LL48qxO2KxbRJO/rVxTntO2F5NHxJo1Mrz1lHGBJi1xCHLsas8YG
d577bNdZ144PrSHp2YVDNRF5ZHhVPz9XGQCU4Bb7GhdXBMmZJesKzG17ROZP25+w
AsMfP12XvS68tpn0Hsi0cm39HMWDa5RIhk8CRzepGS4sgkbU6eYciBgmVHXB+DPi
WzxcMoNTTI5iA/LoDQcMJENlcPtSgy3SWzHHxm8xBbcPGSBUziJE/u3lsfb3HDcG
ihXfo+I8ZLQQsM06PcxtGI+eIvhPTUkBUbHZxKtZL4DbEeSpIze/IEUHAixVjqmn
8IrlyIeWJbVZNZo/8G9vzO2wJHpNKQk59NwOz4ndegsVaB7skwvP0q4RQb4jefU0
XnTSYDlHvH5MMznwl79d4gngMMYbfORNBZyz6ZlGZrNG5bySvk0oLYnprBevK6jI
ks/ed8lsiRpTDO/lpNPUgroKWqmk1JtLDkx59e5Crh0yjxeTSo8bsLmNN47coNYB
hdSMhjvlfbRvBljB3JHRjZer/zufe2/QHR1iBosM6+J54fSAwvueDOt8HkDHitlg
PAvd5/ca+MZ25XSl6KK9BoMRQxgOXjtt0/ay0Eup99V1sGxvzUM540lItzAfwo6d
v9JUwCsd3SpPaJQEORRdrQDHSN0UKrhsFhTG6+PGcTmEeVnbEUExKRe52zq5FT3j
zhtDN7edqEe1PoOvqXEjVRw87rQNvVcsSTiFSqXGeTzb8MewppKjTJLJaPatB8k+
RWlYIGjMFfj99oqnNpDR5PH+kewacN3xb/o0/7st3SCY+EkmiOm4rcTUbf0JVqi9
PXairkp1IuAnZ2fMVdWl+oIxapOLM8boM65jYPg8/0FTzLMD8CtwlBQlnrIId8c9
wvM6RAvyB6TRcZr+9WaulAV30x2XZc53KudeA0/cFuQqSY5zPvWYmIJvXDFuPI41
9yzOUmkg/4NUtGT/1ybZw2x/t8sdBTeZe6mJWEDtgO2nQUH3tlqbKzkykg003X8V
HVoePUWqlIym1YtRrwfzgv12lvf/xlwRtO5ztFrwaau3ub2IPwLAIFr5OSESyWV+
aZJkULjpLKXmEHajUb/1PU7caq6P/trPmvOjKxw8B7bNxbD++AVPWrhL6ewo6jov
FnJpum3Xl3KY1pgzizwVht6tNxArMVcTAaXVLDmLUXPkHkYjfLeZl8xR9Wdylnwa
8xnTAQr0lP/s0txrVcWZD95Zg/7PRWD0cuT4rh5RbzcOy+Orc4dTk1tsAqhcsbh8
KmjYJDTRkKEAe6DhieoMdkdJOu7Q9TRQNZbieZtNKMmyyCJ68/eZ7fzoVYB4lCjz
ua2HegXsA8ECB/Yi1fwa0L4nTFGm/SLfYm3kmjiGxDzvtFCdBMJoY+LoqmvfJK4u
8NChz8F4wNAwGqUZP6AtPf5x4hkgV2fHfQOr9D7bs70PWNXN1jwUmoYEdHS4lMmD
JZ+OV6RycVCSOYb9QDL23g8fIXqXvF4SbXrI6FKqtJtb3hSzRtkWkEbzNKxQW8Xf
4Yh5X8PeDN55cGqEJlXjBow0Tz3nZBvn5Gmny+S4uupvcMTwCmE7mjI5coruAxgd
qoFJ/I7PvHfDoiSYgZe2nlxs7LizHJJawSFZflYFwrsy2TLdrbRpNXVy1WQ8CTG9
NSG/9fUs4KubmDDBYOc6mV791y2yLRfhBrrtm65UXiIXdRr7rhouLHBt+4RDPK3g
ycrobLXtGk0F1D+4YRhuLSLmMPPs/I0sqv5pyWVecA9tgB+pj4NvaTQQZ3JkPjBD
M/VY2z0Bu2L4Q6DMx28pWLHHwINoYhQjEg64z9fOyLomgETUFWmM85IxlFq3v06u
GnSesw4wCwnJo2sevMWL9p8UKM1SNlupYibAsRHJnKZrMJxmv2z34tIVscIhuQEb
M7299+cXQd/rd3F5aAy2K4+IXX/uUQ4lbUmFjAMGIsrrT5zit3UkOIvzu1WuN5ES
KidxeDpbxXT0MqDqjq4+XO/qJkMBV/zubr2GziPqbMXGDuP20T06spD/SDGzae5M
u9UWFhOezwIL6julfkaAkJY6w0/z6WlYhrDE15O1XDZ3tPkZ1oefIW21E9CgBW57
vEZoTegq1qKseqeHEoSKNcsJw6SYhItfOmfVDzAoagIggRLDV4kLylqQOauIv8Xr
M6QlZk4feA2rcApEqDxnd0UhI2/BNezf0LJ314HTYrt36ZH/9gdouyCfuuj8f5/2
mD/dOJtSjqLr4cw+dThrqmUsUJjD5WtGSyGFDcIz52SBfqAwaxjf2y6MdE4VYDbm
UxT6NjMSe2J3x+Sea+fFW5epxBgL6Jf+DpkX5+WfyxyxiONJaXFkjHriKxAIn+Zd
KUTrcHPtU0q+tDQtMBtbxjB/ehQVCkhDdudGrzmy8Qu28CNGfPfeh8XTdiQZxJuP
EDKc5fX2HCr+NkeeD8cF6TaUZiW/OZmsIr6pFSci3ecm6SUqUDGW+42F5EGzqjIc
QiszERYyLuBpma0jLwIxLY1a5If/XAmd7xuXHpVmEWcJIee9hYyQtJIgOBXrX4NI
Ckh82hg7BNHZymLFHvwIsSkNaoOc16RbGduw19tpsiIN7XxsmgsU2caIJBB3ykTy
62foU91nelxp5FOLoGfSWflfNaeSrQsYDaNwW5shK2TwA2/Mst3H7cXjIq9xB7Dy
gzRMLvkzdWnFjLj3vs57x3uSusLYL0sU8Bvrg64rszRFL7pIATzg/Bebh7PLua7g
goVz5Yh2ZcrI7BN4yfW5Eiba9ktD16N3FrTZVg0pQ8nj05xmXWtNv9w8sfzOYXHU
QEdwuuSzbMFPzLf7CUy6DyKaSHGcE4J7y019vCry1qfOgP55dAmUdAPMe/dPnNS5
xdXmbq83APV/n8Fso+U02kyWLig+v61pJMdHn1hY0N9J+WetzDXF8E6OisNoaeqG
U37FZnqGCtlm3jvii/JYz5I8CcOETbUVabNVC7d23W6g528XRe9oq8gV9N+XTabu
zmAsfdZWEz16vhuJYD1dTWh7vVutxVsf35Azz4oqQYFFlPgqnfCCOk6n598EiHxI
6196RYNJkkLsmxlJ/p96KONX8aLl0Ql83jRGyxa1OTDkY/Fxs2GkFE7cBWRJWlJn
oTXiKQ6eU4BM9LsfwgJ1aaGKQeyH6VSfznu9rbDpaiX0QO3GT2ycKtvYn0qApnqo
frrWUkQITvzzSh03Nfqp4xOzfusHNDEZy4FBwAy7Wjds2xgg9cy5AK1fBlAGAHVE
oP50ANqFO6y4bNrPnJpz3kDSLgLhe+9veAtXrm+g1jrUDRpgTF5FYqovG5CJA01G
HxTfyANs2Le21YlebmXLSrEnP9XK3/Ms7yWJg0N4J1y26YyJkBoZESIun6Hv11XO
7UXTq0XdpT+r7aWbZHsdf8E9ANHfI0QOW/tHOwbuMTVKf+8nXueTgCBC12gG2dws
6Cg+m76IdJjacVIh773EiazuABqDUaiXM0WHbuHw9NrIWGeJXhrGugZmgiuESH/W
wJ5ruoiHwB9LWSjpV9pPBlri8mn1Mzyzx+bFGUf5s8LTMQcblFkUcJ4nlPJq49vV
bs+FVJvwDs1LYOrhljqWS+Qrlom6Okf5TqwbIsqTRajU2J2LBEfc6QYQMvp+DuRu
nIM5AY8vOJQlUhk0hqJXdlxgukLwtHtqw8VJhcVDZRZ+SPBE/yYiwfXNkGzG5gHO
uExjuc3/fdKQ0Yo3jlf+D19SWd4RUOn+xHDWhZuGdnhzumt8tvfRziOk4X5uyO4j
fJDs/n9Jcej9iUBML8H8D2+Xwk6inAEOnBjN0btdQHLsSADnP608ONQxsPY/p/L+
8HEeFTZIcy/Kh87+Jfzd646rEvE1oHuDj6gpqGy+SjMpnk8bwKG1kjY+HTPJkkWa
Fkm9pcj5ftdRHYOXdOhaBBTyBn6mVcTyGKzr6PQv6k97wl98psg1dBgSwP9kODzt
YmhNoIRY3qWWI/LyMXYqgxKCvsCnXwuDK9aXzxh3Cl5b/jMfOytyBoJPITviahV3
iIqq3Eb5GSavgJ95WZ6yP0nQXKsdLkhTFZpiN2Rk0+2gQVsu0fM6NYtO+HeYFyzz
ZwCMEdG9c53ZnWbcRVUOg1obz8KNEz/O0oaN8mrEpwNKvBZSsgsAHJP7zLmWvugd
NLrXZtGB+54U4C1ueUBy1OADN/b/IepsXy+WJhTYe3/+wURFsonsuth5ale4a4Uj
Xmg41xRkFjtrdNGV8VD0+K5AkZv5AhEbDSXAr/JbeA2YMfU72n1YTa7N0eBxhnP1
FV5ZL7GSS05Cm16QVSYk3qrcTLtJlqD8ELbfF3zNckXshAG4tfzed5j3mhXMbRqu
04XbkPmcXsbW9uM7xlnL/jlGVp/wHv3qjbZ/TZYnEfl+0PwaLaiR7tDItkpnXMuV
TO7zc/ilvBILBZQv3WntxBe1Rzb1PLmF51hPH1HVnFjcHEvpIJgx51sqPYTfLt5t
C+cnBwVkCPCnXS0FVs6SdxWmbI68QLI7vere5EO9GB8jjpD3Bq50kN+lJl/F3KAR
LrVFmPffZgr4QsZB4dBqZIOz0bDPIF7gDl8QTZbH3MlkG7tVHsrHxzQ7goQdt+b4
LFf+RwOT9HyRpG39InsKcZx7eUFLeNU8AdjGjCTpd9n6PMcnAYxFWwjAOEFtwU2I
xwH8dyrsZjCJxvQ0aCyApTYLZCwrRRsvYWrxfbok1YB6Cq0BeRQxynaaWuGR5FGr
3Dl7D18VmLBZgZazEj1G1QcY1TBVVg0b+gtE6Os1bG15LHdW3yQkZkjouTg0G7xq
ukzGkLnTy/nr1mVjeaRQgbLHvoenkVz5LktLdnX+80Ao2fxKUapeIQsyoFYlYj4d
XxJwCoHWYFbD0vdp7bsMumOWBui3y1lYm+DJa0q44Po29VfssFdobKFg1ZrPbEmO
ERkbYjBDz2mdQWP9fWgDhiju9mBULRs9N3BO5xqnOVbGDo5LF7H0w/uonxGsqBzI
H0OE0WxpOnCBfL9MhdxYAcmQTMvHnZbyZ402Bj34uyos6Ee6ttlvYeT54LsU0+20
gQLvVhy1b19cpAlDm6Dw+UFGyo879XOh7gonUtEuHayaxJoWgyJccIBfCjTlFHs0
CgEOCBbgMVugC3IY8/tKpAKVrrKFEW3z8v7dH56P6SSZkOIuOsRMPY0sK/GUgEv+
tzh9tWNGs3hugxAuzsP6nbzhQypQImpHFcFSev0Kxx5EVLxcM8l9rLI+4Pvlub6Z
8pI/uB9vJ9xjEe+GYfqElYuJsVuG1oUrIEdWcncoLGOqMSV4fdeVsa3+Tjlxvi7v
Ptvj9IyshmyLW2w/lkxYugaetDOrcMkTZf2noiQ0ZQTscwvMCJfWv+yynDCxozKd
iOrYuW0PHJ0eKqMj+zc59l9gDACKQwhQMwGVdjD1zWjJy/ThYYtFRssAmpZryH73
S1gHIBLb3NptfYoS2vYX5iNBkxSfRBVAd/3KYxkobOk6GMCrleS+EakETUQUuelb
Zlg9DlS+8+ua7C+Fa9wvPTbb9rc1PRtp+l+hnkPY+uxFvIQHatbThCVrJhE24xtA
CwZukLdoGeBmT9SkFCg/QiUsd7HJQi0lLchxKHQfcHnASSJ7bA/USn4ygU4unmYT
J5WDZWWvTm/SOD/LTX4YwkSRSxb6mAuRhLE2yChFNGSDcQUxjyOmM1oXbX/XH2K+
kj1rh79vWxS9jYyMcEaWI50BvAdmMp44+jgJa/Npl0sWZyXGx1ca09S4HVcPEdkk
uOdX2j9xLK9iR/syXygjMXn43kiN6hB3QeMTt0VNpL1t62GNIgLvqf8UX6xTsumy
+5YBsjFR2iTHNt9bRjGHiHf3zTOq7izasc/4DQdmt7ugphDq+mKn5yygWemsVz7v
bn2rCf8PxdmZk5Oi5XUzdWwK51DZXiBdLeTa+H+UkB1LZtgIfHPLQMvePG7vRetW
skB2Cyc75X2GKOapfqJAvXqa4QOAzMjgfI/GUUTwntNI4h3a5TrgM517VF2YSG1q
kScqm5QvDzelFFe/lFKX0gnin73CUE1g2nlvOowARmeddRJs4KHHrZMueo3BWRHU
r0+3l4QWp1KZMaUHl0y8sTu4c18nlc50SHsNF57XyvAuukXgGPlH4nVKT6KCmAVN
aJOM6CSDvN7roT7lNKQp2fXRcH/DrSfOf6U2dTlXuxmOBFomYUbjYUR2ny9xqLqe
T4CSxkfYUVQ/K5+WKCW/+KkGcLtbKNLKUDuIJwepVc+ujuLg3PTsYewraTSuXq3T
BblzKHg3xWY/Tt43TAJQ1cQJoJPABSFeUJEByGJqXij1G/HTbkboYx0L1B3jLFq/
8RRo7ArYzgMoUVCw0OJjVDBsl3m3L6xZg6ca6YXM83XmshJ+UzGU94q0LCwWpsyj
7cj4W8+xxajuVbL+H6EEEWw7JW1UxRYr1X8nahK3PyyM03bXeC9ipLaexWw6jN34
PAYUBZw5zqIMjMhSFw1JSYbsCv/A6kBFLU+7C6TRGYNrD5z0uOcbIVfUmQWh+Tmk
69sQC4CoKOQGWHcQYulLCLy2OniY2JmpB1M8t8kI/rPwvb1JB100liUa01rY9kj9
za1k0ob4PheyTS1R9FYOxb+nU0xxGn8M+w+CGqO2AjtiTj6z1Zac5T8mTaicl9+R
V70Mup95HZlXLPwDYr64xzY2RkgaV+YPQN9uGrQA87KfIEJna8o09xNUxD2WAU6+
OuO2KeLp35uey9rKA3PW1AWaFppInDqHGAxP1U4QthOpkaVn8pG+dof0u47lPQD6
K0fj40EvYH021vLghqUvwGplJrrBYi9Zdf59FgppskGl6gjvPkpq6Cc5+/OnmkGc
9LThErQxy8BoA+JIPvBc8CxuWSmU61mrTEPdEXhBg2PCDcZJrD0ast69tQcgnzTr
odJCVFmtdd9rwRtiBjAqzphozMm2B4iZwJftslrFDsI9h49vGS+FP5R98LwgMW3b
pKfrLaCfs1ocfVFUbF7B3p2A15dwo6Gmi7QBtHrsIvSEM9gw+VtLpgTeVrpDg/UT
pce0prd56Iwbhw66t0NmgzSuT3TDn3mbli84S6df/OztmKRBSzaZ5brxX2Phi9i7
3nMxoKFLPoGpIgLjcnLYJG5lbEFtOOr98C6V8Udt9UVSJVL8x1NeNzBZinOulX1a
2stI4/iZRe4DDRPHEA54QJCMleZYBz9tUDkVDEu+CRHJPh7FdHLyaU2P61kqcIt2
snBOt5vSqhbGDljZBQHP/uZR8nb1S2TTk6BlQef7IrRlnPhWlJjjA5ytyxVGqohi
jSZxz3s2LAak9FQHir+rko7eU3gXYHWfHFs7dI6laIx3jTzlQc78yfClsys4iD4e
aARzu5gUv8gssihKupgGYCi1ff2iRdgp602MffLoLAThtzMFm8DIjWqvHnNmjGBG
MPm33Au6MUTHF8EwlmxP9xmE5eUp/W8GdRZSOwpZdaaFk48g3tRm0FZdZazWvjof
e7mMURRsGBF5KRFLkQR9P8oV48MvXW09HN9ubQ20P7COC0ztcvOLFnoi2sEQSPiH
xrM2vtnM7kZ9GJczxJ45heo5CQLrbtEXehCa5QNxxfPM6iIlUELXEMCatQxKZYH0
Xv2ZZE6xYjYfHa41H84IvAbTJe4okkqz2iPOKS48Plmz1tfT6Bn0bXsYUzst8bAT
Y+zQOlOLPQWLTPkeV4kFPRz+4yHiXsPysxTTYAvly1OVopYuOmrPlZYYqIb3HtGC
BRTpxFltHiADjFFyS+NYLiwSZI4WIosDWNu/lIRhj8y08Rx9kGHMycdkxuEUE2Tt
AkgbCoeV0fB+3VBDcDMi5tp3CHDlc6ZXttnycffE1dsDlX+cHxmXVjzgQqOxwszr
ng2zgZ62CW40j+UY3V0iW7M2avQ/hYNmB6LUyVu98owdfY30ZV17uIDkrXLS/3hJ
I9YnJ5uq8a99i178+herIi/hq8XrZGIDKRVacEX+QiK5NvJoAgh0LW0lwtfv5oik
Ji5mZyeLFRIa7SyswrTyWqJHo1zbV5rvE0u2dbGjINXl02rC93f+hJW7lFLoz93g
QIFGeevDgQz6axl9uHwJTyrrLinQbLP+LAmUHPaENeZavs+hFqw86KfDRaRREpQS
iJYVQzFOQz/59fJbXmp30mUXeEIHztVu30uN8e6auAKW8z6YiU6kr0B4EcdzCFT7
vBqSkEVAPVkC3YCRKZP2y7cDtosLwsMlUiE/nC3DfgW7x7m5Gz8TE7Ar05NutKnD
5s5gJKdkqtzCXhHP4LOuQRR4bR3kyJ9lwh9vI2YXvzfE9wvOYhb+l6lOJ4CX+apS
sFAOtf7cBy9M+9LYb72wM8Br1zw9XOn3D9PVvIOExkjArUw+Rb9kG5p9mrgqclzJ
sAoTvN0TzT/KWesQlTJVssVDmyscn525A5SOjRJoUCaiyDcHkAj1oqe7Km/0q3ZA
4crVBCQyD5PGGJ8D3iy/mQvaHzI0Yah1bsfquaNTTsYnfdywWoIkJUEans8hoqjp
qOjwpnElvVNU6sLymlI7/GjS67oNFrwp7qOe8VfmGOt10UHOMI0NQGRditRLpade
iP20RsQ6oE3oFouScOeleclMMKe23QCLs7u6oMOC3VqfK4S1JcmR8MDJDVmU2mZu
NqbWTFg06D/9AG0a2e1SdIN4gD/G4PLPEAFTZ309HHY+yfq+MY70S42F9iaaFR6E
gZQWk6ffaHJ5Yvc4tUECSfdSHG5sr7UiCvIFyJ0elnYL4Ukmgq8jf4nuF3Ovrqmd
bJqfvmp3wtMMOZ3Lx5x1+zwnSCNwT9ywBAQTXqGZgmP0cAGCZMIkN5+C+RspXMbi
FrT8Ht4UPtZcP91LSua/Uk4UZypRGA46QchIxICZ6DgQSoCa6o+NMqgPYdWygFb7
JvSKbzp2kukZFxKWa0kJ62adnESkOrzbQV0KXres4gysbO80KMYzQmYcweeM8B4l
P7i/kqb6109rGU3B9hjJKafwBgh3FH4i5ZWmT25tgnkzyBx8UrTdX6WHIM43Lbc9
W4VD6JytpP623+anFx0lGTKRn2SqQDeRdIr+WcN0qlZvRXCfeCL6cd6eniiLucML
A8+48vgoEl0ikVGEz8yrLGso/a+RII0j7wT607fnWf6KN9CuBZB990HxhEK2xQf1
13VCwWRRLPEQQ0xj3PrBKpdy5tce4nk9sDU32s42AypN5GTLXBv9alA4e6uZuHj3
p/pDMe8gxvTPpU6BUpPZOK++sEGXQPisZnbjnFCyRf5pFRDPUfeFnqyc50H3Nj4x
57nya8j8wMQRim2x9tRi3aPsW6xeVumLuDYZ5f5kczRnSKSVY6kKOsdCdXW/lHKs
FgsowfEiIY4Q6m2j5+QW6FrFktgIlnHxVLIf7CrVHGQm5qpk2Ib+ejM1yBVnucRm
P+ITQorKBtPjsz3MuT7zuy2oQlgj+cXwgGC8BF3334yZdn2+ydtYVVLKwgf+9A6J
KsmpuN1xI3jQg7jVOciaW5pqrT+2BNSgYK6hvy/XfIAhRaQtCIY93jfJtj5Z14W3
2wLI6vUlrLUZNPb/IIs8oVsxOywpidZLlTwLryii9G8Bso4R2Y7vMnsU7AjigJ5d
p46DJVX5B2OzppKjoP2Eq8FXyAiIlX/ctkSeNnBFVksNO+zHXDs1YOsbLxLoIHns
RG5vICqCJuuVkfZVMYW6bifzUE25OQ1KL0a9MBlx1CAJOF3UaobeaSrBo877NJDc
hk1KnuHWWjzlTV0pLl2VDsnUQ4cWhEzrOLxWU8DB9UdmTq0Ijry5Xf9oxqBOx9hZ
nAa/TWRfHWcNI/dWzpTu04xK33dhiEVh5ZzrNpBpchR2H2Qc3pNV+odDX7WaN4N6
QDHXdOH0Sruh6eqIRpnv7rreq9ppprXjK5w66RueiRuN9a6XXmA3w8JkeuAPJTu/
XgDjmdCkCE+IVqf3xdWLwQJqkP7bfD5iWgtT6pSV1YKkjBhqvJO7sGs0Cu4b6R+8
SeeuPc0qc5k0+/uxv0T9mC24YvHJ9eeN39C08qv0k6RSNR6eaZz9bf4ghLrhVp5B
AVECDiQr7yf4n5OivJVpoYc31k40Io06282Fj+oh20tnyLwWePkEfA4BPYS4vf+9
iyYzO6qhJXQzOFv1n/2peqzvqIBJsYlBhZDgAvzS7JpGUyn1xUFzrwLi/75yfigG
gm7t2OEZritFYvytv+ekxADyDiVFSWz91v9NwpaIgaFStTsB1g/b2SvWlN0cNZfM
4CFldwv3lQukxH9uUDkydxg/V/ecB3VFCdnoO3YxLSeAyoQEyrhlbv2w5J/Y5gl4
bVM2LT/ZBpoRmFrbV0CbSUWNY8okh7RYKvuKKy4JwXZ/rRQrJf3yCrnd6uez63xw
vv3wTGim9h3rD5Y/Bu4YdYCEDLJ+so4C62IbhO2SieHKnYkpqh49aVf3ZWoZK3Vo
4B0aHVRVK6dAQyOL7iLLGyC66vcmkzam4uxzMAmjoTTr7GmE7ha/nQh1Z64783lo
IRXR1Ka6OA2KW2jDeoOhhdIGbUAWIyW4i/miVj9cADCR3F81FgB1V9jiB2HgEjxr
jATWJXiX924iI/LuyedJqRDtehMiv8nyHmmw8ViUTJo1u7GS3aQbqKwra9ADDbgG
VpS41B84rIpK3P8hCUkMJv0LgPnStC0WVptKwsoxqpXHKqSNqplVrJx+ehp1A2qd
0dz6IvkBEUGjSNMxZ+5ot8JQamZ0iiBMq60LL3BqgsZneiu4dzPP9AuUo/Vu3eTD
GLbHdOv0vauNkrfm8bBd8d9uo6wzoO8iQW2Z4OQ7qtXTUdD+coVqB0aJrDqF4bpu
u0XyDcykbc7UuW7le5R22kQ0q7wljQ4FloKiXvwh2fUZuYdQ7iKFScFd1gOJpPsv
lZUetVzacuAn6CTOqFdPJ60x+OoI3cS9DuyyYNIuFBHOm60Cx8MPEAHYnxFjqTTv
KqSvlUvh61SVforyBcmF9jzGpB0AX85FqaXNuqzfx+xSZUNbFJ2zr/VDU1trynUX
A8Hu7ha/A/0kEDdKTBr1g105ndD6lqcsTW72X5AL+gMxew0s891g6HLyJ7PGf0V6
29v1JpAuiRUMh0ywCRp9kOXw3hZZYf6N9md7W8s3iezPNXaePs0/dZm3gZq+da78
C2qGDoatoBJvr5MfjpbS7FCcTFt1+g07wO4nRAil4u+nc2+3tanR33ZDJ9ll8kjE
vFIzLiQCkRS3+pL8dWKuMpYSE2IlfUwD0QDAg3mNS7Ttgu6L8jmaQMf7ZexoKzNX
6WYaxFU1+ZT7k81kFhi61mSU+pxF75bIQ4CPvB2Xt3+koorHoNOsJDz4B8IfUol3
w8iBY7CZxYHr/eLv7DljYu/OLAnUODuwfgc3izeVjR1cdzpREnaBSKPhVHXGLOce
5b8g4QBCs4YGyQrRYs0WZheT3t4UJzbZ4dif86V1Q6HLtyWjFW+FNN7MbKSmNUP7
6X7ZS2sB9OKFdiQq1b2v0Z1s1qIDxVCBkMrm0/23SLxggH2Gy9GZDePopDtw7keV
AtF2Axi6Keper6yfyKbBnp1Zynnji8WtTF/pMNFc30NVVV+raAxqSFGe4RMifbbb
IeMC7twtPUnTWQ70l5/OzAkfymiZ+99kPWopTnuSBkUSALT7dR1k0c8gtDpaICOZ
MPQ1qmkSs8dGKscJCnom2o7m/hSj5m3xirtZBZHFDon0x+2k4WM5y2ZGhaPzHKu8
QU42i++AOJ7f8EuCB5osHIM7NS/SE7Hs0d8IMYtbZj40hDGeP2CJutncY9ZBTr3o
hFA4TVenVS3sOs5v/voCH1wHVaMqQ5S2SWlR9zFf5lonkOq0WCDEpCC8xorCMvzG
XvIeTNoa8AiaU4g5l8wiSWWj0df8F/DBvtJXni5w48u9oZBu/+pj2iSxz+FWxtit
NZwcayP9egRREFbXb/d8iBdo4E06ixsHi5RaH0IxaBYA8VpmTq9HSKARvclvl56D
`protect end_protected