`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
ddtXksX2+yylW5zu6QL2Lhnb2d1sD00763mmSITNX595NcHTEkwn0zB1Dry37fOW
FufOhVzEJp80NC5qZ/+F0Vk7Ik02dIR0elf3clrjeJRK85K4e3Hoo4xn7YbFUIms
l/8VZSb14+JVGURjfswrIyCUotIzlzVYZ6gzoZwDXIi5gQIBf/gI+KxNXPaKV+PQ
Ufys/12rjO6aI/pPlqSm0hCvftmBcnezN2hk1UeXgOIuKZnogjOsf0iJVX2aOOWE
6pD/psybjbnsNB6kH5uFTA5frkzIzkzl5d9+YDm9OyC+k84E83I/7/j+rk4L2dah
QJOvksSIzN867/4Qt8qYTQ==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="MvBXkzurAa5VTw+1JJ70nePUfoQXBvZOku/SMmg4TwQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
oRtzZL4VJ4iwysPsC8SXYCzXS8Fw2gtZTOskLcDV+1B9Nzn1zTyNtlo6lNICRmmK
ZRVu2BmCc2G+fmzynYlNTnSa7C0Cuel6FYpxCBlOuk3OF2tzAmLAuDyOH3Z1Yjzk
a0aHuoCdIRKv7BrZCdALt03JeUmXKPdOmIlkVGFl8yw=
`protect rights_digest_method = "sha256"
`protect end_toolblock="Jn9CQpRhJt4rnzZPRk+dOpzAubz7omckX1MrFd4p81o="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 2944 )
`protect data_block
gD6l00tciPUa6pDNTk/+t0OO0nC/UTtBwLB41d4inuAUA3i/ALrNyoJVcBnAmEQW
ptbcNp5fxEUJjnOxnedyZEuEBxWRieZFQnkRdF269oPUbqa3peahIDOCGRAXtPPJ
ViTKPaQtQexHT22Jf5J5Lt9UaFIhnf2+RrU2l17Gs4e+a3W8N4vALq5RaffZa1P2
9qHHcCTa6jC347hPzSwtA9QdDikJrtmFxc6yho2IZ0Z5wzodeNq2U1B4aCtjUGne
4P8sziS+gv0tBaLqBb9KghuFOTmgx6twm69i/7PVX/WwUzzWy7HJcdZPlSzBIFCn
PLyKzyokAzjAQEJ58oU+CJcqcg88tr3In/NxxaFSx4iI3pDwYp/vcdDeUvrD4dFB
vsaM+ABPlaQu5ixFuykPFQBEr7fbndTXAyglt57HgxEMJOgTnwKj4G2E+9Vk1SjA
KsQGdrrVRuzdFoaPg+l46xLuMgMth8uykbds7yeUsLcYlwcCLBkmrRzFV3an6fV3
a4Tphl/TmVROciFYD0JZRoOt6jskzskiN3awx5nu9E9hVGh6s8DLYBpfdHJyQn89
EGBMIwgb6MNnvxEkXpQN2ohS/ZBzYqTjD0GXlTQDUrULd+xKH00YWCYHbs1GX+iJ
usOUMrZx8HAZDppA6m/LBR3+D7r2s4dCKrozroPjlXpW971ix/+siha3hMg3zWPm
MEz9ADL2p9L5xlV5eDEj1sMdPvpZ8Z0meMKauTlEsEf0OXsGZjxN+PujvBfUIN94
TrxgGgib+WYycFYIJ2bbV9lSZwixaC8VjgEHRuldJiIqmczIj8kD0nSjC0by68xu
KBFNhSPqalYJ7CLJPZemsr0i22ExRFBu9AQhC9ZO6eunDkIiBRXZiEQCQYjlYFq+
1W3gnSCAp69ahP/xpZanqH7bHbdoKk7xGmsqAUmsVXAHvKtscUZYaNmXEFnwvi0j
fyF3yQQHZkBJQCPeKrnsB7TbtA+teC9Gf1l4PV+130Hkl+n2ChIwQVpyQefdhAES
NA1qM/AytSrOaWW08BI6eMs/VihI9ShgOr22NoB/NfoVDqprxcsNw6MXWqf6y7m4
Du2plpuZyjurzJfbU1jwtMRp0EljHZ3ewxl/2cDt78o7MhzPw+MEKoBBk4U1xWi0
xVkee+AC6sxpEFgxQ5qV+UdRDHHEkaMpJNnFGJXln4good/W98cg/OWfjT5ym/TW
ngCQ51ZiIWiVfwznLyvm8J2KvLnWD0nS0CRDJTzwy532jjmBxmux3bCKtVsdXSo/
bmdKXz0+sZxsg6ZOJfsnfhVahOj2/uY5ZWe9QdgrHd6hVvrmnxL8WfUCASdJfRAB
+10GktWRyQmc5VQG4kpAW7ajBOREQBh/KQxDeIESkmOUi19vy530O4xkJwfNOfO4
P+OgKA+LDImrxeWmKoQC6wCETnFvjp2HCtrkFRhf8YoL67lvXEMP7esZ2fVrdRUQ
JkEL0oCy2j8jcJy78MZSoDffwqaRiKRR5S/76ToOMnRq7yyty42SqWBn1QCksJxR
ArJjqwd46Uj3zD3ZxBEflaSyUKX253AGqCB7JnnI/oGYXVtPf4N+bYKl5mpQ4YZP
kjqjsxWAUOJ5O1y3IF3bpVSnObYKTqQBB6MJuCj6Jmnejbq21NfgNYsVieayg98R
tBFsy3/njEifEQIwGIN8QNWBQaKViHsY/kEgA1n6AdoaGB0mUGrDi6u1y5gg3Fgv
8I7TgW+9MC22FMa/2PxwCt5mlsO6RKiNCPzqXJxi2xOpZSoD9CmRFOpKvU5p8bXa
CI9BG4oJmEFKYyY153GMQLQxg8alCAALW/GD74wcBLl81437zc++j4jiMrksFomN
tXn3+Od7Wg6I1/pG2en4+5zNqb8YEGseAb6I7jVnzGHrmm3mk2rba761M+svA+xz
YrAoC9Iz0MA8QkoAnWjE7hf9k51xxFuGnX40mEJ9mTI+pFi35HjRfL9BBkbGnOgx
6z3DdG3S7HOksrnf4lLDXSLpQrkTrKFGD6YLSFh2k37SKaUAVm3FM3ksZFc7h85c
pdrsAVeHCm1ctxGE6VBvev5DPbGkUItEXUklmmsPWT8q5q+T+mz4g6cXculX+ty1
PkAQN6FEk4LvJwdE1MP2F5SoZSVdE2ZIIDh84BF8NA2wuvSPGNGEv86jjahUjyzY
1aQHAK58ea9olo4NYXxbnLHEeF35gM/I45ExhtXQgBVJQjpZYt9IzUxuDN3mBasB
rUPdB6Q/AUk9EHvV/eAWEd9rxpwO6h3iF+yCco76VY4MDpmwpwCNBgrD7myOar6a
jVKG1Orl0pE0+gcssVKI/PTR9IWQH8nBZi75W/0yO/GqSEV7UzR0OH+VuU5pfWkl
Seh3XTRdvwYSb83vlrVK8rsoeKpBYg/f+s2uD66d6y/o9drEGRJyGi3zXlBWi9jU
H6LlbNpI8GtA0ofNRofc2zORFbq9tgLIRhHSzdJe36FyrN3IoVu6AW4IQOIKoGRu
sxtXg9qtJ5cci1l5V1lOfemlyjdgamOPoeU+Md5VSlYW64yAe560gqHSVFIH7ljk
hGhxCiwIcBQ5euB8MwTP/Xw4R/kazeqP/RWmhWjVZOY9DbgQNNFAU7bz6ahy+kXX
SHpoO8nLOl4fn9sSClTtpGUSFG9+1gNyrD/vrKdP0STlY75LPFuCDlG7iytKxFHu
0uix2iczAL61fwaxu1mGwejx3MQe9/Cc8iT2SF9PebP2wlhD2h2xusHjHhq6fqdr
xIK7v3kuPuW84qDalvXRmQnVCwuB6+ltWtyplkcpQv79Ad0qEb2vOkPw1cX00nmO
NHFUHBRHjIQVE2awYxl7ZyQxwu1ASO8iygcxkgT1PH5jBEuqg3Dnp0TZ4VxwSjqO
rCFeXazlfFYKvH4MJEdnCXkctzL14pm/xu8FHDpOXtNsbgfNb6F22ULI1S7G9Jqj
5hUXknrWZklBNsaBGGNqX+9tS0yUhJf99WNEBJ7tLtVVymzZ/VHKO2brAqrdY3iL
XXjR1Z+WGg5r892WmhaZr3Euqe5xzZDD3VXQi7sQ+FokufktkYPq9U6AjHSPV/vZ
jaTQfo9WOYChSwZOpYjzoKbmuc5aAnW70omQdlYAMmoHzNTfDRTBsEcLiAk+Ai0s
D3QoXuc9qrhytBdUuJyFpLqZ8JrmrshS3YLlqMbjL7iH5G3KrOtEpGDmO+kD2XtL
JD7v2YlERgdMya5wXNqjhVxhR3QpqMD/GI4grMJYoWzfFy7u9oZodqRKMRyWjQts
iG4CGdQbHimxMYno+2WpsIu9vOupv6hxnOY91/hh94aAJdGPG/myNEY/OVKHFlLv
XlvE5gJJssu+LUISSZ1TRjDx617kLvnFCjSOO/4xoeCi8LSVBz6vtNyDQBZUgVk1
Jo3p2Xo7y/U7FaDQ/i5iKHbUhZWhRf7B8KR5/3O2gB4WyIxPK0wiVtPy9E+ft8f2
1Ks5mq4Ob2T35e111rbH/vXtdqtJrjV6NW2oyCUFp13rz5NinABsobXcXe5A1jLA
mo4atH1lCSet7mcFwC/o1X5MSfIcP737ngXm9W8N6CzS1TdRU7X+8DZdVSGwpm2X
YE7YZ6xqetDITZpJX15KlfaBRnbZZlPfpMkjzLFZv7v7zGEoTSE4+1nT04sduTCn
BH2GOG9PzN2Vhew2kQsH43D1/qloedtdM0HvXyV4/QIRpb41dwSkG0w2LuTORzV4
duav5OvwUtI3w+xteINUggI3WYQPYja3G++VaJ++JM6aocUbasqvfLwdf7XUPYET
C4pxTgSHkd9cbLyrf+1mJcjlaUEnNp+NIxi3Gs/T7b2pcP9CVxIxvFVyIO5yT/xD
CYrRA5hi6hgOUpF2EYsdye2pGfY/bsTzKqtpn5619HF/r6GAb3qApECWl80C7zzO
1PBJVLy53peANk+fbUmnOA==
`protect end_protected