`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
ddtXksX2+yylW5zu6QL2Lhnb2d1sD00763mmSITNX595NcHTEkwn0zB1Dry37fOW
FufOhVzEJp80NC5qZ/+F0Vk7Ik02dIR0elf3clrjeJRK85K4e3Hoo4xn7YbFUIms
l/8VZSb14+JVGURjfswrIyCUotIzlzVYZ6gzoZwDXIi5gQIBf/gI+KxNXPaKV+PQ
Ufys/12rjO6aI/pPlqSm0hCvftmBcnezN2hk1UeXgOIuKZnogjOsf0iJVX2aOOWE
6pD/psybjbnsNB6kH5uFTA5frkzIzkzl5d9+YDm9OyC+k84E83I/7/j+rk4L2dah
QJOvksSIzN867/4Qt8qYTQ==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="MvBXkzurAa5VTw+1JJ70nePUfoQXBvZOku/SMmg4TwQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
oRtzZL4VJ4iwysPsC8SXYCzXS8Fw2gtZTOskLcDV+1B9Nzn1zTyNtlo6lNICRmmK
ZRVu2BmCc2G+fmzynYlNTnSa7C0Cuel6FYpxCBlOuk3OF2tzAmLAuDyOH3Z1Yjzk
a0aHuoCdIRKv7BrZCdALt03JeUmXKPdOmIlkVGFl8yw=
`protect rights_digest_method = "sha256"
`protect end_toolblock="Jn9CQpRhJt4rnzZPRk+dOpzAubz7omckX1MrFd4p81o="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 9728 )
`protect data_block
gD6l00tciPUa6pDNTk/+t0OO0nC/UTtBwLB41d4inuAUA3i/ALrNyoJVcBnAmEQW
ptbcNp5fxEUJjnOxnedyZEuEBxWRieZFQnkRdF269oMJL+7bWG1NjtSmAPCSnJpJ
1auINm8wX2GQKBRSseeuWkvymvk2XYgLshtdqOybO+MYTr6i9yzeIM6UHpFgiVaP
QptYKt0iJxWvkmFnkePj363n6L5KlPzo36oH94RdSC0dCOz4rpYo5LC9WMfYYHIV
F/vBa3dbgHFK8P/U2v7gWWzdwoUJLW7ruxYxYzI/19CpsQSeok2Q8UrPbNCGbMMU
CkKgbXag2iNG4HTy8YNZQCZmMKs4eN0miVfUN8SBZZV5RbVIAvEXfKYxrQ7Yoe3a
MChBJaRA33tgk2kUXXqtnWvkheEM+Jcz4ISsq6Tz0lZq+2IsO/EFaNwsiNwKyMFR
HpiQ/Qb9HH+7uc3C7CdEHOGT2Pw4LDlJ9pSyg8ubYCTDz+idPQlfHOUcKOEUEegX
EsKEKoSdSIhN1ZXlHdSvCw58SS3ffzdESg6fIlCuj3P1XqmMahKpBwroPVG04OkE
nMegyAtAvEeWBp3aLL5lufjIGDUkUQ4T+HSvvE4MkUvVGvGCC9Rpfm0pvOBfAbUq
EWijhe4e1HTea+X1nv4H7FDbzl996aK6aT1klPpF06jOjDjuIB8QV6PRjbtAI+gm
dGB9yyw3I+6rgplz4HnHviaECKwwisX1dzzKrYGbVb2FTFgBODtZMLU7ptNU4JTT
t1qraTAnbELuicBv6xdOvAoRtpSd5kn50BO+SQWzvLYWBNb5jLtyYzncz4bjwAeX
gfQNloMzWLWNVf/Rdp34zY5w0j+3o7/87bDprpn1xD6TYT4kF+q2YQT9AKJv3o1q
in0UvFQn/P1joneB9rmxDWrOMLZLcqR7TYZvRDafmVUgd3Sgfk6cF16UX/hL92ni
/MMRN3xHYy4lLRkyYWTCKTY2KnpdhJM0kikK1LIc4OBbhPMrg0NQgh+G6CEhCqG0
BEJGVNgdggPPtHgHDUraOfDDJgaxlZE81Nmo/O6QpHmMy8bhrT2S/sPVg0xjxA4J
VWX8DxoIUIgAF4c+4wRQ6FiGUMRAknVjKBT58tLoxuLjE4KJmHiZi5R4vpD6hs00
RGzqVepEz668Pwot4mIeN/XZA5B84flNN/tmUV38u/m3qg49KOjeagDbSRirTvVp
q/OCG3C4T46wE+1zDtNP7ik0BekDMUCz785LAW6o1IELziO9X6JGUGBO16V8tJWU
Xil9ed5TqQTPwNHCDEGn3wGiiV7OxCn/P4uME+3Aw2BTEhm/M7xw+WIcrHsxLmB/
7I8Ly/DRdKSCVds/4Qi9X9rznnb+vqhs21Z55KC3JBiYjVV7f3OeqmKCtoQFEyHN
u0lcc8NdYtwC896qqssadoAF5H5HJyT9lv/01p9vBak1vssqPJ1bx+tysHGYsBZ4
IssjcvKeE5YznGuKSsYpyM1gECcUhGU+elcuTVrgQifAVNvpIUd2fSiv2Rq+Xt1q
AuNWMNq/shJn8oSd5Jw9mr/KhfCOl9JWb6DT5h6PcTWg9S4NcGXMu/gsRxoPXb5X
e7qqnjtexNBwbYozwAeB5IKmj2a5C15PYQBQS10M77XHfySnA4prm5dyKRo9ENJF
QL35LLH8NdCrpfdIAy0tClZpF2f+aCVEchQOG33kCjJ5s25ttiIVuJxgByMk8p97
cLiOo8o3qSYly4/g6P8KBW6zJ0Gzx/dPiOdN37q8CBy3Sa86OSKpOKsHlWZMdR+K
DnhEBd0S3zpQZPQ4THi29YzQf9pN8phKVQW8/g+IjltLMNbU5atkHdimLVfgZoCB
QEIbk9RkYlK7cKp9iY7uZ26m0G7P9OjRT4GjlK1jl+awLYVJqscDVHCynVqjp7T2
AFAEq8mQ2CzvgRBCuSH0c2ZV9cHlntpWREbjaqLEcLAy/fAlKjNkaN3kmuHMJ/wA
D+cz4GsrwaN0Tyaxko1QYD5ISSTLsxhhffyVd9nivqtM+yc1aaDMPFlt6q0xH3eZ
mnMfERF2mqwUuWUK6KlNSbzErjuKV5W5O6yghf/jOCuviiP/7JRAo4pTrArN5lcB
1k0ZSG2bYmYiDnnGhib9GA+HYSGkYmCy5WRp31Wyyhm4HGP56WhyuWbwylvZdoEF
CNYgeGABClbt2Fwd4+By13KVbo48rhn8HNxns/DVa++JQNNqrC27cuRe8hpX/G8B
10AkwKkltrvWLDiEMawwYtGuSiosh7pMGU2ZSyNn8OKkIlMY1ZBBSnB7yw16e3l9
1EHMCMyJwhfQZHSluzKTyjFPDWVg3L3k7iGPiCQozxhXczPNtXw5PYUKfgz5VWfx
4WlcYDLq5byBcYvLLOootGjyCELfvNe627HOnAU4K9OIfUvTsgM9t4J16+Uz029Z
a439uaTJy/PHBUpTaNMewOIq/JtfV1yNEck7KhFO9w/JE5gBaOs6Omnhnz9sQ6HI
zurNPWrAYWhxmhcIvRezZMFMhN9V2MCS6GaykNQIenuaHLIFn5StwDgxBCqaUPXL
jKWrxS3pq0tGHj0LIGvRxh+X80V6g7w35Dp2AhWFeZStF5Rk+NxyXPKsb0uZ06gA
OIf9ZmxylQek5EGKhotLYHUO/rRprixPK4IrKoZr0qs2Xh3SxY6f4eRLANMVWE4X
b5zNx9IXyMSc580+hxP2wi/Q08t4wABlIL3QQmb0AOnI6zu9bqIt/Q4KryYnfQ90
6BSSAnRYzZvbaHkMFVPZuJWG2xOkq9goKyHJq66mzbG6q3SCBKFdBwQcSIO4Ubcc
zSmevIbpXMfxW2fM1359UAO/LHNW8CoORB3ij5UNGp+uhSXQ4ZDI548nEl35kEeH
s7usEtgIosmP2p1WgSNRQdrjN5sLpLToomOw3wytehNQkX9rxjDO0nJ2AcSFtir4
e5akb1nfatSJUCovtVm8LofNGoWIEs+3CcmWLJzK9Ao2b9RHZwXq/YRGXFBSw9Gw
pxAFxRQ4x3mpCweO/kQhKW/9oeiQuWpdz5LJ5iGP2zqQ8PFbheZ0ka/ofKDA6jqJ
RECvXLTX2j59CS2tZggXv3wx23Z2JdvSxMo/2VK+WXrj/bnuPqiZ9jAR8zd2tTLL
JZ4o8i3qBUwSkhDUzblgsUVw8S7Wpgpb0pKsv8JupH0wOoAPdn6R5WRUEJ6tzRRB
TmK+GUSfFxmsJvf/rLvl49yUrzIC5K/+7gKPTS8uPYsInpzommFtITvEAx580Wrw
ajSutfcHCPONziVZqtjSf2WMK/mGruxc/UcZTRa9rESgF6T7yfRa6OtV9h/nds4z
c0TCTILFqV83djfZgMQs7hBlm0tS64z2dNvo6gi/RNSMpN0MgL62WHcHivp8GP+G
zX/nYoOMTzfQJmwQHKVx2EGcR57/VfEWfT/UCcrd7LEc0SBMOPlttzVXZLHgFmlg
P76xGHKtagM39VKEXjJrdZ704vy//Q7F8qIVO7SoQ7J45xZwJQPIvF8GiK+2pccb
9tkNiZUYqrgLUGoDCEtTrc8qb2tnLIftGsl4A+9S6z0vYYpVTOdFBb8JwTqDKTku
Jjs6AWCtI8ZliNmF9VE12ULVaUe/oWoBB/h8wb+vsX0OkJsSVt1PHSE/0dhn1h6p
79tc5QCkbF0vDe63uvpGY77cxUCTTmB4ZP3XF5DO3xekNYF41Cmb1bnntlAtnx9z
rTjWZTP6NFzHrwBMutPHKnDO2gMG0b7aLW5rDYXOTsK4xO3O/+6LA/SMoRNv3xEF
0I5io8PavHfo0Q6dnwDXbx2/ePYZWLjCvdIAiPzFeTTAsi06D4pQwKFcosDxUpcP
6740+VK4QK+60RM6mNxELpyaozEDkdtNz5VzE5FQWLO0THlJfJKTHc6RAznSLSyb
0rXo7Re9NZffM2s/fV1k0M8gXPl2inwYafMNkX7h2ieTsGhRliZ5mS+ncy5p+ZBw
1ac+ZxvxF/5lU3kbWqs20yXlzaQQkj4Lw2Fi9cP0NuxSfBtkCAkE9jOBdisUo4u6
uLZPU7z39f046ObeQ1ba8Ihz2gdYKRMZkaq3jWEuRZDoJoW8YwMod4W0XNDKJ9xY
3xmg1eZZHrUCvz0sdCnhCG/LK/kWPNJcsnO08+VDH5lxHDdEsvEW2Ag8EBGqPiMT
L69h0e84vbcnvrBlQHQhzdY4uCChu3EFFmSZC3dZTyhOJ0DwBS0FwnotZeEBknG/
NwB0nc++diSPy5zfoxIWwmuevxcElvEjdZwwdROzxcBYuVtdwqKbWT4QcMAs4oxn
bW298NRkZ1BEUUawyZVp8NE/ixzkspzK+68W9kPmEvWvA9Q/tSr0XqLOtouVrXM3
KajIpx79azMxrBzj5LVsfL7DRCQ/oNgX+w3FllaYOEPx+Ujq6U3T4bf9iClRs5cm
h/A+GRe9jofb0X2Eo2Qjc075a8pZhFVa7I/GQFEYx7ZpnmZLdQVwz62x0oLoBL5s
wXxFEK6D+PJjp+mj4jHZiMwR2VkYd739iacV92UdCBVKYceIBeVImdfpsFaQwuib
qXBYIIn5SspsnRFG927HM44UuuJFY9GQ5dwt1HyEaYnPlZ37u7NIEE6NWtyiKioS
PuWjtbn88SgVmU7i+iOPtS9lFV7w1LifkNHGQYxmAo33b4knLSoQ33bXYCGxNWX0
ldfvihhH0908kYxp1nRAkdF0n5jFh+0rm9pTgT1fOeDcHsH2/nrsAwvHtpbmv9Gw
sTu756YiZ1jR/rCrnHSdKZtan6BjH+dltIhwpUI9rC78RAtb5xlw4ebaAENmGeKE
ZoxnxE6gcnl5Cah8VMGoQ1PkkZFqknwrktdDOIinwEhEHyExtvCMv9pafTfyIKhd
EycFhpJQxx3zOC8gT3rQkhw2B5ttCBv7//aQJBHWXbUGoQV+j18TXQKL6BPGoK+n
LS64GOs3Qc6IHqJaxMOCOiKLvYs7CmSL2U34QOcnmcMH/Cc7V5X7CTL4Zs8urcl/
f32MTqmF0+qeDrVusVWuZ733hJEgWUCcArR8SlsAmV5IS58Wf/t8w1pfR90y+4QR
ayB4XwG62kIs9frpypNULyVx+9r+uVRxVrSRPBzYMfjjPwFuPKhLoEm/9v4uu6bj
5MJn9+Sz0mg/7dVPZ4u9lY1Swao7WEPzm7k7dC4bopvc5jxb/fwFyNVYTsVj8kQS
hPuHvpU1vrORBr0E6hFzvXQC766mWv7Jlthejg3B4nQjuOI639ksnLowOtNZObAG
x97Fvor1Z2rS7rDgAaHehCICkl1g5I5nSRYerYZUI24GEpd5ggoNPR72y6y7d3L9
RBScWAQh40zpS6BQQEn2KjJDSSMe/GY2PDOIsjle7c5lwjT10Y7e7lQbALWiL0bI
dhA6iFxUAxRrxp+TKnMI9hi4ljv7s7V24xd1LoZ7VSdhiTFPYs3TKmHA51crKSY2
E+ffv8VoGvt47bE2wO5125e6ZytPqW+596sUHILcZg4P5yA6BkjzFP0knDMLhNg8
0q5DZSKt1LexGgsz2i+PVqAetq3iL9eQn4Il/G9mAgdmmmqxH/TB1120Us8ViHtV
/RpkX4BGB/5xn8qcqqW3MeDYr3mgBC9y9xklyuYrxqeOoEh3apE7eF7CIqG9NrjR
XwLZUdsDRcYhPqsiBzt8hZ25vb/HsYKWspuViX2Dz5HGT4gw/g6kl+c1PlqOsQ2U
+Udycj26KptagoYG6fphVpZIqZhmrwhaa0b9MjPJa4Rukfz26iWt6VvUcfW+/olK
/9tbMLB54meBd3l/XOPvlipPGxiZpYtMTwlG/5zSOIF8LAKcmamFwBhMJfj94FgR
tifMJu5J7xiFetOyBoBpcQGVULRmsm/0CUEFfZc6lKYafkvxxM4c/73ZiZq+ApfY
Kqyk0lb3zvz/XHmfwLeQgHqVYeJH+DSFjBuJZm1FneYonJ3fhxdgTE9Ud7bz5WP6
IXZXRZ0VbjkssN2ov1EGk/oLCJDtxH8XycWsySxABmBQBsX8R4W5YUfveBu08Lb6
jLQBdtz5Gs33yu5SToQbnY3pIRVaN4b4hhWSn4HZpEVvhKWCtF/Avjk/iQ/jBirO
/2uy3Vu59Gv/Vvbec444TaoYhB70TxJOviCNcz3Z9OtLH/IduHtstqL2z+aFTd90
TktqtzP4bO0KW10EL0RTFeJL63iIne+VH8m0yYahGGTQ+Un7/9EZzSFcTLVI7hWg
nI1bvTHZiwszxFHhhSpmBIGVQtq4TRtF6nTx36GPPJ02ebY/ElCP54puO+T3Qhyx
2IPC1XoLfeV6bcxJBYy+L5DmORd4JtFfrwuIQ8Z6pAJjwqdTn7+pvT/s90R0NH9p
FjybHl+J3adQopU6MDZJ5so9No/RGl4sqphvV5Jhn04Ir70nheSC8nZeGcwfzzvA
egJ5hWwhn78WmRxUt4ZkQ61pUFxdhxIu6vrt+p1/DvhphG0YYKLL2tAWdUjX5R+3
ZatFzf8IbxBbz8ztktFm8bmihHXEE9ph1utf/4E/WStlOZkwvxWTLENu4kSa7KeC
1M2LuQEYeQgp7uEXAohMwpgHUysBDwrl/E6UtfhM4nS9e20dW72xvKnPGrVljo8n
uAg21cHC5biNZ1AHV4HD27DQYvZwrybA56+WZbdRPZLiHy+QjUCpexaEbbIFN6pB
FlIvRF20EA+wN+Z2YMEjqT5x5WRyHjMCt2IZ7K6TGi2mkkkI1qpEpjgHWj+8buSz
BkiLh4bgl8Jh8B3RkXsLfAm/0AySHyrBuw+0T47Vg/QyH5MNSPn84XsDCc5mCm4R
bEdZlhZAmCqjLOTwmWaSTjhEFF75FbH4fzRYVUEeeEN8QAHPfH9AlOotJDVb8kui
Z+bXYibFvgPpk8gzG2tmwq5ppgDWFSK14PzmMZ2gFds0YUb7WxivEk0AKNikCpQK
tlVNu1zCKC/3U4qAqeHg4k9Zpd9JLXJ+dyoW9knGtn/xshoyjEr1LkzF4pfx/tPD
tKYYgGcIYP+umN6f6KeTdxHkud1KU+6mkoh3AwkimGM8c18Yi76ipuMUYItmPRuN
oLtciwxaSVGPWOn5NgMghXD0FglS5l2HnLRCwaiCh4nHVgZE33LeA4AedHOX0X9k
678b8S8yoMVrZ7vNdv1sQUcVvCoYv9E/Cy31Qc0/BB4MuvQcnDfLCAGNioyqXwYC
bf7EpziZIlgY0UuEdqjn0LFQWrhHQTyJr9gDBUXgrvsxhGGqwISiLqRyGO1Oxf+q
Xr53d/KRk/kob8SWQ5J3PZKxkizgZeaqnOIKW9TQtCx5VDtobBHukUwOyxzhSveN
0XQy/Ahf+35N+tDCg64IjF7Pwp0e7/tGOTR5mVrz4dAZ5q7S3PhWV50/+JlCSyjQ
vrLakCadDzQSiOertgVJTqAGa73XFY1/oqrotvlAvf2kV5yQaMk7aYQ7DZcUUiCF
rMV/TSRszuEgWPmhuTbF8eUYbqBuHxgxEqb4AEVCwHuvmCP5q4bKbZoD4bvAUTt3
411WR97847jNS01M1jhZdQisDCNO7D0nIeoGFxKrtDQDuV+d1JmVIQqja2pNbh7G
UVnRG1wQNyK2QxpzzMABDrZOfRGRDy/tTu8zGOFQR6AyShQVVvTFKy1WgPluc2Gq
mQ4eSmUJkvIjt0GiWMumUHTtydmE2tfmeXS/+PppcnNovkYDWvseYp5QhnF4Bbv9
xKwmPBnQS8eJlwUHKIfKS/Z7Rxwgpp3cWkVsKg4dervOqYil64cn37ZDrbSauqOb
0Z0MKGXPTF2Tb6NDcSgREKs6cCbK/xGyjrgnQAX/zmB41dw2YxYGFT15jDrfhnuM
UmYS1qgYDAty2wisYfDV++la4ca2d8q4er0j1rQl8ZH6iMvNDjFIassoLk0UeJZC
k4Q466gIXlhQO7yUVLF6582tZjctk0tEpXilW58MxMgsoJMPC1twZEhSsXkgUVdp
l3s+Iw8uJCqFca7o96zHOF/C0dwNUlKAKQxavlOZwN+9ML5ZQ5Ql6xNBzv3LWPUa
GnE2FhCwYvHkM1BA9j3Q6dlJRJ8U5NQeTwPu1J/7AHQ8gxuFAkyo6fb9N4TqkQMN
k18warptfPeKeF1P1jkn4sLjYipSdBwbLUa3kBnQiqEI9L5Qdg6qpEqETtT35Reu
MKP9cgzWElYflhRtg2CjjBP1tL7By0BuM1kRI7377i1BrZx3GCmTOUyMncTR577C
38bI2gA1n7vODjEexfm+3O+qTERpR5bl8JTKGuN+4MEEugRkUHWfng6oiG23lQr3
gDoJb53NXYvSuBSXGlS/JRX1zjUFsw18mBO7rCpHqIXeUZs+KIXXDkbIToAhH33A
FCDKmgy24xJQ08A5pJXr0BD+hDi9VTbFtuNP9tM6M8/MC6j1/zLblpIWKOKW0OhN
9bifKjfgGeTiWpqSf/cR30xW4B//O3OoH1+dw6/kmT2i10R3sgkICNtzlVtoeRTA
avngiyKw9K/IMsSqKGcUNv66sY243D8H9/3QV1Yn9dGM6xx7Lt/NRdfVU8eV+ggV
CRby9qi01WWpYN7qg8P7G2SpQpC+4K2deoRkpGw+Uj5HKSz8KKRehzQQUkcZrS+7
0BNCVoW3OfZ21EWo9Q/LD0e90rg80CAHTGGSW2+uWglMaY3n6uu/hvmOH5in0w8n
DcZMB9wSo3njmQm8RHVsyiItZBJ0X6jPxsdelzYen5JD4RMDfn254Qj0Qt909KWq
y/KpbvvnEt39E59lNO1oiKbluOks39O2h+o60Hhb/0KtofJ56TApJEN9c4mv48iC
qqvfplV0YBxJK0y3AdVsku/MDIxEx6KBeyUYLJSPxcGzdGsXUm0C/9yVIWfU3WJe
PtXczEHTZM/hcZ1b/8LnGsTvCh/8a9uWLk0TPxmSXUTD8f6ftoUiFCRHlbR3U3xj
z+YxQeZY3ggpsMXVyvFGurAqOCZFADTooxNAGU8wRGneHW6KdbmXHrGD8GjRbzGz
2GMownkXEjnRTtI8UCuIHivXkjc4bHR7P+h2kBKL6onf4i0vl/62bJVDYxoucx9Q
2dfPX3AWh5hqhO/ncajBVdLLFZjdkz3rkwq/ZFpmUG2D34qEdZk3ZC5jMXAOf40C
GqlJm2lJMM6fYKIymM/5eas0U2RiQAt2FEPyQHD34uHeMinXnZSg3EMxWEppXqTt
qALLwKhLnhlOirkd2o0KP6Qrypf9hE4i9E0DOffI2Zbyt2joeURSVUvq+nMGM1ag
kEWInRpa+WvCmdC5b1d1Vzj0qUHpAr6uvzpLFmuv8DIv5reMkqNwvHH2a+6orkJ8
Fp1eYa3uDUZQWRhEfprXfuezjdb75FO0sNXZm/hPsRIakIAEzNZ5cEpY+CQGQDtT
1XGXip8BGmHQajh4/e2qT8/SZkloEziFshDSJNQTlkNVZtjyMspZHvV/sTKCxPjL
zHgsErbxF8IaW7AT52r6BAEZVPB8y/HrXXXVCbwQtkS+lm1Jq8wRWHbaSab/EStC
n0RsM9NQuLn9DBHMrNPpi+gzQzyxWJ5Ak5JIXaqCbpXaKg4rhg6ywhEP1D2wQHUY
uVpuodNR4f0Y3knmFktyYiy4U6d39sccbevyI60/6Lut9oSJZmPSkcHz1W06ISa+
s+gE7BV0nFqZLt2T5gyfaDTRDWkG80iXtR74jCqV5fsXpeKmMbxviDExt65Ylijn
jl2YXIzoGtOPDIf2206ceBtYlZxt20opjFcX557vPFQMo8fv0CVlCXqca16jlK9F
JcLezXhrpfAgo51o+TxRAJg/0mS1EKNrlRLjVu07CKvUdbKkWhVkDyeVNqem0w73
SaLX/hqfLg6/UbqkzcY1Vi9TnTMa9Q7yWXBkEDdICg1cB6YEto9qv11YoRCrKi0q
29ZEt1cihIIZzc8hK15RFZm093gDNdrIrkiI3FBTYRGl3Y7xsRrPCKunntZWCbO8
Tpp/vhiYc/Un0koQ1dx/kzymmZILXDUHBA3geIyNMRQSruVX/hmhzsYzhLzLReMN
2cgtgxubr2gsK8jLIodeywzNUJOVF7PxVBjjhsQsDw9ZrD6YGy522iPdhqFrp6rZ
K+b1u6qc9UKnPbMDpndy72hO5MnUF+1hBaND9RFEEm5Q6CPIIbzOrpGbCeYe6QG3
sN+sNVpPzb+mKq73nTM/txoVtFHLqOI9ZJfgjquY6bDNS+OmXSaqj+jRU8BtUueA
GaSyqcMuo+731m7EH8MAAfDW7YRrcVuAUGGYteQOxnKlE1GCCmw2EJgJKVGki/bK
UtN21izhol2wn8UAbHyZBy+ne5fzx6t4rlB1pXX5+CY9mby/R0tDzbWxj+lpusU8
UpyRw2zYvEoJtwDl8xHxth5IoVpM9eZ+Udv3mbjt8YvCPjZr+cW+SMvhDka2G36Y
o/Onpq9rpLT1pYPF+w5rzSmQu3YA+0NHxyz3JzaKZmE1hV1v8BX7XWUWYCP8H2g0
Jec+qny+9PuVGMH6fHcWRoN1SbC7SkkzUY6izBAuGat2CzEu4AFCz2kK36WobGsP
5GP25+Q080EHvqyF0EVguR4v1liUIwXNxEL9TTUXA54Br7+/zoW21W2HA9AyEjLI
kL6j1vKnXrtljRAqCCms86NnOKAG9cQoD+wQm+FIFqTnauND9qA2ejSFvE4Z8hjg
yU2Pcy8Q8G5z1F2hs0+1w73MqXUeAsAB5Ls8po2jeKDMPn2AIk03nKrEKv1/FL47
F3xDLbFmQ7iTks+SDiZUYIeSumfuiS9qdZg4QFAB/+4HlpOQkQosnxH1NhanPGN4
bM4tPGBzo1uFAawLvzoy8FN70g+LJpSNohz1YkJN0X8sZ7FmX6cgcJL8kFmu7yuF
/imjcGBLdzd8xVnSrENlM4hCtih/RIY0+JnlaYybV6WWJdd72HI6rK54qj7c+/w1
rvm+6UqZMicIfmztHJUCSpY/W7aOEPz3lbJAymT+c1qkqqbiPL3Q5DBGGMTh5ckl
bwaT6ljxDPHq7Qbgz+VLoXtEIcLDaF+8FPiOE1uNpofoJp/hixQJvUTrR/VVsJDK
VgxFw9DlrLTpTPRmXHNEgUW/Ry44EAPdY4ziXXrV6mTUo+hHgR22JgBU00eAazMw
VKeWsl6QDCY3XBE2jP/nQ8CKyLp1fKpDHHuEF71HyIHrXgfsNXS6xr8t0kWVru5c
u2a41r5BBBB7VcA4LhivKkN07igD5Ni3EhwM/aoB5o3QvXmhImIyFKqgr8DBqCP2
BWtqK6D2JkERaDfKFSZDabAjbphP1hhpb+Z1JtTZaSoix2J6ynmaM25Ty7YO45Jn
PsKRdD5YtKUSas+mX0zTGiyEf8EyWnxOgUdMd7uXzRtFTDGazPieRzrvdp13Mdqg
uWAxRfG77cHVtuqIkNFrRlxrBeKjVBFld9EBes6TGGB52slm2aCzgIquhzI4k40V
sUrX6a26fT35NhmUNvG5OwQCcE/BOB77qWvXYOxh4aU8shUb0JiGHcazQuaOKiwo
UAAbbhDWXkTd2lToo+v6gjtjpdu8H/fx9LGiRU99nFsu5UYQC2k3bpHIzKPthA+f
ffaAw5vKbI0dlPyzovS7h+mk7OrOv21UagwRXOBL0fjMCYShHpuhCR9PX7Krtqza
feVKJdBsEwWdX+boBJK471/FaLpJELnBoxpzzccFBsRkcUYklj6Z2c77VTHaBBRP
jQsPY+lG0J333l9Wx499rauYtual6f/4kfRI9KE2lriUcV4S22sZOn9g2Apz/xwP
q/JSLP9vbsT8dxg7RpVUh7is/j6O0EpfHS6Sh7LYPHyVe6HkSDNMgkZwGM/HZBw9
zeZDePiYttCYOoUFiwqdgTkKmEDU6yoFEAaGHABVPjq6hjezgWKSfUb1BLSTfdSG
Fllm0Bn+64QFb8QejAD3VlhltlsQN//eVk8YhCd/608dYSrKXWjgMRgsjGEyRz++
CFX5Y6W8H683wBz2tVAtGgQW4MB4dgl+pGTlgWdEcMTh8JHVJpdhUp8+DyeokTqr
RrSsmdJXr2lgo8EBGGVZnQu7cyiBbIGJygY930eWSXXmhnwVo2olLfN5pZy9si2y
hfFmgyf/xugKoGok2ooQiLQ/sqZdiS20OOIlJoy/nNDw7xSG4jmV8AjfZRL13GdX
fjDlzw29GO/vXIHKsr5JXUQx9V9o2/wRvTUi5uKfa+xwbj9Cmf/gm4TC8/jrJ2OA
1U5OLNfxE28DhdBlDm7m+pDy4EL/skgreCqnsexMT5SDJ44O5cVmIPWjjvHYhs7L
ykrWlftZyNTVZgfCo7zo/ckYdSaV6jPymCroJW/LfEVswbil9cqUZ6RhqzWlArLp
y11Zi3mkzmYobcdLOm6u5nGACFvfIdKpAjAD/n2urF5fgmW0hfiw/bbwx3rswl5d
yPH1G0FW6X/bpLlsmXWcatTszk2ngBZUJ9Wa7lLbkhfL04RsgZjFOby/32bJrgbJ
5SrR4OoWnaPSBBUwV144EUUaYjQR8VmFgtAncPJKM736x3zQoFWdEcvEuCKM2CuJ
lpZyGKQtC/rKDtUX7R24FT0RehdP2qvjDEJ/H1y9EN5MSHxvr/yGazeXIQtcllNV
RwP+Gp5M9laFc9HuurZdTFzefH6CWVtjVZsgmaLGW20r9vL8WvchAQmhvjaLo9D2
q92EhhDCZpabNfyq1agwamikvz3ayf64tuZyVq0iOTz+F95U2JtNaNNNAfllVeFw
r8PW4TEVKBvaiIYGexbEYnIK4GUhi6DO8fdqqMnNXS5mIi8Jyrl8WTzq3fnuoPBI
b9awJrTipsctQPp0U20aUKr0e2vKBeyC9lKuEmIgGWXUEh9pejR1sejVdhl/QiM4
/WTT1AOOHZAs1ODG9720hMehMq5h/+ef3iWEuDYaCgDS1JJ7mRF4eOAn6tuYa+CF
WaM2w/6yRzJiUOeeRc4tSFOeB/U3fwikKA5OgG/eEN0Gozppk7vhGBBsI6PVjoEb
KyfoU/NzI6wWXxgKsU6Kmvlr5Fl9sEgFevkkK1RNMFw=
`protect end_protected