`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
ddtXksX2+yylW5zu6QL2Lhnb2d1sD00763mmSITNX595NcHTEkwn0zB1Dry37fOW
FufOhVzEJp80NC5qZ/+F0Vk7Ik02dIR0elf3clrjeJRK85K4e3Hoo4xn7YbFUIms
l/8VZSb14+JVGURjfswrIyCUotIzlzVYZ6gzoZwDXIi5gQIBf/gI+KxNXPaKV+PQ
Ufys/12rjO6aI/pPlqSm0hCvftmBcnezN2hk1UeXgOIuKZnogjOsf0iJVX2aOOWE
6pD/psybjbnsNB6kH5uFTA5frkzIzkzl5d9+YDm9OyC+k84E83I/7/j+rk4L2dah
QJOvksSIzN867/4Qt8qYTQ==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="MvBXkzurAa5VTw+1JJ70nePUfoQXBvZOku/SMmg4TwQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
oRtzZL4VJ4iwysPsC8SXYCzXS8Fw2gtZTOskLcDV+1B9Nzn1zTyNtlo6lNICRmmK
ZRVu2BmCc2G+fmzynYlNTnSa7C0Cuel6FYpxCBlOuk3OF2tzAmLAuDyOH3Z1Yjzk
a0aHuoCdIRKv7BrZCdALt03JeUmXKPdOmIlkVGFl8yw=
`protect rights_digest_method = "sha256"
`protect end_toolblock="Jn9CQpRhJt4rnzZPRk+dOpzAubz7omckX1MrFd4p81o="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 13920 )
`protect data_block
gD6l00tciPUa6pDNTk/+tzLxvdHE2s3DQL3/JqqujQBC/Ei+vcAB8wM3doqg5vTg
mdfn9XB1bLOis2CVSfu295W2DNwHfMSTc/8BhCDRnTlLIX0UCJs9Za0+LoM0rMrV
T7EjVWppbP+Em6PkVKCwlmIQ7JKaifJ+Y+kjw9HCGboYo5074hY+K/CBbfsBQY86
h7FrhVb0BFNFA4lVvsm6L7ReLMHd0r4LMpZetSOEmigSTVH60SJCHOaQc+lrSn9w
TDsPvIKSj+qxxfzxo7bQJ6idGzLr8P909WdpnM2cdkisV+L9T5gZ27HASCARu4fI
yHbSEt0cHWft3Ku1YlycoJJ0/5+eZao3guzWYi9UiZi2I55OFWC8CVhXl1YB6RlF
6pD7jW4QZ4UMGQKmha+0BB9tml0BbRRVTJJA4HVVf/ginlwESfn4BThZ2ZJF5kg0
4LBr7WHDVrvfXVauEEgCas3Bel6uiksJ8w8SkUwBeVyUyV1ugnx8fgyH9cT9vYHr
KrwuMUPO7pIdU10ozr/rfKwPSd2MMoulb9Y9UPyfrdsnddMU21Kj/7qhW4Zh7lbq
5v2MImD4u7L+36PX9RjhajFgHRVBmAd/Mp92reBBdctypoR8ZQ3Qse/aJCSbNFW0
u6lJKt3BLgDw1Ekk9e20vOuyRSNWw36RQYFY2lv8Cxqq1kTySP5kVCVGAfUGApmt
yLe9L7K/J8RsN1hAlqXfoQGohTCymTOPAOpx6KYr1FzthtvcM1CSJNJoMKE4WlmP
VwaoewrVg8ti6e56Kz0j3mtag9rkA4tuvMw2+wY1VgPHA4Xy5s5pGw4FziHatwN4
XZF/2jNqYrjMC9QhJDqoq17yRA9UOPLojdZ24cpHq3JC9HVFW4Ybp9rUSbtvvnAH
U7tUo+/1Wk63j/AMCcl4nFpvCiZIf/pS7CRRdZoTqeBIyeqpoYhrzpwX+jQ5GSvw
1S6umwvBtUIDdF6GwVfnIbuQz/7TXoLW6PA4hPh1Y3Vo1ynCkMr77ZRConsreReX
XTuzCTL5p1M5qYQ+pexvd25YSoN+Lxz41Lvxpmivo10IQkvzA9+D6CbHrym0qCiN
3iRmcdvU3eaHFJObTQSa/L1+AO9kpctjfO7rFr19oG+yCeXr1dO5UoDXn1PJYffV
y/zXY/GuXIVhq67006Xi5dQto4iCLI7oCBYj6DmLI7rUB5IDqIAiRWA4Yq7PsEo1
XPKb/7Ot8vLgGuhJcefHNqRKxUwfRp27V5n5H6/sDOHiBVsRLkcx5EGlRl88DhpQ
mnTh2tzp27jAjeg60S+GSpeUGql2YjcWT9FqZcF7cIP61EbeSg5CG1s1jc9FKXki
gMBkJFOJjWbiwmY8ujqUumaUcGaDPoU7P7MCLLkRQVrQI7rmE44nogVOujWbHC51
tYzj+7Bq+58g2pauep1QX6ACz+6c+K4BgLl742SA7939AyR/7ISNW0Wagf2/wq4u
f9ekWtD9bq9WW84OWbCypwSwCW3loPJC/cz6ywGdfOrmHWfz+N5OTVTVxk6kSkJd
icVF2ZJeS9I+nBSiYLmH80EHgkgfJ15fLM4RP+8pdw4kxIFCoBr9BrbNGVxoZAov
lDyjnQ/gILPP0jYSYvqLF3hgkV2yUJA/zb5TSStoFtJZAq14saTu2+qjloAYIoWF
50jDcPJhR/TwqG+/BZgRE+sH9NgG906kSzIQmIigCgjew5HNyI/AdJArv/3rYymk
2EOVI6u0BIkP+SsFEqT9r2Rcv+HrL/kGYNg0MGcWlqXncFLVbg24ktDJE051EjuN
cTjKcKaZ+dotbUrkbjHBcd9bT1xssCHasxD22ttJYL1PheSLT4C4YqCap9u4kDyT
qSsU8DY61JEljHEGrijVMOVqVbLmZh/1yme/UXgqLxADBPmXFMonJNGDvo+Y/TKh
zWGD/X/VL/0Q4/CG1vjjgmZ0n3pJOWeXnvs+FkLs9VH6Yc5zasXRhU4wm7B93Dig
y/qP5sud5lGAY8vx2TJ1wGWVgjJy6Rbo04zofdwwWl68crgmszqqdOLiTQnGPW81
FbRFoHWwaa8poF6ktqo8RiJTHz2V4F5mgajwQV1il3z5ATIcmtswkAFA1lASnKBY
TanvRVY5x3SSiD4GYQV4jMw5o+A/oY2pZkj03bAf5s9PgKTXivecnspHoOPoqSsQ
n4yh0FuiJWhH+olBxIdiIgoTTe2L33AseFiMgGAlg6n7meWMDJq0dgA+QthxmEOJ
B84l7lxqFjhEhag2IqHIZLQkTmLn3vyvJnOo9GjO+guwOp4Jo5okkZHB3lDSxgUY
pxOXBN+iZEOqdPqm7bDtySkxqinso4fNBtK9/CfmddtXEqgO9wtWtb+KwcP/H63D
HQgx+QNOrZTwfZERXrWtr4RJI/aE5a94t8wAwGRGNSWfVXE8uqovTuCdlDytKoqU
pegJq8/Qryy0hE8R4wSe+iWZKrduaL3c4W809k8LG/zIU+wtUmevgXSlIs4Ci3qb
ZP5UbLJXgJPTqqbyy1NxzPwYwYeIUaI6LQk0pFRT4u7zMicrsX8FWGdrUNxWccON
SBS2jjVeLeb1F83cHrYbRV8bn57IIAbVFcKgheJoDzRLOTvF42G1DDrsgewOECsz
siT8bjt8R8z7arxf+ppQ2wRRZAm5bKe3QqQ0VgX2ZuX308KrUDfeqQnBAZ5NgrOZ
bDfgdNoByCl8hfWuN+1+6UEe5zvtj4FQp28ixgKIr/5ymdvbb39CvMGL5CCAZxmW
V47IH/MAiAeYRu/GDgDhqooLYtZmga7m7ze5kDfRtqcQli8pY0G+PAW8RTLwuk3W
NEaeJ8su1OcEYZgyhnmoSTuUss2VueqhoB6ik+yIg7oX5szoT1QGR5nKyh334te5
hLHHDMlpX0rJgjMJO9jsxMbmft+fqR++8onYjs5Gg9O1tfXkBaCai7vbzL4m+oSE
WFrhjHKQXYZgvKyl3mmkLpkAYJxSUVU87t9inph6H/y7RDmmFvsOggoefQjKtVhB
jTSYx5djakXi/ZfMX6URhLz2cmdJY0etJCZKahCxfT2CYF2YDXRVTB5VSZf5y66W
3HUB5Kzc+sRQCV0xrSYhj5WtU5mN9Q69xKWsBjLdn4isV7CGnVarbW8YHUS+H3Mf
LtAIO/c6GLswg4yu0+OddpwJ4tyXgJ4c/Sm+LLfOO0iSGWF6YE6pmtTV7h4QlMNh
8qufvbg3ldmFikAlMMCuyGL8zbEXjrpIUjxP/74UxRLcWC0KZZKk7WYZp+QzFMiS
DQOT10+SzV94l/H4iFDpKO/EKh/Xm2vEHHjvI9TyEhCvwcvcHnzNxh092R77BwHB
HY4PKd23WBz6eKqM2U6dbR3GHWVEOSQET2MtTgbh8YB9y878fFJ5pOmOKIY3aWxZ
SDzwsf572S1XUGCKdTVTelCpOUEBmd2P4f6Gjs2qZKW0Zhi2wQVec5LwxAfif9bt
l8ADCZOHGaF5XTzDADGpil9msefxJ7vKMxUdNOZ8oh/fwry7l0ann4qTs5BVRPq3
d8YEUj1Lu7ku4YSPUcm09iyS95K74vNyaT+7jfPH6aX1zzH2tSQNGIXl/7d24eml
2/vBMuMzZ2J42g5mBCQZazticRp+DMlpYIDdNZnqnbYMZ/+4vJkaWYBG8OybY7p/
wLsxert+e2Gm39bHP5edHsZ+0expuGSdbv743pVAxXXkhKk2Ndy439MPlhup6TAL
mshbgJz7UPhMFDz5lO48fPy9pQFfFxOtRkE/bpB7kv+wPDdW47Z5tYNvbZr8bop7
OStMrv6YBQPf59IN02tQHjcJIUE/2BnWWFPqwmsKRT1aIkQ1z+dkrH+uiz45/em8
kPkqBmHkOMeojsbGQHH4KCQ2XCp/We+SaK2oZYBL/8/ABeRDkItwnwKIF8x6Ur9t
Pq6/bBmy0xFHousN0pnzazsgQ43ogaj2bzaKrGtHdpEgVy4GQEV7dpBvMiubpwFy
TxvVJ3PHsuGJUFGWaP9iztAWkJb3CdsVk8QIRUNoMO8GSJjNwdJ2C5Q1HUSKFFc2
NQ/zFY9Fsmh8VNOa8CxLII9/MitxUzZ/7NhIfVT2bOc/RDrMpgXlfWhl6XWLPj6z
DWpq9FEnbYV48X11QUuk/y4TF9Vlmu+1eEiYYPhXcPqaTBesWeWhR8BeO35L527W
PvCxufvhgYArSXbsXb1wLtSC3jvzE+HUy1ExVctogpypWmaV/NRFq6KPG3Bx1lve
/HaJkUylxCxsqx6PG37gv/YbFHamFWWKAKuYmjqQFmfkq2KRF4o4dnuFIjTBAJSq
euW7xXpO1Rap/sR52Im+8qN/WlmPxOqozeG7zkN4N52zwtHSQvDbLXQcYDRgoCrL
Ov5ASkTEJ9frVefXcYwUm8iwqEy7h5d0rMr80lOvb9mzKb/cqPUnWQ/r5GfSsz3y
tb1QTGagw8OrR/qHQS8yQvjKJGebYMg6EpNxybAAE1+vTNzAk6jkXZguEojNjAu/
JSbPitggX2BW/jo1gynqqk6AfjtbwOnZ/PwrPpo5xGmJsyjiSiUKUDUZrk/6OrTD
EBptR3uZ3x0sb3cWfpoyYpElPWojW+/TIvxTeHytl22ixWLsJJ2/c8oSMedrACFs
A+7M9VjafSsxNzEeI6JLLUzfs1dWWwad5oEJRAAfWjh2lc7JhiyV3yjJqwwhu3U5
2RONIqjZkKTA2aEJa62M1GKR2wX6FeOu/VVdCPyzqS77BEoLc3Z8/HMVSH61YNKX
jq5judYi+ZWA9fKFAWJD5DzADv4uxDHFOCiqeuD/lK4E5ApvHvdtuWpTOqZN9SNy
Mb+SEDZkLLQBOJgP1A1qUF0lpLoEc8tksnbJU8mx1P9NwlWxtl83Cb0zsPfcPFe4
PPaxdmE5N/jrByc9UvSk/QhVyxx+tIRtU3L2hnz7g/YadMJJGzqSbFn/BOZbdMKs
Dz9FSXI7tCg3iM6y1tj2lq2txZHFi+Z6Q5FxoqR7YO9q6ZYuU/JOWyEjHQC9065C
EbGk+tnhPHHVABkTL8CtV/DWUXCDOoNWX3Xv9JEqUVLHt9gkEZpfsUlCZRT5DsHb
fclbwkTSywgwVxeA+B6GI+kCoo81ZnxEXEx7QeBdbozk23AbNOWE1yst5zJdyzXJ
blqMWb8XspPA9qz3eFVC3ZbLPZd6fZRWPp4MieGrhOIX8OIurxkR1qxsl1KH+CKp
8qum+66Gg64W7lMvY/IIAd4fV27AeImDcDUThWoK9SY3Y05fi4nQuSGkpmIzD63W
iJPGjMh3Kkei/wAbWl0YmOkNQ+n7kHc8dBspaqx55Yym0by5lniuJ/vhc/m3MeOe
IYynKftgVfG5qD1McNDI08h0ELT6czvB8zE5elSl5ME4m/FFifgaBIz9Q+7n5QyQ
qnMNbD1L/PfBSGPkTIP8qdSqjI2P6kTghNvd41rvXoz7Ig4HtV2j+uSJe2sKuV6K
50F51cZC/72NgWCn3CANJNRg+MrqJta3utoX+fp0fMNho6chPERp6eIHKp9QG1fn
gd+EZ/rBuHqTHsi3P8ENmXBTNOzd6DhBvid/03zwDxL810el2+sTfX0VcowBX4vm
mCBkbEQfJLjB7hi9H1IRDaW1sjzEzq6U132e2J2bbEZsUC3a0PDyr90LG7oknirn
LqSjpgK/6+/5qon+MJdrEomQqv4QMLAEElwmaNQP+sRrfheMVYjMt6Ap8lQXMN3E
s5fSkep5YO5JAbF5SBUIj1SlJ75gJ4opAYopuAKc404NY3IQhzTx8LyEPV3RtzfH
cQoUXwj9PTlQZSjj9TeqtQVUXLWJ1SVM04n+E4lYKI3vbHC3a2C/2xZWdNpsw/8M
riobQZDt3lG6uRG6S4kQldgiBVp9WMyYt026eWsTOY/JNgZb0go5SOG11hMEEsVy
9zN1op0UfHOcYFV8DNhG8G/EHY/GPebuWrNuKhUomUrY9KhGARGpYWtcPYLuOqvR
Kdsj8qmWPLBS0mlLzHYFG1/uFVeLCJrOqRF4MBaglxJSSD/JSFRjGzVUFvjGntKz
uP1/RDjN5EbBBH38s9ic8JnX0Q2hVZgv11R81C3MTQllg14bNTt0XI9SErSXQsuY
arScaYYPYh1ihAv+x8P2F+h5etG4oqqgAJGdVYAmXQIMT2MiCTjmiEvTiGTkTHhh
75a4oDUJj95zdLa9i7lxHFPgstB3IM32xz1s3c/0SoTZKLLQta8GRPfsMABJLtM3
jQ1pyTHDvJv67m43rUNeY3Ufw8IyJj4UUzc6M374g/+aEgLO4f3HoaL0ND2nX0PC
2uWAc5w7hqKphE5WeW1wighLQxQTlaqX6s45Nv2Vr9bHj53EU9ovafx6yQAeHvPj
5fuNxT1ajC547nYvsc9EGj6czFhtwcIm544Z4FxntKZ782g31y4MZSPsFJ8tpcc5
O2hJ4SXJhLg3AmoizbZ6qdXcRk6+VpBW1jmhIlJRf6anZ8Z9/E89T98+wYkyeI1Y
SfpsBNDQjr1uwD9ArcRn7iAyZEZ5lJqItIdgjYP2XZucSwR+GI58yeWppOYihx/y
SMYAXSfiih0Fru1HJQRI78bwkSBWqKw0wR7FuFn72Zv+KvsOKxWcQ6Yo0qheTvSg
TFvxUvlt7tuOnALp7HMVl5sxX/Z8R/SJyyY3/bOY8biLnMVCF7M53MOtogU/wUXH
SWONbK+3FzJzL2e14xjwD76XTjNINlRgqZ1MdY+ZYiZ9Orvlstz6tlHmo4UXXHzH
80ch9QCY+Ei4rzaA8YD6acgXD/+LVITXr5DywzmJodbAb1k1no919OjZ1wDJxJLk
XkA/ngN8RdKZ/j8Nt8mfT7qRa3W7htrnSycDEFlJRDzZvQBfpT4YPHj/rcPT4GzY
/QATNLApfdxDJ4ZR1ehvD5Rzc1kU2eNQUBzUGELUGBHhrPRC1ls3FHoKmXkd0QDQ
UFEcZIdxWtUxXuA4qpxOkhFIU/jc1SE1fpRvRB6rICt69k3HLrwSXY4IZaZUIbP0
Ph+fksqOEsOprKrZC6ue3CKE97cY7zMaeuM2po3OrhglGYLjfuk/T3lg4MpJXUYY
sheG+6gWgZbFdmYOr+VD1rMs1oSfNze7G/aiKF9aBpbya9hsGlYZ0gVKLszQLsNo
z/RJjna+2ve0EGJDY8HH+yhs08Y8FMXcaUoLscQupUh4XqH7/dD/zD2THHgH7+Gv
pTUCz+FBnixKD53D+gTn0bXten/ME3qUmt89Hiv1gHeI2QBnGRMV9YQY2of0OUF3
S2MAlFUV40yHQrtUvsn+R4c5Fl+QTNmTXkNt21gzWrK2KSUiLRS91dPc10SXmlCt
qv35Jgkq4JvdJMI+lF8lUbvktfAUa8WJGap8eBYznPEXJM54XZyoDlBXBuis5en7
IMFxHB18LUAla9niDCY8XQ1uYslYdDnQenBL5WWqZW5QyT/kdJVRVipBrWBF4NTQ
9nQdcDh38KMethnrS/tTnGqwZkGr4egBUcFsJQIhbwCwhRuaP/qj5VE8P/llzNq1
89sqkhNdcUYkkckNtgmWnjX4V+K4PtrIaJK52T1ie2G2tZs6ZMFE056nvbJ0kqHn
em13prwOl4ykfRZhnK2mUf4pnk/yvKk7FmEqbBYRWJJzIZQVxXRm4A/HEwCPfNWl
0ZMMSidnYJwEeUyrEZS2EXkD3uL4+lnoUl4jiGRohBBLHzdO7Dn5RCx34FOR2xG+
f27X+LADIY692J6OK8dg1wMdMsbxU/LKP9VkkOgXQuTmpW8LTAsP3HWJonxTV2Xk
YnM0sOmyCm+LXlo5OD1hcsAqUlP2VzIStM76O58i58uqL0mflJ/UvHNy6+QyqbGx
5IUuHYFbPwbMlGI7qvrbDG0NIw3byS7Vnl3EZwrAstog42LVO9L+fMZb1aDuEhYj
0JBq2SQ+mD+ePIVL7J22n2avLoYr3JMhX7/1FjTkDA4TvEGpCh00Ybtf+7Fj3XDR
Bl3WBW47V8VkI5nAX2XCc0RGVc9hXIjNYsiEs0R9aHz+0IpKhedT3qFPEjVRQQ03
QDhEr4GfIQiT6L3RkJ1Eq2MvahyqbaF32PSrN6SfnZUcY0VppzQoZvnTmYgR5WsN
xnMUZUwpx9p5taoJJ1d9ULzgpFeg48M7eVI+5mr4yAjVBp0p8rVH9+2bP3foKA0E
Nue0tweNgje1h2yPW3tO8yIJ7e1QdW4stDUMPolxwmrNwAveoHhSoJuMikx1OVIF
qjQO4t8cLG8WSqlLH2TxRRqqupuZUTTZDoJo/RO9MC3uruAEC16BrqC7FbsCvq5G
eOZJDJwbD6voEdrVKmZ6/S+gARC3kH6fShvZ3bKTrkvcG78AZPf4n0wG2iBcSnH1
ETA2+CHAKlk7f2vZSvJbN787qgk1sme3qbstEBinpmaTqONZq+wyyGWWSxgF6dRL
IlZ+4hA4MNoL3gLaqa+URVdHaesyA4KyPXyUY6PSL5Boxb4sqi127Ul3Wt8/r/Tu
Lq6Du10Rtk58jfODHV+m0+ZIHivya/rsC/O6ERL2FNUMDuMSujPejAlclAiLclRq
c/7At9DhRh3CiGHIbw8VMA6txEWCCd9No1JH4tXj9jN+PC9c/LJ5dChAXEjt0toe
sW0UtTw0oxYslDrmfbSi6lsy3X7yNpC55ixhxKWeId9GhY6cLc4a5KDygRrRgNiF
JQ7pq5+bVAqSc5FS0eSr/SEZ8qbUU4IatdbyXhJjgNKtZ9APhQ/mItNUEqgIKR6U
ZSjbtI5bfWRsvc03X0A5ChSKu9rZ1Griic8Pm2YsfwmnX4HRzP/YnAPoIxh+DLAC
5JvuGDFrvqfqmU2bUYEwd8x+N7HMML74ngsE9QzlSJ+wWGR/rzi8g3FSBaCNJ23E
SakPNA5k4Pzqbkh2PBp9TgRcn2nozOipY0BiGVhOILECCfsMe0vJEUOKcwU7XxoT
pcPJaWQ3K/dOQ6aflpCwmP9/OIfh9Ii1zruqAF9SZoK4TtQmPIe7s3Tsbky4vZ5r
Gw44233EcXnOU1x4sqWvsIxmV4bQO0nj/3R9MlGqxShV3+oJ6Mq17JUcVwzC5z/S
Zzd9UO402FLSdg4LcQZQ++o+cHcHY7ngBlHIFO4lkISK2FjztOuqFsnNULSpCI8z
HeIGu8ZVWLtj9n/PizyJh3zVMbJV7vihx3A4CuqINW9y1nTFnqokGwXkFJyeUt0D
scd7O7RXUah1CHes/Uzq4d0y6+ktL2e5o5v36Ch3psOrBMBbr0Dn4rc4hVs0rzgk
M70RffplPeiQDianf4rsrUma41PJmpbzKG0NPrd73oJqbaMleMilcthhEs+qfssM
BZHyY1uzmdtLrX9apmvnUXVycZKhygCzaV9R1Cx7AYqx2v4TVEjjVFn29gy3Zs5C
NdDFys0/5X1r0UIAVEd8TJMQVLMc6i0c5S47kpdzErFrL4XhXfi4OsJffHzs6+8v
fi7qxygPe0WBfuj0RHntYPnhLiPLIiTAPMhrc93fIz63t+9qlUtDRgPUvNmwPmO9
UpaQFAR62oBFj6/y4BS5Uw6H6lFHCoqEQk2806+6IGllgaEjK0AKpo2TEDsLAmUT
36ldVeYE8fdVYbXXucw3kDalxRX4H6M5lFW3BrdwFMqv148Kmu9cFfPS8mMG2xpY
HjdrzXvo4e0yeIABSfJliBQC5VVgEH4H3cQ9KZ4/PZPsqNjhiktX1pa9OQkxCvx/
ZWylOslEvyG2oiAMaiEDRdcPOQstamqv2Hvo94l5K3L5CmwLByXaCBCZ5WOJfAeo
z5U8vXyaOGtGB1awcPG4Ic09ivDGim4dR1PgzVwhW9b9gfT2iQtz24Ssh3NFXCfl
YaCXkUwgLa18JyrdzyLbAD5qtlkORKgJzprOMvqdDUDP84ZNUcobrTw/e8jRWbUc
SXY777At75knYpBf/BO+3j3bb5lWMM9Xj3il9cwEzS6Spi6oi2ABHZatLnjLyj17
PKpBqklbIy/whmkwepMem4SC4MJ/TBLcXMOrYouzpWhsGzce3tWvpZMf44QaKxCv
oB6pE/dVcOS38RyNpal4mcLWm3hrtKBB0zfkrKp+pXh10AHWTdQwk53eFHeygrES
j5cvFPpltB7v92lbFKw1jwePGJOR+jjMbXJR4ZT64oDWt24HuJJuVnszxWmV8VRK
HPl3SUPAxfLC7FBBPFZmnKKQ9cuKwA1EDg0JP5eILrk9w/HVCB/R3UInjnQZMUNM
+gJfMbGPsOonPJh2CpNTef3lmRutVdpbSAHeNIAhJIJwv5E5ybaJmnJt6RclQcOu
o/010QDWB4jMSybotQjLUClrd5kRoyJADE+h+1M3iIsRJ4YwO1VKE0Y08v19XEZX
5x1aSgVTncWO6AyKXIqHn5gJUBVTnhaZS3c6l19EIFGLIqzeD2E0Q+aSD80l3M+E
oU7ggxQmLsuKIGO8FAwMjxr2DSwTH97XAEF5vwDuWAvoeXPyUVMs4/a8i01n+FK8
M5N5rkU9Knv0+EhqLNJU08cUVHwyoo7vVTWsSJsepoGmKSjFadoxcUcQbhG+B19w
GFPEweKWQ4a90plE5/z937udLbN49bpMf7DfibKKbHx0N1DdQptGeuL3/cfE8HaI
eaAGframyDJGmIHYUT9saxqH2q854ltvEx//t2pSJF5jtM9j3f/ANJIq8jG/eKX5
UNOg3iUxbMLthP1ye4icjMa7oH9IVwWP7yYkM0CU063e4FGJPCkkzC0Qh51lAp/Y
Ym+wKOHFnjG7DFeJhf+CNhnxCGMda2jSbZfUunrIMJNWyRIUYBjuUGKMN2ZHxx0Q
VWoV3wVVRpRRWYmVW28m5R1rytgaimMRhHrRYdoBPQPriF+5OyXrZtcfJYlO6jOD
F++OTo1Z2P9TdoLHeJqb4WphN/mU+z2Rc81pcpHXpdJRsDPp0nzNg8KreqnPpWxd
HkxdGpf/tLpmzs8DnPwlh/8mVlIQELR0hzZQPEw6JkjLW9pURWECZe685eKpUPzc
Lk02J7sVIhWsKWjLH7pQ54HEdtnFV2RVl82yKSSq4q+7tjEh61O9ySk2uCDcWeeU
p6Spt010YocjWItSf19CcRElquRqCB1W7ZhW0uSreqAVUL0xSeLjR91+xDygGvfy
kooLXhhgSYpfNN81wjwBOhQM2srd+uAfyv0a2sS91Tbc7fu5iJ6zDkdkdRDNrLDm
0AE21vzGsWmdDuDNTxbSBvfYbqIyip81qePbRYs41ZmgT7vfkTWlOLonHpkW8MGB
P0AZtnGbfL7GAKWlB5DzmdAcxJj2sYoIbeXJ9a9/ksAc6db9QcBixUdvort1LCzs
95e3v6Vj1TcNK8cu75kjeV9ADmtJif6BF+kgKzdLB3zVXnKg2NoamZuRyA4RzvN8
NMQo5Nx73eWf6ynOq5jOcaOTFcQ5HRpzDtGAq1WeIuZK7nFd0RPMoR4rJW9qjoUQ
AjVxvaisaU4XVgJPBFnqayhoC2iQ0I5qVDHPcDuhGQBWMXY+ZMsx1mdOooB3adN0
w+ugljLgRdRFRSvFgRwYxLeqRoPqCzEIBCZj6RmmxysjyI+soJcfeM/lERJE4K9g
je7JQbfj6Cd4TtPeTxuHC8m/xFbb2c3s4zHXBfQibPN5se8PUC0jxLQvEHftYFQd
jyPMi+NiprHEK8KyZ5BIjdJdM/TvtCVXmkbR56Ys/i2GTGu5mGA4u5epsuyPYGbm
9PjrUaxml8SOoo7HxmhU0e5XMejut9Ak9k1Wd99kjEVQtOhoVP2TAfu6CpjLLq4h
KLeeOSjlGIOLWWH5kx8vX9DdcpOuxMb7fF9jCPPT+IAYxa/xfFtS+SgXXhYWSL5Z
QKI2Q88Ccvtox4dYYG8Uf9UcQqBbkR/x5EaTf8iScvB6dGg9+v0wZ7fL9hK/Z5cS
+ElZkWAEa+Pu2WRGOYHtgupA4NGva8sAWMgE6hUVnGEJVjO/u/G6r0l0/kBIkaAp
AVMiFUTjLQQL/GRkxM3bjd0ZCltZ6P3RgJVV+mu0RSj507pMR2W5b8whZtRAHXov
uEnxw5fcGkGHqf+QUe1kLQNmlCUOmBBciFvLzsWuN0Oa3GeFzaKmWBqOyuXMValh
NEuOhf+7Cfi74cSAz45HZQv0Ib1FhhZNNGuWZamWO7QnqcESgydHjsVZ23yXUJjV
jrU5FD1E7bWhQMQfmCiBhCC9jumSadLkwJKDefnlsH2Sml1LtTYtplQcfrePgz6b
c5TGUtDjjAbx5B8oiQuKLdsAoYzkStPvudH64VYkFUNhOLQHouWZoCSuTAB8nLxY
g1CxQhJPLNrG3nUhUoDI4f+Qduae57QIiZl29t6C6S4NRQaVetq7lt0bGmlz/be4
LneMXXVM7qJPN+mxpbLW0brEkDvhW+U3a4PmrJorqBS3fGuropTlwG4wY2kntQxQ
VNfWHty8H0WJnCAf2EMtikVUVIeTh5hG6KRcVgfP5on6EegSyEWmjunP0tNXaLkZ
xfkOacr6//7HsMN7wrIqk1Z9nddI1oskVdgF/TjvG18gTWcBVHBCxfIZkGgmSFEL
HxJJVA5YNIu6F4U45F12Kht2I53PEizx6BJAlyszTh44bM/8U1UmQ9GGfFUKvhhW
fHotvAsM1SxaRPFc5Q88gM03amkAe5qrdnB1obORPvwMNIEW5dqnLLw7tcsIFuwG
DCrgGt0qsytKPSOWztGyfb9ri1VJ9MdajxgGC/jbAe7REjNeGPotDK5mS9jH8+78
H0RbCrrFvmDrB2qtaIRz5j76um7bBLQGCQ5rRaePTFjUWNXtEGISgJw6L2kTmjYO
v+HZWQxkhPaaBut7GZnTVZ3at9xpk/H+cHnETW83DqRngjv8HujaMr9tIOOcep6x
KfBsQ2sDmg4lr8rQc6FI1YkaF5XSjy11bTpKDX1Ms7MRYHtVQZbURwdAr//OOmMy
5zd/LtxxKu8TKSsURVmb86D5zrHkbR00xqgAFuwNukOrWAipnXmhIBTW8RD2RHqF
BsUn9bDiVRh2k3yHL9utO3UJC6GtOd+/Dgc2nRkHkTxwZw+GJANqSi8K2UjujVTp
hkPGfVk++kEjbBfI/tXTQB3su11vneniw2wynMZHGNkZsNOtJOzRQRZydI5ten6M
lu3WiJw35X2ECAkzg5VaE4Xyvd+jmrqmKYMz/LPTjWme5ws43CItOwUbxfNIeX1e
V6HBFwC99KA8fTsSKlwQBVDN2NqGdeYpcqD0sGz2rlcSoqqSfJgUfUrto2v6y4aG
zmHtItcTq3W0j1cme6t5FspgwqFhzbbRP3+MUyXJ9DLJKKbYHQ6dL0hKzQuh8uGw
nipCpj0ljdtc6+CKy9hluVnpoZ0t4SHD6gVkdhahZ6cRvVWiPOjGMugbFrpbH5Cn
Ig65qp2ZEgVKuncsOEjH7XAFphvPf7HhBRHVkHfouci7m1hhNMZ7zObKwMhfgtvw
bY2klH9PHAjX+Cmne0vx3dVQWVOY3h9lIToUIkow6zOSMICHvXclkTl1xtshtwKc
ffA+5i8VQ4RkA9cmKJncOfxjtLOlXpRNE8C8RZzuAZ8HOyLZG0uQoIVOFjprliLq
D9+to+Iq0dwlHNG+9BtB2EhIfJxhh0A9q018efPJSV6+qItG6XDfk721Io4LiDXu
Wy7J0nMInTs0V1i9RZR9GTYZFOgsXIUhtlEHwdbC02MS4moyiVJH1ijv4rUyF4cI
kTuTpWz3YweI3YUOz81yZdNVNO3vb/CSkr+VHLzGl6+N5uz7UwTkOrDk39C9J+0E
gYn8eb6zY0dNBpV6SAyiJwQpSmSPOqYxWS1+G42YTwGJzo+XqpeY9KCSNTRuMKXO
6d6ejK95fbZBuEqQc4l8sempezQ8ceh7YeoXK30fWKdQRqjNgYqkLOUwNUwrANj+
GtiYm9rn9Q/1j/mrEaTT+ItVQlWk8A2tYzamxQLAdyFeCB/N6iMKQwQATgncQKzd
FX48IVDZMcHlYUJ6qsTnEJlF0OBDHcxiWjpx7nXO2nyblgy2UO3d6ExGkD8xTPqK
/uxJE01juGRPqfEx3hDL4QG7V7Mm/jmpTUzyhwBMvQgtA4zyPDpWb0Ew9+QAhUA1
PlBiA/PlSX0fuYGC4ud839zeDiQjkyKGySrkn6FMtx5MdWssYQQv1a0pX9Svu+dr
1LMXmgpxHBqsko1Aokps9ah5X1bTDWwMSV+aCuBqHvqy316bcgpm5q7HAyhhFcfC
EBFXpxHrKbQh9g2K8wWqXJhSUqbB1OUDbij/uLOiunAUnGrg9Qsz33CSMUgHRyID
KxGX3+uhYRQeX/oWKjScbYyjj4r6mSgOCATv8RPwaf0z2rUv7+6kJYP5PnEM9c/k
CnkGCUSdFKqUCrar+7mRphj6wIA1hq/n/okKuPv6CLUhTMpwhnyJLORfoYpNl1dA
pDRxyMvebmxat6Wzd1P3xOex/q5umH7f03vjC0nDpsEh2cBJQ5iT3mUiRQyCTX4j
Vn+UGJYPzy6v+gYjCZ/7Nvh4MoGZTwnASPgLSQlnVYFlDImnf4wuQHy5kur7k3m5
SlzxdgUuNvhuYO2neq8IuB27o5yH3UGcgMQkZDq+HL0pwvDzeC0BjxKrrD7iMD3J
gXh9t/FnqBEsJsxOEftDt3rvG3gbnSacbX086a+/pZGh5JAQATbtP/fZzDm7H1Pp
7WBz0FJK33BRieW62RJ2Jbcics6QJlmSNf9h70UiRgI80df4G1QnafKDgNXkbjDU
PhIk987rNgZUBVeYKjmou5VIUIhqPpx3qvoE9lyIyOATR9TnYsjGWH5nNXFyph1l
BVBX0Hs4wn/AJ0x4d7akCCjeCE7SaFl7nZkUTFR3wki0ejDARqrI6PYhFyTE5cC9
v/ojMlb2PnwVjDd3TmbFTkPtFRgBx05zrZ7ynD2OVj/eV5DB2s1uqGMXpKIkWRbL
w3kb/inCtCMyQF4TUTjYpe+B7Bx3fR0cAmqvOJdcdcei5zWyAtPOZtMQ9wsWVcYo
EVnvjFDpXqyota12v10juiwfd20qn+dPaqWB4VBMDHY7NpVoQvJN4x6GAMCrZaQ7
EoqWf67Hu+2+uX+IA8BNJZ2O7/U3f/HtBdCKmrks6/2ZqP3DvFC8pTfO706S6h+s
C8tYqg5fRA8nM6rtOVACOoV2Wrm2wPU0mj+EhYCCi/B2tZQUTiJlCCFHfc894Oyc
f2yFLJfmnODadRuZSLMLv70XaifOoC8nZ1nuhoDzYk/iOlj1OuwU9DPrX+VuqRa8
p1/iaPo9EbqYy6GiD7uYafEVWTcTGMW8dgmkQWmHiIQJIUegd2KPJe9HGJCZBGsA
sQacvY0IRTBZjQ4pCXQr5SglfPs2CnTYtfrSZw6ZdU93C/pqG8WIquq6+4d6HSx/
0gq3qatH1oufwB+2ZvwMbHtvnWEa9A+1gsbb1mt/adTiL2wasFmuPK7psyNSpaEi
Xju982V1Ak4bH0pyp1oGhAg4ADCxhAmVE7VM568dTQWWskcHJpjR0AFh/c1hc4/i
lm3dtta7HRDHW4AvClgnf5ZKPTOxCNipNz3jgZFydhpgdguMXRJfd+ScZIrKV2zF
0itOcm0iHZ2PN5kMra4A0tLOCSUPbsYrzWXMcDBxQIjsQNSnvBn6F3Nbwy5Atyxr
0AtHDqD3rJouVui30jWK3tRyXkUg3YyoHkBYTvUbRFEIzJ98AHaOYly9s+LMP3IH
XaImG9Fd1j+YnoeF89v/8XKAM53y2pO63MzmaNw4PVhrnViySHn7poj6aZZ4UrUO
TfXD/bUlcnfHZYX0hLrv5kYS+fkB/1sn8KLO2maBG4Jle/2LXbXG/avPJz0+wpsV
2r1C9qDQWCoKBIXD55+hljPbOTztcLjskQHDj9JyTX3EX5h5UbML8Ycu3wa7UYtA
j8/QGxlisqLJCiVtuXEdXOYo0yhfvUgV1kDMi55TvWJDheNcu9/GnX8ziv1Wh7dh
LIU5f5ID1Tqmpb8bb4r0OIRjcnMN/plwTnDysBxFNGpYNY1YzZEL3ugKApUXudLm
UL/i+15jpvJJRYRrABIjr6zHZ2d3T92lQQKCdMcqLXDSfbU/f4+XeNM/F2gcwSKX
4T2lmwu/w3Ppj1CE4H4BTRC/UcotralLf6Mb2dfWabAlq8eWvNjGj5STCSP+07mh
My8mqdwaTnUxOHj2vxapS6CRlt8E2oQzr+ikcD4cdgumi45PqfIRCQ3ZN9CfcTND
/CndVWdQil+wvIHlMwqhORCALY0GyyrVwBnqL03uSFU2Ocdiw0QYC+qmK1lriHzt
0WzVUWYGGnHjQZ9kHfBRPegU9hhlY1GZd23tREISWVGOI2+o19BQHO8joObcZv5W
2GK5eNrnzV3QWLVnlpx2HnGFB02aB5PHAQdVCaVrFp9yFwrNnyJ9KX+fT2Q2ihrv
Zx3o6JB2udoUdyrGwN/rKW40snrIxRIho6sc//nJPnK5qjPaYbk6RITT4z7KhIOC
znQ+VfK8UpfrONk07jIqnhANuCNNT1+KnhfJS/HB6/WkZ0uFMdUVaWSEuYPijCsl
rnicZ+72jOv7GB9j9yEeSxU9Y8jliD4DD+WDNzJDR9NRymmtCfV5s7dekbK+LNHr
T4+kLC/5yHUDsCamOCu6qIeA/0MA1/Ul45Z/uKLH/K8aEOSnGhAGiPODnyixMGjy
+NAoB/tYXpxRaeSqb96nIaSgcfYUtGc8DhWXKJyqRvWgkOA6INE9z8LuE3Gv2iR+
jflfppZaoY5+dlIa6UTiK4lLbEqzMwsJywHIWe8akDADj1Gqyjqdr2XKi/IL8096
XW969IgVlPzizgtjC6lqqBY7CyB1QSaNIDF6bhO8kq38zhc2wZfse+56ctI/89Uz
kWWFb8cDk8l8eCkihpcDDs7FpqhPFqXujQo+wDDvmhkk1sgpmnEMMaFdbC9O14nZ
E1v2LTwziVJfSF+3IjRboPQP4zY/EtwyqRMJ+pomS9d/97xc8dqwf7V76KhxgDL3
QLyZVeUzuUPeX31WBlUVKaHYI22eF/kApeuoZN8BXkMsop0rUQLmn9mxXNyl4SDQ
i/1rQY/gkC5cBMwt4foyAadS+4awXaqemfboQukCyg+aj2/rH4s/6Twj0XMA6g8S
ttQS+SHJWM1PQToHKITfGNGsBKUSYWcPdv8A9d9SOum75d9CukRXWXBIKNsCKxVD
N/VimRyFX15uUyKQT5dpPQIL7sAVN72K/GjLzwGTyaVbEE1vpSHaT1ZKjPmPQIh5
AQtAFOuSMNBq0ez+ZT7pmDgbHKkC4TGeDgR/ad1NBF6j6XQjYQLB25CvMKjHZt2F
I1RtssWt6rPmA1i0y90ep2e/5068YntI647NPzgVIz75WCV46MjQeDVKsiPjuCiB
ZD5yCpdPdo8RKOOvf8p0THNqLooxsXKxty7iYBDxuH0WY2iwYZO0gvQEfKnbMcej
pWbU1qKS7gbzzkwqE5ZoTbHuxonwNJi7STF5UXtpR5bUbpaTe5x3CgYA5MVwVpjS
MD1EBcnhChFyOZ2o8lgdnDLXYIQ8PrwmbCQHvCU4CFdJ1v1KC6lZ+rLkmEBii+AB
gitthfBfL/uysDIx5Q7rupnT3VizMomHDVQqWKVBvZrcbBFIXTilY6GArAq/uEub
hoc9Z7Vcc88fU/NVke4AQQbAcD8sTSCp7Gd1+Ow/6RyRaMFruF/+OzF1Re/s8uf2
6eNbiFm0pyzNB/0WpEm6S/UPO+4XywHlG1/1UePr7+BkZoEch78o7HsGG+RTru5/
flkT7HHLmuZr367tI+XEEDPwTUYSdzflnEOFInCH63LN0z1omtC511+rFibrb61R
eVKyRgTmDvbPdvVIg9dmk4Hoc87GCgVYWFa1RGxywptXpw0WKOdylSZdR/cWRUwz
CmN42RjfVayIyDApol+Ku6l0xtk3Qw0mgAozDIkNumjNumsMUS8KGTqNr221EQhy
3cTyUu6Qg2xRO0CSA8Fxem4kUlmZVlVVWEmWcS/J8AyDVZunviAavfnHi0OCqNkz
YTxGL50FkreqNc4c1CP3PiYrsx8JDo0UhSRqGoj4LUYh2cEvQi92JN6vX1KHIf3e
sUWR1zndTyoMTpxNlWbJx57EkDEyhfpafZ9he5MuKw232TEbPPrWho/I1uZE59cF
3ZEqGMmtCTVZn2zlBjOiB9pO7kUxjLcnrvLVRJRF8klc7tWywNc8trl7u6NOxzxl
oQRDP6ll6koQmsEztOYPYnOLET+XtWQTxa19Nyaq9I+jNp1X4ZzjSnSpesxG+vHU
uIyK86AGI1EOCO33Kt0kEFpWnYDhsFqLPqvOPsRSSs3n1zUwQOJe7nXKnJiI/GZ0
Se16EoyzO+W5jZ7QQzGjUD7gOf8Qt4Gu0y70U06iSz3QEbvpLADwDbk2eyxZsuvQ
8E1qHXgLewG27Gdi+YfNbeaCCkHbp8nNXCGY8E85Gm/mdeb2O/kYulOkfRh5pf7J
0Dz4LEWbfdgS2dlOzXT0DriwyljJRtEp68Znsca85SApv1JEK/z0OURQpnE4VcT9
l8vrfG/0P1Xnb0M7ib6D/A0MPvJRNFZOkOifXeGOkjfLWPeJeeq0KlIwQVhyN15T
1iEYm4S6iGfSZE3drTlKx3WvoQeiMkT8xe8/dfEGNxzR8MqKyDB7aPBMXir4yOOB
`protect end_protected