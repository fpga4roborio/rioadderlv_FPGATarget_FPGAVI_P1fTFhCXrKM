`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
ddtXksX2+yylW5zu6QL2Lhnb2d1sD00763mmSITNX595NcHTEkwn0zB1Dry37fOW
FufOhVzEJp80NC5qZ/+F0Vk7Ik02dIR0elf3clrjeJRK85K4e3Hoo4xn7YbFUIms
l/8VZSb14+JVGURjfswrIyCUotIzlzVYZ6gzoZwDXIi5gQIBf/gI+KxNXPaKV+PQ
Ufys/12rjO6aI/pPlqSm0hCvftmBcnezN2hk1UeXgOIuKZnogjOsf0iJVX2aOOWE
6pD/psybjbnsNB6kH5uFTA5frkzIzkzl5d9+YDm9OyC+k84E83I/7/j+rk4L2dah
QJOvksSIzN867/4Qt8qYTQ==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="MvBXkzurAa5VTw+1JJ70nePUfoQXBvZOku/SMmg4TwQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
oRtzZL4VJ4iwysPsC8SXYCzXS8Fw2gtZTOskLcDV+1B9Nzn1zTyNtlo6lNICRmmK
ZRVu2BmCc2G+fmzynYlNTnSa7C0Cuel6FYpxCBlOuk3OF2tzAmLAuDyOH3Z1Yjzk
a0aHuoCdIRKv7BrZCdALt03JeUmXKPdOmIlkVGFl8yw=
`protect rights_digest_method = "sha256"
`protect end_toolblock="Jn9CQpRhJt4rnzZPRk+dOpzAubz7omckX1MrFd4p81o="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 13744 )
`protect data_block
gD6l00tciPUa6pDNTk/+t0OO0nC/UTtBwLB41d4inuAUA3i/ALrNyoJVcBnAmEQW
ptbcNp5fxEUJjnOxnedyZEuEBxWRieZFQnkRdF269oOvr+qtuBZ9SJfd5JEQeeYK
k682knXsuPB5ymVtRzEp/lNtC4EnHBkJ9Z+SkT76MsZ66ZdCDDWQ+02GdmPZsXri
D6qe4DZ6VLbA8e/ZJ4AmFWzavG1H8iWa/pMh6EQcta5cbMflQwP0l1ohvcLBhlNB
wYCAIoUUSz7GF1sqHHVXkRPz6ZGooM9xpqCvze/NRQDmcsmRaheZR/2DkxC/Tc+i
SVvn5o/nL8zVAsJzlCOHYIDpwbgMH26O74T18GmygLvccQoaedjW711erFyY1VFj
BKvH/croaJ95LvFgZSRDHs1ORTvv2LcStpBQxaziI7I2G21Va5RDsSQbXv59Nsu/
3ZrEeTawOqTwuDY17MKZssLscC9fGxP3vj39Hs2v3QT39DFHmLQnMpWVCCYWmhpn
WbpDfAsheIGNtzXJ3XjRMCLh0BPbJA6qn1y2S7CL6zLgdQQoNeiP8NFJSrKyV+zt
Qs/tQSkuVSkMyhANViOXHYbjRizg4aF+ChdS2aBmYw1Vz4M9m7rPlVubVarR0pVM
jyUFIpD7Mix9amYgh5DM/VzWeqrGtKvgI3fskHcG2hzIeKIeX99XMkC07S9jeT6v
M8hGqGrlfViwQORULlJkNeKs7Y7ScU5R4l/pvPHZXOWfrFiNWhJ6QGrUGyt3ZzO0
tzAyK1Dzi0hEMeLk0/tAYCiaa88BVGD9/uuHgHRHZ/Ix1cRUqBWxYJwu6k1sLJfE
x/gOJJxRNbVh2++FXTb86/DDWwq4PzhWiKpSlGez6IddS91f7ZbUuOnJeyLpnSHt
WonsHdWsQ8miSO+vzDU4uaGJcGXb2FfH9UYjCYY1g7bqGrGd8ELq91INAwKvkkgg
7/p0S94KYk/MeNMQWD9Ym763fARwACPXflW6KIa3DcEtEWM1uOfPKr7X6LcZ4ctT
UZTzU7fvkSkNRN6zrm8kCCcZWwtDaSXoawKk2KuWF/zTgoTN/c2gR6ZCr6iQnNgc
5ROU/Wb1/0ueu9UQdTazgD54UvZixSyUcmMhmAsKhwsrTTzbZFT4jIM1KIV+RoWB
2awbsW4sxG/m0EAh3mKgU1NYvTSwBFJXQhEMdVZFQuBOC1bg9K0Yp82+5rLijfsU
bPMqCap3JXUTzdzK64dTvaaV8wlwgfDdE7FHhM+8cEfElLxWcR8ZUDJcpQA4P12M
0XULsmV4wnJm499/kkdKdj4Pb4IBA6N29Jf7lhGOS6cT30DhuRqSW200gJTmXuZn
bqTDLZXfP3e8agzOMA6ZGMbApsNvmVKZcilviBGiIu+6VSVdW+V6ECz/EK9bY/xc
bUBNyj71AEvt0fpwhxEMSLyhPh1qwnu2UJumUW9s6ex0wdUVpQMjRdaXJ2Nbe0G8
497xrtOIxpAap5Xxy3s7HjlMNvfdttHP11/5YcWxMsgJmi03GEitLhlDlp8Jokr6
lCRei788RNnHpzgP9uNVLeFxXlXiVGY4pKz9HomaWOvr4OB/Km3e6n4dg/xuSsIm
dS1sv3iUb2tCwzx4J5Nk/QGRNICUuzPgohXW1riSlmyQGlzVj0DRXBtDTBPNzekI
ipeTVZoTEqV+JOJhWX0zAheTXeVofwGtBTsyJQHqHRzy3FS6IpW3FHVFopRDrwrM
woNyzD34eTpAToaJVcGz19QPpo/d+JB6J0Qq+RsTYQ/1OCC83+DFoRS9u0qD50gD
JrU5weQaePR9zJSpRNDFwee7WcTqP1VQXSQHAv+yl8toHoe/TcidBRr9SLnUmab9
9/NciSZJTePTm03tcjri32F9q3yoN1u/RrC/K0RIyoH+vxvRvgWpiloE+Mo5Vtjc
xB7Fdclghj0cW1T7AkdQGrHKztM7bnKMGgi+VU9TGUCrwrj9djKZUwoDuclBlIva
wEVmrM+u6A+O+Q/Za2gj/iyEcG4+XHLLc4j92MO5kOxLD0AkaSL63MYKFQ8mkkjB
fe74l4MLbtDbuxtmwmKnt+5wV5BAxWxIJt2HIy4RkCF7iFwSOf5/qXgZdUs7YVTj
0pZuJCRwuUpxK8Mude7Fyd7cCEq6ttsTxnFjas+6WTutn3WR3QZI77c8hVdyxtFk
XX3c2wfBU33ZeDsMBnC/IPxJs4EV26Jf3LU4ooDJQTCLxCAqxt1OIaequc0N/3uO
LnCHNvWS+/qEBRjlgzZRa1sUHbGcvwWo8FxthDpWqabB8SmsdwovaaaKevV3THX+
EygYkkl3nf9pDZn9aWhg9qDPED25atHjXbF7r/k+KzDchcOyQHS7hNqIJ2Qldo67
zvXWjQBbTbkRl4aTy6R6TBMe7PE88ljTFxZf00e9ZzUmzBgWI/8/Qjx42ZRR+nZ8
cdA8vtHOalQN0DnzUp579mZAoTLePSNVYaDoaxsdynYdXHl3L5Zq1PVMVuUqhmx8
5eFMXMF/cOVAIe6XlCgeWF7HxZ1+ceL1xsNDeVhTynje8jnRqC546KGANtPHWfQJ
OkaNkOsaL3ciafADgaUKqieZuFp2DUdicqmbUAoEQY9K5BadXo7w50ZkcXuU7WFg
894yJMr3oTws/B8ehz6PArtBRRKHyeWrC+lJ4qQ/H5wyfi5EWt2dWIiNFxldlYPT
Qa/NG8SzfxynPZukEN9MQ2FWkY21wOFKmHrUsHdvLMWJYltvQyrXHq1AHw/I8zxQ
fGIpc84g3o76uZVwFc+wq3leUR+YUsCphFAm4zvxzloOXvodsCC2l2rUBCfZVyK/
aUK8sykLGNDHrs/MDFvdlk+MXjFsecf3IXqvU3Ia2OdjefIf+afUvbg8YcpduK5p
nijiGdiRKoNxGEVABJt2tKlIyBJr5ZO/wKAD6kiEegwKZgyAR8dy7qYxXuMpw9CM
Bigybbe59y60iy5e1pKWgr+dSNBvu/bi+gV9jNNUe3kQ/kSNpAgvs+isGZ3e///9
no77TD65ibEGfu8PY8OfqmKEdDBsRb7IeKXvh0UDT3U9BFJRBF2Ne3dxeUFXVavA
2Hs7i9IxRnIyK6zxVZyHBbV1BgW3kSwOVN34Enoi1aWswJ5/pcpyzrLtS+0MCxbX
aViOTzF412rqnwd1+Rb98/GiUgj7MDHqnMPx9VdAhgnE1Wxt7NCQeBYg94CWKRLD
THMhljiSEq3/fjgQyCQGJpepucfE2Xi6VdfBfaK5TyP+vtFXJnryawsad3s7QAXS
RQL8dzWy/jYv/A42y8HWRMQdKpmixN4ZBqqKNQ+U6pEQ2KWusXTWKAc3atIQ5j64
43osHvF2u3rLooiOnRrYlQrMbxN171CZl55RKuxJuhuxehO2IeCplv/b3svLVZEA
+0/s6s539KstUfPUCzbBHMSM3atlqSHC9WoK2PkLqbUTsXQMpa5qm2oPEoAiEhJM
aD0PAUpCABeG+S3cHnJ+Q1IX+9AifOY6umlQJduDgFkzwuqxRwIdOaVk4zX7S1Zu
yH1vjYE/zlnRdH+dmKIv1RN6eTjBlrURYYGbHmHqUcM5+tAxxGya0T6CAmzioFBz
BQdTgE+o2vZf/vyc0pK15A5pPI+yNVDk1XhNs0aGgQ8xt3Xn6+3xqwVUvWV4ccnf
0ZWcnB6YfMb6gNRSSgpcMWQZE9GpG+Rcpb46+Adhu2yqS5nS28BDtKc7LsnUnpLV
zxOP2wkmQzNFvHzRj8vZ9zrXFXIk0Zl2hwkaRRlTJGwWkhU9Q9GNns91HJW2ZXH/
Clhr+J5iIPI49LyASUjOvywHg0ifhNtfRtlozuhR5xY+vrMc+Kw/VbbcBhepaVW4
YfogNLTgNL9PbgDcKW0pMGkR1lhDpdVr9bJfWNsui6fhDuzc9tCpolPL6i09SP+c
GIMzmlfPoQLwkRheCfdhsBQg8+nTGZC0/+5rRHesZw1mI83dEmbRzPrHTMiXwepw
HtFCy89kusvcu8Q4hRg/ztDHcenv2pUQazpH+lxPsozsVTq+f0UAist7UYbjtWFT
YNGdW39SXDRpm4hCAbWuIAII3l7uFploEZSVnae4yOoDeAw6rc+ZrppeUGZQLYl1
1s/wzmlV00+wnKbSmGH2RXh2DPDutNmgFRusrlcU7thhF9bP12kv7JsvmIn6BHHK
/cxMFiJALwp+rd5IKJgZ4Nk7EUYm6JEEKL59FZUama/18RSExOTbFOTpmZp3b2tH
rFfP89nG87JCRt1b++hmALPfdGwX8KqV6oVGx9eizgTnBtrHA9aXdxAeSlyx7ZpO
7jaVbhcUl8ij/dCdbz9zk5HbcH4zV7EgWKyKH5SnMPGynZ2BUJ9x/Ww0VvLIS5T7
3AyIebhxSpwSUJnIbbn+cxAVh5ZWrdsYhCbB2bZidE1QSOTzrHqcv2IUT1ehsE/p
MV5NC9PCVUCjUhZWrdSI/ejMFT6l8vFwVZVvYb5VBgjgYd5Af7/fHie5/j/aLBx1
DIL2rOQT1XRO67xXOZVdESEYTf9ocuNAt/3Tfd4y0IfcGzkqBfqwiWsJ9KyZcqTa
KEsuG5iMCOUHAPBa/jL8JHBKtrAXdGF0sdzERQQMKQchihaWFaH2nYlecRJqnQWr
jqpzg3sYtvbtpRYDK+ZxlgMz/DRkwpE0kQwdl9YCYVVzjo0piuqqubJAUw9uUMwm
r5ftizFpcZiIdFiNgoJs4ovl05/zCQnAE8lW63cSBt8sGnWM1vTIxa+qXR0gQlgu
a0v22HVHqnkbS477GlEsVq0/dmOdWT65zNX7pP8+NyBMbCjkhcVXqljCkRR4isMe
71+i5LSJJ+l3Ph7N2KELtJMmibDEhuZQsmysWq5YY146so+sUIxl0sWnW+ks95Ih
Y8fjGtQG6fLzs1Lrq61gNRFDfnIsxeIxiG6cJTD98waC+C9qZCGcm3f24VhanFvf
Go3zgEASlQH31crncgeRzZ7xYf0mbFn5L/uLcKOCFZ7tdJhTGGUCWEZwuMBs7AaA
zU7SPwh4kDksX/0J/WO3vSd9pNNLselL/rKRt0aQysGr8R3Vn1pwLTkFAa58YnpJ
as0MAb/WDgUmsXFgqi4TUg2kak/I8JhB+7+aDnJXy6teNibo2CeJiMvcrdvJueqF
QFxWemkNSAzT/1eM4D/VEuAfgG/IeghWl9vB6c80Zs9Q/enr9Iwzt0Lgm7UNa/ZZ
vSUONJCgCiL0ER7VrUzwqZfbPg3UdBTBQeawR/qJLVJE1YrWDpoHj97QJflvw1Qk
4Ryy9yNdSOx5zS9UJRQ0dXmHC75OROJ5py2XkuztHyvsq9SzFF/95XphfnRNzTaR
0UQ1LNCEvzjG2NEC1L5kzaKXID47/OJPOVvgSnjua4Jyc5ibN1VJwZ6KwnGIuBYM
d2NrQYpC3rmcJGikU0beuKTvjLPQ01lkePD8bogvIP/L7TCcJcr8wkzLQf7ohe5D
EpNJZWvRQr/Jutugfpt8G5rWcZtnI/huOUVLvvtAkMg1MJJsxoatFz4bQRJJO+1B
PCelfJNnQSJ8ojK2MKFJYLAYhWAd8ViMoLiy8Sfv1PZGKqnm3l0RVT4oy2LZl17+
GenIfsyO9+3gGX9YDk/RRpX2g8rttUZaJ/UDBjLmRT70n27huZlaAYYKVus8E+/W
fYoLU7E4YCeaVK1FepC8SoJoS/H3CTjO+5HmtlrlmMT5Xgsiuz3oeP+sPTDMrDwi
ub5Y744shXyqYeXBy6iekDZsJX6EOXqXHABz3F3KDsHDiJ4FGDOgUEuRmgXDPPQI
WR9Jg3f3N/YZi9h/8PQ/3oLZdrsXsRjIE227qsEDKaO8MbYxziVzTBXOdihDNh+V
Kr9Sbn5CisDGrRX0q/ZXdKWo6kz1U5NT5/3VUVZ+P6imj8Ib80yYIxBWEq1bI/vz
s8u9TLmieKr0nkJDijnxZ4kKhlblMfq2W0mx6bRlnpKPptTjkxHmP+qYsDJTJUsf
MIg2BdXvLOgWIiFKlagu0TK0SS+P4z+4qELt9u1kQCVf5R4qYB6IhSMLUwLuUhCz
yko0JC5vt3ZEqmzTpvnquaiyGEnDCNtYfAE9cEbQWaDH3noHksKAMz2zlKSiP2LI
XK6qxjk7tsvN7rEQN8AqElio3cO4IK3W4yBHZ8s/RFEpMQ4/vMRPTMrMFmK5PLtR
dJnKY6PVEFbYaMyryVMEz1u08nnRP6mFW4URfSm9/qNoOHVJzsUXse5+L0dp1fP8
Tqpmq5QYvXjpioFloJXGj+TSjYkReKj6IAcoVShhg1XuSXU+BRv7gkHj2W4Tj0es
ezH2Pc9sN1OdS+iEqbCHG9Qqycb0AoPMPf5aGOXACl+TxSXqdhdUaX906EK6xd7D
+Wxh8x6nf9W09Y6tA9HRWpQjlf+oUdr4DtOyQlelOZYdu4+oarhpRjTeYfslm+5k
boN02k0NyyNqq8fqQC39zZbnBJzzqE2irdcarljsSsvEKx01q1Itvj11sEaMWN/N
+qtRbaR6LDTNM5o07uxK08Si+wdunzN3pg2QgBmecpkuXKb8bfH2ZmZIHQfe7aw7
UxMDiZeotc+KR2FfGg0NeuIZMXyEM+dfgjAdLkpnxbVduLfX8Hrwg+V7p5UajyVx
Nu17bANuiF0PpYWiI9SjWcKVoSHjKL968xcG5SmLy/fWGBtzjiyObCh1Bwz/EvJn
cusW0M5ALDqnH3yYhMNd+RuuEG1HC/sj4vOeh5aycp4i6L2Qe6nW3+GgQT+5DKmP
T5joHAQ4G9HWCfitbUQXNsBPGMOFVeU3AzUX5UgiJQRts1ullG/W48GXmItf8e7M
RoPVkoo9h/f0XEv9ASmAD+OU7BQtF0CNwMt3tMMUIj32NMzkCGA7+FMC7ap1bwz3
VcSV12HaB9STVBzytAFBh3uhC++JYyE/R16zzKRaD+ZslPZWXMYVtg1SyPHMrXPm
pMNZia12GtpSvGblhwBRvSLg5DKgwT6ahl5FwbU26IgVXKGcKvvqaV2eiFmPm39F
7vslh6+UoUAKdHldp6+GW9F6sXCkAX+xmaK6ylwl26dGVhVYFIzBK1Yv2c+opo4i
4wtJOKGWkbyqC7JS/wW1tKcbajao2tVAnEnfC1v8w+L44t9+6yn5uFOnP0GSPJlO
MozwaV96jBjAWY7pEhMtz/mvQx3ra4BcxxbuftrqPN4Ky/4VSBJdFTXPQJqaJSq2
xKRgjXg9sYgY17RePKe7qAaqipS+S3n57B5+zjDwtu0o0BTS8HUGGpPcdzu83YtP
18pyFqvtAs4dr/RuAHiRQoA1G0QaThGWJia2Azt4Cqcm+upnk+jldGODYvpTEPJz
bZK678JZ+x/cPeUX9AfJGt+JG7TprjpFQGa7yBS0pT08iR4htyY6Y67Gnwt9y4e+
nXNBgtTlydXM70cE1G9DZdYClt3DAT1qShJPUmTeU9GFCvf0nBzuD4S8+IajWJga
5Aw+JrG2BLAEZPf3fouj66w5eNp/xWZYisIcE5l//CmO+6FtyrK2bqPFV/Pcw9XZ
CsiYAfyOeQtF7DsG2WtTRrVHPrwNSJcyQiFcEp51IkP52JdGPa2ZhqY0gx5pHGL+
XwbbFRwzbf0KBEBIclDfV7+oDpuc8yrJx1LkodPF5fsVJRmaSB1dGrA3NUDWFahR
kO1D/8g0VjrhsbDhpZTRKULLfRevkOfmbadA7wDYqEnc1xk3vrJ4NHdAHV2nVOEf
eIQIOZT2HXMmxmmch6SCeGk7yULpZOR+/7WHEHErPQmCqe3e5/CqrY0VSbC2+4Cp
eGlvVQnVV6fgJNs9rcK+cbKay/CrDs+b7xSGxLAq9ZorGsCsJ4Bmef/nirZVX3yU
j9Wr1WMSZ5ty42xhECJazwknvz1plBR7mqZzrsF3i6bGKhhp2jsixtRge1kPx70d
WKv6jMC3+QEZhpHK47YMrMDABQRnav0hQNumpx02zWQiO0ztGZcnfsJxLCjDCOBp
i6zEe60WLxGfzCqBW9o7aNnMVwwrCApcn5TgRoFsiibwrP80/iZHqbNcOF8adDcD
bsRyYbdewEm1dVPJedsEwU3gVO602ufL1EzquSTnarXpAN+ieurem0ZnIuc3jPbj
z8uMVebOnppWcgnl2y2L3oFVLwnBPKfwkRWDQddLEn/vsBMkt4P2YPnjDpmshXoN
eeFFgB7pDOfNQ2uh5SUNc4IEuJmfmr65K1Fjec71AiZrNpym509gpnDup9dz5O2n
Y/IRFO7n/7abEzhJncPGx7Gm1m2ZjK8bvdz+ClcDL0RZ59Stp29gMVlU3ptis6Fw
pdgcseuiUbq2NLJktWim8ByYjD7N7JUwet+aelXKgtKRNke+mJ2Hci7Q8LA6PDVD
6dmBj9hYiYIWLgIVW8XM55cbA6t5B3nT1TTbDkrO+c9uF+uBoXN19n3CpRT2rJ7N
idsPr+VWEe7f74vJ92qlvAMNJRZndKu+4vRFnM5DuxwgR/FfuSxq7wtgjEC3E4I6
afw14iHx1XPjcajfQoSvMOOv5a8yj0UGII69dU5XDq8YcsglDEys0RiC1k5C32PH
ZOyEbKqvQMyAbovaPwLeg42qF0154Hr8TaiTg7JuDAIDN24q8Poqr/GEQeGtcILZ
TvEdIU8d1aeByLbnaRhB2qx824kkUHhDfbGOq1NjJC8KR2LBRbpsbtPKAEQDvkPL
wSlQvviT1e2P1WK6y0m/hhQ6ibgzOKmjO+IW1J4OhQc0HXglw5ly/7J7FLOLf9kp
fdf7N0wd0uxW2aQzVXiYTG+gr+gXylzllZ4ShLjsq/xyo4Po5/mM5kDkRz9AGE9Q
mAz7BW1H7WNgrQetbFXNEIx3r1l4boGyGQOBoiNsyyr41PUYj/+DoxaaKfLZyBrc
nnWZJ5rLexl9BZBBwy4t2Fd8wDwZl9aK3b0AOF3jlyTTlgGQBBMp1d/FJDAdvI9O
NQ4sesEgek3xgo3HsVNuHA9pOqzsKycO9DiqIuAQTTihqmJuwlrVzRHcsd7XQmlE
gstscaBWwzBhWBSP0MXqMRTVu00pLSzDGvgqer9vjfdPIYDV2dy/qoJLNPGFTur3
9zMJL166QWK4JdTavCXLS/riLyjeixlZkBJajVPNTwwzOGH3MTCx3NpjRlUIeunG
eFL8bjTpq+Dad2HXvJRFjj442sUwILgEeIP74NBxxlXl62xnpk9uIDtRj2+a6UJY
FS5m9hIK3PyNDGUFt6ms7Lms7ye2JC0Y8pNb2Or0qUJL53bp4oz0xZpY0FFxGxJi
aELkr45bkq+DjO5Y2V04XN8LBuvZrPh0VNVonaE0lJcrLmSyBpYEHfeXPVLGHdO2
Gc+fYftTmsTrtC+sH6R0aBgcoUWnNPXPic/LqffV8mOie8HR12MOWy/JdpQWgndQ
Tu0y//V4N8NwEz0EXpzu7O0ntmY6ZbPtpmkq9CrtIFSLMolws6RD5TuQAAxewsDv
SLMmWrfL2/6CLISGQWAgdhfxeTUw2iaC+PB8TY9EpgqT6NTRzHd9SoR0wiH08ntJ
n+p/CNt0ciL03SSZ9s0lTX7/xlnw+p1aWz77+8+FH0BtUshTV4RTLwf6A1kk5q/l
Khm8/cU9UPtQT7BQ9+ZK1WURj5UFVlB0PYPkBoQQ138gSSuEvfZa/oonG8CKCcm5
zym2IPtokux2Y8YY3kcEjb1cdBKwDF9xAeQEVjpf8QMzROndlXyacH5tRHKBnrmW
NFKRejuMVW+CqQEbrYT3Fur+M6ty3+aY68EUwFGSzbt2k0sSyMuTdLJSIg6LMOjl
iTtfkWxBlzbGGiBR6ssW8uXdqXV5jlW2NDgVEEy67WBuoGDD39vB9LsScA4m2EN4
+1R5x4wcyBKK8bcqJZp04/dzyVDlAavUrMcIixK34nnytoZlsI57FqnH9uSKhypw
LtLqsdtqQKQ2S0DHYbg2oRDv4f8ZbTsB06AtBg9YMktoqBqF0BmV0j2nM5b+loC9
jWvqC7k24wd5e3SAaM2+S8G+8PMZWmFSLy+1PciKBG79qksoctsjVeFR/+qAzsil
GapnvmYBhXKzDXfrIgtP74oyXe3Fc0lw9jLsyv35P4rfKpcawoo3g5MiDtcCaVIk
WY46Wq7In8BwW8Hmb3iLeNk9cLoPaXo9T8fTUtViJVjdQl6vgINdu2r+0KUxiahv
gYzYlZj5UbflpcFxw/P53mn33adg0aC1SyWHL9yKaBJU460+F0LfxRU0tYfag/gD
/lNlLeV5mc/C9+gGH9B7FvB+x1UPzB8kk06HPgMNX6TZmMyB5ObdTJArS6ZxyuPI
Lu1wdX4KpYHRQHRpM+jhFZisOsGr6hrL8tsNrDMFz8zCjPRQa3cdLMpkoLtUvluF
JGPO5IWQZBF3mMIhpLrKetktQBjXbDVZWSOneYLu7NYg4Pp3wsTmEw8NE9dQ1o+a
NkxJf3fKPaCHt9E96dIjoLh7lAjeToSLmfOIuW3v3B2aynm6k66zIbwV5CTvzqPS
GSF6lzPOcsvFdW43CuAe9iG5XDo9mjJmnCdHTnI7MsBS4rOXz9DefcYMzeP0Y7Wh
ujZGaMper0bs6OhGTStXsFzAzjolSV9te+XPc8yRinKE8E2KN8JI0ICPl5lGkU7k
SLozjPnp74FNXrG/kRweLdimquvwJB3guBiZsj5hxbe2lCUl82IrJersPxLWse9w
OHbqUdBNXy5bWJSvYRuY371i3pR+Ra3a4bj2KQCGqRQi1eRq8xqUohU6tH6H0ooc
FfDJWK4KrSbTFPwrLMX5s8uxlYknK8SvUz7vghxSYKqcTS3C/gTR5uWyv/+J6/kk
Nga4hcRZupNAzjiaxm+h0r6VAvnVHLdWpiY7PoIp0xdj1sCSMU7AZfa1z7Ho5Xll
e88DutGZ104j0OTUMOJ84hKwEH4bVr5pLIeAIp7I89q3l4SBDbVV5kQo6K5atYaI
j2x/BJcFrc7DcWQJ0YBu2OXAIttey2h7zBeZQXtRPH92F1C4PGgWYpIZMHXDIv82
2WvA/q8G3eHd9ceINW7tYX9N/6aw8kzP1S1kzHdiQucS3czdZ4Y8rUHypQ+syq3B
NYdArwQ/LBaBAMHooshPaGX2PbV6xOl9/kBuTsId/OOsA30zcFWkukFHcg5yOdXF
/YlkXtPDOAZexzO+CaRWkriplIWop8LqoRkiatUbeUnWTHXVr0RLZ0+2QZU7ECR+
nvgPZlZsBx77FbN6obtCfdIaby720nrBqpLd+nk86a6JdD3GCzjmh52f22itl/92
L/nivKR0WXR5/PBnfiKAvrsDxRiAWRs6Cv8w7fBJ6g4rSbow0WKX9gXVPyW/d7Y7
hTwQ1y4rsVVGbYNPJ8a8TqEl0tMbW6PFzkSWI0Zbw9iJp8GpU3t41scQWgaSv7p1
hGkAVB4rJ6QX7Y/YYJQ7tkOitTvMTU8lIDeRfRAS6qbQiwZGROgET9GGFep2m3jr
MNKM7zSh5977DvMLkLOoO8eCgab3mBm3yH+5p0bH2fzwHJCDj4hsj96WJKIo2Vle
apVjXC/9kKZFNTXEvvlJzBz1JvSPMiVaeN1Oyl/gHLgPhWjIYKntotGn8M8TfX17
Pfyspyt/+c9t6jQBrVpdhByCgWc8vaLmb4Dcaax57oclDh7j4bupjAnD9OHpbkDt
ozj6ypMxDucZop0PixZTinYtDvNAOfAbTamvZeGA72DS444NsfvX8N75y3f51ssy
oQ3nslCn2llbvEwKAEyrOtsjRPsJKXTTgqGx+3CLgzOmY8n6FzP+H9a4Imf9D74a
51OWzLAF5GjCiyfgJHHP2tXukgjwmtEMFqrNXaIvFrbUmpbuDmKdtUDjkT5m7+j8
iGw3Iuw+wYIUAgfO5TU4XvQ4RaH8BVnKRgmgU/KZMo/5UbnGlEPipJ4arMMhJM3K
iKQKifxA7+xTqiNTxczPbRd558jOis9Y5opCwhL7mo+AArpYtutE2GNCwy+XZhFA
NRq/L1MaJezm6qsjAGf/+Q7xaLgP5q0JFo5rNUvpI4q4IQ22ACuzakg5Pc3kKASu
CCZR2qq1GwbQmjc8QBSMCX1j98ztZ+Cm8vyph176nOmY/aMEJVB342tf16gVtrqX
jQxJzCRC5vVVYkwEd4YTEt8N0IkjFXRTeD0ADXBFqxw37sjswyq9THnsJkFsvAJ2
YVVQllyNoTvc4sqrn94BYCKHNu+OlIx0pj27yW4BAkU5qaPWW98IwNmgwvkAV3L0
+trQuJkCGw1ymbDPGGHnpqK2RjiN7J0VQ0pQ/bU7fDHCzvJUdrmzgg6sdFhdg94o
uteWJtt9nNSjlohuzWKrV4LGYSzhFyiETMcoVTrNTdbefbB0WsXDxhE3w2CgiqdW
XOiF1hOsS/lz4yQGBTNVL+d+Ru9Uh6oos8ThqO1+ZpiXlRSO1SwX29gTIVmy68OW
r3G3hcwKqXP8178v2ZfKtsolqQA/4RCTh5TUC4G5J+rgd+oJRnFi+x7F70ZGfC79
Be4/LQV40NdGN1bcmg5mt1OYVm5t6rdzjds8TuiGA1PgeHYZ0ICGACkb5bglaf43
johpFie/DxY9RSd9Z9u9g7u4+47iJD2+g7KF6CL9QaI3oxnPB32BpoluiR3nIq5E
favHrSZ4fm0MX7k5M7ivfeDJi2IjtfWvPKXM5QepEYqkZJfDd8fjMlY0UrJ2cIcx
WwOyHoWey4jH7snsizdWCguxt8+UvNMvcM9hq+VGPf+i4bmx+BzDYmDl+Z3PuYVs
q7bEJAt66s0VtyAfoF6Q4PfhMgyu81fCfpZqeZqUx3677M1nF9Hjxd3A2jHM78EP
pOyzFYTUPYJ1z/RUW4SMN4JF7GnuLeON1VhzTWIaRzTLHX9sec93p4vv02ArjJzi
0lvHJLGiMKNL4wVVPpkBxOLK5qlBnbLU2XzbbF/04AqFZ2OFVJ2i1xLC/z9AI42C
P6g2KYKoKkhp8NLlrrtmGjJSJHrotGR53YOYOw+zIrWn6mjs74kfH1eoSMsGsHAP
0PIwkN8yJiOV4Inzl2zPCA8akdNfzJawDKPhK04yhVpXlHN9CY7vnQuG5om6qr2K
5zBZ/FY3ZzGkdt22DVwEGUhmYYqwIR4/Ftq6F9SiIw7jdxbovXwXz3bo4VqeKHlL
GFiGjjezlt/2Eoqj8IQUkWTX4d6DMobHbH19hXOdL6JMnVFul6qyd212pKL6Caos
3aNtElPeWhP3CNd+06YjbW8OAVLIWlp1X1fTeZhqj1LOuuqGGw+DzVR755jmKspQ
qUBbtecewHuadRGJtslMiM8PNOBsNCRhjOZEfP1KmQc9K8wXGzJJmQzZdHCLIu3V
JUr5Ah/lMSoPE9RdMNGoMztKHOrf0SgaFkUBph+aZZ7y/eTZsKKviP7lS38Xlhaj
HUC1raxaIDWT8NTJFWZbXi6UnJNiymNlG3TXFfky/j2sRMm4X7/tEK6HXLyTCDXQ
oABzxJF4vpI5O1kwz4bGxic6kjM+VmEr8Du8rZv1PxWWFX/uu5pQ27BOYA+HgK1p
QS3ifg77K7TIH/6hGrg4OPshszpjNw6fB9YE3TKsMqzEsX4TpMX8mkos1gv0ce9G
/YWf66/9B9uR9KfTvqBOqnJ3PIzH3yX0fP81hYg14/2OxB/ROowU/op1Ak4TqMF6
RyW8DKMw3AQnfF74jGbjEyARdxR9gWPIbg3KRYRx/YepSSduy3xkizQpiQcKP7ya
yYX+9DA8QPTi7Qaf38S05bhXSdZwfPVUgNnBSBFOqNTBM0fcFZSrTf5KwbJIwK4a
QZk5Y/lZaYxMNHtun7EsDnv4MHr/IFLUv9zbbvS+wcUoeR8FC0nRtt8RgzWVRWN+
180BSoAkpvxMk39X/cstM5naoRCzLdUZ/Y512R05QDLQn0iellOkka1cx58GD68b
7r8UlEtI9G/VlTNLKr5WOkUtsp6YAuLgI8Iik/zCNcOHWLbMQo2HGGOcTMnR/O99
sVgcmSwpmwyYcqxsuFwdx8CjkJz8LUSkBe8isr/SrudYT4/TXzMsUpRebemDvEtp
bJAFY/tq/cBlNcMpPg3lpOkXlhc8KAZVRiABYMhffoE6DpEmCRU0RvGhlzc96UOD
iCfMWRS24jMoXoZThVFvuIKPHbiaCYSGp9BD+XTDAPrOxdQmUdsSrDIRtcGJCX1s
lyYNimj5LwoIR4bCV2NY9C+0HsUZi8JQxstFJNFaMEwZ0010jaLUM4EKn6N48On2
DiUrKzoRKCRB9nOjUZPHDeKe5KLDb+TjcWqm/tXdORkvN2FiDTxfW63vAE2S5x8O
uoVdYAXEbsS1peU6/Uy5gJpDg7X3N+8pbQaK9JqnoptvrshXIuFYLt2bH+63ohNG
4iGAf9kIEk9I3xe7Sp5/JjBgh9EzXlbkrc2/XZ2S9DamSTiQHsmQbRZNDi8Eh7L6
H146yI7nxspWkd3dgMKhw3TZC8wMN33Vg6eLjzXdV0x5D2/mIz9BcOSI8fXfGJp9
gYOQ0cVLtdjABKJ7yzz++DR3ZJWV0E95fT3he9TH6nQqAC0ity1jqEbR5nVnOfDE
JBldhk2Drv3Xt9BwKPRgTSf/i1WuylqG1pvuRyPC4uD+XlcOh9roj2F3R+BmP6u0
+tegz8ntspGXl8JfL2W9Pamydegua1PFaXYAcgVfhdxuYQzw39cTVC0zMJk9n9Wf
dn6yD7VonEMkLk/JK0E4Zx1Mq2dDDGc7KJsqJuE252mAJgPqUHECs+jN8amW2uIw
7i8ShAVGVVUJSquPWvjFGdCsBH32f9x0pehU6BZ7fA3/Do+ixJ6GnadLH30kaDZZ
d74yK/cmsa6aJdDYiLDLmFW5FkqUfiP9XjkQHGxR4Fc351oerNoUnsGzl3TkugNh
2MK+9cQ/idYvCwRPOywXPStaYEm39v+/9n7UfHPG+BM4hRP6ZusAHh58u7ag6FcM
3iWFDfgVSNnZJv6XGtd6eGdGdlb1TfA5rwgDU1AejoQYOHrZTHdm4lyhFo+mUwha
V7GYUD2PkxYzlNK8BvO57ZncQUBfUbFwGvRFkN5EzNclLPI8n9gNcEsJlyb0Nfbv
lLRL+7GLPEO1k603kj3IOmte4EwAHN7xZg++Tzisks9rJkJi+oL6WV5ADYRCw+su
gsiI6h/QgjDzEjWsdWGF00dlkGeok+xs3GWEb2Bpyy0C2wbl/5lI44Plqz8oED7j
lpVm/Rp++TFG/6+/T517taPhM+oVrnyMM0YOrt65fnN87kD2P7GuuYAQ1p37ShPp
UYAqseImBv9i91AgFDFvZKK9URFKuK8ObiyW1F1D4JD1m8VVFq3SLIgMh1pCBwSF
DS4KAvVMXEWGc7OZ8BFpvopMVo/H4twj3h6VUOPphK19+mBJVJOXiLkMQeTFhlNH
6Nv7Fd5uyvx2s974hYJB7S5P7XwaSNKSEag/gFYA107MEkUjQM5dE1K7O7t7CgKa
UGYirWc9nGrckIBgoISeD7+m8TkYu8ec1DhEWmZmWMcC6Lgm+e7an+Hb5zPUkZf6
BNsZ+foIL/VUF2L2/U5iytJusGOCdO+V5BZ/TAkJ/3cDY5I/d1ZD02jQJB4Wndw7
6w7km+DDGjDZt4jaMgI86FeOfwMCOQ3BkiePKGOYWTL1Ene4iep5W7qI3EwsRmZv
wvrLD2g4l1x8L6qZuc0O1QTcwIpyzbCKxSWzl6MBYTH4aCg/Rvv/SFMJsxlufb7Q
L1dK0GGKsEb+BkXBtTwHQfrt/z3O3WuOfKdhm1aSjIY4z/HkKgcQWQ/qosTcnt8i
gtFy1347Clbg0oNGn6+meHvV/ynUdCydZ9gMsafgzvhGu8HlSfUj9zA14yqtyOXG
r8F2TBabNfXbnyKkSfjyFqqBBmxFlmFMwchMVnEyMx4SFykNIFHNTXBUUCWBZzlo
Ya/ZA0WAohVr9gNEMak5fpvMc0kAlLAFekOyRdTkIJLQwBUy6nUGyPL6zEMRD0ND
lvxXTDeH1giGV7gnZ+EvNSglBAyxNmoZJTASpibCI5w5ZinLWUcJemtpMnCA9mb2
Pkv6Pe6DjB+GZr9f+N/dMOMv3fCoh2v2IkEWrf7QrwSqOIuBTUKl4E5knYijJ5Pe
2B6XRJpNZqRCKWW5fI4fkymRqhqxea43lx8em4KJBe5mMNdNs2JdpNhuggD0oYW5
8mbG6IqvRWGNLfsUfS740QX9Omg4y8NhEqk/pu1Ik5LWmZXSZNVsmVnqijm92vlk
eqlMfsuwisTzOCncSi1gnw7Pc7MD4IN8ybwsLhYUXTHEj2hIl9+ejuZ4IvtmvLSg
up/gARkTEOkf4CM7DbRYnfVknBFStCFTrPyplqxLLMVEltxUIkS3GWNZ4HUcutDJ
HjWqfpBNiw60sNFd/bEDjSXfbsgUHo44UvbHfqt3YGvv7jrOVVFIiEjDT8DPUnEH
q1kfVCh/+jjngubD5SHEsOLyVIpT9Zv9WTpyqDQRMGg43juTAG5J3yBROoh/ioP5
qKZNjuaMWPZNfZZTvNrSVEPrFWl2ckqk1wvhv9gBOcdSXkkVmAzUshSMN2KKKilb
RN8xIsQjbNZFzszI71aDg8NhRhcQRuuxQjEEVM0jWiYcFYWM88aAz1Ix7GpjI0om
xLzjQfv+kLVfqOG3z6Yny1XvtgLoKY61gGdA7hP7yjZpncbGexQ8KPRHs5sVxewS
OtBCuXBd7eKgaBdI96YWO4r/xLduuMTlUBao4vmIb1V0WpsM6fntezqqk0swjif4
BHpomCmAo9t2U3tAEyeUMpXwXJA/kjJRQ0QlXlYPnygynaYJyITeiz3U0V7tJ4lN
vtBkEU94ElHW6AG1A4hdbqVm6HnA5elGvl2SRMbdIvudEnplmK8YhaQA8WFYx1bA
P7hK1z7rNfrXX+p3wfmSfj/+QLQS6c7j00dZ6C2DMSPbJaGjQXv1iuZ4JjF9qSmf
K7Wb3Pkg8YdUwpjNhFbV2uaMArtUy8cm8YNArbN8IeVxLxyhLf5E7VRnlyPBl9LV
JOLNravYijk1vZjig4yqWH0hICFiCqN2UspBcDQl+mBiREtimeDS6YB3peSV83sf
cCW8PVMd1u+AZBUmIDSoKHG2QUAsn2G0jeEKHv8Ycw8eXuNElamFjQbhk/+BDVxS
vBar8aZ6FX15IHklcrO5gJ0q9r+4mAh62qGvQeob7vQpLgfXzFRX0OxTQwnMKaYH
+SMcrY32/O2msepU/b4Sb5hr0AeyT8zmU/zWmGratVF2Lod4g3qSKt3IScGYVQby
Un11jVj1e9W/j7jGYDgSXWIQ5LmNOQwgl2U4VbEGuBGtImIScMQ5lwTM9RGBgtJ1
q9pXL8RwoNkdImIZuymFikvJ2WWY2n1r8QS7yqs7JzfLLq7rHg4AgHzrehLWIAcx
5PTixKgZkvoxm6VYLow/09k5JRmKNHanYxQoRPU9C4hsR7II27Ll9kIxVgsoPRDv
rUsFSCxwy6pj6Hl3ep4E106RVFFE+rBFyd0pwnE0ll63nW/rVIAoGYmED7msrqGS
1RB69+2+QdpGRNgCJANsMXKwrx0FvuImX7Iunf/CEHiTboy++rgcYCW1F6M56dEa
ktJLN8Qdqo4dek+FQwzJaJgfsYGrqGDN/aInYCfYZy16q8NtO6qQGPYQedhmAjvP
O3x7AISoYoghIw9h92tl6gRGV6TSu9W6iMOmAAtdvVq1d4KQFiWPFjJPQlBuacG4
iH+ghkczgDv7GHNSc5Q2XlIyQKsa0cl9roW3TIPCXjyFH0XYIjMiBGmL+Bok6kbj
0a8DA/A3v1nAJT5M27fKcDQM/+iPeXZFXyFc36Rqi2XS3JmZDxLJN2jAaIW1JAPd
ExNQvqBlW7aaQGrL98vOqbKPdhMCjlRBd3jFw3Ht+L9OmWcz3iltphRINdbT5ppD
yfnrgN9BWYP/HcZXmJjxhzM65/9KucLqjNjxNIrGEUXVED1f98gBMVJCExrwjj7u
wSa7ycoKejiV07tmv3M68pi4UK5WVEJzE+GxVKKx1aE2Ph+AwE2QCXQA2LRdy7cU
EnQBR4R5URzKvV9eIJfeXM1h6tnQalJxUUxh0lngzQEnujwxvTM8Mxtnic3UmP6p
1756TONKL112m6LfV/DLiy3jbKAcU5nCG7/QVw2fKEYCw+VSIBb/Zg6LqYAFnQzr
W9BDW0uNFr8KvzZp1s1ntkwh9GVf3uStSlcCo5g/y5lBWW23BUJOiCobj4dpgk6d
rSIADncKPnOSuQ6DjshjHGcAN3inVguYrSI0cgqmqBeVIS2YBIkDl/gnVVhXRfGq
IHSZkIcqZxOLXxIZQyi23VDYLRDDr8/GYTI2LcKEM1I+IXm6+2S1dxjJRs7knv+1
GLx0V8XEpsVVEknERhJ2WQuy1zrsHtnVnziG/AJfr3QY8DRAgOitUQclrTrQ1tvV
HuE6ErdBYrun98jMTX/NmQ==
`protect end_protected