`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
ddtXksX2+yylW5zu6QL2Lhnb2d1sD00763mmSITNX595NcHTEkwn0zB1Dry37fOW
FufOhVzEJp80NC5qZ/+F0Vk7Ik02dIR0elf3clrjeJRK85K4e3Hoo4xn7YbFUIms
l/8VZSb14+JVGURjfswrIyCUotIzlzVYZ6gzoZwDXIi5gQIBf/gI+KxNXPaKV+PQ
Ufys/12rjO6aI/pPlqSm0hCvftmBcnezN2hk1UeXgOIuKZnogjOsf0iJVX2aOOWE
6pD/psybjbnsNB6kH5uFTA5frkzIzkzl5d9+YDm9OyC+k84E83I/7/j+rk4L2dah
QJOvksSIzN867/4Qt8qYTQ==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="MvBXkzurAa5VTw+1JJ70nePUfoQXBvZOku/SMmg4TwQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
oRtzZL4VJ4iwysPsC8SXYCzXS8Fw2gtZTOskLcDV+1B9Nzn1zTyNtlo6lNICRmmK
ZRVu2BmCc2G+fmzynYlNTnSa7C0Cuel6FYpxCBlOuk3OF2tzAmLAuDyOH3Z1Yjzk
a0aHuoCdIRKv7BrZCdALt03JeUmXKPdOmIlkVGFl8yw=
`protect rights_digest_method = "sha256"
`protect end_toolblock="Jn9CQpRhJt4rnzZPRk+dOpzAubz7omckX1MrFd4p81o="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 21040 )
`protect data_block
gD6l00tciPUa6pDNTk/+t0OO0nC/UTtBwLB41d4inuAUA3i/ALrNyoJVcBnAmEQW
ptbcNp5fxEUJjnOxnedyZEuEBxWRieZFQnkRdF269oNPyYAFw44nUwnNUpmeXltO
2rube8WDEW/nuYMVbq9pOkgZLnnLoWcAw2FwiOIDzWQrGuXdNxdXc0uRfy45oOGo
STzompN31hoxgssyQG9eIX+bZdcwY/WqclVNd2/1/EfFotPGga7sYzcattdkkFwG
/yy1UvK+qyue4l/Z89pL0AdWeGieJXKtkY8JEHx323g/G4WJcHSX+E3dnOr2UI+y
YGXQqsOtjBjCfros/LwrjZqPolUiKdZiA4dkDUvxpryd1G9skEJjnur5y0nXbtvZ
LBOQlIQEHdkF6wCwFsxalpLWlvIr7N3GO/wSEY59+AbfxGsIfWs8vo7dpoTFLeZw
DE2y2Ctnmv7avbtLoZRUvTjUZgAeuyeimH2oLSTwnXmrhwuLapl/9WoBmxwYOEeC
WwTsRIiihvZufUjnr2s866bKah7pyJCUyP4CuAVATfladI7F2IU4TnS6C99qBX8B
E2h0lHeY6TQ39M4dZGiMk2avJ9/xzVXr3KV+F48jXQFtP+ODhH0A7/LvZRcbeBHh
LKpmN5kN7sBg7SgdHaSVLFhuqKrouzuzbRQUDegWZTodd5IEBz/toRFDw4w1e6V6
pqZhNcTY/Ki3rcTM+zGESdy7iipGxaMtUoABl8lYcpLRQ35tXY/G0Cjy08FyZa1r
A0MBoA/wCXMgP1XJLM7o6S6r6G8gaQ0lFmQOOAsY4gQjeiTMGNQmNDovLgrWSAyZ
a6Nr2Vlrboe6Jv9zW3lkBL6tzhHiNgbdIK31W992Ga2cYS+N5cM/0fQD8BFjgAX7
AFkQ/jiumn1mSz0uqSe+4eQHYcr4RiZA3qhW6fqHnIiQcVWW/Abvci/sDXPSrBc8
cRe0qGxkr4UMg4N3etzb0s6gKQ9wdj1VGCru7Lk5mWtZUKJMdLR2EjH1+g/E4c3h
T2I1NABHH8LRbSG4Zy+3tMmQ99GbM/3CjzmZ+16yLAykX0ZCYLVRYlJW3WCyUK/j
EfUkX+eAhvN0jsQI2LfBh4bkc8Nu7FPF0jZg0c90B6o3bEnNjQv92wOy1wp/vokz
1A73C7bv84jtz4EXaApHFrbpfzHREgh+rWpJZXPISTFbkgBLWjXSu9xwMpbD7V4z
KmHGC870CPpFDWnH+VwwQyVH7i0jcWmymZUSHd3K+YgQFCWd4DWVrNlGaJ+70s62
5T5OXzkOxRAMk4+CmFJiWfN9cjp9Mcu4hYrtk221YYgKCiCHHFolOM6GUnJIkfuQ
dDP434YnRxZEuGCXV41Goi7JUuR3M8TTFvPAC8r6aJj4xweF35Ju0z4C6j9C+OXl
qTDsKR+RU3o+spsizgiLL9wDjeKpHN4F14WycbGjcDI0I4D/HRh+w8Izq/cGcIDI
qTgLsC+/1RCbE4JctOddW6WirZDeRq+KIaQjje/xExVSAJItfLOSQ+ewr70YTmgK
1oR0cK4694oZhQK3sWRotBPp8IKZRwCzslCZxrzuqFBGnRo8o7N3YoPBp8yLjC7u
2FLQ2dvrd8Eg5IosDqtQICnvGnRHJ9+cTPHmVzaKNuMfAO8j+CGmAuRZTXe4XQ9w
XNQqj212KaMACt1WFTiSWbivxttiC10T3wUehxuBNbgxg8hg4d+pFB++Xn/ydVYE
1lpKSECDxvLMk0d6VrdMeSnda3G8lV+e/YBaNiB1unyF4RaoltIEMkc2DxaAcngC
eKZE3o3a6w2pwKBuzAr2emTyQCO3IpD86vco7grMUMbHnq3sEXxIoDM3uOzoPmWn
lb3aXy4HZkZ0++ah5PJl1kakzFN60E604rvW2PM1xM2ctz3RXSGXFvRyhNtAJpBD
U8DoQ1V7FMxxjWEhlr4lA6qRed1MhNmMowj1v4ESqUxmYaLrOasijSpvBeuO/Kob
z6m0Nt3aQa94CaC2hkOpydwWCz76GaES7+tWz48/6shp8dM1I/vknzMvf8ATXl2p
2TTNs+V96IHFcR7eH+kFkmEcVEWnR5TQopG0qGDw3Q2I2Rzyvq8X+USGv2axA/Uu
a/RO0ol+XXT/bA1Msh8wfeC3Pdhx1iTNxA4jHzaiztQ6awGDG5/FMS/JVEyyOgYk
2T5tSoyGFOzyiFnyNbjIOimSML8m3W5U0vd7Hg7OH3L/ujDZ6qu0XGy9FHAskBil
0U5AqGG4ckF79EKlhmddFSS+pDMi4hhnJVdryf9PsGIaBum59gULAtTaJM/1x1VN
BS43RmZDn32e+CGeVP8kRSqJBsT8z/pV/xFWbQrKQkZ/zCpv2GZqri1R//GVCuk/
g6Pqy3sgRZs4ZHcv8+nfQxtp3G5g14Gx/UQHKIS3y+jxDPMBoSWm9rMlrf6yAu69
r91RSblcrp3ZU/PHcxcysNxURq+hFxISaoeNI0urcZU88CmQ/M4S6YyoCxLcsByh
5rShfQAPh41kv5aAOne2PVRKJeBcnIZPoF0xkioXJ13cbQ9wjYYU2iacHMkJXm8Q
HKqdgKNZXZ1+mwT8hHpXZaIAv8MTZNthA8jV0D+shqT88Hlua6tCwO9tV0mnFnsc
Z+V34shEeaJoX4JogS/3jITKX22yQNlQZIqEt+kJA1iVWbMoIqG5/vP1BS56p5du
MdBQyaiU5K9mIE2bCD9pF6TBlJRBMkdMTvV4EEj7nqClSgI60bynhG8KQbo6+HNN
k98PJGQXN9auTPiDXyl3JSScTv6SQPhVYOP033FcfZRJBKsZ/PadsL4sJldI/IHi
ZW+AOzWZ4ECngDuv5bgT+0V8ZPP8J/S81iGEtIdzjN92RKlkKVH1hf3IK/FTEACl
lmP4mD7Qsc0B/sfVAS/sl50yABMR7vPuKjw0L/GsDkthEJOWnrUXv3wpm0ci7er2
pm69oOwjD+C4bP4jTOGDiK1Spe1V6vjUyQ0aEz8jghytvab2olQuDcDi8Gw30e5F
molObT8VWIEjpHr+qn2S0FUE4QGmHzVecEu7v5xqgG/bV2Ij8oorcgBBzKTWAVLw
Xm8Xhtjjn7wNMUPSh+4dZl2LK4RFQrWDk9BKYWnqiUgymjcUAobnW+RoywzSC/j6
Wt1URFs/gurQc0GI+SqDMr9loKGYQSL15zOMNKqSa835CVth16X/lip61IUGX6ub
fONIoQ4BQiC3mzq+YtU+lBOdr7/9u/qHdkhVh5NVZ2sZupZRTsQdkeLo/4lrRChS
gq4Lq5m28eMvo1QEoDfvGR5pNwcy6jUwtMzy6c16G8kAuE+fGJCsVhumk4YbLKmQ
n5aDTDkC6/6sLEQDbNlJFICD1hVOTe7DcNmK/vl9SO1QxpTJBTDBrBW/G7RLwmgC
N0lUfpf7uvGQWtJIZUeo77skhe0MupLv/Ptm09Nb6wAFJkcQShFRvifrP/NX3JrI
gCXpsEycKaMRvpJ/i+TmIW4qN5fxX5gyDWpQb8YWEitrGx1Xqict7y0fIViR6D3O
TGzyUeNLF6RnQgJubXMk1aqeMBDrh8vWTL6SS9InYJ/Nb0cC2wi/6FCevMiMLqv6
3pHS4YNHufpn3hZOw4pFRKsXCGm5cngEnX48UP43lLTdAqd9Dv5DTgZkHTX62mH4
hY9y/12mO/6VAbV5s3QaugaiGzfqAAlH/KjOv92xzXap/hHhX5zdic3/kVSWYkcS
5csqI+Ov4l+FLmxzSWa0Bt8HjRvhFQ6V3Jzhdvbh/jhNmzCB+/Z1vRBBsSgwPYjf
LUp/HRJ9BSjgd+/AXW6i18ZY6AgD4rLIcFg3KwRc8EbHgjYlcRwVY35b/sxMKF4W
Ps56ILhrlimT3CG425SFixin7u6MQRUtxmsgTOKxFUCxw0v46Cg98oMKal8KWyTY
SEJNRUMI2TPq90LhrxsRN1Ei6X9f0cww8DP/58cvsCJQnT/PtejkLlpyoyzxnk4d
wuhtjCVgHQxbg/8Xcnk27jMRcvKA1Iu/sIgEjz9YH/QYOc8NTLjYFCQUtbjAz+Te
l0aNBC7ES1FYfm4QlAf5Djx+IklfWa3kziYl+PZz//+tKf6Ql1fU6rOx3Es0yzMS
Xeq4zhRwJUakej6cje47G3IFT99aCWOL68IJ8Vl+ZoEH+MlaI+kUoKKYARly1TmB
a5Liq/O8XVjQMGzxik5UdK17QjoV23td85SFWmcqQQI+5kbIpD3eN01BzY6ymo5l
yS58n47gUUIX6HkqmLUdHg1oZDtMbPj7KB2bRnfBOzCQIUf2aCpIYi+xod/JUbOi
iitrfeS3GTJQnwhRH14llZll68wWIFh+xqEJi0zw4InDVCH5u022JDRn4pOmaMLs
BGp6KoF7ZxeApd1kmg2Kxfff5g03mBuyvKj7pWHo+xpIig1v/Hd22aFRWzJ04lD7
eEnzEsSHjOnlmawv5RpqL+BpQsQIxazReaig9j6O4XSlABXziDKjwPzsdHsVmrpq
/VnNCNsmW5cey+643j/yY6OnLUQdx+3o2yyxS3KwPSMVD8tqcqJnPh5RrJFveqxY
2IiD78v/HzVLApLfyFpJfHx7OszCNTs5yFy1JV3kaqpfw0JUc/fu5wHHvOjb8pM6
tfTfw4Dk3pjDXJ5ym55mBDrJoGKELZA2l3V3Eeq3keqe0+UHLtrw7ukSwXhwv9tw
XFCmRH8ni9VmUE4oovV/LC3TdXnkXahFyoPZP16wcnMAqVNYh9jW4nl9unlb8nit
0sbEvV9gdxuTdL3LeTWSjRq0/nfXYMKdvMdOmDttlNatUZ/JL58uUMUmS+WE2sMT
30DWNPUTlCU6Uy2tLDH2FWZbcNaiLVYmvTyTefejuhTEY8dv4D9cTN+6w1rInDXc
aKYfQVXJiInUIre7zYeHUBOf7AimWW/8+sovyDEzpaHDDvpbsQtMwVLLRKvDs8H1
In2nL9neYoSjZWUNZpqABBCUjnAQw6gdTGNU6SCWFEFrgKlVYPtNuDbH6/HWdt27
Q0QSCGGxphqdaJhWJjWnCmpFcKooBH+eIby9j/+RmdUm9/sLrgTkHTFJY4A5lCoj
7w0HmKGp9j+os5bb3WB8748k1AHFxyjaIIbirbEKuiLWevBvHxQO77ZXH27z8IjZ
Wu+3kcX/RIGmfY6BcLMzzaYLQ2egDzs6fti56LymqfZ7QwwBN5I9auKwoEqAIAAa
wj3lAoBZgF5dfsSIDWQRqbN6m4lhfjHeEP/mR2lMnBliInGDg0yIEQhpqs2sdqTc
rq4BRiV83tzYTQVg3x5jGZ1+maSj07IeQVyPgdu7154UcpBfcVZs4zq0EPY8+cvW
KTY2YLlJ+nGXCIT0QSihMzhc+ovX2l05Nteekq0adNEhmTTeES55Yoo/I3Dt87uz
bdZzMZVU5qEKXzdOX4zSTy7HTkDhESb5NjWSHDbVM+7/2UziegFvPFPJ8yh1RARl
4z2bcL8BlH/A7ri0hJCSSPAPJy4Lz8EULQAsEQcvk6e+4D+lJFvIvvb6KQYIM0u5
YTyCY8kImUJN2kQSHyAMd1nxgL4q4Zfhh6z2MEcgEVMVX+VXcJznK53g1bWYJsOT
zEDW8V3utMjRwkKQScldzDxwzoMGYxQCSxnUGCm1w/8vsL7Fv+IGUTXMWAvz3d1y
lpeEVx3peYGr2aLeO99ETmeGPPGv/3Q1gTRtZFOWXBk3kktxr44VZcrQQ5TkR0jK
fnLYkWybcHMwi18uHhtwnQ/PGpLVADuT1DmlDwZsIKalrT+JDRuY8issRIHD96yG
BfG/Lu0eUOcT37FeT5Xw2igC3Lhke2KGhcObHSpdP9CRA0Ej5mcLG3E1ZNPCqqLH
9tA6Ofoq2gbX/YvdzkZRHc3ExuwfOlmsJtf9r1DmHT2iSeajGbhnI3axvOpN6tsK
boFJFwVfWoa5VLJcoYuUcQ4RWVfRE4kJmgqyTzWBl0VzWyv/7yWcNtgtiRJhCXyw
6wj9AAqIjaTlQ/5pW228fJqT293rgr/G5dqpdHY6bULpt0DdGSYzYFjFK/VI3CW/
2f7mx5whxdeajZkZZjVLxF9OSr/3uhd8uz1O5ZCkQjrgaGFxxo3YhU9CxW45Kxp+
hIRp3BTSJ+51TcIaamAPWNz4AXtKu7p17mo+qNCX6uLmqqx7OeBNdEyyqX8gUwLs
4lWxOLuwoBuhZiweeRNV+564MLofMH8kU/t7mvWgO3sycH3QV2fw2rcHAf/xcH10
DydRV+VydpyN5dj1A1aqG3t9/vQsv+sXsuiubzr6y3ziFLOKBPKtYBcAsNpvH19+
McI60xoUn25dV0LQZFaWvsJgBBvmbU6wCPwIiAKrlfNXI2smsDxgDHOO7RT87XI5
s2PCYTlw7Wzeh6Abymt+CCjPc3mmE8xuO5qrpbmjNi7GcolAInYzMyERjtEb7iKv
iW2KsRK+E8IcczrhmtOZEQsDuzclzzhlrC56Rdd6FOPkQy4UFqDTTGI9BYID6v4c
DRRdX1UfoVpFLs5/qmzlZfEZm9tQU1Az4S0sW6rL1p1D/gfgw1b7VFqht8RXfMbf
zwf1SkxYdXCPgj/zqjyV3ccvOVNEuBLiOpXtDoCkfAV8k5sUmX7IPN74VSSFaoSu
81aBw+Eam+xNI+1jqBtbhpxxp/Ya/Tm/RMycpprTaXe2NXLRgR7JKiqjqUQMxBLI
v/oQakuG4WhMYddTY5b/xchQ2LGGfYBrpdqLZgBNrMxHNqedBnY7jseuQTXYJU1j
zZgmmSQ+ZPdXnDxllCld5mqBiFL4YM2Tu45iTbfDj3pV8SLebxDDg0dgzrpLNDpQ
J27MWHCO1O2cfcXLZi1M5+7JNWETp+XkU8K/OGtnpXTiujxkwhwKic8851gQrCm8
zCRB/7pto1PZXYAeX4iDKASBimMbsj43rU9cGUlxJBRh+xhN0Fls3ov0V2nczjK/
qIhRVuiIm9WVyjGBx5ZZ9EWOPdS5lIH7MoFZs+tb6zPaggCXN84rKCSV1nzM5arg
2kCtjgO3ZC3etMU1wj7EHgix+WZ5yYa9EEYxp35UwoIA6hOXc2l5CkxyMjKYpnfE
S6KHxB1E9eh2TBo95kMoTyQzE73nC4BWmJGGVgXuxiKnUMWw8ppFjA1Aip/5pyQF
HPrHaXq3jBEKToyqLrsd/BHy/+tjbHSGaqYbdLcnJfaF5E9Es8lrXmjTY9RDhaXr
9nca7yR9D39MJ4XYYizJxh0S/ecWCJmqPBJOd4bYipNPpfVO+2ChZpigexSoSuu8
Gxt8AXLCmPJpWsZIOGeNMn3+q0IeIrPK35pkzhO/8fK8otschkZacsYkOrezBnUU
bwTteHOwwiV9eyxMJkalRnCbI9X3KJCPNjVXaVicbUcU0uk4wh4uas4YqmbxqLYD
dTSJoc0+6aH7RM2+L51nFimCQQhhCIJBNkmVKpdtyTa+D9+xWnzXyxdYv2RDGKNM
UDydNJkzgyuQMlxZ2Q08GpbVh59CWOXEZQvC2Fr1UGbP4daJKn2jDmzUduZbYy/+
mPl41vNGyzwHGQCKVf8x8Tr8DDYvTfr5Xe+2vi4F8tHcLBHxAJWXga+MNR3s07Pz
MfoT7Xa20rlyNXaCVFxg4v3KwwyLqKIgAAJ/vWQT4z8RfNA3hTKDQJa1exT3tkKs
52hcMe7TMUbryzjwKtU4YPnqfr1litMyNOxOvLffFimK02wfUX64+F3OXti/0s6x
dhzWDdvnaNC/jaNH0gN5/bbZ1KO3PfSEI5DDinykwzauN8b3tmHup8eXahXYLVFH
EFraU7KaQrE4sNplEZW64sQEwBNxhdkTUQhcTMCtDockMmsvukHTWOT0Ebwugm9I
BaDpWqUO+u8tqN13p5gfbvI3MMIl+BOqy2IxOweaTrBDsjK9AuachNzYA2omzCuE
7ICpOqEYW07y4VbzwNr+4wiTPVxFhJc8v2uKSHUAN/hm41OKVBCCvoOZT9c4bmrz
h2quPE2I9fTA/5MokrOJ3Rdcb977EDTkn4VDun9QQgLfzJNODJODaqPFY+DZYd/A
uaOWphZRS+Y1w9n9azwGjWyp6bMOFVU1wYK89vfRkayHqH8KqcQj9X3S9EuOc0YM
l8U/0faHjcWa29Nhw0Gn1G6Go0ovQZCTeOktNHA5tgd0W1GoIOtM3vfCdRaQb20+
Mpkt5lFEiBPrZRgcJ36I49mAoYzL7U/3qhdZNEMemW0CkW3O/Hg36EtmWq/aX7QS
OpbZjYYH3wKDZ+skyzFBL0xW4ZVRfYmJwpBHyAjovvAYHkkxQTsBqaxSBPh+78gb
mC4Zvyceo7bXIW9afMbX3mG0MAuyxz+zoUdvBHrr+7M0tR/4pMUelsqbd2NBwuD7
VU59SKyCvQ+OB7Ua24UuZWunSHe7esubWDIJOLoqU/WGIgWyd6dA83a0VduONIZ6
dblfLD5uAKnTXNHgwsW9bH316nqQ0Y0IDyfe0zb+D9Z/1ODlQYg5leZctT29iL5T
zZLwCOxKjQx/V+hE1bkddBmUxnjJU4CTmDsrVHryj7lf4A2VrU7FVdZuROnKQUiv
IVLL+FTfCnlfsnPypJTjqwN4/bxOwEDghRQ1BGaGIYx4wh8nRi+9vuz8OmuQikgO
tTd4838n8zK+J4v2t/afbk3Lx1lj3S9mkfBH2NZG21nc3AY+u8AQGcP2M9ZrTjfU
5D+oZrGqClmPi2PTH8yJf2WTxmhg8bfxGLl5fYmaHl0cMplBxZUoqpnjk7B2uBFF
tF1OWNUuJwSLS18iXeHUFoQAwijnDcCoilVcj0lFqYczot/en+Xm9D/9qbgkP903
uXJTHW0fRPeX2WDK6gQmatOJokK6CS8YwzfFVaz7IGp8zTaLzFHuU+qN3Ud2Qjxx
8y86vW9hOJCQs9fsd/5EY52BbP4T9cnn6OmWdWtJOt/iJ+xtU4Jewx+XHHEKvTI0
clscy+YCL2CbOlj3FhdXaMKdIINWEPHs/QR2ynoHQWZvJIEI014djYexRct++v3R
W3rC2sCNsyWAff2O639iAjuUa1ptkwmnlIak8kMqu4ZDBmmVoCitqW2MireN2IEP
Uy0tIRmTV/Yzp/VkDZBtKG64HGes/vNaH67GQdouD4itU5Kh+H7MvMYsLycsmub5
eG1MMSw1gQ72o6Q1iE+ehY5HCsvVZ8bvBaT+snKeTshJw0T+YTa2K97apPAO3blG
2Q+Rd4eoHJejU/0m1ciuU0/x3hfS6OiReqpAyb9yD21a4GEI0XiXpf1sKP5UUcL1
zQm5HRCjVXntZlc9afJgFdIMUjXFap37B1qpFTdh4JReWsmihPLwGfnwXNuYBql3
BgARB2XUDzcrhEh4DcK7rxZeFDEjd+Zkbdg2DdYeI5qLnk3wIb5gXkcxJ96vb7b9
nDyJu0N/zSXtJmm7zusPJT9/EMd30hCHi+UpkoRp8ErGds//Bh7EPskQt1Q/pRmV
5b6QVt+8qU55dBxJRPbKmBk+ewPn94+KiSaVm4Qv/ZTEfP6wEDzAlYLx0JzVOUf+
gZPS6lWVKzWfaii4SM19XetWBPbWVnueZyOmML4W1lFLSNUXpfj4GV1r2UhN8K9o
iYRGi2XZGKHHF2sen5p7BdB7A34vlR+DX+cJ0VGM0BHskFQA6rT+kmLh8zegELUn
iXi11ew+TnQQUwroPp8DsKnahBaBJrhFTY27IFn9lJ/cr+rs1zoXTdq/YZ5un4YY
lgxnvAvwYJMMBRBSDxOkQYw9Udu+Rhz2W8QAICtdIcs0ZzvvGVSbR11pAHx00icj
+VXTBe4xKGFnDOsHPaU5zm1sJbqal0CJxyQAX8m0OF1FCcNydgQuPkL+0Xkh0v0C
GzSAIIr7jMqzQu/0g4dD4gzXP36spJoBwb0IBAfDoT8yo1S9fMxxs2hHuHcWjiU8
6hsFIXkBl4gl8Tns3a85Kw3XkmAqAsTnkutye9A8Cxeittjrl9u3pkx1/lP68CxP
saMQi0XW9dYIKO29aftNMI0rTp1pTP1WhCMbluxQBHCKIpIZ7U2f4GhreCOyfwtB
pUffPJgM8jZfIaLmUbhBdb57GjjhOozN8hcxsvbHrdZuZp5A4IpNUQJLRqa08DYY
0VJq1AJIjJZdDBJyiYDJZhVyGbTX8NWAdwuuy+25zQ57zwoM/AVMXhpKBVgtkmpm
RxGCQP4KQKlRr/cAkASxGBjEd7llJrxzvfTaQCGqMSLZ+SXBWHbXmGWLxny0wAVP
cZKFaxljbS9EdMK/N5YsmVEXhdM7SjeuOjr5pKbTHciYsM30g8Xvck36F/I76id3
izvIiY+9pDwG6RXduGdTbZ47U8xjs5hgx4rqxXjjVTTS7SEuCduIY9Y5L3WgZq1B
Y9MxBq04dj+Ij34w5wBdIWeqKROxFnN0PSUelYEx2Bwm4KJ/WvQu06KAS22uEUiV
lLHKVRP4CeneXDOsCYYB+KlqJOLesOUy68STXMxuvKGVS5n/S32L/bNOIoR7c4VF
4+qau5OKAm/NH6UuKJ7rfouWtFqKszHtASlRz5CeFxfL72lHQDAdc/uNtHKhf9dv
V6jPXu+aZKJP6AO9emZcNP+9e4FsAS71lIsdU+VK76ThzObDjeA2QSaDxG4pSrPo
XzKkV54TKeKx8Z6fsVmaLx3PifOsOliSeG4McjZqKJCIIUCwZZlPwHS5HV3H9MJr
2QuhVpq4IKhkVEkb6B3/pVj4bAeldecIfsqVN38j+PJi6Ckf+d8/jRR7osO/6YLy
3BENzOOHpmFkqKVPNgLM7fJlcYTm2/et00+RrP4U5D/MTi/iZKCe/tCWzZqSxLSo
7mFE/Yu/dkmfLTeoD4QxiRCytUEScs6U4gKpvTQNUtIP7nr3pPMU85DBhFZ3vQ6E
fz/x/rE5oB8+8dkqu/XKRCR5ZMDqtmpmKG3tU1YsdyqPUEVBuebspyQuv4QFcm+9
ZbzC5Hv4ACURqs4P6UHbOC3lbtFtuR4ouAMA0Xo297U1IUZm67rGtBCxJSjMKljo
GFcqY9zgeazZoNuqrc5p8twLJJKHVPyksNP/DyiRMF6HMgRZNA1jfdBERS6cCvhS
tRRk088HzM+9i2lqdjJUdjhk8gByEQbEblz+6CJhYYhdkQo0Vdo/jyx/faKfeC9E
eFB/nSWn898ZSfkEBlhQJbS+AheVx6Lt22aHOjO+Phl1Zkq0Ur0ZPdKGGkaP0SHA
nY2jAMUP1ROfult+De6Z1ca6K+MZhL/INGm3Y64U6ocoxYZK7vyYTP269vS6MCUn
4/Cg/TwmMmkA8MwfUV+skXSK3d1NzXs5T52rfw02WQj1iuP/E22l+QQTGXSxea8C
u3KvKsw1XISSchdKKrIIz40tp827gm2ePKjD9pVFoVygi4RIESpAVc9nitCa3w73
zR2eaH7EevhO66shO9cZRVqaVlaR40qc7cfNj71iFsQSoFI9bbhdeAnrlOAS4nd4
lDPZb3A88yikMs1phIheRWUhQ8dRtpieo5A1lvVo8XJ3SGMhKQppN7Os1YgJDXR8
XxZpvgjF0OraSvrLXj8/qvnA4mIoTL+8iX3ljk5vQFr+VHskL+B+ppHzbZOtOXBt
Tb2smicgM4M960d9M3QEGchtVd2TEqhzv8WbCynGkDm99014iSGF2c57IdHd+R7M
xXQ7IgVoR+0Yi7Vu/w3xGjKA8u2W70jGtvq1UoBr58UBgZxH7GaS1waIB5T4Aw5u
4/x7diA6l2JmZjKuH9uuX0YaBb8stXCpgJaSno/2B57gY6JI4tnkVW3l09EPh3BQ
Ja1Oe5dmIMDEC961z4RIGryxzjSR5FN1HFc16HmXj0t9v5B1fT+zwv8FevCR8p3s
l6/0EoEApPLNZZUr/6qGXAUgUxjOuwrbrZvxZuPka0n8/b5vPlZUUecKdtDhHWOS
glbBp+Rwe1T1CGW1rCuH+kCqAtOZwhc6vf2ItOCNZ29s2Ky9Xc0vfZNjRNuT25h+
FAQ5i2uz9ivZwpHqUnSzartNw6RnU+4K9w9nDa5IJoC3oWzoM3orEaYlU8gz47P+
ry+HDUaWKYC/QKgywJgPV70iS5tnyLVgw0ZP2Gin3My3R+6G6PKIVU4AhwoXISMr
0X3lwIKkXh3IkRe7tkauGzvyJm00sSppFHwHdMXOzDwgeoJhFzHHklib9J+6h7Vd
fR9TOoJriPwdThsAPsKvJrr/k3GiQ3nzNpbvnyl+TBfuwGuXOX4LMA7IxN2we0RL
EFguU0FKWPEUMXxCDfYbWE0CxnLm7OFuncRozlvaRl20x3izSehB2D/J8aVcL0QR
zvsb/yx3DYk/j4KyHxiotfplYID0XYyYCry8GHfVbQ3/EfFcRfLir+lfx8apNVqC
MqUyN/nmaRUlbVsvUvD5CkPjIACO9ld75qDJeJvvDp+X2XuSdbwhjmhGnVMmfUbs
9xsOFCyYGdgULEvkERMOE6jVq9c4WrepblmWOrKLirvdOLLHN2D93DdHmbliO/Wd
zIE/9hJHuUtscyywJ7xaCCMqyGEDnY9N6sJ8iy6N/Ec/xGHYTBwNHIxpqon8E3Y1
QbEL6+oe2Ipoui31JkH9lhD8K8Rtaa7Q9AtKiZhgoBTlSVNirD61ICQSkla5WoWt
a1mp/fU8SbT2lRW1wPgO19XyJXo8i2qxRB79PlB7P+Ydr+zX0ZRjQDHlrEbs22ci
h310KLY7QdYJBRueVf/vZPxFistwS2SETM3T0Fa62KXYAyYmv4a0nW3bO6QoWRTJ
TYKTno5/u43A13C/gab/8fzj0u21QYarf5+E5vhx1BCBNj69rArzbXbL6wbCxE3T
fgKuqJ+VEfVMGqkn/2Ah4NOqVIz1+yt1O71+j9qgQSymZOPpOtcNRODXM21xMQSO
SovNiof3zvFapvkDTCJYvBs2bOq2kNIMDqExzrCW4kQ5NmkDnYU3eZtit46CSQBm
LziZEmRZMGpOe30jZxMRk+TDDuPXUpbJgkJhA0STHoQY/yTO76eukIWZCWr9Y9fa
DXqyimFQjZx9iRqOp2LRJNPios49FDlGI07AfqHmmbHePhOxKpr6lBxeRN5eA11o
VfiHuhLQBlvyzLVcD64zyfr3y5CL6l3k+C7axmp6zE06Td6aJKlwxdgFJPmO8nYz
d7UXQCDo63GKGrc+399wuLCGdLHTBrxcEfHSqG7fq1wxyA1YlxVO2Ql9Q2xBvQ5s
gimB6/E3kKs45qIgmoE7qTHsnLhqBoS0pc7feGNNcTns45tfk6YbtRzCykBTdnnX
48AnVFZOwRC64sJwkNmEeM3YPc2bXeZnhdx8htMUh2Sg2ktf5XmjjI9NbP/iR2V7
8n1sN8GEmzLGkrrezBunsJeUfSrrUJW3NnAaUlMm4QpsXWLAFp/mi/3a4m+vAZfr
BwrqS5ahnSNCoVlUiyzy2ZeWoaAyQFB1htGNIPLbRniWE+DMSQbaz6PGYdQ22p4s
9fXbLLxSkRhCOHuaSCPnUQnerw5Ni7dRJmB7G4rKXZ67A9d/bN0Ud1AfpwjI7x4R
6gJgd44Yl47nh5Bsq6rJTIyjjqN2P43yDxp6Vdc9E0tO9IwlOYIlUh3+64AyLxxT
dHrn8BSXudhrsdyZBctVlXeNC5hyVqv2rn94I/jZS4b4g147zPj5cBmXMLvEfrnS
xEm2eHM1J9C4SkGJ5hP0jdGtqBaQ8VYnpsTnCkggA83aZmKQdF/gPzwdTqH6j1eH
1VhTcfioyweSKZkkIEJlVkChkmrMI0Yj2RhtsYfmQ0X8ifA1SlDSGtpN7pBSwDQn
kjnin7e5lvMdJK2M6cEZ9q7J/TaBrWH7BDh31QK+0MUKnIuA1ZgqH8YpET5I1B0B
yhS2n1+j2OwYI5UlGUoHglPpfTE/KIE6C4tySM8EJYI0L+DHKBSilyfnRiz9r/CN
5yevIXVpklTFZvbG7ZJK+k3GoGMxyn7pn4uleCHsSpXvCBI7d3yhrSrm6ZBk8OW0
LM/WHAQQPH/g6ITjh0zsToAc/OLFIYYaLBWSsAEZHL0i4jDeM7bSET1EfKRwvrui
WF6foOYbhCO3LxVAtdWIQ9F3kbGhaatuAjGAXzypuKFXxiDVbk9Bef8ab60gNfq5
xHh44+pvCSrrWBTpbanG+YoAfaWh00Ksqr5HtEQkn5V3Rt6qrJXWidMrYf12d2M2
OczMIWzhvKx30nzJNOVqkk1kdG7lpLDiTnZMF84bfadY+6tgnX9h5v5Hal5EvPVF
rinCoJy9ACGfRjmBcbLqgJ1vunYfqdzeO7BlBXO4PPV8XS8ir2qK77cmgqhwbRde
wJeiOXECKHyHBy9K1PVtBVWijq0dVI4EV08TYQy3Ce6srOF5oB/Jz4p5IxsTbyvk
yHkdhX9MRjFehawzuWktn463S+xLSXIj6ewB0gdas6R3236z262xxNGDyAh6+yza
YTGt2yXuQHhrxqIMGgOLCZCFgS9XO2y3AR+nmNJLrA7j+y/hTiyDFghS0JKkMwjv
PEM2I+XkffzrieTdf8F+1hXbTrbB5m+9Y93DX11b8Uv/yC95KDG3QdvSUo4NtnI/
2CMBLYOHmLtwwLpQMO3ipKluoyO2CfbQh4TEBriZDi8ZDEjWIk/uMXmVtMOnTE7w
ZwMJTG2NFDfYiHAwI7nS6CZLSMrMRrmyRtjAxE2bwZxHNaC+DOJIZajaykUomseD
9e2HjzQ2O62j6v49DYupUgutiWmdUiAs+Olo0mbOmzsiUj4ZyOBK5Jhfmt5RL7p2
7RLy2VOQInBA8XzK+xx+alNWi3FfG+r0d2rWxd5ZqbETANeSvulvgrd6/Y7AqlY9
V/5htybXw/7y2gdMy7YwxGmelX0uGMqI6qjVbvop7kqkQnUPq+DaH49+vZvLcRKN
XvjncX30km6TEkKqe8KBSbCZGTVjQoSkiX7it7OAwwkHpW11Qu/p2rmyYIe6/VM6
DDawFDAx+IOXukp9F0TrihZFTUjQ9LT6dQxSvuDEolaMiY5jl8B4FoHF4Dp2g8Sb
5UBbnlKT0J1TcVPxjSDCnd64HOg3adO7hrCYbOtHERvOh2PpOT2tcCGa8ahZWfLY
YP9DYTTa9ivrT3tlRuDeHAq9mviRx5PO/NJiVCSYoavzFvbC777hG4RxuCJ2WVxj
P0ZQN6GPC7k8zTcU1R+JimAnRu0Ndn2vX+Wb6Dn5u7EwUaVfLhFcRzAi3bRXXwKR
Qd/LPOHf8JqIi45TJVvLpLggNJ+lTKnq7x1mf2jm98SFpfJBWlKF2SSlgsy3/Qxm
6FEw8ce9mrXYmMNPjEn3jTXNoISz7XnZqRSkL4FVdorufYUkyv/urlvtknhCC0MI
1sXkaOzO757hxr+8xYSss83fX3d8Asfx19VxA3KF2kodHB2V2u4Ra8VfFvQSgCjY
/yFDNdmcV3W5fT202iwZBRXVHjuObinMsPBHIk6vzOBG8vJvqPwMg8Ss8oU1pIJF
ku9RJSNbMFtIBx1nwVlCmsZiGnTFITL0N1jc54QMwRc0XvlPwLEqQHzowNF8rk9t
r5+4IQTHnVKpS4tQwjYaov5MCpGtuQrCMJ4UbC7ao5ZqtWhXwY1rbdbLpoY84uPj
+TaxCMe0pzEz6g/JIjYdATI9u3FIM4yhcTVM5MpMsQbluqhrtiJCfOe+2ZMGUhq/
kfbiplDDsDhWIrN035O65yrWt3EqDak81WAZeFspaHNTOr0ouYGCbxr7zM+3zUhD
D4e3ct8wXTUg5gOQ0Gy4hYI2EhvlDD7NK+89kZ+TVPRlN0G5tehWx7JdvL2/KckV
aBRCfIkAkgv5hwivChJGJY3/nBLdLnmq5Ot3yAn9tTwkiYeGpi0WcX2KHv2z5zcP
KO1CIrBgl3daKAZw0x/akqDA0a/XC4+9iBUTacZj0i67da/PbV0X0h636krQfXcr
vKPZKeLXURW2s/i+uckoiLpCgkznC6bsPt2UCPWBdTqIftQFxOV8S4QRgHJo3sML
7ilWC2E9oZg+M1mKFDKfmwC+RIiXmIU499R5O0ClM/v+Zpuc9on+kqkCsVy3viGc
OJz+9IS8hup+UJhZ0o4tOYAqSwJ3kj7nnVLrRTOctt96uXXKqOALUA1VV1mxwzOR
YHKmVfMUolssaVUT/CkzVQMb94u///g0KbMs3uffE4BDSZfLivZRbqs1eNEzYgJh
ckLmBDmuRHkmGVpSaimllJzkVqodmf/ODxJCG7qVf1MXAA60roT8JLxP6RnZteaC
76PT9pUK3pibAKIJ1G4/J0s/x8iJiL4WtI76S3xfAj6nYREhUtLFdzoMnG6ZIpKy
XEEso6yo7EfKAGjiTx16KYmlHCPqxWRtQ8a1OJvIvOmnqz80cryhvMYwiLbN2dpa
XQYSktWW60RmaOrQyv2hXtMIZI5G7DxXGHMruO7qLvm83o4+QekpYkvruGcAur04
JFS/rNiaSr+9sOdw8DY9XkzkOhu3JjIYkFf/YHF1aRE5N5/VHPyaRAxKwRg+g1mn
oYgxhM6gpxKRGIE/eOOvvO+KrxoZfpVPq0w/sEmhJFvpjkb0wHS+HNyrLt1YXLLq
mesGhGIe5uxXBHp7OyfB/HhFszKHRWYn4viYWVXWqzKOezAzOSOBWZXH0Sdpr5lr
nqFjkc6HZBS2FRXbHo7L/8glwypLTWZkcw85I/CCS28a4GrtD/7xqDfI8e6aHSke
HqJ0zFwF99gL6C+VYCUHf9E9HICPCBorDqgE9fcJWXuFfrrndiKSr6IGne5TaeRk
UgJdRpUhihjPvsPosxk81tqPAdlyQXpgxstUvxoVjb81DqrRzx9IeAuSpTGUdPOQ
F4UqKCIT/uKSrCy7edm1m9gwhO1x4pJt6OLFrPI0x6HZKPxmcO1bxelpEySaYfxI
UHdntn5yyVaQvmThPPE1xxG/GjYapQyLy5yiccgvwLRnpSZdjsSbYOKrNYXfSLtX
bcgUlwHovgud0JiboaRl5hBVpSCuRAS5HBt5K59w3zmmiSx4HDNkADZbVzceN/kH
+qj+6fQgCd+iBKMgR/BP4dA9nfty9APpid4ztBPb/muWVId6QgRY86ychcvYBdTB
04kpmrU2n5gCqqr8W/mtakjFV+PY25lJuwv7bNPnSsoLsZA7BGgLJ7uqPOi4bwG4
96/KB2Juprpuy7gSTY6fifpNxAwDXdbQq6xLDwlvaotQmR7GLo9TTK6028ESMxkW
2Jun4e7PBaIxARWfQyStC2lTl/uSZKBiPq36u3hz9oKJQrseMSL2lyj2BGJXhomh
pb1Fl/PbentpC2KwAoCGWeilPHF6QX0KU+ZRMc4KBOgBA0o3Lm90EVRyVdliArsH
EGoYrgL8fi/T/0x8nJ6LI/AOVSuY3FVdgBdoYxRmNzflH5jdpgZrfG1NiestuIwZ
Hgq9lVhMsgHPhSRXLsdkcluMGNnIJ+6mtvTr8QsQLd0OELIDvPjPLwl4sKLYzLWg
Yd1IGOwJav+D7tj5vv+YnBadQpqGkAEuwiggwT94OT/4C0usxlxyBBUyzua1BdYU
pMHU0raltjFnKS6/LTN2qTv47QiYn04ZVz08HdPBlRLXn8Om5+8pKDeA6i++dCQV
O3XpS9mNEJwsLWVorgxcKgdIqnLrc0oScJQXmuRzH3675zKjAHhECRePDyJNhCxh
UOSNPZVdnSXU3f8Zng3Fj0MK670nCHrl6PhP+tvQFTsuEWSKO43rcvNs5RphkGal
a5Pw2OQCpACyrVPCBu5eJtDBQurWrAisNM1rvwwy+gQnTX9yQb9ctZ7LTy0ZZci4
5860IcB10OYRiFjsEK7bohu9Xnr1S/LCiq7qB3nnSwnFFVBVBxr01OwIBQLAMQyt
qP2PWLJQIARG3Bg+zEELIJwlLqCc/Z6Oh0GklUHmfiVoLgDsl/V0lUkFt9ieT4WZ
9Q0+9STWr2SzmzP79lyL1/1VkImbWGC1bVJ8Iud5AQlOHgzlHM5qvSMD3sCX+qFu
wrYxExOK6fLHP2+IRaNi5u+cjeFU8eQislBpUbi7a/RP9IP3J3Ice7XpivQzCsQ8
fJ9UJ8lIacjACzp0VS9KdqGTAqFkW6a0gAC2GB5MpztF4VqNRztlcgz02CykM+6j
KHnbKXQNec43g0QNModXdmkg2WWewWdwINDRqVtFj36tNYr9CJX/MQs7psqQFk2O
C8CwIOoTMx9rYxu0MN4iydNRMmyXtnNpgnABZmOugYlqxzeVRwhrtrijSuaxwks1
BpMWEFNDcRlmuj+wThDrvU8B4yzzudvgFQHlXardT2ezZgrGc3dujqC27y0o0EjC
oajWKcIYeQrtdo0+z7Jf2varpBDHJZUTbRmpNtsdt3OiYjMHg7Gwsaku1SzA91KH
ofHtH7HXeiifLHpfh/ohqVdIwRJ1U/CsCCFglFEu/cW2CIKbsDCdbtHCNnfSIxR8
cy7jPYDS/k+ICi7DrsCQTb/QU87u5HCrhpm7clKkyASvQJu1iQgZB/PxG0kICMjW
axoPiS2qns6bWyTKoDf8NARNloXGhOkxwIX8ChLurgB8oU6FT8+uApSSNjTVRl1N
xFA/XBovtfgPmfmxxs3GCP25cOBBa/IJCbGXYjzubNxahUdIQ42rz5WmueJukF9m
yfLEguPG5smi7KMW1bxhgF48j+qaUCOW+etVh+dc7YMclPD/7y1owri0f6pdy6bB
CyuWg5096PL55G39681sGTZEmKeWcnVSBoXJQ0JMZk/hhQu34q5pDPS6KM/7Riny
+sHUlEVFPhlJG2cST8DdK66tRgoPuyeQ2HQeGt9fawptgiJNn2pgQKpZbgJgBaQq
HxvlFzQrWntWAOKXaILjDh4oFOwhHSxkx3+hbBUjF6O6Q+fDoAqWpqKLT6Kq34j3
XpXeQJa95t6ko5W8cmBxNaIGMeqXvWVb5Dpnm823Y9SdWrLy+sDIAtTEnF/NuYQr
TvwbNyJMjoV7FJJY9cDTLqeyt+MrAkWXwd43Wny51i1hTZD5A7IyJcRQgFPxApNi
FPy8jjAhyFddC1/Lfx3wg1SmUA2zVfDKVzqXWLTkgsp9y4qwwE1QOIJizzCCDVV8
qoUZVrQ679aEnBGKBt/Dzxq9yb9F8cT9mrOA1icYfK2fXxjnNR97DUuBb5fCPK3i
uqbr7iAoLIJItwI9XBlsYdCKbMf/Exl4Pahow7NIY4lvja54SwkNe8q3hcHG3nvT
eYo8W1T5rdNdi9FSXU96TOFVaWi9TD/7W3KNPIIF5pgbeW7YsN23TaFutb2RW6j9
aSyVROT9U9G/fvKFsr69D6PzZ3M4AH1BM4YDsQeiYaWGl8BJRoTMu9BuRdefi978
WepVHYrL6yfFTp6dw/CBQgCu+dQXQb1r0k7vDGIjuamph/QXn+puXAIh+BkwCy7g
evbe6Nh9ZTEKjl0AM0/FHm7viHGxDp870wkd092Oci4aAJtlK9RVgcE8/DnIcqSg
dPTZEHEuAlvlhENWC72JQQKI13SfN24Z9iLbT/VfsQ50C4ETA8zJZ5/9GvdS4rCl
WyWtfRCu0tr/qB2g3dJ1HZ4pZxd/AQ8AnzXVyaY1jZri++IuY1qEo0KaKFgBtkk8
h1aRKaaHOX32N31gDRM/4jykzH0qTSsYyv7U+PyzlNbKRDHKDmvASd9YLX713DjM
hcqB77NYvblA4FlKCL3WCh0FAz04lh6GVmOz8r5sVAUWZ6SjTN+5myFxDqjbX1PE
kAzVWtyiee9zXzr5RH+sD6lfRZnGvagx2lfw3zUh4sPw/XgjkiAYPf7wE/ZSj/FK
RwAQPdB7LkQpu0Z5O3p6SZrnaIptrXWvW8CZLJ53ctyC5M7/rhzOBklR9quajEq/
BpETw6eqm9uLpnvcY2yGkhGNz/0bmUaD0+2Oau7Aai64bIs3wxShsTZXZQ7SDMZP
b5woE/qvRqGvqn+jS+LwM0LdOVLH7lQmqDRCRsIkbyOE73M/wdwTUfgUKM5iRsA8
waelpNYp15ADPSW3Vb7pqgd0Z/ta1VApg3DfROKn7HY6yiUhnysyia+UTG3Ogui+
mY3hwJ9rxM25yP3ikRVQ3IY2duVQ4HP9DS7KgZ/M/qxQZ3MaFbOorM7u9t8TfJky
acK+PLPUeNNJRBwmXhpi1+uefrZDNdstwoVPsTnQBhlUXh8M2xv2+OMuwBP9Cabp
+Yb0DOY1Jqh5pb+kIPwWttFplI5qJR8OOuM4ZKWZ9lV6P+q16OOY5BToguma8Gtg
TAYWffObsEfXl2Brmk5ypUJI9Jy1NlcffYeECDtiUgb7bjSrxsCRAl3N6bRLZLsU
/cMCwFlZn8dBVUZzoAgPr0Hi5VzzIofWvOMxNnxea32UmZVpZ4ooZ54hlFEwclzU
32EN8SHsNZeY+d8UNtomaR79vZ9DICGKIFulYJhRmZyKonv3iP8Jmgyf7pw29TlW
CVtLm1DYRhAWM5dbvOoBFRerQ16OtzMv1ubBNUnXiTq++rE4mjQjy3gz5kozOWHg
/YmhQG+q1gS2AkA7Tz3TJByHOJDx/cFGFZqADXVtaPBNT5Idciw+O5HMUR8sBUsu
AZ3yPs8Xj0s8ESaNDlNaaQla0FgRdJoh0k6n5MpE6KaFS2Vp6ZikmdErmNno6oW2
zT/nUE7J7LrbmcLggue7sh1CE5yb0TzkDDdIihT75gMaRTjk1p2u/aIbsYwqsVUe
i/besLCv3MEqaGAlcD7Y2mM2AEQtQOgXgR5xU/IdJqT/zRW+4aOdPxStzI3Wz5qk
GduqOsmXcZlnfkh42J+q6OCLNLCfAjJuo5x4yOI4ln5ZPMbQ0H5uzLnrQMwZg0Jt
SEa/maD3bsYcDB17Q/Fy3JV2+Se2g5phAVre+GqMXk8EHwRfsezUPY/P5siw8JJQ
AChT6Y6c7Gb/s3gadaPw6TGmxDYBr9tNPr8oNX0owdY7WxcpvolgAACt3w1KWv0y
Ucv1bDrC8jHQZtRwSAQ/mhbcExk4etbLrI4p/jGBJiJiv5wBozTccUnDxOHm06M5
gAFkDH5x3Kl2w9iHvuQeXul6qqbAop2napBRFA47xECToP4RsOmZ+/0XzMNu+g5N
kOF5b88u2U/CEoQu4vPCopEnzXrKlGE95fh2vHfdmEToeF8c9ZF60COaRnbEbuVD
UvIcopnlDYgJwqKVVhdgrgUhCaLg74j19DZ1QxLa9Qp8VN/KSTIzg7jtCMNucyXK
45IjUObX1mAQCbBzJ9qKUaZW3t1ByaZcRmlqeV4edNtc1dFn2KsZQiKKcmY4wUiL
pF/YQqerGEAZjVD4yQAfDxh5Rws+1PxU5SmhMQ0iKk3EfNotUm3bFNQVX4Ym/hwY
PvYIQQSTvVxtC/z2YdrJaKFjXx5bbq3gEWmPR+FnbhmLuO0WP8mBkW/brVz8TpNV
iCA64g3Wa4oVx0vooNdV1rjLqGht9ZpOGwuEh/JNfN2TR5EDvndLwfjh2hib+IkP
Cl1zHMPmdwUsR3kEXxPOnDqWqRCox3aAyT9SNzo+/uyMrQsD2q0DynLuShgRAEkb
CS0FQ+PiOyBzXBXEtvQUKyu1Bqc4oTSQRC3CT6cAdXDNdlG2Yq29EWvfEvJLatzI
6GbwQCMjZ3CZRB2qkjQpZiykZPyvkJJvNUzu7zkXf82c6a0xjogthsVt2TYM3DCr
m48R9M19wR2tVZv0hBpv8kBObAeR8X3XYsyoAHqvxg5X71SGD+VtQRBnWMW7yuiP
QwHkg8McgR2A4BNQ1WD1JwWYiRtVs8FsoBBt6ZhcARoIDF6LSUfm+giY6u0NI0YA
TTv1JNFjMajw4cx7TVjTPpk1hrxXPLY9Lf5S6eecdFMjLr2mEJkOeZ5lr83C99fh
W5BQcDS030Diw2MgpaQjnOs/IWwjab5P5MHsX7F5t80kSt9Z4KWnc1CnvXGiOi3B
l3B2GOW6GVSxJOFgWWw5h5GsfcXFI77EGhixGAnUP7Ye0GNLAO9BVJ44mAWbdauu
eDujqFvEPkpsSxAa7cgrCnYXh5YLkcP/OmNUlk+ekQyU0kRkNjRA/Vgebs48rvT1
wJ1Bia3aqtBTQ8ST15q9+zvy6b/z4zSZW50ZEBeHkftdUfsBxtWbpF3n7AOyG907
miC9LmzoLFjF5bdEpr0dsztA8Mp5ImYSK5IIO+JOiuoSC+sqcGgxYs5xT8lDN3cv
oNZg/QXmLzAHrvM3+Y+fHgY0gJ3Uxuw7BrkG3vcj7QBpoRrX3qqed+lgOyCSFEcO
seRrwrwdOxLHBKZTJSkpq3jfsjBt1doPrLgBs4ByPrz414XVY7mSfqDCw97Ghxto
0Gp8zkogOFG7fzfOyhTF6Jfiih+nWZpsYYmXAs2N8LN03IhOat2wBVKTxOUDJCfl
zStRfRDAexY2qjl6FFijgOQokOSNVtIx2F9HIXDj7dmkKcHMpdXKs33l/kFAW7oq
t00wUn/i8Hm53g7UIhRnyKM57/1r84pjTn1hJ2fPECFaJIOxiCmOSDEu4PapThqu
SuaKjaHL0fHUyb6vlVcSKJtGyZ0J8PSDgeiAl1dDKmstBp8eS0OL7LLm91xnYPh5
qicj5fG9f46iLnHoo4dIUu/zS7C7Ll0fYek2XrlPXs8ALTMFsUeWFnC9Wn6fuQ2i
/xUmVo6WHrP2+G5SrHuuPvJ6bxCdhyt7xXhnwKI4SklxwDjbVRZEwBjJOpTBuM5y
f/UinOCK3VulKd4shgRQ6o49dyFaBO6CcOBkhM/fwDpsWq0lSDfDOwKKVlQuTqyQ
DEqzxApQMUVnm9wyPEZU7/zaxiNWOkEVKCVQZLoSbj61hR381eGuBXqTJ2jTQqYo
ZsnwwI1cggoTwjTnNgBt6mtyeiz/dEkjuc8a1I1CIKdcFhHgW55O1YLvlqfSY5pY
mK3Q9noJyJ1wU0+3D1YurXEW4PC7/DVF/lWVnYK3fusTk4G/ORv5P3fhgKtqjo64
8WHIf5hcTc/W++04sT0LT/6f7MUbhfpM1qnw0/ojU5p7ovcixefLOkSbGFO9IfxB
2IFCRPYICJ4V7B1Ux75KhFT9VWCH2ym7wwqKS7fKbnzZv6zB84ekdIo3gKUGd7Nh
O4BlTJJ1IX1uM5E4MYCI/qmGVXX9LhMMvunn4XWbeOkOQOWsmoqihCwvRs2woCVE
aS29sLSB6NZSCggyigl1ShUqijiznzlCfBcyTIjfZToS+4zEGoRqM/9Qd8atNl7u
O4mu3KsMXLRiqwUCP+0QrWMXlUIwBpOpBdxtkttbLtoPMhn+kNbj7IIDNrRKnzaE
6sPHPMr/Yn26acQaVDVwMA9/W4Z3cuyKKStNBKr8kJuN2Bmq8tjIiTYLgD9NwnYE
8cn5b3vNVwoNyJhEXMhsW/OuC/zpd2sNhk4NNpyKqgpvRgoKxUsKYlELHELUewwB
ENGulgSfegiV5hxPztiItrG3LYSKtumE1hr629bO29P/D6gJ+tgilWjDt+PVTjbM
mye9EuPQK/WZklyQuQ3Drub+C4bdM+43MScWJqRXhjHmaB9ZiU4GbKHorPmkoWKH
s68SCoIq7R7jRNDrx5Me5jJSb7Q07N1HPuXJyWfCX402N3rZX2jfr5o5HMCpuslL
Dqy9b0p/crpTiPkMGyHxdug8W/8AyE1E8RClrtuRtNcTXGW4JFW9NwTeiBDq6Hoq
8jWFwYxq9ECoiwBlcyw2s5vEqXHNTZkeTTvQxXig8m6CRKx4GxZdFOQbq60pnaqk
r0C6t1y6MFp4xlrR3So9Zm41FmFeZCq73gRjNs+q0O7wpkh7uAndGVjMMt8sfmnF
BY27NeR1LCR/jNv9yOEGxi+UT9yn0RLS1GAR/OmRwULAQt/lGIoCOgEC1x+5ZqQU
ibzC77xjixCp0aUZC/CZAn/AX35LAYTcb2JHfYvMp9o9KvFnaLYMpHdSLv/oArIO
N3RnXk1/3hpePgCfXfN/LtiS9PS2e97JZOuUhH29L0QHPFlzv8TMpm5G491ZmIO7
9YVLOmaqOaQJmt3FDetgRnsqnsbidjv8qRFrfop2NVyGBg3uBHXn3MfYL52wE+zR
z+SeXFRkcFxRyyZ8Uqham3ImUwefhEQ2DcNnw87yUk0ffuF6nIx8WlhViDruM+Xh
439h/K2EckNgL66FpJxHYPZ7mX+6nJnxVIuHX9ir6XHQEAuVTChRm3xzVjTg+m1C
7akE/Q+kW6XIQicL2rMrXfjziEPvgo9+1tTlBDTwTacTpH1E499bRvbVXU4VnI7p
LK83Z9/FmJuEDgmAVhEuX7tQ0ptkU2FjgBIUuMaCeAYGqpkBiiXIILkP5xrfD7Zc
SMfNThkSCh075lvNYGdrdIFjak39QH8jn1zTftEFRm5fYkMfP6kL3joaS94XdNQX
qakHOWT/PJ8Dy3cNvXLE1dVm0XGTlmYqqKi1/9rzPDdVQ/+mW3PNVH2xcmlRR0f4
AVHzeSUxF6CalZ45VdQYQXW2zoU39ClKWUqd61ek7OaDdQ/hOZlkXagsFvizSCXe
b4X1kU6MopRK1kz1uefaPEcxkE1WPFh5xIuQQ2fC+AqyJFG/YWcBFgU62NPBITrV
KnO7ywvQrbyWrr9Kb7fI7497Ie3m6MncDbtheap0RE/Eaewj05vlYQpinPsdt3Ji
uy9PoBSQ9f2mL4q2SxRzl4SuxWFn0dWRvWDY0PQ1bE1/7XCCivPtX1Oa6r1CYhx2
IpHozVY8kfdCrpnX2/HSdPPNzfWoo/2gWo1QnVo0LlSzrSVsrkTFWbJZG6WVxKia
VNvmSXMyqQPhOAFzRGsrxCXXP6y3NutkKR7l3CRvTNgHHy6pBoSHgiKng/Rwp8g6
miy8JxG76ryMe5oktb6ZwlyhXTRzEukf0ePjwSNdmi7szoMj6tAwjDADa7jFBf8m
8TKPA/n5Ey1pWuQUP1wqtdba3nM4pWqL+axphNg+Et7gW1z4/5ggsQH3UvoGNDCV
HImwqpWFy7GHmYZHvK0vPE/lZ2Mok9E5xhfBQUozz7neXszZL+u0P5cnBxXTNWWu
S15Lc/3Q9n39m25ju/OqaLItFWcvew3kaIcTjZk4pAz/OKgv21/j3/N28X/TtPwI
gZtMz/J4oqZDwEw53qk4ZOhQean795eB6pfOf7Zf8LVajCfjUTwEvWqph9YD5KZD
1zVBxgIvC+h9JQYEl8/WoztKK8pAXec4lHX3mDmYxq91SZ+TdgbWhtUykTijqx4K
xd7BCEIEzgDNBHPAxlFjDRYhTFA3M/wHhVjSoW6lPxUvgpj2dRG4BM2h9ltXKuRc
zZU3DivAO6cQ+xfXl46oxaUlxUB7vSWzOz2joI5X1d/CKBG68pJq92gQHlx8svVn
VwyhUAfYpVEsHoDpghN6ExXkc4DkV4N+rm1X2Td1erDbK/1jA94rq5sUoa6gSfUm
Cqhy06ca+ELW+aJ9C3mpfB6w1SpkmlNsCpuvgJx4ZnGLq4K61L7VBTHeicNQ6dB7
bLzyQpSTkuOGled5PyCk8VetJwnas8lFGcXyqAGA+SlWSUyVD/W2Ro5Sbz0J8gyw
N2VUtAVn8dA6cV9PdCRo8V3mesVeULopyZMJQICUGW0rdGdrGPDPVi1IQ4udL2Pi
NOLxxOT2s6u04w8X6brzmHriDpym2R0hBdyaH27lf7wysHwHFpzsZ8W+nF2Q5FMs
T692FlR+1r/yiUO+eOYk3MvfNJHcoXOwfY96mrD3VgBJ7sEctUjUM4CyRSzYIZMm
PSv5tBWESZD+MdCxnFIcy07Fx4x1jGejVXKrz6KGcNOJxB5+jHigP7yuzrH5Tf+C
7OZpZAUCJD0qX5STLZNH81UfT4xNZOJm2fR1cdZ/WtvwKS5Xk1NRh91ww6UdLS1W
lyzkbXGBRDAPhS3C/xQPQCs+axc1/1ot6VvCM9XDQ25y7r4Dki3kTVyIqGGXxAJV
G1q8Jhc9zuM5fbdJi6quAvb8oqvthsHHabLJ7zq/mGTjWwGAR/4iLbahE/bB7LKf
d4ENRbWSZGdSA1rUVnuLpzrhYMWtROCUlpCH/c4YoFZw+DEQTzFT3Pi2HfCJA5mQ
UVn/i9N4vxObq3Li/bEMfFvVxzRcgJ8K10jLVSqrp8G3Js93QXwcbQwK+slvyuSI
LKbFaUYIMH22i7PbxqCJUWuzP51dIRjlGfIrNUL7EecwtLO2c/5lNPlmYMofmTpl
ArUQ5kejI51+5PfukeWMGazoBP7AemYLCFUDzsbe8l2g+mGhHdMkNxZ42GdBVuJs
p6c24aalJt6iPdZNJ2WLNEZ4xG2TOBTfiAznI2mbzCqzefFNp4Npu8TZIL306ILp
kum9NWv/LO+gXbUNcJnIA5C64UlmIZzgZVh206QySQ57qB5hRElitrxuvncYNzWz
62to0uMINVOTjcq8dhqyxLoSIn5ScrWtaR+6axqS+wmC+R/Ef4wC179rdWtlg74o
4Xl0RYrFBPUYkpMFGeQl3nC+u/+6TD115ONCObDVlwNXF/+3twSsgCgf2SeD2L5S
PhYYlAMNu7KDCGuwzCSeSzPbA/CMMDZC7gTaAlX68b1hs/ubcm0MfbQGwKKbmOsg
PnLAbUb5QI0OJHP+jqk0CZXRF2iBD21oXP8oXGjslthBNLaiWjtBiMRmw06MoIcF
OBO7ued0Z+9m8wRRGz81FZowzPGeG/hNifjM1UwJ1N2sQo/ZJeUPoEUku/RCHFTs
9Mr9EhrzUwk1Q6V1bjIhb8wUIQi8J5T0u0B7RxHhbl0UYCOUCJL8+M7z+KaMfuoC
meEssNQ9oWWPRQjpZQFY2riTr1GlzLBKAlhrE25p0GcLVYbDZ3++5ql2/6UoJzvc
JWlxB2qr1OGdEAhpzAiAYJBiydIlkBcQmVqzl3bhZcOFWTnH6MjnaG1f/Cuwa2x5
oSidnRse7/EdIPzYaAFaUwuAH36NpGvhkbA5ooLbiwEBWGGZudf4qwCFZntQZn+6
vMmBDXfFa6QVTcAdma6UEeBfMMKUWsqOcmMgA039PyNatPqoP7Jg/StTM5CrkY7g
AnrJcojaYmAskwGXh6ECRVUtT6BsnS3CrG5Z10c099WVU7XSVc7NugS1GhhXsszv
7EOdW/ooNld9CfzTdYNL6V9wyHpb+/aK39G7Oh09Dr2vQ6K6RqwAqb3K/qyEgjUA
zAfMAPRvlAcTJl8DwMiqVcAylAkJ8pjkfZJ3PqaYWDGKwgAtVP5iQVfuOE7V/veb
26oCQMjf4QOJoFHkWBYO4Pmp3S/kCQT8u5bny5DqdWDUN0eT6wSz3d48Z5WOo6BS
S1lqJlY6VfdZBbbI3M6TUd23BYQW0SW+GAUtwAlHUHoAV3zZfQuepX99yGjc9jrI
YLmbLX4OlqwsdzHSo/kaG8eS8DV2EVPzkwasuyWCA3zjAt4YRTq9YjjSBb6qmB6/
MADco7f+KFYp/GSoEYwOeoW8fw0LLwmFfsKTF0G5cJYXQ05Z6BoYYckiYd9/QYu2
fa0l840kZU5i/iVnnUemIpDPlw66KbSzvxaqBakbr+h4LxmOq4PSEZNbz2hqYomL
OCkCaNSVU9b7hLiMRD3n7m5Ecg80S55jXfXFGUhaZ1qV1uya8CK4k0T1Ip3MEDaH
FfuOIqcsmSyaMu5nrIjFNjFxCsqR+uZuYHVWm+JDmw8iWoQmXQO9+p+/1joCOHSw
cA0IsAQTEdesFTQ010RnV0b6AWIQQux3FfK+k4HLT/l1CtaNki6vzNpbNi8K6AsL
u4dv4g11KuJ0Tf2r4aZ3YbpVJwEqS705nZaHp4WjI3JZ0YZ8lG5b9eqxyN4QWKpt
1Rs+PFm0pAemZmQ2Ikb98uJ2ErP5gVKtRADUtrbRirzWOwsQoUYQ+VjbuIbz8s1Y
2ACdMX6vOzEQmATdkKP/d+YuSs+zAA1A1/ZYY/KsUF/XHZ5oUvJ8cDaXanwVehxU
+VkCGnpml0Oo2/lUbRuvuQ+26AxKX6RbHYyNBDBgEYtjYvEebaeq4NcGWwhwpfZx
BRIcC6/GEQc2fXfQRnHBjDll2BGx7zcq/EDfAE0k3YexOGn28SJCN2McjaL1JIKB
6SOVGgnXEeuoOZgsKCKCWoVE9r++gpMuRtNuTCWw25v8k5CV3HGsbgLuIbOyyPQI
iqVyrId0eUmky8mvJ3pWxCznD2iGZnXm1pJpM6nsG0yfxSWnL8FLCIKz1mdFkH29
ggV3OvjIn3q+cnqx0B4AXOSEYZjzV471OCKooSVRQ4oeDS/yVdzCmBNTPv1Z4zBC
LxBqjRh69Lk+j3QVCuAl2A==
`protect end_protected