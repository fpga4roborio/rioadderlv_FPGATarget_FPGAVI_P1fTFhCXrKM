`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
ddtXksX2+yylW5zu6QL2Lhnb2d1sD00763mmSITNX595NcHTEkwn0zB1Dry37fOW
FufOhVzEJp80NC5qZ/+F0Vk7Ik02dIR0elf3clrjeJRK85K4e3Hoo4xn7YbFUIms
l/8VZSb14+JVGURjfswrIyCUotIzlzVYZ6gzoZwDXIi5gQIBf/gI+KxNXPaKV+PQ
Ufys/12rjO6aI/pPlqSm0hCvftmBcnezN2hk1UeXgOIuKZnogjOsf0iJVX2aOOWE
6pD/psybjbnsNB6kH5uFTA5frkzIzkzl5d9+YDm9OyC+k84E83I/7/j+rk4L2dah
QJOvksSIzN867/4Qt8qYTQ==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="MvBXkzurAa5VTw+1JJ70nePUfoQXBvZOku/SMmg4TwQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
oRtzZL4VJ4iwysPsC8SXYCzXS8Fw2gtZTOskLcDV+1B9Nzn1zTyNtlo6lNICRmmK
ZRVu2BmCc2G+fmzynYlNTnSa7C0Cuel6FYpxCBlOuk3OF2tzAmLAuDyOH3Z1Yjzk
a0aHuoCdIRKv7BrZCdALt03JeUmXKPdOmIlkVGFl8yw=
`protect rights_digest_method = "sha256"
`protect end_toolblock="Jn9CQpRhJt4rnzZPRk+dOpzAubz7omckX1MrFd4p81o="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 6544 )
`protect data_block
gD6l00tciPUa6pDNTk/+tzLxvdHE2s3DQL3/JqqujQBC/Ei+vcAB8wM3doqg5vTg
mdfn9XB1bLOis2CVSfu295W2DNwHfMSTc/8BhCDRnTlLIX0UCJs9Za0+LoM0rMrV
T7EjVWppbP+Em6PkVKCwlmIQ7JKaifJ+Y+kjw9HCGboYo5074hY+K/CBbfsBQY86
AyoN0MKhsIx+eViNgnWjA5Q+FYCusm3YSaY1max8h0b2OP7xr2inrDDCiXZzxKqA
2NTY4A7shKLpXc8QI/up6S7eiJnPbf/cpHGHCE2LnfcIG7q80Yso7kRxZlAwr86S
1x8MROhCzHZQehroS9apYeZrLeqPJTIOiEDVazcfkLVTdG+LpJPuTHJISsi0N75f
vpqihKU58duWmH+9inhGsMMSk/7aYcFDubusbY5AhuUI4ZfyduT7tK+5QeivVx07
cprwrdeZUXptacOmApxQuhh8PKivSLVFEs0m8S4ngpg9NuE/zy5oRckhXprufTLS
ByT2seXXVo2QnA+kTrEp6r/MtTXplT3G8Kr7dv3V87P3L4flnI6tpkiQ2jKzwqN9
7kBh+SMg1BA0HHsSR6ymqEXrKRO+mV2hPCwKLFNiD5SHUh6Ma7tvn1WQV6FlW2Es
MngkxpF9/t122/F+IIy/BG9fAJQv50jyEG34ii9Fq8uOyZZbes9MQDahuKdP6qGk
r0riZm4W72+XcZYcdQLiVY3oYl/yVK9B+GfFJzug8HoO5590Njtx9txxT9CV9u2t
Li5RrqNTQ8+qIO6dH/sOgsQUHeJbJz+HY19wwuVzTva6Bbd4nwG3jOolWZ5uYLpi
T3JDlqUkHIRDN+wCbKFtTDvbkB5y3u+yURPttOykqoCO/8o5Mn6+x/jhD24hfH8/
C/7fh1SC0xUnU4QprRF7y6CKBrXNSXXa1ebCLZXZ/eTKNpajY0D6sbXGvARVXmGP
uo0SAJJJ4xWTBKjRiwhqjUAtGVkJbu3aQkqgEIMOsrTVK0IgitXwfFB5k9eHimD7
2M/sH6yZPaJKUULy890HsP9rgBBD8jxtbXnGucnKWI+Lx+O9iqwNLW6E7r+j+j6z
E4UB7Cso085kEO6aebsfSDqnHou5/TcsKA21TEm1KtCB2Y49WcwCYFGuS+4jmFkZ
TjXqibS9pPNKc10gMfwS1qKigCXVN+55oHs52YtDgtgGW92kTJgBXXj+NpZCh+Oc
tiNI/VUi0pS3BDYlx49FkaxS17F6PZFP37sNgcoFcLNgDU9v/XCjXJzLz5oNIffe
vByH5a5TxpUsiS6OPhpxr/cbugohkmMzNa+fd/oUhpmWvkE+l9n4m7XmMKfoZnC6
l5VW86d3IuPEfrd6OcML6dPbf3XhS6SYS/Vqrcmf8ssStJIyrGQGYp++IFRkylGC
F3I70q/q0B0Kp4LkL6Lgv8TjLPQY/2QYHCr2R3R86puupwp+qA2afz2Dx/bdATU9
LsJwCkPyCbeGXUzvJq5XhpZr1P3eU3uCHfqzVKfEG3CckyGZaDWMp07Mo8LwDmIT
PKBvpa9SCEe7TTAUQzDH1jtDPovSzC1LtTHpAWfnHZkPoPyZBfP+kYALgdKiod2g
zx6d1jdB9v+8ejGitJgFkb0cPj3aMye0YYNvHIzGwGZxZKeQ5OVJbPyW2aO7DfEP
cq7Bt+6qv13nAiFL/M3u8MQUJm55KqglaEsH+c0W82WFOb86GUQR76Ol3vrPi2WE
9X4AODzB+jypxvdDVo43NuGF+p55puwq6GV8JzJTIlVEjLTHIucMhJBud4N7Wxnr
svxoM2RygAXB9BYqpz6YTdlg+LMEqAGHpp59Gozmt1xFmfKrlG36kYZLe0EIzHlC
sHntkLzve0Kvs0vO4OyyIjXEmB2H1b3iSYF3O6rSd2m6sLxrRm2HFXMUt3/JcpVk
EXv8wOdC2eYVxHbKHmeP7rHGBxPv+ermH/PSlCgfvvrahxWfgb9u9xVUdKk34aes
1TM+TKOEQXlLFcXrALxGwjpEZmZMaOlJ9tdJNweJmJmHpQMV/gb4VLebmZ7LaSwp
c4IOmDSCXyYqeKglHeap3UnlKLcGbT2onbiG2JxPjQqq7Vt2azealRx8bxRsQp8k
zLXaaHWN/oIC99G376lqJ7X78uRDSoWXHaFDkc1nzaDU/1kq9PcwlFRWB2Hk6N0v
mZZzdG+6SWqLC9wdZXmXMl/VL2oWNJgUcBD0ZcYMagJz8fXdthE6a8drRj1cr6Na
tOiKqAd2c9KUppJM0Szzpq+NKBmCB5P5K1mhzBg8UjtJ6juhaVcSx/y3vylteY/Z
cOn5AWWmUHNShVwp4fSW70HaL4/JFOHEzN1b13PgywAbSL1QznDOJND6Sb8OUAd9
DFJH/hbbDp+VcfoqgCKMG00wEj/TtFBmo8T+fLqA5orPchwgLUkPUHM1Ksv2nhJe
mcEPnqe787orYY5SmrNxJ8M1eZQcCaRI55Eev8D7r2GUJk2Bgj2qMigT4YkIKSyp
/QOypiRytBlDaKMQ02JS9+u71cMa4B9hziDGbi5Fa9Tjbr3HOXtQNNA/HTHToEkx
e6pbDoJsivhXMUt19iCq17+Gu3Bco9cqeRa5qj+db81R5iewlNZtNKC5zlqqyBG9
pWegsjytYQLMaqmAsW5tet0APK0TCFrVm+nWsQEwUS4iveaXUMfF18xoAUIGClow
yuCrxJnBdliZm0qldJg/aHaxYclcldQKPs8ZYKdEuLgRlYboFMNnuRyDmj34SbgA
YD3AbnEpcfLvVc6OXiP0TU/qlO5f1MuYLALglznZap2rDm5dWJyTHVHR4VENiob2
FxMUl7BFMDa6zM6HpRHcBp1Di+X+kBL74fw7owTrLRqE2w7ADKbWfrbH/rBbiR1B
gvuc/4Rc34SgvtsiP51X+OVeqvB9a0UhVeM+SyJ3o0fDYxvVEB4sW3lMZP6EHK6j
bLEFn8ENxH95aCYLDUnvrJitRlZ9xFW86K0p4w+Fs2PQwTPr34x9bIqHXmHWJFjC
F7VTp+p5dhIhXIXKTc411vrqImFs7YLWKekkD4pKk9jZJoqdlisDYmowus+YoXgm
hrwyupKtPeIXWUZG1+8l/auQNjxemMNMy3cABfux6TSvRbXWfHR+/wnyo0Q2PY+A
AlKOKU/RNmS7YsB4Q11tgX8Za7XTLbWasZ8i/risEHjxWTRUHJYKgsv7PGg/8fS/
HTeEKKlLnYHlzRqjrlG4TEL2EMV2vTCHDlmleY0rKrH3rAq3ExJTUxEkp3/oGyB7
0tgHYtbCrWWDTfK9NGjgVk7ijrqpEod2XNqZJQrpn2AMiZTccET9wN6w6rDt5MQf
87l8CfkZrWZm2M9cZpHobXfR6JEWwbSxoXcAXkG9LWKCjDXPNWXeyrV4qrutoCtA
McJ6WeEfYVdcjPJ5My/jAx6lmznZrIy1hAl8cVAj0M5iu7om93NkkeC5oNY4OtQI
UDgXQNS06v4u9MtPKkAMNO9slskccQhaxMsFH1Q33qmYMZ+UXh3UK3E6/pjdjs/y
UsTnlTRcoc9yiaKpYheJmFbrIfciZhdxC8cZ4l30skg80R3K4P+MRWe3fSSI4Fdf
f+i1i32hZhbALYWwGpyKwxAolgBnwrwwWGT+LbTZFQoYczUlcB+s5lC+vYBxsUhz
A6Pur2tPy6CnOLw2nnWuE8JEQYZGwmxQvY6xvMbJwW69AyU5uSJZIc9w44B1WV/+
JPz4r/ANa8u7yf9J4B+VhCI68QX3cPtObs/dn+X4WoOM2ZUJ59gWAs+osCklOwx8
G5q8QXHGjK+YMXjHoQDiXAHSAnK4CDfpf5h69YXIsubxt3W2OQ2m7k5i3y/KonwY
VCBMpZwZ4dOxXCRYOMxAB0/tjCoR5zsqb/UpLA9uBCVcFmHQFxgYCKrgs9EFFRnd
IKbH0mqt/oDQaAgglYeUV9Yj6d4Tr8JmPxex4Wg7f3dqPwtjo3jLCBtC1+dD+vMh
1doQo0xMQ6VVCeEwPmyDvObs5nZjYMLcsJxLTHxIzvx8fpJUjUWwyKGaRjQ+rzuc
YrTRExCHz8A7QweefaucFK5qQA5mi9J/Y7sj5UcvLznAcUSfRPX+xZqNLKFL4x2Y
GKT/5KUQ+JcQDY2ZBII4zhF21gIdZpdW9pAt6sOpXVXuXMQvgevS/cs5K7xlM16q
y5od8jzTCO9fClMXkOPFpOdK7LID4N4pSF/xm2Hga7ALM0pMmwkqCzWSfurQPGWv
IKVj3b9jAa2lFuqpaAGPSiypxUB5h9jEbOEUHrUDOpfCDbPRHdeyzKXEEIPelthh
mnUR/Z4m1aSAB7QXT9G1IwFNYcQbOjgD4ArVrgLmI6WOQ49U9bKdxzNwhHo6SGCR
nM0UFF+Q53NcQi+Wk73B4gWU1El0mhffDSs1OZk17cCnXXLtXdv7z4XvLkO9ejle
62XShe29JUeu7AUDjUYnmyjtW4O2OqL5j1gL6b2FqCPruFDAMFs0tbNXzn91xBCH
llTeTLAxpTVT16dHmeXB8s0o4Ev/DbIF9pTBhGZQVvyAjN8l3yRB3DJxpfuCaxgs
zrEkFFbrhTJtHvzbd0d0abjZdLP4htHO8nbopZ7acQ/5hlyLB+qo2k4wdPYo6JVT
G4nxEvX5ALrcBxTKVsJEiMe0FXobmFYYrCJeDGgh7XHV63ILZPT/AUQx3hJDe8TZ
M/wJhQSQExmhb+18Ujmg/gVB70rBMOtMd8GnlgKJ43pWktwBoM5/fc2msahLxCpL
CkFsHNY1+b6B/KXz9+7/B8V9F8qQEkirXOnbImjFb5GOqOQ+bCFrst1mePGQzmmd
UU9rwmMwlGGdVBcIq8TP8k+X84YL6H2yqUL+qg+xYMtjnw+RQbKtN19MtcOMlUif
2qOXpFDJ/4ZDsN+ShMa7o9F8AG4i6xbsMlY26f8LVcB2kmjp5w8BOFboJn4xEZ/6
WDo95wNhYytULEsEdktkZzVS7F/qTVK7lhNzi9xiQfHZCTk+r+bG7H3YhTRfsMjw
p6l8JPwR2JuRwZGpnpTgOrQpkq/7pVSfeRk2pEUI1ppq0+hqehz7Q0LSwd1daxAR
WAue1Bf4w6OCwRMeDmimnv1hLRWnJPRPuGLzrfxCkrYnSd3lC2taSKk0rNnioR/O
oZOhJVKLzN0A6OxrdB2xscFMGaLr044qKjh2WYY6RuvuIX+5w27qodWqfzJgaJLs
UUcJWBe5CRfAaF0vM2qXoUx6nX40v+BP0OaO4tI4e1RPZ2r2fyUXbCaPiSpWIOeO
2M58afvPT/JreeJ5G+znipWdKSavEcvunDOjdTl2RI1T0ucrmxb6Wk8iqomK1B6o
RhsnHEOZ92apgxqbPrImXIRm0sTmCH3GPZ/dB0u76u+cZbDenxr8TrwRHOvHsDtB
m2z6zjLryoDdd+QlC2gwwPcdudWlkfmyTotI00hEW4bBXwL75JJb4vIl1RUKI8Ex
ar3Ql9kIOqkIl+UYD2ZMJp8g0mFf5E/R2RtHLex1mVHCXkTa5Ie6nVXmUjQkjkmg
wv8SCV3bkg6uN5r0TCXojo7RkegnjsIUgABT2aGyNv9eSelPneacAEb7+IUBKurN
poHt7+0m+4/VzRpJXx6DRMltP9uxl7NGJ+OxD1NSKzMbvL2hyGn9PdMGhQtMnpAG
fSpDzMNH3iHfLmw43WR8yv4eSwOF36nYWaiGMnVqaIAkJGr0/7ksm6MZhdZWU0Ln
zKesJgLsBWPBQ15SlHV8FzjOYb7pl/ecz36dQAw/8vqdTYUrvqvZoWlGHTB+AA8Z
R/ON6UAEWkff0uR3Wkuh/49bnyefvaFy05fKUPs+dq9S3ZBXKPrTBKHjT/iKntBB
UeMx8nyD75ln55r46pkfr5Cz2NTJADSmYxGuCFejXj37cQh2uRcgxha8/hzBccfI
W/Su6ho4P3mR8BC4/my+3z/EWN8Gq7HowvlIWvTkcGmQ2jkEu7HUx3/ygejxleFw
DQWu4O+KwHH/xGYHvC+BWrEkuc8zD8va46Yg93HDW+fpTyUs5CkdUrKCE+zd2jcE
BALAF1eVssYHL7pz2ZZKS7hpe/AreQfGxGERy516eDxfaj3LkenQPlr1bIvmQZLw
e5PcVV3R2zwgUVTydq5PILGpSfiUYF+WlKNjjvHxBO/NuvvSGPKQEiIwOmc/06PE
MkefOVP1p6UZSJMW2dHOSOYPMDzvYa44usog43ffhjhpu84//vGDq5Nz3as0Xy5i
dJA29R/qhtghhR/0coGODCIxxdAJrQU3MTnI1EWSeOfnEvIrlRDivt2njrkHso6i
UTk2UGumssvD++v40abksucBQIczQYLZpvx4OMz8xMzW6OVFzqFnsn/eIB0vgTug
f6BS2s/vhkl26RcCmM3atV9nq4on859wP5Z930zLcRtU/id6F6SWXJzT2bUUVni9
gaWDd98DH7YfXXX6tGA0CN+l0LvOZLQAVzBupGI/Ftf+gxTSATcruOuSvdZhmoAQ
VEjRJ4wy+LNUkFkAlGDQxxPtUp25MyUuFTZDtAPMJME2R0HcTpQ1Moo+/9vXHOin
HZWdlzDGtLqHbt8179XHHzcGhwz1XKTU0UxwzKyQsDttj0DRShvpDVgOn1tWwmFp
bgDhkrwMN69VwlcHJfLKf/f8O1NIuI3oadGMcQQJkNxaf1YSyauLOrneAgIOXE+L
7ADZBSLMXPygS5waieTVIfVJzv6lqZdqnS3OLqwFlEYJe3nNUIGiquZlpkSfyTFS
kTD8ac/2m/TV7jr826PpdqaDBo/ca83skXeMubj+DJa005IjV2WqLFzUFAvltaZb
NR12rteAMkJJrpjr5cZpOk1E9THbl+zz2fGuxGq3MkqlDL5Fe0Io/2BOBdJeEafJ
IiK4aHWCYAIkDdroZ4NeBEMwA3bGVKT/He6OQJQUTf1mhF2MUp48Z8kMVaOUuJHw
Ctdk4H99ce1MQoFePtka98u9oNQq4cGOHFwL3irdmlGt6eeZ4EKKU9yPHStPEO8K
FYD6szzT7HYuzijvgIm2D29daTT9Rw4au7yK34WPVkOVzhiPg7hsnRb2S8MFl8mS
TL0v1nRQuc6L8BTJbmPtBer/396ERzdRKeHd8dTAe2Pi8uJ/nBoUAWZRQJjbSoLZ
kybQUxfHB2pw34aKR5F/BUM8C10kIjQiOL8rmAqlWPw6J7RInbWef1QiDLun+d+E
MsDK0lhyTc5Fp/UQO5V/dwEy6fm4rQpI9TSnlFMOPN6vTdxHjY/wApMYkgr93OBi
tRS4RLJrW7S9UFy0sxyBFPCaXvt/rkUmBLwcLsD587Px3gx2ITzf6tnYrKJ1vw31
Ia/o7ZMlt+PEreqxG6W86jfFlT7MtxnA6cgLI60oCHy3uhFmE4Ac4i39YonikpWt
RZiMzsmfUZWBmjp1ngL/5uzTbusolZVO2mRFO9dXyIupJbLk4DjrjbG95l5vctal
CxJIsbkBU+SfgcFAwGVTRSR4vt1wGZ2LNsV1Fv17EvsNgl8wvxj/q3CvQZXWQKEW
qTEufdUUfZ7JHc381oVUlzBLYkvV8J8VhlqL3zzAx5fD4rO8IV90V/U72VHIxF2d
jtOgKNbbyjEqi5PNf9iPlv+YghYkcckBjlS76oEllw5y52mZF68ltFgdQRdO7phJ
pLJvsWLe2xei5wYUcbiyyhHNutiNR5qlcYTebgK88QKIy+mJI/uOaVGm3F2Ye+XW
DUdfeG8b4B0n6RCg8UhWvMS6XVYolAL6JovSBsniVBuw1FoGhCJ9BNzb8wuj2YhN
IRzA6CaD3qiZHVsgz5yF5pwUHs6ewd63lFZNRDuja0I3pOnEKtsLJpCavqo5wC1f
P7So0jW2N9oYZcc9Pl27GVv+csXugDydyRNMvw8rNBugn2wts2XBkXfeNER6DQMr
ZmDkowdMChjD9BJqYJoD6Ks5RI8GqeYTN2TaUecyfjnoTvfISoLlglDmNw456MQY
vqRaAnsjprRtRBf6zdM5Llf3pRbnkiCTxzvivtb7lKPElutdFK5qktOHQSqv9O0C
m4f9gIOD3ieGh4SVnD0CWh7tBsBGYJi6VJWQvs8/WkK+j3nRXSWODWGbkSVEy1nB
MX3G0wjLqalhaV8LlcOpwUretrMmG6SKWi/FTI/eCXZ/vmtHx7rsOna9+cnIoUJH
urH1McMB5G126Yu4Gd0nMT48sp4pb/IBdT5dUZw1fBth+F8wE/NTwDIykkWAWguy
EVWQ6QDxsFmG6ZJ84NhXEvoJopwfwbW64P26znapLlYqJCjk+7/ILxPZeDGiWPwn
wlelptp09gQraHB0Eza9MdaOCEB3SOAlWN6SwaHjXjI7faS/CJYb6ssB0L+0ifUi
lM8iBKSifLXZoDWYpWiVpt0hrZlMoIKcS4r5KBKMxZ9R9wS0A+zl2CHxwQpdPkTb
dVG/fxBoaL2R+388j4Cd77pVoDALPXThh3zAVb4/UIAqm85lIGpSMbSiF118iQ+H
d/vNz9lOb8+t9JzJUxU5gWV9bzawIBozfTNsuhK/tbPByGtQQG6TKi8b1DrU/LTE
IM3dbN960e1Hl4NFJWei1TJs1Ok6T7o92O5emnX/hgdg7AxB6bzW4pYWZ9OIOd/p
NfUPBn2fj4ingdIk2r1vHgFUtDFgbXIiVYbpr0DhLgiAqks4Qa2gjViJcYOvv3Lc
MSdn0RzAsMWco2VZoD1DQ/7Ol9L/fCqEkrqcEk6dViiZq7cZ8E3YigLTISaNdPDX
VPKIezuBCZkZnyJgc3mTnQ==
`protect end_protected