`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
ddtXksX2+yylW5zu6QL2Lhnb2d1sD00763mmSITNX595NcHTEkwn0zB1Dry37fOW
FufOhVzEJp80NC5qZ/+F0Vk7Ik02dIR0elf3clrjeJRK85K4e3Hoo4xn7YbFUIms
l/8VZSb14+JVGURjfswrIyCUotIzlzVYZ6gzoZwDXIi5gQIBf/gI+KxNXPaKV+PQ
Ufys/12rjO6aI/pPlqSm0hCvftmBcnezN2hk1UeXgOIuKZnogjOsf0iJVX2aOOWE
6pD/psybjbnsNB6kH5uFTA5frkzIzkzl5d9+YDm9OyC+k84E83I/7/j+rk4L2dah
QJOvksSIzN867/4Qt8qYTQ==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="MvBXkzurAa5VTw+1JJ70nePUfoQXBvZOku/SMmg4TwQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
oRtzZL4VJ4iwysPsC8SXYCzXS8Fw2gtZTOskLcDV+1B9Nzn1zTyNtlo6lNICRmmK
ZRVu2BmCc2G+fmzynYlNTnSa7C0Cuel6FYpxCBlOuk3OF2tzAmLAuDyOH3Z1Yjzk
a0aHuoCdIRKv7BrZCdALt03JeUmXKPdOmIlkVGFl8yw=
`protect rights_digest_method = "sha256"
`protect end_toolblock="Jn9CQpRhJt4rnzZPRk+dOpzAubz7omckX1MrFd4p81o="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 53920 )
`protect data_block
gD6l00tciPUa6pDNTk/+t0OO0nC/UTtBwLB41d4inuAUA3i/ALrNyoJVcBnAmEQW
ptbcNp5fxEUJjnOxnedyZEuEBxWRieZFQnkRdF269oNfXMBxHWN+xMRZiCBR2tLM
Qv/Zls1PSupXplI3/TBsxJenY/DantRMGDISCloal3wh1m9OOYB1cCMdK5UGbAUJ
Ux7WnaSq5M+AtNhuy+ABJH4xU+rWPQXy2rcVhq8i5pCpEQqtDd1LaA5t1SBguh+h
3ptJTQopY7RkwiC+0Llk8X4ygn8yKnp9DseYWfMh/llrIzZGQlXZfZq0e+8LYaH9
H7SPzwAVW5dO7DYqabVo7THrT0NeN3l3QzNsrJ2bwcLn83yPMtCDxi4/P2NjUavJ
UwK0W2zTG8sOU2AbHzsBnWqdqSDqX4HayyrmEWYIwDMKRJnWUoZ1eJkkFuLd6PwL
0Yrp7ELq3ozToq6KF7doLvdh9cNadD0YetoTYyyKs1ZZHS/B4BCWKN2tyuVAuPHw
SxoOEIZeXh0BneEdNGqjjB/LR6ILOJMTnSFPQ1pxHwjjL9BFXB0VR9vGr3zm3Ak8
2uD0YAflGSz4dQdR8B4SA9AJ3+zRT8tYvNUEFmzcy0hA9Sx5gC0TkOu3untCNcwW
ODV70pxtah6N08ruTeBoEjh4mEpUuO9bTS25adfL4WNyDYHJjCtqHB8FMUnel0Ok
En39fwv/nzHjJIhGB/9GiepmTFIKiLjMtf+oR2QZHHjMZBX8WJkTaBbgyqsMRZhQ
vMQl8nuLYl7T95S9D0IdJKpRyInAfF4F7pdDUOK2HDY86QP/JvgIToXkm6WquI9S
GfgppzKCfYizmPYrqhv6FpFjx9M3rZETBsEIwlrKV+/UPRDI4VOXY/SeNJ22F4GG
TePTChhguLD4PRsM+lhMfj7q2k/PdEVlRE3ftidLk9JuQnkRWP9nmnrYofL9ZYaM
yuChiDmjIycjoMA2qOXcStcuYix4RuU3SXllcB64vST5ZlqR0neOLv43WTcKIAt2
cqD3p5yEimBJBRQ/wECzIr+HixLNEtBTACDL062hNPoReSABWiQslZnE/i3MXwBG
FQBnkFSTK9lgrKizSPrXMARYPaw3vSnjDqIzhJ383XlD6sdivT4HoAgqy0NZNsIV
Ldyms2pEATQZotjbl0MGZdNl+k3kvMTXazVKcQdr+nnufxikywEPx29Y+8s4fRdK
frxaT6MXLa/CwyLCsqAHN+62ca6x8ACF1Ys6QCcZW1WHKW1hEAbI2a37A+zrMryq
azxO2CRcNRBLfW+f+ARm+qVmTZtwMQNXL2p/hE2JUgM0rpH3TbeSF0vEsuQiJcZV
wlKxGs21WArcYObqZr1IZ1Ps8IVZ66poUGqVGkQYIYyO9ccapiaczz3d0jPpNIM9
yuvDv7VvP0MwNbMZoU2wjajpAFl2vtVPmqa5B5zQfPeGzj4SzrpeeiHKaPDq4ZEF
TWzn/E1r2slNQMf740jLns74K/gcjMqjyRP/DUB6KqqwLUbX1EZyaAw0MDU9DrsZ
Uk93q+xRCSaudacDnM+On6y1Zx6zrAnkDvlBYI+xyE9rzCfu91DwtCsSk9Ln7MRF
W5468XGwRTkbLZ4rPyArHw1Ddgq6L61TIv17J4MlKNAmcZBwICMmDwFD4sE8jkuq
Qb40p33cTasTJbYAnGTZQ0tguRvgRw9J4tU/JhTCJq6j/MmfeQY5T1vTiSophccE
hNBLvpBOZ4t8lq7d8+uq+KdSQM8MUhKK6uv+9rztNkdYQhUA4VBOCmggeMFU3AQc
cQyT3ouvWfThWjVtDHV6XR5/7sg0LoqrAy8Ndf9J6UDu80Ld3Q6Trt44K5cSAumf
iRkuIxwp+TxsCUB/N4lH8IZ4vwSCPQKudVJH1SUJ9KhjlO0JobBeCcL+EHgXGFlE
mfT+AvLdE5xJDoCxw5FQpvyBdxRLAa4AwJpTajt0vrZ5SRxDMkssZDPVxI6iO6zM
yvYUcgJ3J1HVOl3J/H4LkpPJb8cevsbEvJP0f270jGDgG2HswV3WBLsURy6wkfA3
RE1gfdLLw4WqQxjESOedy87wzkZx40b84R3LiRhzra4FC17D2VmpNFm5AuTCRYOC
dFZQM799rtrnHcoSz5w6I+nQ89LLaBlECmcUe+0qTnALN0pZ4XqxKr0abljmhNoY
meaB8zcYGqy+C7XaefDNI+ZZI3ewngTxb2eQVzu5IOZQCPOd+Y/wqT+CtfHO9WX6
bVJ37IP33AY0guxwX2H1EVTcM7CsDflashNizP/aqp0HxykS1CAlK9IpuIhPEZcf
N2JCxzuiNC3H0MUtxysi406BefTem98v9lWPMNnXg2B3IjfWipeYMBPeP4Y6zLUc
BGr9Zws/krPS6lm2Aw+tgExW4WVWaaRhuPoZvJ17ZIFGfn5iINfdTvTDMeryZHKX
HYH1Sma/A5TdPbbBYGsR52Y3/gwDaPNLlLEkLKOw5CUWwHCbkpsmk94WqR7hJHxB
gN5tPDnHL2/5nK2cpOikUzJYJ6mgnbZOXHmG/+SpmMAEGZlReRqAMNpMvLHlz+r+
dHGiQuGbcLagt5JknqjFiEFBKRAF2q2C99mYDS9V52PQmXReB8rvVovc3Cs7TlwN
NJb40iT4U9VLMOdoFyGTw/yLCWydrqXuuV68hi9aEkcz7MVcC3vLZu2+vM0AmgG6
bZanp96UQHjBC5ndRVeYb2lZzo2i84phwlpH9KAMf+jTXhuh8r6jaSpkyawuQYUz
Haq59cmJzdj3ArAqXKgtbn2R3K0xB75y5DyNACn+VHpwVTeGxamPAGsLx9Rrd/qS
BWFrM/gN0GUbwCai9CyxBRHFkVYNGBPQB2emwbTuLeJLtyAoGNqw7BH+Ue0GXblJ
QPtlvf9147NIGHdAHwjI155crq1cIzI3CzTAIh+vArMrO3FknHoylWtHq8TksUqK
fcJ7/V/gffF8YFBjwlClLj8zZglnv+AO9Df5KyUOnlRZXFYLeY4qsRWP/vaM9m0l
rpMwSft/PKOCOg42Jqi13LBZ5ljfNzGXMjxghlPGy6XYkk3DSMhVLeUJQTGf1Pyh
ukr+Ncrt+yCvch5F6Hv7w8CYTXwMErB7USojjsaImeKe7AmfqCe5tsJ71BhzYDZv
JpMZn6BzlUkSnIGFOGmk3OmBulnpoaPv+uaM6q0rOYrwq2JvGeb+ZOd1tRvbv8Vo
o7fMOfW3aUEWvzrwof52US6lzP2fduiQi56q5sUHstMMHCi3vjU2C2OySphxm1FT
LuEpdWaSD6by8BM0xkBCeUF1OpTEQ8VNXLeeOQpwz1yUbUYB7mir3XgeU9UHc2IV
VUO6IvFfDky8z1GDu+DZBRvuZn4H8KscNdQTLemKGl7gFKfxCqhreEJV0XnKJCZB
2TJaz53x3wgSaXB0BjYOIJa3NDoyZ0w5c6qOi9QqaDkhUBkmKsnm+iB1l6NcRoXj
v6hfcmB9ZmH3NP1Ya5W6BI8rYeLUEjgTrWaI5nN8+yYdcKz9CHg3ML+mkQzBbB+4
AwrWxRmDHCBO9suf4cJY4BWbB5LtlZx3Je6NIlJWsbCHtKDOe3ybLzuTtLwc0016
WMkFTEoKeQHgifCmSnVOTIRVcezuzg4WkxnRacLWj3nU/Dz6v8LQk6JBlFTfF7WJ
LIPMfE3cOcjY47jFp74YM8bh0etolMPElYCYGbuhGKxKUw+tkYFZsPNfiDqlJY2q
0ERacg1VgGJ1DCpFyjaEbl6bIMhR82SPTzbPGrpu9GrtYBFRJyVnyLm5tTW/Wt8Y
G5BjvjUU8fwQ7XStqVBqX8dcEb5Io2mP+1FsHPHVrDJ3S/itfe+VF8BQ3Bokies1
CnKAeVIirIv3Y3dqSPP/vXJNFY03e+fAJwhnS4UTD7JVEWSt/6RJ2Z1Yw49VZ28g
dvKrjidN+lYKtpKGcV2lmHYGoHP/2ATsHDDtKRIIO4ygLvb0sEb1f7+pGj3QiVEo
oHvZ+1a68M7UQvgrtNj5KQS79McsOnOf7YWLxjx338nmDRfwyZVF4YVUJzO/SAGz
Nlw9GW2VOXBFfC3+7D8ZMzsJSQNxHvCinlbOfnupTYlfEmRnDAh/i9sIS5swTtCD
elkc6xjXVCzYOZ5b0NR4pS0yoKIvVAk51IoP8kclX8G5/FnYYZ7b7Nc3T66p/+g7
jk15AmW1suYUtweDbQ+mkdo2EwVF2F8pBA18wUvUX0WInUXOIxPCCfU9GLlN2ILi
oTrc8mRBsXKHOxEgdrggg+rvjNW7J5lml1k6vBECnWTjiEBnml7Op32+6oc4J84c
BA+AncZTdUUg1bfZj2FzGUy2b3sQCHLEn49fR9C+A1AMrcwzgoaOeWKDGwb67qh/
66+RDB7BS2vVLOruXBFNCj6FzqX/RIwCiGQX5XZXvK2m56zjR1RnueYp7ICPClDf
3wdq87uriQpD3DsflVUZgPe9fu3bCcg2wExCNhKIRXIx1kELHSnrx9ONLJyLtxz9
O1JwuAfXhoFAbzT5i8WW3rQRro5AGLd8WkJbRZNzi8TbsZrpRZC/QViLlv2332y2
GkV7uXy85pc3eXgXahiiVBruTSfQo0A9gesdf66DCGxRRbbaFbjCKyCad6H/BIkU
fuI3Mh9lUF2DpCek7kRSzRsk0P4vR393BAsd1z+3j2h9sdG5Nt5GoRWyEyTk1ZKl
x+VscFgVr3aCoG+xFhXdmMCQArTP+EWuvgQIThdFQOlBctqajYNUxd29jZQZeEV9
kYloVwCu2ZtB9xhqqjLEJcbih1jarIvf+3STbfwkNWYE2EQnvan5Vfmp/RbrEyGi
jwAAn9ouaoWfwi4sB3/IZRxJqssS2/qhDskyT0lo+9EI22P9KWbVl+O4Qpep4dE6
Th7eJ8Ny7Kw30KIsRMyt17N1JHRsEl/HFh7ckoXI9LarhRTu3VSEaUudfYSfC4DG
qm6GQLhuCKQ2bUcuTCACWAPrn6i019Nw6+l+0voimFah6JuBR1eUV6Vw7p+muVX4
6PAYR3ej1Wu0SxBjlNk1nxam5zqZF2unpSMH9ruw8VUfms2P8a1BMxRaSTJPnCSs
CiDG8Sw5DG7vBOx5hs+3MhpowBLPOnPOThqKhue6y7pTdy5Pix/q/BiZ08T1ZzHO
J+52w0rt7kzH/9gw9Yu1cfee5vnP8Kby7WDs0Ehc5cRdWcuI7JWs25STcVLLvbIl
05DP+Vjj8FDPYnjE3Xay1TkqdUPlIMSQBMDm3srzeMO4aYijWlsPRFj9fPViCyBp
jGLgv8TByylyR/mXAeZrvREhLx92m+W52GO70+98XYorCiX6Zgg/wuztwKe6RVjC
K/FKyUIL241n5LgzDE3GNOD1pgC40Z8gqXtmj6q/Yi96O73NHVNxjYj6AdWWzK6+
R1h3odjtXZ2SEoWQ3k9f0fkyAauiuMbiA+VhC2mSm9LhD7YuUghUQL+ekc3Rzc2W
E1vVv/ULJF3y1003sUTno795KaDG34dPvt923zx2STEcpvY5uQioeu2JTD47og6Z
LXJYXQWZutdEh4aZOqXy5s6hrXVLHjw6eM7HOimEAoFA3uyvczfQkXb6apBQ+G17
oEoY7/obgkTKflDDdgyxnE93hC9lBLACOzttdT6yV4Him2QTzruzWBBPFsgnwAae
ySWqVjWzTUzQaCSxpk0nP7tBghoJx2flUaJkhpBhqsPsyve20NcTpSyBqjGhA1Ek
ilq6YH2fUltV2dhPqihVxdEd29LGCwFMEmIK2AvApUA3UcROhOzNIQgVER8ULLfJ
jNag1028UxG6BJMRBPRrFhmGVS/JbnpcWsXl8s8HctnEBJlYDcNsDUiC47ZU93Py
O7wn3/G6qor6wTXUVxHD7kJJMd4+Ff6Ea+eS+lUa+py94nkHW9vi2hCU1qo0wpB+
RrE4ZjcsfwPX1dttqmQsUCopoT8iB1vhEqtov9khuMgX55H80KIFbr5niMnkaqsC
VW0xMoS28/5tFElETzefSA+2Oz5jQ9ORZTsUZQkDQTQJtlj4AgLU512FtVpLvuG0
wKg9/NXr7DsTUwW3hdeaTaSEeZ47WNDSic4QwcV7itJV0ZKckjI7uMWxEsb1RsZK
CbTIBdyBmnkwxnwTvdeFA21LeDbvaTxWbJFz6X84bninvQQBuGqxrIlXpDNgtPhI
0CMIN5XAVb92coKkPzvxeFiac8H/oedycVwQRQQLBHGx8+WppyNh7jb8i18nkmyd
qSXsklHAGuwF8GrN1HH8gNcldckhfjljyBZNVDFNs6r8rtKQb3GeBF79g1pnT65E
yTvkLBUqepZ94uB4rdXh3S1z0j3Wx6QMrqOW3wqkAy6e4l0ZFgL1tMkJp1rk29zI
F9DUmCrfXiGk/4vpUMPvNIM/55w2GGfnSjivXxF3md889dSQgJMAclpmg0RrXd0a
apQVJL7GUBzHvOhEdmnG+HEZ4qLLECBEdK/2V1oFaFknx0GkQERDCRV5xkpRemuG
V4oPsJSaQVyC0jV54qXzlWRRH5XOjnOO5tFUEukzZoBX9s4noBHxKtpa7h6hY6oR
vCtdX3HrFS2CyRymJCubT8qbuDxPNpmrifRFbGaZqLKDHqgNASyWyOV6p6fUZtSR
pr8VaPls52uX1kigvwkjSvM/XG/Kgkvb2Kul1AMlQxBScGK9dPRN4QxgYgX2LJ6G
9cYRC5n6wLLBY4JgYO9hBDOjSwj4T9Ptxeiy8JW6RKvnJf2y7WFo3KBg4MpVKcLO
FyUBxcIonU3vZWlNdp5EKx+yG5DMvDLRni+EY2BX6atksjUaic0OT8YA9IxJoE4k
PYAGrNuaKrlOwK+3GbVJbnLlHJgWYBkwUzAtk5kVz5+ltgX9Go/jKo686dztZ6yw
uj0EbbO8IopVrms3a6JKo/DrQqj9XwlbzV/sx8PUudzh1a9iY8B6lQTDhlLoVkLD
Y8gnNn+BcGvJgbZ47UEJHKfGaW1OKcmU16yffKlKWoN57UWnCFDkuVTPIjYS6M4k
nve6XNwsjUZIHOWFqWvxYjYeULwWMODm0mAO6bxdV7o/Ll73kT3EWYFcatnXT6UU
Xz+qZi3cB6OQmQjPSXrA0x17ZoKWia7G6YvsmtvU/1Y6Yc0+SNNIgdQEs/xqEB8S
rbkDLSPVnr2p8AdBiOc2c/eF65jfKCPzZAQY8vceQlUZbELqhODudZafn70GjGkp
HIL8fjOUCBaRI/CK1TyHVr8jtWTELw2OkTCI97LEQyag9quWvMsM2haaDcMNtnml
3o4b6aACXPtOi0Tj78drraKT2eM4JnL7ldVqFDB9ipNVsd5v8iCFOjf4WfP3wun5
DEoG6tsMLtdnPx1eRkN/yXN4GHhxU1Gto1AUhFQbvFVvOTooyOGDW6M5Tv7u7/3B
2K9WoRbsfXzYUqrYoznCRyhiw658r8tyaqB2hZFBXz+qV/IgpyKc3wuzunQaN17M
AD4051qFgfPZ1LvleSYzUa03FR98x7p1F5fQCoJwc++hjToWFofjwKIUWav96riL
8o5PJsCtZwH3vFN/6UO1CNgYSRP90Fy8O+xZnK5cNoTqdmJys5C+MfgRwoq9I11D
PbmSPPkAXYlC5inb8jhnsfBIpF/89Jsse7tx4WYyUfX7g6sT83oMmUPqqgPnjxXd
EAZZQ427o3JLjB1PdUo/rcV99YpH5harhvrcoMD2WY6gVQAlJk1I/xIuT3kYVyya
97MIBJYLPUr0BGE5aS+D+k0XSI9v9lQnLlwwjAYsSWt9ds/1FD43DCK6T5z+gSC8
1hXTSzTmUkYw076Gi61T0j7+kgoGE6XFWAnfjevl1xHfqg76RvnXGi8XZ0h2+YnB
g0vJVOE168zrTzunRZkEf/DMePx+lQwtRXiIKzcAYZ3BgwaT3h1R+QV7M2oxBj7d
rMTwKYbrjLS69WDoCNQcF+XkakgCQmqfwlSzRg2b0sSjTq+avLnKzCtspN++wb8Q
oz1RUjUoG3ZVX45cXJQ6JqgbfU3Jm7nblgtCGvtXt1pUsxyXWfo4dNS/KOMLrFQk
AOS495p8CZn9xGmsFk8SSbHAXMvMR8Neshnd0abwRvIuenAGfFku3z04LZYTjpxI
7/njE/ufDcYftjAaMZHakxF5gRYggdUE4KjvrsnKJ4PfXOtOHJl6wP6bxEoWzepn
fYiLf4s4UiQOqeMO3OkSf5lR8hpTO/xCZtto0Uzgw/qq+F8pWOZMHvLJie0wTJsm
gIkA34MxPC6EaE8XoQB9jTcjwiJSn4tqKMvIIWcKsF4LfJYzGbtowpWYPgBNzkcP
50gSi8CbZv7EvdFGSMa+KYn4EPSW6uMQ3Tg4JX8mZi8i/SBZo0kvcGZ0lxH8uT27
P9o5qOZFzltIymtbZ7QaLkH3bVdWG/UZKS97ohoVKNwoX7cs72NLNScYeqYJK6M4
H8ySzQTKC37FQN4QKptwGnQY4O/QwtZOQMnoyMGk9l70s9v39TOqRwos0W5rXxzR
7pb8N8NZEBRXlWw7rcjzbdtrnTJ98zNv9OYAcP6i4uMtNrGBLoV5LeKXjtZgrX7q
mBzD6Bs+dDVDukxW/A6qoiNzHZhk93e8OJSdQQP6WlLdQV1Wg5w3uyV8RhHktkKf
T/pe6YOmq6UiPrlovbwzPsjytfx7rvVtW58qckNxqaNHCbW8yC6vwbZWRktsremg
BYnUkcJEWlq6iycqS4h1I/dkc5mVxVjK/NHb/1nX4w+vgm6kbsD3mxvplfOCV/VZ
YHJ24HnUIX2pUK7rRgRWD8sj2dZwBeQsPRDR0nJ03n8gBpCHzdW6p1QD4VfFyw+q
rvO+6IBhkD51QCuOzS1kd6YTA7QT5WnMNHSnwp5M9IY/4TF8ae2cB1dPzbjEQYeK
AU15j1FSuaqpNig0KD0zXG/CRdqFhqeYdxHISS7m7zqnQWAHpoTDFew3f/r8XUc/
3lRM+Ho9pskI5YmZboiNyM92udGOUyKBSsKwlNMnjaE6AOngc6Ms9sH1kYNN3ebn
Oy0Cxrgd9YC6uKYHQCRhNBzvhalA3HgO02TNx2QoYHBPGtEeJN1WWBDFC/Ll4ejq
dvnzkF++gn1puCSOgRGsGfbpfDQHkp17kVrHfU+R1g8eDKkmy4/iXcJP7YENIFc9
z/JxUdqgiQE/PRwGmBdYHNG359xu6u+S2xkaiVfRTv1YAuCu0CK5BF1uRIweYKwx
SVV4GEmvUU93dNq6RCkctth8mSFSsYCSpfA9wS0iDs6kxuUkl8WCul/0zssihGpA
gi1NWglr1EgsXOEA9z4mU++DNbvZHuwF3alQ+Did95nT++lqqJIc0mwCcf9RiLdO
TWEijXYfkieeTB8UJXfpBPs6c4FL50qOUNOFXeO+2gJbIjeWnD/VXU8upjAUeJyl
bpyoY32/NvNx0n0Q8zIBo6ncYoERO8opSAZtWJbsqZ2UIKrbayKO73KLSIVl7MDb
6OicdKXs1OTEkhFdxoGm+4PaClQ8/aL8yCI6qS0PmRoHg8BOHO2zDnAmurZJy93B
IL+ANgMJhUa0uUKrdcK8zjJh3Lr0wy1hyuxah83+vlMRValVXGq3EwT2wlPfUf4d
8UB9+FGuheJRUOWZ7HRHl7Yk2U8xRC2xgewmHzxb7YsDiN9UV1v+y32ePpkefX3/
IT7u6yQWLOiAyA4OgB544DqyRr5pkmZKDZqG3II6iZ5DC/mRfPGrGZyHtHvHC5hX
mLWnpltwj5D8mEC0w/cA8O2gDf0buW7IVGkMWqMC3H3NmhNBGxUDdC4l4CMfLGAH
QcSaEX05MTkc4WqOQGlvVWeI7RhD0z9Ahd9ivNnOl+g2lvqYS0oxUZEHmWf7ubXR
tQg2MqedNEFgABqtd5aM04pgmI2lQxXl1Bx61DPMP5P2waN1y/LwKXuCBe8k75x2
s5NL+gc8e9FJ1tJkecNm5O/4LQnzLfX66OjTJOTdkn2vkeW1eAFZrKKzE7guGatT
P0SO2tD+6WKe1xWMQNfrgTfDy/poeB7/AZ+pUND1NMAr5qU92s68QQri2udiLt2T
KEJAOhuVmgs1kp4heKmklnIxEasftZqLKZ0U/21r3WEJsAG16Br52m38Mkeou5fT
H/4P8CntbruYRs7Oza7LWfCr9TCy8qE1tcQQPsD7cQj8KqchtVjqARzhZsRGwcBv
1MVCembz2sybB8mzr14orhm2/PURlM7F1EPnFZPH16yAdYHgf0W1MWCqyUgeC67L
AhfoDQtPWU9W7h20K2ev8zLec/wSnBJn+n76AWvDIY6ToC6fud6MNbywqc2OWtVj
cr49TeqYrNBYdXaYkAwHfjm9sPNxEMT2XTpwGgqfACubJrIogsn7iSV0GTPrmt5B
ztYhGs6x56+d62spKj1uLnyScGm/4sTQ9qe2rIPjBB48n6gwBEvCwOIdSMKV8oh/
eRrUcv89wY8uZIUWngvx/oz8HpxLb7DdtmWxo1jVsVW5u74Jb4RYcr3pwMxGvedP
tc8i8tOr4U1Gpyx/23B/J9kOVOfKcoWYqKsfsEsKuIQaDt7Yk0FkG2VZ10mKRX1g
cvmJ0Rqyh4Mw2Nn4Obg0wzo9qtuikK9A5exMG3EpnTuzx9DJcRDN6/i3VIlmFir+
tzDylnJ90tZzp2yQByEtNGWe6Ci97M3PJ3NSHk5KY1apnsOwi/MU1oOUxoQ2cV8P
Ouc0sEr5OOx2PpxTCMDgd/ko/U9W9TzwGM4jXLupFRiYbKRYv2fmq9eZhjnKTn7o
F1+CL+BfCUGr+J+P1p0J2kpsn2cfbS9h+bKoSdFumzzd21J2LdtdLRGlpJJNqXtA
8Ec5Cadu9YdgAJTl8iTKmYvJOEa7LqPzNXFmL72Y8r988w7pAGIrRNZ4CYzIumN5
iLs5QfyiGt4QpnsuL5DedhMZnTDi9YrDZDs6tBZKknwSYt+Mla2ANJZZR3XxHBLN
emxnV++WrLBalEhcKxN7nR5Pndkxyk/loudOQI2OUTDk6uWFL4rWUWQfy3l72Si1
HZ7IPUIJ1EB7FEfDp8KYDrNerhsDWEIYz5TQ9BsBVbVrD22jS7cvwrAFvUu76OYf
LC4jm7UQc+iU7bL+WwHhll2t14qP8HpNj13VO48DIgBLsQ/g+bHxZQjhxpj6Mb3t
Fn5ZgTz/SiYrVpZUc3NmchwxxiiV2XAS7hArmqB2F5vEJTTNYyov8mJO2qFqcAx1
7CVrNQFCmG9uUCzXEQ8TVuNgoAfwLKSmVKHuF+touZzz5INctcd1gII2E8M1zZLx
3RlRIAqAv7WbXisR9Vx12lMmbhEgwhx4VhI6DrJCn3N2MvCxn3j9TOcud0Sb48JN
y0chMOoPhxmJIrgCEk+dTui+moSmD8GTcUFgsx15CEtujnnsyJwK7MT/VkBSl1Bq
BQo5UHGTW5UERJubP4+o7rfbvZIHhO7LGETrWeK/uUZ4oQELaXoVzmvRGklIlis2
PNi3biZ6zuyMwSOQJqYM1sFHIUfqObHsqk9GnRsE4LU1KHhI0B2Mam8P6WFF7s9s
7/BYihHvDQM033CrrxCAjLIqR+tAoIDOqsY3ZqU9H6rzy5Lgyct9B2Y6xLaaZEur
0DrOH1XPmL+gTlO1oUkHXcnfwKZb/AWP4wzM8MHzA7IDXq1Z4aFf9xykKf7a8RlB
niwcplacjpPkMNz3vAEzDP6JEdnNTK5KbnYgwx7WKINd3ZZvoyCmGzYizt6zcig4
aazysyH81wmiC3rZaq+DJ1P1eS1ZcxUydtZqvH4v+NOhZOpwt1Z6DMFzjLy9BVtw
3bro7CAztPfAPT2i2Yx82fvyWNa6lrzNLyl76W6kke5Stc+Yjj0ain9+Ucqo88HJ
UzAhAJDjOyaLD+RD+FY6EM71rhFvHY7/c4QdHXLpfNrWK5LfnZ6PESCG9R8AZ+dl
+qhxZfpr5NExVbDQOH8jRxSEqhDwo3nzLg8FdW5aY004gx2KQtso/hX8kplBsM4R
5ckdNcdyIj5bQ1rjK39Tp42R8Nkb8+4vS01Cgqcdv/qfoDbwG2hLAJOwJT+g9fP+
sDV57H7xR3KftL5SziOnHwNRF3aM2YU2vcZXS7VyvY7ekU8jvVlPb5G3NMEKUVmM
OTo8J/PNLHNXeXBB++tePvNpVaqqf5pJOtldJ/+28Rdaf3fQ5icDxr3wQWNuFC2b
9LhKHtySKyl/luLaI7mc9X30rMuAekjZEzUhtG3goKgl/PC9B1mS05qFOFAd5NSo
2MIsxtxXrGSHxZL1CHDKK7ZUJxL04W99WwkKjgqQeYnKZSoYj+t4Rs8voFiobBxc
c08DRUZHLIruoxR4q+lFlSy1SkeSceyHcEkrVA42DiR7+WlFemwkg30mvn6JqeR4
nrVEFZNnAgbHb7cJFFjAUoQ7xL0L9nm8XVlCuJGf0VL/eJ7D5GG5oOCNr+cOuSKQ
2HHtdqn+kUPMvSAUX5g4aMIkGteZ/8RBAgxOBkwYLRrnhsXpcEYXAwZ6zVTvq1Xp
tJAqqe6H4RmanMSEfEi27jm0qz+96kvnWvJjPkWnjLkIskh+SPtMSFhZFPL+CiUr
xj3tNCucV/4SImOHmo30wHU49gWUXwnTl3hIJ4a9ddBLylVwwMwcP5bJDo62oc5A
wJ0cxQ19tIDYoBPE9cKBWopL1H9Let2j8nrxnB78jJKNkmIfZUa+4Cz3D2WN4OR8
/TzJBkr2xZgi/PjMgnXi8kyaxHi+BGJt80jvVJca1S6kXo82PVMVwbg47cKAqBnd
FAvGen+VPTrryNHqzdN6rtBW6XmqVIjB1aYd94KIytKaDt5tekdNsRQTISpnBxUf
xXZpAmh4P0OiCkrae0ujwidmuTcDz/RbSWQnTpQHryef1KLIQ0sg/HSRufsN8ZsS
yEguvEZr7bje7K+jxJmrPdOBWszLLfhyZkUbfwx1dIA5j3vOoLeT1pg6ZttGW9ka
oOVh5MPoPvFSy6y+dmAaQwhgNM8IjJr6FM2BuBm362D4tPuN5S94gD8QU10OEeJS
rtNaB0WuUFeLmGFU57SomWJgrs630bdxEKKyyX68JVsJCKDQdNB9QlIGNnSoTtbA
klYMOEAd20jnjXqmB1P2L5UGbe51BL+mEWvY+yQCUrrV5npTMYfNAUyg6gyR2wvl
G7fyVbI5ruL+K6QsWoWFGBiDSGZQtqNtHfDTNw6V4tyrfirzy76jgtrtnSZQW5fj
V4uTkPAVjytlYhvqpg3OssCJJXOtfKWM7P1EcB6r1QEcoqCHzI57KkfYZNf021p4
Dn4asQ4nuWK61Sxraln0RumRV8TemWUelAIr71AkFkEpIPBPLP9w20Vimf/lXJuj
DPvGR8v5AdxxVXmEmXS184ChoU0ZQmfQHAaxm0bcfEddQc11ozKWSo5YKyzO7tny
0jFBUmLEh3wwxNfm6Lx4e3oJcbosrqqZVtWSeWHPqcsU/x/qYa92XQdYLxIRoen4
vIqTvWnir6gF9MQ3bebAEXESBI+XZtNWeFHLuhV/UExfc9xsMu1WI0xE0zc7HRG5
9Nc5/7iZgrcMCJYVbjGV2trO6AXm6JtQJUHYDQr1xQ2vyESB+4/KkkGNKzs58ZBs
qtQZVQilNN0weBNtbzJYbhSZphrzqWkO9gEd3C9Ov4AI860dWKuK8UKHkk60I44z
QMFPOGsSCJMAVjErhStlIENyAt+1a0+1zmHPfjJdm0T3QyYV4YGSlmIXLObsarkD
GqM/JK0CYt/V4InKhEhkSz8NdDkjpVGz2S1H3xUZy1LeI5iHzdbR4mwVWL+UrvjT
0h126XBRlSUUxtlS3U5Cq8XNthQP0v98ITLirmuIHRE+N0YiYh9AJO37AsYxiUit
TRDVJeAQkUrCyXvMjYl4OI2THovDoQQSzlM/7RfMbZu7u4y8dPBZUHC3PsRE4j1C
msdu/EnRCmZ4kOQJ/VIbHqk7m08zZm38o5TQnxpjpDwHDnzqWJcOlAlWUXrARsKm
P1xdc5WjokQ+yzl1jaSFxxNKgeZSbkaDKs4EO3a9bHJR3IJOs85RJddcMd1b3fI4
wHD/IwjpM4q7iDUOxjelZmGy88QYzF+cvP4BHniuQmtDRGM+UZGv3ilC07dRvft6
gppc7UAnCXnTiC4NYeTX1mb0RuuVPP4vitIIz87NSaXgkT5WG+PgXPhBJj8ggG/2
yTWzE5OGhy5mFodM7y+/NcrcoPK3vzdHHSFNrertVUEyidRjlmrgUiCaOTDRI/3L
YJokZWXUIlOT5sfvTlB0G6LWPoVF42pO7n6eTfRwfe503oxgFw0D3LzzWoX2qKZ3
i/m8plS+JsdgepFUwL8W6nsGDenuwt/rEyQwZR+wR8DX6FmpdizvX0KjtFxrBBK2
Iyna+6bdb71sr9b2M2x+/1ZBOF7uNrO5ytut6AfP7pnypfqDGt8OwINQsDz+ByiF
xZxL7rE14eIMGqwevxzAO/Jqz3JlBiO6iWzDKxau0IRH6awjDdy+CRlx9vJrKEHy
sWwqsAaNHzlAtEk0aHxz2Sdfi3v6QmbOjCduilKaMKMMRMV6HpCZDeT+PFOSq3OE
wxgmlbNk8sxkaLb+8UD9Uxhr75FZXgbafZyMhA+A/XC+g0pQ0Y3dEStzYutOAWVK
HIGEDKdTIrRFN4u5DuJRhvNuBB6Y3AGyCHfX9gw4OEpGox3Cu45yVrM9+dsP01hK
b8dwcmkq+yxE13xrEpLMRPKwlkrrHYnkTGImrMDUFI89hzkTpe4im9UR9z1lfpAX
Mh9shvh7EsbUb/Th6C73lIVyxrvxlMdBr1DjguQFs5MfA2vbGTMfitfVy79roI3h
NHMX9Cz3az0k6qBNfF66mj7leYWR3/sX51BIOOsp9tAnz2u2ReeVBTyMchq57p57
ZPj9xbaTPvcbrmL5w1WVlXk3FNGk7D+aSI51fnwnhDR/RhCLE4LffWJKtSC5gsJs
aDiLOBzeJ9w+bORD3Y+Rc6Yt/tu0AvELrQNjEcIEJDRbs1KZgVeJ2tkIf79vFIeC
Ko9IGBY1GE4YrqIjZAA0kuMTJzLeyDVzZwddzrp6GlJgnl1JbulQSAg59RDYzA91
Aaj3JoMVXrj2g6J68BBz2h9XNEqcE4jaikNG46YuHyjTm0i5iIA/XrbbcGQPK4LY
OoLpoFOMGOScPiQvDQfvZ0e5blPEGD5CR5SWTZJ61c0zd0saDjSTFm8oK3SPUwXU
0uu4Ddff4XQnHYW23XvTy9BGCylxQ0I54oknoo2ytN9fho0cuHDEX4s/V1K24JTa
+B1IRujtNk79m0uhNdR/x1vaeARC/iqDFHTNMvSoW0P6NmaKiDNLyEibxAMXRZwD
2fT3dNi8cazpaslNzroOngeGcGOW3qdgUb6eYTExAzqp+LtShENrj5rb4NIGH84R
YoHPTCvrGkAfxNnuVMPZ9APiVEqIQ3tw0VghWVtACej23rSn7V5JVyo5FQzWT23o
xM89diIW4KaWmUSP/XVdiDoWoXolfj6TQ3uyhRlGjqrd5YKmNorpZpl8fBfj+i+x
QhFIrSl4W9RJsI9S7uRcTHDg/8sEDpljo1yu2xSr3zNivK+xF8kNgnqeUhVg1uNj
wWbCr0rvSbUZscGZVfpFvkl9zkTTaco6irTaRpmWp/U8kK96hDuJRBZrMAYLcerK
/zoaVl5i8PIe51NbCS8R68qLxrPKPnNfOvuiNXDtYZyatt4zqQEYQtUnwfHd6xK/
6Z3Swmc19O2NgdYAyKHoqSlnwKOP4rAnZtAvwBjNUbx1ImdgGOs9QMLvkMawP3cJ
a+k61VlJp3L6LWCy/yYAcsXvak/6JztfIJCPjE9YiVGVpnG5kc1y9uRKdcNvw8ap
bO6uh2czU1hcHHbOWNqWYo8UQ17oJPOCdb/35TVQMHr/MfipGXHZk6LYM2LZylzM
zNB/QfONTM0QRBbhCYEZWEXqpjQCOj0mNVDZ676zChslI+UX8Zw9CsFj9ifEeJwS
DPGNASwi/RqpXpfUhkgYm696hfL83iF0gS6ykWk2m8U9lnbrtPudcs10Efx7iVyW
46rmHwQoy83Te0HmtKVjUaQL8lyAXjZkdClsdjzNbAlLf/mDYYdJrZE3axOL6q9d
RIx12r739+OD29FEl2HUEThAYA4iqGg16ug2+DKKdoypNueYUEhLFnP5um8sbDPq
4dSRQDzBSJ4YY3eyYsDaUfAv7hSBaBd58AsYPsrBo0ddUsj5ua8fDF6dFdSFjBBe
P7w4zOWXHxvaE+FBFigbReDrTEgoB19h+nbsW0m82u1vv/zk68oshJK5mIaPYZmw
R6WyQ/sOiQ5aQtHJeSweF3ql0/F10FUpLjB9yWYiY8RW5NvMhlQOtcwaNJgl635b
6qGjzhtLEJ43h07K2Hj/AZD40vGrGLQXpqf/DCDsS+mUshuBI8qfBRk4CGz5jYhK
yN6An2cQFfCjga5ARhvIyPzT8Qhqrb2N0MTR6l26ko/3RK+fWN1t94S2502hjOqI
NgzukJiX7IM3m5y+PkvjGvCbmNj5oXbAxG6HHcBd5Q4MruIhelNYzHlQed5mPoa9
Cu/9IisoUDj5j7CIyVKXhHAwpFTvTC/7lzfZnvO0ZVlvUMK1/CPAuRNO7LUxJkUq
FybtKImZid9jjAlOoxzWQ5SgVcu1F5V4q2ac0QFVXm2jbEfz026hXQDjgkAYMbnH
JznZSnU2ObjdOrE1IIXmK4m0uih6gOM4cB8mtoCWHVRDl5SrTHjmMcNaFE2FIu4z
jKjVz8mVERaG7F2JRU15tKxrshGFMSK7WSlLx9mUIDVwmDYAaJ8uN43Pe2WAp7Wq
Lyi2zaS3XnxK1SeMuEePhS94vLEGaFfxW4dZY4kSDsIw/zJdiuVHkfGLmAqwL9YS
rjaU+XuawhJsOCb1b14M9507b0bsep+3ihHZy6tMP7Tv5uZFExf8x0VYnETrb3ZR
WoXNlRDptEaVz8Un9rvFXmYRPpq5bqj/MZ3Gn0msvy7pR+xwb5TVUy1bUq0oSUpq
QA4C3eN2pTNgdjX1zCDQ6aADgtn93NM1eYgX9lYP5yZfUOiIj48BoTHTmaiIccJk
JtU9UaXYuVyPqadR8vMcYg/SAPVz9gNSr/bNSS6I3rVoZ34QJzllhGtREMTaM3Z1
/JFf9+XFeRuV35p0o5tdshuqrfgMvCdMc0qDe0QCrjmhjeCjEz0VplbR0q/RsTZZ
PZZ7PjONjhuNyAf25ebwJUPoMd6UDikxaOHdfsV8pDupD66Bn9oJe77LQxjIAfGc
bbAHhYw9igRSsIRAoRx8ABveZH9bsU5yGpKrZHKcaw2CzTLy5522GfROPhoY+3Jz
XS8ocXjIvbv9HRylNhprCb+lzs4PaXaxhGvhTvddvFN/8FAGHx1OeWInzd/fK6qd
wk4DKbbNbPZPVC011FmM5LfoXLoLYJ4ODowEaQ4/UOi26su2950ewzLwadlYXbPA
o1TAACGFXUkyk4Bm2GcERW3Fw0HMMNhLQeLEI3IVNEDG/fPUuQKNM1lfpLiuh150
D/FH7MVXVmiyTiIrJJJFeaKjn2l1DEentio2VpY2Gvm1H2BpURCUyDvxJUp7v2eg
ClGvG5+9BqwguDlh9rFTtcHI9mcCJSQqg/AUJk1yvk+yqBG4GMD60q5fKIBrwh6B
a3rlhp2JBvyDu0cnIrBV3PP2ajOZsue0U7/VqqCkrdqJAsDO1/QU0kZzG+Ix69Tu
+gt8xwYg/3hn8N0OJmI0AtI+je2wEpmMjqI6vpvMc68GyeBdWryrThWnFVoN8/gW
rHV/rN/v0hPSlSWAPyuyRI85dHqv5z823NdU1/MiJ3qlsI8LuYs6nmtmD2jlFD8u
1HTxwsZpU6Srfcau9hsOPaUoGyFBZLbg5vEe+LLvf+fNZZzSVaSsFkr414jXdswP
QmNWo2q+yeHwvo9CTqCIb5c4SUSPY8R6Ld933q5sjNG0aVrYkSkgzhias6ZpTD0p
dQhPLIbndGwRsVMQTeYQtTBZm65yGtaJj4qY4UfDNcrv9/8Eia6++sTgIwAr8nBw
e2Yi6prZcChco4p0RGkejDYo3brS2H+K7qpfvBzR7rWdEhOasDmeDQzfggkejr0L
u8b4de6S58v3Yr0d0VOCJryq2OCOU289TnLUpFC5ll/TNb9/SkwW/oaj0ZG+CAMR
jrZoc533WOVo1YDXl1VYj45QDWUWylo3uHHxQ8FeqFXbiLF3NyzvlFB78/3ug5jw
RGoS/TLK9hBveC89dWWHbpjLIR83b/+F7Q0fjnrIR2YNONHVae6EBpl6NKTH1aTn
WoVeK5vqO1uWogUZhsRYfma4bGXt17hGNwbRJS6eAyCoP8JuwBIT8Hn/Rj7ZCn21
ktMgvAd1hAvG3AcbmWlPxeyBRp8DxqFNUgsM0715gFKr/yKgBVsM0XYMyRcg+rQP
wBjY9S8GQ3HybjWewcwpGgEJtlj5maJpz7ziVc/wvvs6L6SeRbgY18g3+oFCN5hB
DOwOs7fvmZhAy8B408ajeKlbMp84DPxH0D6TDlzD3FtGUJul6b7OozQ1yhCeVvYC
RznLU3Rg0/0oYcD+cy3i/NvBZKFNmS06nOii5qR/6GbU7vyilFmgNIMwNKW+hG0s
0zlDEmaROw/NcU6bRGiBp3EtnsB/r5NCWmHe4a68xytL2VhHt0+UKEZxjKXPL6Q7
QYgShr+pnHTlP5tkFjzqyzyIVxrSYCpapJqj4jpXBrmaBF9l4D9FKqtHW9+UdwcC
Gihp72l27WHZCOuxEKDYnKWfxCA7k+uskb8TQtEPDuirY5NEIfcPQqcQQlWFAcdt
o/cL18DxtdUQ3UPL8eurCfzMzGbe3cmuCP+MImYAkBFIUc/oMiugKLr43HrBXqY5
mrie6VxU/dNemjHOKxThjPFiEEILzGhZAcS2esr+OD1/LDZXc0pLA+8r33VsZfQh
zWSHMGrvDsVE01onFZ5iyc2N+Cn7iPgAnn5KUVoK464tRsSg7kOiSVM3xc8nZzCu
EmvVryIqbmra/HYSnmwZbeXIoPA0sDr0lVqQCW0eEiLfzrKMmPCM6KOGacNQGgQG
+q6ypOG3+XHfz1kehVV+c1yXxET+5MgpJLSClXg23LzJTgkMGJs73coM+uG98BTP
Pz71lCoUAJf87+hWXTUJ5abM/n+zj1QrXxPZ3Kgoq+Dah4qBf60pGydiw+garwIo
oItmoC8M9EceYvZ7kzlFpgVzIjVM+63ahplzAeXLirhUjJQbnTb9E0fDOhMlQqL2
s2GsvYtj2NhhssmMGIITZG0aghq3/wfjzG/NJiJxK5NV7Ww0Mt3qSE4vqt4um8tO
wBV7Q02eQw1QiyS14JFc7A7AKsAvHlUjiFA9EKVgiHrqAHjiYBVhmXNSciDMqHJ+
R1xndF1rf3ogQDB7U4nmdAA/hPcI6uOzPFLfLvY3ExJnAIvAgimUIPZr0Q5aEpK3
lmTN+FyMzsW9lX+1Af030o8JsfuWE8H0iUjUIq5Cv6bjaq35zvr2C5oz6YypIy1a
k+wr3/XaUi6HU4+F7YYYPeXqhtJISpAXBJBg0bWSsebfnGJ0D18+eHk97xGT1ujD
iGf9xtfkEQv/N6SCfOBn1gVMXJQ2P63GUC3bTmDhmqT6LVtQr/pQsvfrIIUODxSB
K73Cdgq36Aw1s6N3h/9751XT2okiJ9zAR2xtczAauqexaDl6MgqUI9/5GrSOvB6S
K8I/Xc4HLAx3T8UU0dMRrAyvZB3S/QYReulziKT9uTy3Gcj/mrUlen83KiV8o+pD
FV6Bu0L1ucOYPJnOwbGy4K1oFh8Z92wMqWHoG+6+aj0dOBtJfwYzTA9JHMGl+z8n
cOggIs/YPfMg84AKguSgFLFaKbMYvAlAGplCPHDHEaSQDYHjmWPkcLxanrsIMWw7
UbALLldk8vqIkHqF8nduIGASIYS1hxRTYBWsyNJf3SUQjZ2g00n8yRzbl3nb1ogv
lG46qiAYPuLI4Hze6bBbhqvxHbRbYpTiRgEboHUycviWcCxBOV20n5M7wLlQkxcW
XnBM1pY4MUs3UVg+MWgurqKNcSCBgScH4JOqyY4Q6g+aSazkIBQ816nUyvFUtAOM
G1qnYmWO5CQvoUktYCIpgResPzWo8bHx/0VNaOG3uJ3TAsv8vfeLJKeRyPYYiFVd
+l2ZUa/5ZGfud8rRWELWVXM3jfkiFdha2H2Ur7f4J+bcCpWaBbI+MJfzoIsaYuAH
FPV3l5nuBPs/HIIDFQxQ8n6DuVFwBNouUZpkC9e+pOApKiBLjRRbx8gMpUczodUs
6OHN//nBF+AP2tVvIZ63dKZxMedRsR2EmfP6GXiMh03MDlt5mCjBXxu1gtVBrqQE
LFhCjnATpkq8ly7Annw0eqxm0rAPOT0IBgqyf+i4Fxk4hziF0dgZsquSohABmxsl
DAewYdTPd1pJKC8qbQd7x4H+LF1FMwvNEmNNyQWhg9TRUZwKgjSbXOBKaJ6ss2CD
uqFPB46Q78V+kbc9pvepwsaNPVCnJqYobAv/fLreabXUOjjyyRxALn87EEbocDNc
gu5zCvcajEPMll+O3E2WEVUkzY3ehqlnPeBRsh1EJJMJoXZIhbO/6l72/49t4Q8H
TJbpyOHHWxhBXMfhXyiuWKOtg9H0zobybj6SulaIVF9jnp3xN20Zd7naPQ+DgibC
X9MXzcQtjTHn2aQYDzhkNkttMGTat0GzeS4OXtnZ62Mjz98Hz4KuUytLvdlSu6s0
zPviqzfLlns5M5E4IUBwBsTdtAbQXe8tZvnNB9Y04jb0ewzrMPtJwZd1LQ2tM3yb
rHJq9TZ5BhgV05uhlvxs4xy6/3hrFElfbDvOrE7pCHMEG8JCYz2Xk4pdeuEj9HA3
uQySIuTtliEczIKbV3uJgnRoSLw0lICsnYJ/MlzxlhbT/Asv7NtuQBf3YE4cLWs1
5oLZZk5+AplqSM+FolAwo0O8jMVRJ2Yny7qYkAQrVUidNP0sCkLx8zRIaZAfIvGz
RhZYveMNTNsAfeF9SOpKCJN4s7P0uUdOqT1NM80BXPLac5zYkgNgsJUVS5o685OS
DDTjsZRFEeUEGhbsMV8LEWkE4jiB0UxDkD5wh5hThIcpa5UVsUNcJEWttaPgdzPQ
BBkgfTmWgw5lB8SHtnyMa07EJ7rrcxQUNmhT8vulZvK63SF2QNr04bZwvL7ZcAPT
BkzkelZWY9gAzuAT6/gZBG75BxxjPkK3U++8y3zWC+hPNqy70C7af5EiAPZh4I4N
P6iNip1fQfq/A57hpJBQHKzTnxkifAAfNrgw5BaJl5B9L5cAygyJTp3qLvojmoPh
39Bv5kRcpuzjN3EP5vFgSOjq+Gb1lXzG7gXGStSJFJb71c9QGrGlGIyu+jQZKVHj
M7zFWPovXmm+QdyL6/RcGsfgtXpqCz8x0Hjo+ens1LOhVmvOiUowe8My9h7vEPgO
jc0FcjNZYcWuCj6W0oMhN1g6YAAcO8+nqpnhnOrK+LHNId6kUo3emqgiyNiA8NDe
ePA117U+qF44mNU8vAfHtixILVO8pdb6RzAPzvhnzgt9Zzy4zWUyCPMOW7i+wuLz
TJMb0bxjxkWYhXEWLlQ+B+YwE2ha63J9MEOozcGU7LP4hpOhiyt5Ywo2k6TvwzII
blhB2GoxzebvmaVpVKFBP5ogTuueNIM/FOnZtJO4qVCYVNUzb8sh+3lXgAU7opj2
zhEM7bcaP1h/ltzV9j7EnRs/netJy957OoO8FRevUkf5K0knrVsg/OtYozzDudD0
5rn8GNMQxysZVQ7aHiGFVTr6Mj2Gi4SxWjzCWyir7PSWgVzMu4dNL+Ytiea5mUvO
1TdD+z2kqQrtJxstUELi3K4VZmA4MrHv5HOZ2QvmVFlAlumpuCfs60PyHncDxJnX
B8NASRultTW9KQ+aTWJNQhB/+7xpgCwL3xbeaIPwY7Ff6FyHRHRbASTVDz0TmpTK
JN5NK2clXezFWwP/v5139bmOezVYPo7eyZDugEtAlxvz+VsM32Ae7hnjJhAKWp3D
KCJ3eW55UERDfGLSYXkl71Qrc29INDD7Z7zqh/FodOH0CIQ9D0miDfaOGIRzMEKS
HCDdxDh9CrJeGr1e9rkROUryNkloQFCk8pP6qru0J63Ph19zGQQZQk0yDtR9jVzd
VnbnsprzHjyhnDxmHTnQvPUUbEX7HN2Y1UPevBFS7cxq05/AZlDgSpxia2IdPIPs
luxvU2y01Tx30WfgO3krjnMfjaO/eDOwkbXMwrzr4l5GlpwGKhSSYiuXQZYPXtfs
0CjlRwsjpuVxfesIlVNNSiC3C/pZfihYaDdqDfDnE4k0gtAURUrVo4i4x2s+wGjG
iHDVnnG9kmjBDglehoeTTVYjCq83z3QsQHQ2CZCOgRl3T88mM71Hew1WQmTwSaE+
AmFX/KDHQ7dnk8mOsGus5LjbYTKufT1zVCm6nz75Fn8lJ0NC32qCT0Uf3BedxrAw
1bH59ykGZaOjhcQvM3J/yVHnosty4zBSrA3hDXg6QBvKBHKImqY1Eg7DYQYHvS7a
dBw/LYxnpYEOLkFbyJ/VNjyYqOqJC3A1RLMmt2A9JBp/aN1fVI44v+Ta6Wi/CuYR
LZVJPQN+of1l9fZ6wh5cMob351mp/d0CMU7vuqJTsb0mkRmUDoXoIXTXHWKAFdL5
nTOThWQvlpO0h8LheU2pq5D2n9ByKV3tBksOROiLVTkn212UC9WPvGxIpkRoeZHn
Cidf5IxS2PPq/dXjtGa/N+ZBT4/6qqO7n7Kshqk4xfQRb4Y/TwotSIler8VcQZtC
0beBX1Zo3scDM3L0EsxsuqfZtaJjT3CQFsGrualnHW8loRTmLdlGmZviGVHfEjHX
Cw5Xn0pNazqDfgSn6S84u0kSW6sKSTGB2smpkJyXF8CZDPgDpwNK3AVI+A/X8r7d
qoniP3uRQKwP+JoRzV4Kl9StJs6v9edJGMoMpKzBVixBewrI9jO76i15BlxgLa8L
wBSe8pkbd3jJi7cRtbPR7ZeVUCloAOCOyqNp1evlngxhHQbRjpGWnS6YNznxMh+I
t0ZLSi2945pNUWmlJ1GJaCKx14VhkLgRaEjlXzv/NWOVjhTc9Rq831aXtfsP7oHY
BE6qa9B/7Na3z+S29uBKTxGblXXFWsJIDk7u8wE4a3u/UCpNTSspQIW8wUM+zO5Y
o7oG+R3/+lgVWdKjXcl7f5PT+4YLd+vD9XjbQX8mUDmn5Vpf23PQv04rhwbVm71d
PutIepQ3bzeDGJEd3DrvZELdgsabNs5xoMXn+6iG+lDhINMjnN7kcqk4xaTswOWi
M1OtCbRcc0UGZ9PbzFjP4BYZt/K0gBhr0bfQjwZ/6ONoT8VI+ews3xKZTncU/JkG
vpqG0YbscrtTBZRVyB7M0ZYmVwzAeohueCZlOgFwE74Gek2sF+QBcBKtVKpQ/JTM
zz5Nh3HD3uKsEH72aguJ3eR8jP0vfm6rKYGT4mwPAA+fOyD+F/K9Inu0LKMLJrBv
6Wa28YlQYyO7XLbbDsQSnm6+YCQSjmgiclsjRLQF7WoDTRIxq5oz3jvilRMouX4N
T0XsCG52EcCFBxB9m3xxwu/n3byyYuXB2Ikv/2y8BshS+8SDbs4iWIqRnX+9Onn5
YLEOjosqdnANAAop6nL0KWj47jloyWj6m/NVAqXrkB6CcEm8YEKfl7IjcLD0xqZk
8rQCq011nye7UcPbQaQbhIXSlsJvvxfwKfVoXoxOkNzu5sdSAnWpJbfmN4btpZg5
++vM2GEyPrL2Wmvc10ASnRCQehA8PDdkML6a/shIDAVMg0RED9zOJ5w2sy+qRWj1
jHtBpM/hVpzaM1Hd/kBdGvPkz2bkbDuxSp1hWJ6UFMOShFlUyLoMSRRr0ufsmnC0
QJp7dLukC1FumJFdzjvc8Z05Nj3JOPf+dNy5fE5HZhNLD3kPOAeYA89VOA805zUR
c9QjuZXH6e05/ttG2nHosUGEjhS92GO6ERc4IrAbi/XA9bo8cVffBgvDlKWgcmpI
lmveyof56WrOW+3VkRsRtRAoq9jCIUXCZJMIkmIqhgS9tb0S/FuIILmxdJ0WH7qC
+rotW766xpNSbf8Q1BJaxx49UjWUT73tlwOwOjIHc2JeF6WY5PGefIXuM0BBZWBG
BgW9DnK9Z+4GqXvkZpu4WDIX6lMReGLRW3ueCoKQdHvzXeWtcgAXwszOBxdt3rA7
d9tGNUrwXJLRSBFpTepXXgrGqnIwgNop2XjxudkI1Ci/XNOO5zQ1PXcO82XClxUB
NSgCaDxIdUXIc84E6JDgP4tzc2H/zdg/kedVh1hmFNQDw4sMbXEqtBAx+oioDclr
DtT+kX5M+FoIk4Fg8l2BB62G4+i8JP6FCnv5oKfJRDseMlxV1hsz5Le8VxftX9CC
PUDY8IJ2FKkE+lrEmcg1SoS+Mh9vMpLTRkWtWE43X6nYPMGjPMBkJELgOYK3WMAh
FU2vJQ3VEsmpshchBiRhXWdxVB88MKomrKzkaLvVb2tynkqbCxu9TpL6c+bmf85a
zR50sy88BlVVoMYxxXDC7SiOIVb+gKNaURO0SBlki1XGnpz4JU1cAHtusKhqYwF4
lax8ulMMz8ljw6zyMyDG0MWbdpr39s/4InTXprCWnG8NsOONCVfiYe5ZtT5R4BVE
n23Uuwlr2cOZ2fVXQiPeJP4DjOuh7t6GGhuW4jVwq9MaCvFpE/E4GUAAY+0CWPtp
2KaiwBWf2ebsvOnEZQ9g1CCH5ZM1hsbGALUwFS0ZAZtCqICfKMZEY7Hum7VzhMQt
U7UzMZjjPsJrhntQJS/rxpt6AWgw5ktNMoMu+AkWuE1Tkbit9vUCNcxSUVLCiGSg
y4JV6RBgJeI+PNz5PyTHyFqmA1aFqCpVH44GVgrMWCrJQ6eNnfFbErW96KGaemLe
fWGnvEL+J2tFeG/4NKuCdQBAVH3Zbd60ydMZboN865j9HSAYBdxmUlIWpCZV/q2v
sqe/Tgn+vH+GceZ3Y60e4+uHSteAbPjH94vvPddXUuo9I5wJdXsNK2e6jeYBxYcx
Ub8bGpo2vBL5aVUaFfs9XTNqqE8cMYLm+M3MEsbhNwVJiHQ58vcXpaebLn7hoHle
bqHdsuxnG8B/7qS6ZP2/PfES6dvptWOk2LCrLmZ3c1GsknepfmhM1VIUkkbiYLdf
vVyQliqVQHLOnHjNppUG0ydkNjprsyjd2tABcJUiRIWMnXjmtJRc7XLSFJ3kz0JO
bHhPRWv3fgiAcNTKKfDWUgqHLsMZ8ygEIWer7r5vulDqJqe6YIVX02DLlxSvCI78
+LtwNZAFLzB11D8snQcMKEWx7C1Xv2E/0jhsf2Dp+TV6LczyB34x6gbKWH/gT29H
Qxla9cMcpYSLdgFtzTfmL6Iol3ElrzSL+dA3av/gW/GvFVJf8qrPPksfWbQUHx/1
SCFg5e61/ecNNlrZZc1guWQow02IT3mA1sJluuFgXcMw7VTBXAmW7ssClgR9tt3/
/9d+uOqvCKpgrYDpnMOZA/vvm9CsHGzl/GUuBTR6AwUH/3XA8QUNg1lOMmpBSXG/
Jvr07b+PDp8AndlYm2eZUOBbwKV7DlzdNe9YwBQxa5Zfk7nYAI0mZryp4DclukQ5
AgQfttmchY4kdSKs5az26jqVwlJZGTfr6j4Ogg4zQoYV1Ssx6K3khb53NJm8SK65
eio31Nb8rwyqTy+SqbevMCagRlUxwtkueEiOgLTXfvQEzBmBLIZIjY5i34uexspk
VT/pt2DkIhx6Zzf1LYG6z79OYMTXloQp3z862oYh44Z4FTgHb94OaVnRM4gJf6H6
E0Sr5g6zeHk3AWR9C+oiLFyg1CIKKS9iG9YX1gfUAO1tNFqPv4kCPfBSCdLr/lG5
/kEf59qfpBcdtk+3O2q9ad5Zl73oGW1U1av3bYCygeMn5M6rzgk1p4CTygaQxlt/
p/UqqBVswOyAOAnpJQOMM1avxtXywvhbNvLx9xjvw1XSs67yi+uTQmj7W4mUS9JM
ZaTIdRqAxyUvzyUIs0QzWc65zASt5SjImnVV0DlG3LjWMOKUEeeyVdQAIyfHt1E+
PZ2DodFEej2IrqI36OBAlI0vFju5vPcWYeJ9VoGM9Tu36ZMmM+C8eNT5GDTAXlES
ofDfQqC2Eb1dxUtk401JFcmnNcGTnYGIfCEj21AMvnicXCsWQQ5Wx533n/fBmNI/
7/a91UVZPKZnCwhSa+1bMgB9NViOXSv++uPSsbtcGRHsuQnw4lFn4Qzz20SIE8Oy
64SAfD2eoWaO8gQYP8nOZeHqHkP1BLXcHZELKNEk/SMBIT+6juhvRaxUSA3ibLwK
ParZTsxpxSBf0eG98ooXUZzwvVzGuulkSkAdP/nvotH4g+47NCLfaIH/NpeG8W+O
1M4XaPUV6vwwYD6Mri6AoVBYzrnLQL2wCHxLmFHbkP3pvTYWCcOF0s4IMFt7llk5
oNBmLW+bskOo80VCiDci8G6iNah8TEgz7b2HLUSVbJZCcq4k1C8J+BM++lNwCvQL
F9UkpWzEffNIzo0ddvf33Q3SrDZuLt5SAnqLNNuTmOcfl4C6J02KjCzeHasCBil4
28PbEhUgz3N84/CWVCi2t/elCqJbHCg6nVJWcJ2Qr1QwWlJYgAVBkdyWwnGyPSLn
dfWztCC8dQquNcBh7/Sn/nF5SVBBCfbWg/24Sl7VXySFY7V+XWIx0q1IeGIPjCZ5
3ouDDs9RiGYzPUmRfsEkkBwI3e/DPBDt7s1VN/vnjXOmXvx+o+LGlYdXP8uBIeWR
CFtQhdRDa6Dgmun4Tn2+MALanS1WzQ5b/Xc79wKNmEUISfZNpDTNZv5FBG6XM4/W
GQduApPHbJ1bcbTb6oH12m92WiWwQMthUGcA6XxQJE5Szc4Zrpz2xkhZoaF0LyAQ
Tu3vGht+cyurjHWWlnzsRy90C5f1zdJCwpXP2AmBbfdaTUC8ejTicciZ+q2P1Mqr
8p3Jnp/NJoTEKd3fJuqpC8h2QbAXdJA2W+rKS0UIqwgqdCprTHTmzsBsJUoeBlNY
RnBRoCdIltTDyLY2snpqSCcSNIBtSTnifw3lx3mdSZpHeJ8qqk8T+aOblfgcPsF9
gUWx4iip41M7JGayZy3YtCdHF3zd7iTQ5Nm7GT1LF1Remow24zy6yFbyM8E/Y0SW
aQdXK6rBzUhZavZPQN7fBA/fSxzeIrmIWezJa2GCU+/Rj0xIU1LaYOKdNFI3BDXF
F0/pLJt0k1ut76x8N4rIJC8QOCXlmzv0d8ytLX3RBsXmd2FXGln9G2acyHGpPztQ
uNJopBBY0IMGwSBbN5hJ7U+7svkRh4iNBbJOPI7mmaPdOaveOQGnZ+xmAzJMnTEJ
gvdWXXl9A/1MQdPPxhoGy0od7K//fz9WqVzf0TGKfo2qd0YWBvZLwp5jTB1MvSJ1
HZFgk+jlBY/HyUwpynkrR/m4BLvbuL5WSgPzpgOVPL8d0kXkZy1PZTU421ULwyKh
NiJ+CvEfPkwZsK3DzscAhLTrBoxq1Ow0dEMGVUchL0tu0Zvwju3nyGpw6DyfEF9/
QW9e4f5FCKTLdF3u3485DE/w5gwHuE/C/SSBhL7Eg5fAe3yOprRUfSHXZvo4OmS/
RLO0ddZKT93v5jg53Vq4YUQUcpXdq6aDpPga5OV1xrNYeto2I7/Z59pkGkD/FrH4
z64nhi9HS1G9GVgWZ0S4wZ6AJVXbQJrqPzIbB+RN4JpSHTNbZ/7LMJ5KmtWX6grS
o8XzB/JYGSAPyXarEcLm7rJVBXJhJHadmQPFBAlkWh4rJoWOW3/x0YZKyuCvBGLT
nxReWSGrcDpy3mmZYE6U1G69oMsx1r9lkuhwHIgocLk4viRO12v5mqUF4e25wRyQ
3xPEoamk9XmmS0KdVIHdeLwsVdaAW5y12IzxRvBupoRcncVJGNrMa0VgGBvEYyZ6
IWI2WdCpzfVzJirRWYxLvsXYeEM7L6OEf/PTd78Dhul1t9ZbZXnXXnvgQwOIqTCe
5ZaqCzpk1aHJJYZYXXJoyXf+Ofhs0teY1QGbqYeECVrzhfi/OOkxCBBJIHmCRZ5S
HdCgOlbYdI5mo+vHJ0d3Styyr4vHnjZ+otS5Texksv1vVhg/ixWCOAyLALV6ymwL
aqkrf9A403QAiwcG6xmyth5xfRA4wpMCXtKHzt7Z6ONGEZJqol4gyb2Cf7tta3or
N+0RQOzyJXK54C7VqbJUr7/DXWRqjEAX1XhUJdOMwj3DMXKSpsqCicKMHfT+i6IZ
BxCy8rwTJgXlZ5ZcJxk2ZqTknVq+NCWV5iKbilMQsCRoZeFCq7SdixDOPWitN5BD
XRVNydS+Yy/wIRuxZaEe4VHyQmTj1oEom9iNBRkZp4QBTQy0Bdge/0CP54g7E7iX
YwWbg8tGuAfCAb3aL8pmIE+/w/ddoORqMQn7Timj/l0tEM8oRYZcNIH9VxaLOPQn
UPbvzlHFs8BfNVZ5rvRztzND9iq6n4vkDlBlzyJ1TpOYUuYyn3kzdHECLmwQXD64
INN3bq8y994TOKVFYREKeNquofXFCYqsM5qBuScXPSQjQvmOWji+iSN9kZ3u0CNN
YMDTs4zQ0OmatdnPR4QHk8gb04ZICZ8OyLJWY2XYwLit/6+ZQk0nQ8yUvQ0YEgqK
gn0v9hu480Q3Rj+irPVGzjX3EtujDtMpkslR3f8EcXDtY0qnacF3gQ/doSUNFMWd
kgyTTQLg69k2mSPbghhyFwMInG3u0ZypIF8MyHf1wY8w5p9JZobxBnmLKIPZfBX/
XBaPv/c2rI1HfZ0AbDvHGpAJ7hVieryiSYgzLtGuV5I8NkAASE/Xno9VHA9QOEPz
Ud/WAS5BmfiFaW/JeOq4+cXMKjrr2I9NFFavxZ0E3EAy3oA+/GbMTzknB+zHcFei
rrnGmY396pu1GKIAo+iVGb2lqUUnt11QUyKB4p2Y54hLggNhvAxcKuneMnIrdiTs
+ZI5I24pq5pL7WZWy8JjvUwmbw0clLypCCCR1GDwjP0ktSwAP0hupvK6SyW8IwUB
WFfaQP2TFIzXCSULcrBD11ZrZCG5bYwG9JYLTkB+dpz/RoRm5cFPh2CPjalXJJDR
r8lKa9qH0B9hYJgbfegNuQzt8M9kl3NFZHAvNoQfYWmDJdArhH28764EC0k/jU6M
zQ8YOWrJmXEzQ+2AFTAn4Vjf5OrVuvJkIbwnr8Xffp0foOQvWM/xQtT0+gTL3Ltm
kF2AbdYC0bzXr9oAG0wRx3C0tMUY9uGRDOkxiomyN9xl2St8IsucU9mWScv2VHBU
4WhqBCJtZpF8WlyWZ5IIvZ7djJGLOkDbHkBCodQo0WYvBKdNWyk7a0W1lrdcGZui
rB8m0nY4yTi57QuXCDc9ExyQpQx8tI9FElI7X6Vw5JE8VC2czgpnRWgilvP9vK4z
0VHW38LodqIB0fNKLYixFqpVIiOE0xTZ2IwW+8TsZUjGCu4PhEoXUolh/CTBk5lB
XGxB0ip/F5ziJOmbN/EsSx3RwEF6SksXiU2EU2JwQPvrDY7tYM1IWoYM/w8JbexH
vEoKO7R8ZahsfLjQBcmx77ugUvOd3nQXAwVwpEJmewabiWI7ouNXkoQltg2nrG6H
62yP0FCu4W3YmQvkqwSGVkslvJpx2IFmcrgY0XntLsZMiO8+x7IOJ7Ej1sY3vwEr
w9olAwBtHBcjnSGqDbkb+QfIfX7awcXUtA/SYlUj3Xbmqf7KZ8lV+Wgyh4wg6lC2
H0PfuUCNiC58CesWum+HfdZ41W2nkTMYkvB292co3BPKHq3AW85VkWc4/16sJX9g
vQ65TLE66o+1ObVlvZthK9fYcxmgmHs69LaRHPrmdPAmEm4iFZLcZoFm6oEjljiI
VmeexdOYWxwYVFRnHNGCH7ProfmdarlPb2LHj9Rrjh+FA8SxGMpwsnDmr+F++Kad
nWAr7GMUjAAHxTPbC2maHaAXfxzNieZJk+ssuyTIbTAW6spFnSDjKdmpJgodTCYi
Do3VPz6k55kfoZW50k32PXGyPfwS8ZJIH7U+CYsWA8oxG1FGe2PnS+YnbCqJy6Wg
0QnUsIqq9XDrWQaH4zcXJPTFGNzbmM33KnY7IQL+YCQAecA65zaI/drAJPoL7zPI
p1NKX5RQm6FX2y5oG3AVckQI0li0YYJ0sPiEsQmXu5vqzGgvpCsNVtwAyoWdG6Wz
BfvLprvOrdWotJcA3atRlmARp6HYvjFF+v464mSZd/tPZTgrAs21UG6fvYkEOtdb
OiJggT1f3/hh2G+8hI9jUKmLn7jXhevbUsZFhANp9FNuFtpKA58S+uz6WbdweAH+
LqXbesg1oBtq/3aXWS1FswHGYH5qwA/27OEZzcLTuIbPhFLWeM78JhOdsXKxkv6o
v1Z7QcJcpzGwwvO4v/Sx2XETsdjP9469/diy1z7FVt79EQU+jUu7FnXxefxElHbR
2EKKUu8qAjpV39AZ5uEMuZktiQDrPK2oOaMq8Fl2L9qvR8fY8LRQnKt5X25oXaI+
SFDgCsmdpCJfcP5yqo9bvQn1IzThCEk1q6S30+95Py5/N8coqGFC/HCI1uE67AwI
kv+fEty+u7TIOeo+TXO2IfErAa5RS+ggDTwBkIT9OxiLq8pADNXoMWrbzAqpNSkt
va71RFNmnDRcnSe/VbW2YEK3QWk+Jyyd1N+0EvcKvnjWjvq6BQKtRcM9zXUfx4fO
J1QH5UbbTC0TG2rDMcIyNkuUVUo+KcDVsbvB5rIhS5M6wj2M9/ZMMamauyCvOs2D
HEpc70zAvukdCft+2A5mgRMDMa7WsATSa9p4rW+0XP5ZKegKWi+hf08YJ1cHdWcR
FAYrpu/J2yQAb7ubu+1cxSqPxXEYHaTQ1TNPr/TXW/XJR1TSrKGQCB/6RVA2Rh19
MYcN+KLwo3VPBkk3WpNTjSy9jhyTTtmZBxpviVHjq8UxojHNWwanhHwFWH7tjRsq
3MAVdTerAHS9Xwx6IVGZCSH1OZvO/LfBXFsHXPP76ADMk7WOiCeD4SBK6XE6cEFQ
PCLj5DLepRBQ1So+6JPEuU1cdmFCWbqS90/Cvub3hI71RuZUmb5Atp8hWaVIaH1m
4GWHE+OWHG6JkUvU+rHTdPw5il7ik9lFNUYT3x1tWXuTPWhYQDTyDFMtmsTI7Ux3
WXJ/CEjuhDpUdWIwvOvbBGCvl44ZvlhShj3ifN+B/cIK0tzMjSzGtO1ICNqHVc0U
rsgxCQZTIYaJTRAci1KW26vlMNrMLp7YbvIUptNKqAfxrl4DuW1crF5ZanG9Cma1
nkLz0gJMb8aQQuJYHXfdhLfUSidkvGib7WJVKfxU4WyVGnxMy/LGdujo3jJb0cQS
P1XPcApzU9MHbI0VHlZAVeyejB6XFFJYXiVRTGF5gFAYTnykvqH4oLCfnKrKkQH8
nT6nrUQVaYh4XJslDEagxmevmywBuF8/FKc2AvjeOeCq6qmRUFddPuFaH5oXIDui
QKXg22Pp8aKWXxXLNlrIGchKerVXVWNz9JQtF0BXi3+ueJhV6q4FkiuUdIoYwM4J
UZC2wD04Zxtz18m6/FLxL8e+lhnJMWIZKIm5Gl74xyIp8Z+fTrX0cm4F0FsFomXH
EF/piNJcwZBqCkE5z0Pqqks0gGBtAD5pc99TcnQcvmROdW6NgylNcsrQxewv1e79
jNoVWaMLWgd8InqeLB3LtmJfaM14Pl+YVqY053A4WOo3YT5XvKd18SZJOtMWylol
0V0Frj2pRWLFtQzITVeOO3NiWnt04+qoYn2p171XPcNnBeYpIvLXd1hAEYM0xz6a
5arp23MBIIEDiiiDP+6UoVsyvFOuCqiGmgyQJTDgcDWN+1Uphn9XlflT+HrSa8q9
HqIURcvx+ju91wi2wfLuFG/LYWZ7MW1jHfgyTgSUPC2YBICKGx9lFpvY56v0zCNc
nNDkCkNoN7Pgxe2OilV+i6Jrv4YueoXNQIuGunJ7JkM6uo0/f16519Nfxv82fvSo
ZhAQ7QXyaJostD4dF5BCAVNk5OVYefjR/X4H7d8zG8kvH+ynnVvD3oLFBCfrtxwy
42otU90VQTJL5/X82ScoS5i1GtUwPmqJrvy3+5+OqKbV7mhXhIABYMbK52ORnS2x
FaF/KR7T2iqbuX9fIRwUaXc7aIHPmAcyDHqvRIEDkEReIcShGQixawWGqk+9dFy7
6RjbNXAiVV0PSbkFCYipejirOzpfUv5YT0F4Sv5WYm8Y0sAcHlXWAPDZK8Bc73wS
umawDrpgKRoAGlbZ0YAFpziGLXgQKXnnK4+nAZYITY2UH8NFt9sPrebabGW4W/2C
W4ZWsnJHjQuAbXAkpfYFTyh7B0ugBXMG5cCVPVOIJM0YLlkqI3kW9/RuvLmyn/ZF
O3FWp1cOPTyr17Om6XRh5jyLvGl+/fdPrcKT5UwnbBk18KCf4sCbQGAxGXK6TYrD
Kn/3t4iE25k2XgIKE3hKMV2myGIxI+NlJv5X1asVCc3TIIi+86NC4At0iF6kFXXS
ANnntIlXtZWyc0kzD3jhuulTWzPJm1tnbXlR0490JUI2bZEgbXnXsyFRfygA3I8V
ekLwk+Vto6PgUxJilDYDxzddvnv04smNf/4Ns9x1jW3eDKc0jX0Eq3B6YEVFUxz/
mAyUzEoDfbsswZoMK5KpHCbLGDX48w5pkXAp+XvOOz7AVbQXuhZ6xj8ot6aMKoNI
jKDqIlkyosFN5Ls3H0YnC/Rt/FVy2MkZMhpkea1+ydS0Tf/Ui1+OQJcAJOOY9i7t
h9GFYoPcp9fdNvo79AbdL7Bl3Mc2ON6ehdp+VF3N5gjtKNnvjlQKeUo6BMVzAvZx
Jvpt6WB+dKTBzBtJXT6o4qySQJ7vc25jxOq3l8GO/yBzyUBRuni9svt1nz4yCvIS
PZWDAL9WQT6QEq8mGKTp0lR70eBW/TFWDRhF5E39qZxkVJhbccPuy4jqtvFwDKiq
52wDpa6RM+aEk/ao5X9NXmDqMUys9ngI8RNJf9TxWaAY1AuDhV0TGLMc9M2Bc6vp
wxZ66rdNlY13ieZyWBrt63TSuIZL5ouBlwN7L89HxWwqi2dT6f+jWVlLpguqqEMJ
yoOom6aLLttbk+RQd0my/8wL6LO8sJRm5e65E5O0o+y7CQTrUrEEB+d0O20UmDRl
8h1R+4d1NgJqNTvUUtCdP6Wsl6nLGXryNXc5JAKxZ0PLMSe7kO/TVwKMZxvlbQgM
4+mcCZ8wBRF6v46W8vroAsOBsxG2JwRv2Yyr4tw20v29HttI1F0n5CMkx7ndNKEm
JHTU4RLUH1mubLEk1Oo3tvaAEIcuqLPtMJGeeLiKPgma8q+z+dkdK45FdUnCWAg1
q44GxMIC4TcKDA1XDxIxi8CU/PG7mP2WXc2FMaav0Qiod/k0fP+G4u9uCZcixeSc
kaugZQ0ixWskOfaCJUjxCNrR97Tb/UesNLLlPdYbdMc78n3tjCHnakc69vpdgR/B
Bcw1coxbnIdy4jT/mNd52Z+lSL1IuMDGGzSFyiekMv/bta6la8HbtIxv82dw5p9V
7cDwl1XrFbwhzQDLduCpeZDxtruGaGLNCVYpgW5Oswl3c/8fJoy2tlutWnM9rysH
cGO3E4qlCoL9W2pd83OqTpEhEnqcGlVX5glEL1Qs6tIiLi/e1N2uOOnHAkMsf0/5
z+s5sCTi5OQZV1gq/3bvwURRJAj4nuuzm8ytpZYcspfsHCSJseAuckNc13jDGGsT
vkirE+b2ES024BiIO/JBhu27LO3IUG/etLhJGziCAcXcG3fVM+uLmZXOHMWsesqh
HBGtXrobT1vzIHAxSPi2A1a0BUdZkiY6o6QGJF/n6ferYG/b7tElwkEG7OHDpBau
H7fdQSzYlOrowi18zL7KHAEhSl+fX85XGxkk+nj+OAVOpnxjxXWMUvlJRiWbg1Oj
updiWjuMMxK1bh739XGqBwjDmg4Y5qftFuSpNKuZq1VU1HTWMICKO0xPKu+YuSPV
+ZWVZ32EpgX7FBfLljjqHmMHFnGa67LWZU009IicetL1++//OirGb1hZZoLfUl4W
knP3OjH8gZbpWeImPMk1pQPKR8+ElsyIOiaQvk3vdl321Dj3RrMrLB6l+mOtUlIf
axJRMGGHRvKe4lYYrL4SM3GpvICA/w8fBJHm0EX70/RkqqIdJm9NdnqEfzgWfhWw
ra1avzOsbtdwtes+ovcZghIWzdZXKH4M7Lqh0OK8qPqUUnaChMCRuq8+tohiUbln
BekQFviAhcQX1z/KoglFfQ5ThLOWBeMd4xQbaXGEI6p1LiJeAmLWZmZP4S931NFy
4aGC6lobt2+4zsFyDGGCWMBI/y9J8zHbKfJBU2d0aDtzBMuG3Gci4rnUQLyDRHUb
c81Scq9u1moDQzRGDDiV7JsQEldHncGhvIT4TUI7WwQXE2A8oseMukv9UbjG2bLp
VZ0Ab1uIuII/re9Bt/0nZZZpmVj/9pXgeFzB13oEbPkxsB9lU399c13p3yEdltxN
g1U6qMUdu0yYtOTQ/ROeZufvMNTlCDusNtjh54VaTHTdp2hu4Rd1X2PdM3P8GIIz
KIAVo0fDSLx6qR80h4r9bqA8yg7CJ25OVTxsq+r2OhxsTrh4RQHpo03YSpvkVBSG
THu/M5sHCslBVtmcq9jxZsmOxNf/bEWZ5r9hLeGzUpXkdRFLY+vUd5B7caG9TbXp
/1Z8ejXDZy67lW6rWtEuCGJYE0NnmqhG3qzr6P477VxFhC/2htAdZ2A+tqFKw6tB
xrbA+0d9e9TpmmFPoFu7EoR5Z7EWogC2THmswJrbbgowEQLWYRgy31j0UCqV2bvP
cYNNdqNExD1uFg3gnlXDpJ9dT2wuUXS9XoXMF2paq9FZsb2gsKrvjkL+z+YIYLA1
dUGkNYzjavFn0ovb9l9Y74fsw4NlAkK8DlotQFSXAK5TbOOOWjpkoTQwX6wZ09Fa
y2Ypom8U28zAsV6zl3jnsdJvPOuL7UsDSa6gm7sJEWAeDmRi5dUrVCx+TAxqhDMv
UlSGoDFs4tRMH3WdLwdEknL39h5xnT8oRuoIt32XcradPhOD+EzHS9CHmiOhrgqs
JRdAXW/PCn8yU+X2Y7/j2BUYmGehACsO7waWfZ5fhAoQt1v9c7YeMHCsiL37qgN2
GmwPlkJ2hX3WeYY656Re7bQ1zUqDHMX/KZ47876SSap1KIfhdFKTXADo617fUJlB
2A6kTlHrHEH1tns0Uc3JfiNCBRpar7/+UFABRv2DeyJIzSE/0HMWRLRr6duiSuNn
xJuE/bIylEXspBuzG/wWQ8yaOgThdfQImlCmKJU957th0fTaBh/ef4oublCxUu78
/cZeM39ruSuFHmJ8XDOO6xkrfrUnAD/CXYfYShvCaD9TJYAfAykPMNfmqV+oliI+
FEWrxc6czqg2rDLN0YISuhOaIYnxVZ1OhY05C4EkMi7NfChzW4bSjIX5/E0ZzURi
hrd6xymY9pvx2KgSNNyI48gYTLOpH1H2znaAcANCDOjcpOb6ui36jvAY0kOQzDkM
u2G2yxpACpmdFT8cu4xZGo2FlxHB547/rrzEliOB9oDH1qTocMbLMt7Szc1sl3n8
RzjO5LYkAbSdcBo1DUHL7HFFDZGpav8PT2NSbosvfog3EfN558Ns8a/ZjntVvRDd
teB5YXxnlvXoe1w2SXijk+UVzPETZC628xQTMNjWUpXd8NxfmxQkn+/TYwUDYKQW
66/im2ykVvalTiGOzK/1UWtiUm3oL/Eie0EZDNerfhUNrbnfqAL8GcV4bnwHTilB
MPAz0VrM7y03Qd5aj3MYSI282W98favLXWd69SiXW3gTu9zlW+QJUJKSySre/l0P
LqPJCpBKy6EmgO876roTaEd2i9cmpF0mxGgU5BExCnTcfUu+phvacFbOVotDla3x
AFMBk4crGJge6MG9IClNUKNUuWhLDARq571cSZ6wgmykQSmo00gXc2mwWj7VbPVl
DQAVpqvsGaD0FthgV/7qb40g7umoiHDi1uKcchLjHUw92IU37883LUHDJmnZO3ze
NwC4pYpr8+Y9XunvmsYzEJt90v5idmDXrMACIvPU+lwQ/uBEJpV/Y29KgTkYim46
zUCv+a9L/9dfZHJFk6iAmN9wgh6tJn1hJ9FX8fm8FrmOJOE02wTe1gg55iiziJic
foOp7mP1HUAC1/ZaE0U8ne3KPLLipvMwbyPQOWn605ldCfNkrZXEmQresNt4ENw0
x3UCTEv32pARbiZM9HZ9Dj/RgYsvTH5ZEya6xUkBE6kRMwcFK/By3HEtT3jmTT2Q
5ZVwlyAHpCgPGgfuYBLE4IWdKqkhpOHzwMhrlw07fb96weRqArADDc6VYNzBYrJk
4cliUbbOglx4bklxhqr3s5eewiv5YHTyjdTqq23cA4e1qv3gi9Ske+uT+oGFylFW
mhtYn47IOpL08hOg0T0S8xrLu2EHAOKx6OlYQi06YhP2RkafWgXQQ+f19FBPRhLj
xU1ngxygfjxA2tCAG9FHAhxj8RIeow3cIQk3lkuMVMdNNx4wUc0uonkF8XTeGLVX
9dpxtM0PyVOQTKuw2rxVNzfST5uYzh+3Jcv/KKCbngr2x49f0torWtQ1JwBAn38u
zbw42iRVS6P+DaqY9D3Mk1dO3KrRp2GZiC3eqkLOznJDmxenfdrHDqjz4hi2jXuI
jDh1RlnlLaC0oHxjwuDhYuvyCfS9CsX/IkOUNAbUy/QO/KgQiQwLdQxjW9SIbwv/
HgtobXnyjWvTRxk6K4efQQMCiGhzlbLx/H8bPck0ZzJldVuBm3CZBfymdbUJpoEJ
JvcTCaucQbuY8riHqij6mA7OiMRBMPlWnZsCrAN2fkZ3iIOS8o/jVmDuH9RTc/96
1G1+BdBhyehelXfEKLuKznKXTitC7zpPjkfJRTCm7qLXFbqkNTejATdfa6PTDDLg
tnebxdRBYKcduBaIvEl31cAwFwgVQ/0Fp1owNUQ16akexHiU6B6KDX5MyKS1mCfb
ictaBwILi0gZ8b6Sk/nFOIcsky75SMFXxFlWse7d7DCzkWNI/EkIbxPS14XDFqQ1
Z5busL5VevS30AWVe7FwQi4VEqpFHDg1+dsLCaePARm4clfenZJ5uO/9aZMDtoin
0S4+3BROPVz0SXI+6qAHXKlznGzpVGhsUcOC3g7t2s4pu3Y7w+J7R65b65H+e9uS
ZeQ8m+a+vTGV1YCM+8Qx0bW2+mn9JRuI/U04TkRc0mfLPBCrhtgmsw8T+L3A+jBY
tQ/xEIHpCtY69H/SQwSNuyZcCdRaPX3pX0UeOjLvexoknNfFvKt6I7GgRmBAeDPV
tmev+pZ7s9GVpVAEuRh0N6TXdtIGQKe02RKXQZY9a76m0Ty595Np5Hc8hyi0it1v
7FmeRRkyopPTr/EQAio9IDrbUUgcyb5oWewX123GITPTteLllamqWW7JUP7P6NYk
iePcZRJfexKzdyWdAKyY2W50Jx+uRFxLSqg0XfYHQOYUeZ1li2khE2Zhal/5Q4ho
e1EeCdM94/a48icuhj2W9U6ev3qmY/Gz9Aeq3Cr89gDTLt90xdNj4vODY7fK00do
rIPJCNwDwvO3u+/25u1xJeHmTAUk2bkV15XJwom7hFrkmjl1R5KcQceHNK0FF0Yl
2nt76VGyy2C+KTLesCMewatI/dl3EmgubuC7erLg07o8xGTkntru3v7XUhMpLjLg
6Vr7sBIA1gcZedab7e+7MrdnZd+VN80QjGCFQkOiTIO6hjsf0flLkqscBQ0TN5AA
8pbqsSG9YcZ9/Ak9Bu9ldHqQGWLpvp7zhe2ByQ8aF+J7xPKzMPu4xImV+R5UDYr2
MZ66dnAdEQjfac7KVAoTOQc2uOFUNsSO4louK6WC53zByRjECIsZjxYtw6BY3dhM
tyF1pUVDUQvmHILw5I7ygQ0eN3TwiBxB8GaNk79BlzVSCnSOTBmp4GSPH0Umv9z4
14lAO6gK5auaKnH19FwhTShSpHgYNcq/y03duO2aWBYouTcgNyo9ZBg9WxXmpnPc
Rc8txdlBJ/aR6XISFDXBNMMsejUP7M5/L794uMfPAtAwBk+/rIECHsULwABN87uv
eqdBDm+JVt+H5Fvx/XGqJA5yDejYcRgBtM/skgEzN8hjIFTF47SUkHxZnfzRi/An
zQbPafnulmkWJNmxaeBSGpnYXxSie2Th5pIvCApckwR3Vd6nFQGRnnblLqxdkvUm
II1Nao5F6kgCq7sy63AZFFDqjMKYXxsVtiWGkJ1SRae16be7rRLE3tWYDsUosh15
rF7JY5T/JejVlbOMc2yTsIgv2dvU6ATclSaSTbv851WDbUYXQhi1WPwUVyyC+Ibh
V+zuTiKOGiKJpoFlQ9gX1C4aQIBnIYUlLjDlHnzHxSRsILwDN4g4bJoGNSSd6Zak
9+5pq2YX+e2QcKY0emwSuypxvS0hhe4dtyvCXvXAWrDZnEQVlob/80jrJfJpBhnb
MUcBo/tTVGRwLzdFDi9Gc02PH6LCJHIRl9JS5Pu0wsbWgJJwfMz8gB9sfgw+231D
5o/Hcz3t34LKt+6bcfD/hJwFO4D+cczvzIcZ8PBNeSN4gCxOSEGa7ndW9DSNrcl3
Wy3fWy2vGT8942DmZ6UAqoWPpPz1mY6uDYCo4gq2t0v7IjzdCbfx4XBDvrfRJ7/c
TjUZ0XfK+FcL4dQbV3wMEsCMlXZ3lH/GlBqAkV3qPt3r+8biFBNXgp3pfETgpQu8
+n/qmX2De6N4ekSnEojWfR87tGYlywfgJTKWLb7s4yMvp+yu60BdzrZ2jKVxpUe3
rCsriPPmorkW5iEfs3UJlxOORxQvDYg6YhmffuGdoj8/LRwHi8Cr5mtC88C3Obws
XI8vagsww1iOUErG1KeiDAZ7RkY5msUcxSG6gWMjhx73Ht507q/ovqEAbkrqaMih
zgnTydWCBAS/h+G8ecL3zLLlvH0L20uDSFenpMN3GjGko9IG8jiQXNnhJ3DGPWUG
KzO7IMSjMGl3sWsLoBc2+9Kta0E9/W+hbpWPnQy+94ZTR2rFbhW4tkA6vlHLlJ0i
nDhtQ8Nv/U9v1PmEr8+vNtgZt5DCFtj8Tk/W2kLzQlBenrPVKdjIfxNfy9GFEiJu
aijECJORtmx9EngOglinQWALme/GJAEiYsrsV19bdu7QO2SYbQ4KBRJKA3my+tVA
NnipIL//sMYLfnMQsBL2k6X3hbYdOyddjfur62rv0WQGW8FlHSW4OboCpe6LbvTD
5uJtMbGFHrzbQxxiEdLSfY0UwbZLJCrKhyneTVo2utdRapdEloFdIp7eS6Tcpwoi
n29nNKzYCSCxRX0Hj7CS8+5BHWixWDrJHS5uji1QzlBzMzat7TuxRbulUCchhtd+
ptDNCj2b/DsyJ4dJpungB+FegbHmYRZoFkLPx6ZwPwdu8mXsT8t7d+TabqlKXWzT
MFET9xEL8GMhXYFv6IhdCz5NxmZyBGOYQmPsLLF6tHQfQ1NQI2JsAjePqzNG39cj
D0lTE0xdSyia/vGho9j/l/WDZy4e2/FJ6kyJonTpkxRylRVeiKU/UgF9I96695wQ
3eg+1bKCnKyIPmYwgdB03HIkwXXllv5KlMagWx4p0rhsSxmzgpGe4NOFHddL5rH5
cCyBfH1DyWF6WzDWjarmejPpfvrALySgILemFOerKxAAmzh4zXsYzMapI4ROWcLE
mB/40ApWId/maMgZOYvCMZDHLE+eBM2DgdUIK6PTzf6SpSor2X2byepZnFdlBNNO
hYnH/Z2z8jehVRRhoEsabWUhbb2BndrTZGDD3UW+dzrEMYb3A2mtoTEzUGTwX6T2
KxKfn8je3mUuB6yKTM4S5owvIn2rbo8FgAWtsT07SbZyBUTbICaBnezC83dLxEr6
0b0F0aXIsGiBRrmuGT2MBdco+R5BysnItzrI/3LpXBzo7FUZzZUbGB2kFTWRS1NG
0MCVkw7kSNIODhsBBO94Tvdso7dxDIJXh2KCYzqjI0ur8ZmXX0H5qDkJJlPlUGE0
WCQw+RogDfYBrsTVc+IKTvDCy/9VreihkHlXz0IG/KZTX/SmaR9jloVaZ0V0Z8D4
qQztYK8B9FTBPPiqRj67BRi8Zi4QMPuyfVnXgEWw7zfQNb9sqejUfT3IE/SZUlzF
1hw3m8YjC/8FR3kyXBC0IMDRTIOBf3gNeY3cXfWsZu6Gv3+Deehvi1q1sAZookc7
F/xjlVijPgJnj8uv/bPT3PD5D4NQp7L+6LtkWVxFMbUBA7eVl+7wlsllhsQoQ/8G
5AW6MRZ0v9ZCSHchL0gUymzrPpZaVUlEY/nlHanI/s3T79GjjaeY7Oxux+Iqht0u
x0mkVBiTZZ/ACc3nnH1zJKS+d3zk4u5x2+m/oVLHVUP8TujOM3Ujo/r3b50EL5ur
s7wBvGQyDIEIZDh53ZfjS3HNkbDySPRPfFF21LygKogElGtyaPabVXWMM03Jt770
uvc5IjSsARXo+8EqVpzWTgBpIJY9VknZtIahiwJNvId7L0AHcjLVpdAGpRZfWU5v
7Y3ewSeZfTryoG0xKdLZJEQopu9kMCVZYZNEwilp9fcp46+DcWBRhJtNvvA2cbj2
b2S812X+BaxDg/YSF/h4wFUr7aKABVQLzB40UcuBpEtsR3ZbzGdCYl7/EvQMirUn
My265zlZBJuGl48Jghpn6c4If3TnsLjX43eEz+lC8aXRw3RDrvyiFqU46eOkMTNb
HyE1XzMDIdM0WpZlnD+tGgmPFdqYpArB71gF71dY0PPwxt2p0AucYu5YcUXPDNbU
KGm+UHkP/VMxfoiAN11whT4TKLC4v7SGL/oyoOOveNJbRXlR6cCXdUHaFrmWur5K
OpXaHQWcFE0sVccqJnMvBPKCeArO4+TqrIoke0XrqLS90YQti+yfmQI2bwb01qIt
aUTEMYMYJcya44MOCODcJjKDMM7AZtpz2WEPL8wnXEvPi07Gx+o2Kh9tmxj3aPix
MEJ6evdH5M4rAGJViS07cWXYygZ1S2zsthSk9S9XHylgZihIDPzoF62PJk3EnsUI
RIROcp+qv4TIfSjxRRUGM46BbC9uJa05vLfk4OHuxl6ElO7cixarqg6AdiBxRqm2
e8Poe3CQQVWXxCBCDOIqkL7Ap0zC1I4PArFC/GgWg9zqJ303CYt80t74zbuQ62PB
xoptWGE1g9RBNSkwfM2y4xHlwo74M2CuJ1AvhFoNmkdbxrk1J7mlVyjNDpqHpSBT
ReoZ7L22mi2Jk5nBuHwnmTqrR98jaDm6BaJl7x+lqqUHvNIwLZs+6wb28m4z5MZO
EtVW+qnOb97shX3WnMIx+10VvKSXiuw20CTXF0jwFKgkrEDGwBmxAV397DBni2k6
ULac3Zrk/6+G77ljIW+ZudOVsFhpXFYkttW2QM8ETSaaRxqBYDiEYhbMNvuildUi
6eAUtiEWjQompqK4pi1pR9e5sD4F3c5xYFA2+393ChMgZdVHihaHn8/nek5/kOeF
IPCk4fwFetaQ+vU0dCc8DwCh1hRfif8htI13Rcd2Q66YzzLpktOfcyHQ+jNBzW2t
SDAYfXiCHR9fvRC+nBG1BK/UJsEyHhIReHO5GvI54Ozi00LDU5UqH5gwW2p3fJFd
Z6zxNpUyB14UDGSCiQTa0ARE9A5ZGcsZr1SB1B1ckUp2TncVwJrG4KW4zXy/9OfC
xUVbbYo1Bf26TjBlFFFlfXjbuiLBUNCxDGmzndMjl8vqjw5SBho3FQ9tJQ0W71yP
N2BDjLk7pZXxdFxmNrnC82XO639+xeeoRZv40tV1pGmdDuyiIhrf1ZzYfpjjathL
bm4vlBqM/eYicsmW1WD4w+kX1FNzpAYlw+55xfZTd+YC2ReJ2cY1yDkdFOoYYnT5
bm0WhV+uZIzC6B0qaWExqXhxzW9u0PAIzbjEZFbjclDQIxFCqliGTrnxHrpqNa7N
xwmfmqkxQcnXaVfdeer80YlTYkgwvkSFzJ27Y9i8EAjwRtTN3DRw08OvKWaNopdG
61aIrIkqACejSncU+YGUz+FIjqhKbZfhHMzMLmfh4a2L00cbAU/yFxvSzA/NUVcp
X2M3hTU41wXGzKkA2x9Jo+ooQPd1BPBZmWgzqpf/z3jJINOqQ1w116PgxQLjW63m
hOH66Jjx/BqdlTlHXE+HXzpPTU8hM+tN8++0o39oaHFVjhrBD2vL1RmpaGys20lT
aMGTtTOPs3CrUf/RFxFyx7eaUS6NTIyrvSsWlRanJ0eoHvGHhoKUgM39w8Fq8NYs
kSp+vrXgJxPLoDOpViNrdgJCvvooE9VKXvr7jC0Ve0U7r2vtFDaA9jeX/wk7h463
HJqV6wdywjgcMwaf9ZxETj/uY93BVWGWInsHpwBf07AFPX8wq0FHlKPX18jHwQwc
1KVV14Fu+CSlEk1V20auO16JCHr/QvWXGjLREwlNrkpsmCrP5HwrqG8DqPYP8IXf
uOpNWY0U3fupBzIxuunndkLKsWRyMI+6nLZNqoOWXEa8G/5XswMPYe8RogZAc3UU
OYdQM1VBb1OA38UCUT47et+PGu8AoH+L5qOdf2sjMw7yXjK35ClN/G9GrDxyJP2m
RYYjZ482XzZozkbefsG42N7ev90xbQp2PUCfrw9CzxJmWZ3DECXFIla4o6PcAbeD
F7cOZ9v/I8bHDloXwqT7bIzNCCRJoD6qpkeZsLi7FY/xZA1qi3ehxUgXnHvNi2+4
XiUFUjh/sKkiupE6JgtIt9PtXn0I4WkFp5kuZn8t9WNTmtpkpKP5UmAm4r8Tm5Vl
7j2fgffbLB5qBd84EI4lcfE/mMuqncmTtUp684uQ5aAJ2dgHtteDcAsyiEEpDcmT
fA5q8knqThdWvAj+CUUJYoulVFfWht7cI/j1GYTu8vrel0pquMUR3Wy1TDT4koRe
VH07t5vNLApKxMl9C0Y5HUFCHtuSi6JFDYlXdZpPhFc3Eaz0T8Er2mpkd3zwb9qb
IfRnJwCkVFj3MfMEaPcD4nVXwLbD6VofS8X2cu4z5EKg3pLFQ1csXPDKLo/zpVhs
xG1/tEx/lX+01h2r5o5Lbgdn1tBtCePdb09X6u2gmeKTjz5ktqKGSv5efYqLqeWF
6upP2rOWjDhP/jRVmK3aQUfzlT+1mYWTFXxySGQ06nAhtngLlVJgBja3RN8fcFSU
z9vYins+sXTmtDqwg6wIYR5sodFQA+QY2G5/ItWhwEm9u4IP3cor7nXyGxp5kQAD
rUm7MqacEOHKTTnDWgBbusxXASM0KEJDVvFn9DQI10mjbDwBWyEgFZTfWW9LFUb2
uvX9+/BzKIrYPieUq2FaB0nWofffrHfg1oIO4olfJ1YDeQOz9a2nuXoaG8+Es9pB
vOKqH92uauUyNWwDONBIjIXD8jzsygCHp4QDDXwsyBXewoMERe4HIKrgdW9iX2r6
xErzDZWCAk5UC58/FvSzY3cu+TlN9BtDJGNeZIwoECrlIJgsJsI5wPO4JcmLA24F
oO4gZxNP251QLUJQyICndcXH5cO3QlFGRvc5CkhihsF07OJK3Tuxyqguj7R8k9/C
/xKFRoQEwBtTU7uoJxCWbe1UlRORE7m8uApjKfHXbUkBfdt9e2o2/taasy++CyVM
sHX2YfsNY6WFdV77p9WmSxw/oEqGtw4O3bZWvSylfTKZ4mjHalqZHU2MdomRIgN4
orHHsfl9NTLcD2NdCS2Wg++O0sAz0CvHu4FxNuZtza8P1wQRAcwCdm6dcX+E821c
+uEemjc+KvitfHTxB9IhzBxn5w59/T75OPnZfkaj5MySr/Y3nXf6NdxDzPizzMdL
UeTEeqXKf56UeoHPxG4vN++YRZy2J7b2xInfhDkwtwqxsMxZ+tYg2FtNACmWFF9w
xKlQ2ZCrF1DycOUcUsQWr2DnziX4fBTrMCxT5qiF9qVrF9S9dssnbYANXy0Lo3Wq
tLA7HovWp5yNhHydM+DovhTb1zNCVa/iEEc3+PWGaJCzENXLdBRULJYNpGq6TMor
HtIKCt7EMwuB/s1gpqeavVwUeJriYmVORFgC8R2Xr93UCi7gd+nSMcKjVNDMjREa
1mqQ1EoVFWyyjRXQm7cecNnjYgvs9LVZnxmduWRPav44hZOI6CgOXv85kEj18tzL
SpO+GEtNUpfoL/T1yLcgqFV6Zsd0Fj047U09S/AWbIfXKp6LzAjfi3F8jZGhdEuI
8H/u9s7xrW4koH+RXJhpPYgjEb+jDuz+eb2l/5efX7vsZjPgLuUPseycqwLT4JAq
HtNQN1S1Nr12HShtPSleh7ui0pBcX2v6ogE4V2TGNGlRxxycxxVFLMjtnxRIGjFS
ofWEl397dB3N7E70RbRk4DMP3PUneeTHYXGFUoNYRTVNi8WP7fjLECQAcuVIUdpA
VZgIe9buDlCz4oe6j1tB7KMWHGDKm3OCXG/SMzTRpTC4RUc8aze5/5booO8sA0ou
31g4TwvrUvRDDSWzXhQUB+xlnxvwEVPh1jwI5rkxNN5gT1kuzvgwPQIORiZpZzGR
ejCNrScvNrgBbw1nLpn0Nh1EUDQU3ir1jf86C2hMffAMIfj6FIdh3ruNvmCiFo2O
AKwk7xXPzNWnymEZf9JJyrjJFQbRHQAUvp3JkVpdN97D7AREydMp4WJPTXvbkIYJ
12XDt8keLebH1XSs3MHNOPGvx0kYpT12NI2S2AX4s23/1OTWXMoFiATyerSY5jop
uXrufacSbW9fylcPnfQi4wsvsvBZEOVEMNVzwJIopthPe9gz4E6qwV+CGuQpO05e
SlVOTdsHJ1qMaPMrTiOxqaa9IzPi8OYT1uXqu421PxHBQhOzYrmE16GV2F3atJPI
ahr+N9x9A1H7rIOrcnlqxO7zss+UGI7G3q1R5N9Sx3bX1lS9w4i9r95NNGY5E+TL
zHkALoregN5xj+yYGB5BEH9aES4ibhr6vRafphNxxY2WvZluwsbyn24OS6JiPvWY
cTKYu3le1SatUBWCspNm8zh8MMxB3zftxYs/+xMNUdAMohabHNjC5Q0F0pC1TDYz
uwpBF/uoWDLaLXF/QxYDUbgcnudFAGVGXTQfwqvtb1drS0X9NXSgSSLLUoFTZymx
5VdA3Q2f4MS219uzS+CaNFUevgKNoRItAVnXeetNk/iavVS54k/XJL8Uktabfen6
ZdTJLwaKDyYtnF7XXZBLe4N8c7CHYmYd/GSky8l/C70YiH85X/IDPAto/kk5hoXB
M1JwV9Br9gG5mhUD81aYggUad1At5QPJPzN8hwf7KyHGmrpgYxYYH3S5M4NdZx0C
6bqDYK3kz7JWvfvWZPnPznl0ECkZkFQtM5AoKre5p7vpw2skJro4oWSbYKcj/We6
dp/c1Yj9TmDLoGjGCrl+IbQr3TnAV4KNYMKv0sw8hAbiT8PLvqXeITmCFqyV4Umw
dcaWpQ37q80u1SvDTge2JW79/0t4g2YQfjhfxpGx/yq6sUv1yTRgAwEMxapoTjNL
x35XdHeZkNe2qOI8p9rdIzcsfgJjwuwaiAAHVA4eaCDKNapR6z+61MhajYlf7Nyw
rzx9t3mB9Vd3xjN3cFYtxR7ctkQxCWOBQKeoSxvSvay5Q3dbjtXjR0yFdC12pJ/5
H/HW+bR/7+rZKZrLKF3aE5z1yBCw+N5C1L44lD2bqKkIffb0ggcKruWk8BXAjlWF
70ndRXv7l9XotXjZ8Pitr3L0ilKVO8sjD4y6Kaz72OfZ52s4XR0i7Im3ZkS19j7Y
TqF+VeKk01qmDVkgNpEu0pf+kJbQZdQE3pE1E7WwHcYNFeN/KTJnexeuX5LQxWaI
21xoVCEa4SzXGqwkiGK+rb3WvN5mdJ3f074+/bDKpzHMDqnC3jzY/aJdacHhObqg
MTbUJLmwiMmIr1kmpA3MJkFabmQZF12qfvrVg8oUogucCf1KzhvksmSNHw9Pn3kZ
jsowwoi9jrXU15CE+ShHXn6kbEh7nfkpgAD0EJwODQtBXF71xgM7KRBaBDdpaxOp
pTYku9rZfxG5BEcARW2xb0YUwE0+5YKeQTJbRXTamN+EG8SwSfxEb47LDGyxjnoy
Q1aBkLQ4xt2pI3c/ext5CrusCydB197ky2L7ET4N9bVbnNGZ2RtRbBq651rq0uE5
njcJfGcB7qi1rKrAm/HtrXAtzm48+2tlbhf9veYBjJ5uDIFa+uf9KkSLKIy2Xx48
P8CgrNal908d/+RWI8AegcFnpSdmKTvIyhF5cwsw3ULPPW1vtynjGBvvDBVvkum/
XS5hTq1cx7BtAlDYeCv4G2O6xGmfCFejIFgrsHAZ11gJ/fdwI4cNR4lgZBpYh+6B
ED4wK22tGQgPde6SssBYMhDUlgu83RPoSQzl59noHhO6aYEWz7prQSlcEOB53p9z
ihFlv5QapSFLYQYaRx7loHIZv89CMDH2kNAzn40colT92PwQkhHQe2GQspUSIwtU
aL0NgCKlpH7hjUh3TkFR379lqZ0LjIpERRu58evaOTjfRaYzpF+guM1mAj23z0dZ
7zpPqt/wSnX6rGlq7uIPgLtz+mn/zA1rL1OacLAqgiAhgP9+/j9vlKmerPVdK8L7
gPLF4l6vlut6HMixmw7IEjHuBzb/k3Uk7TWADY628Bu+yGL140CEksXpcH9EG47v
X012fARG4Tos19UUs+fFXeB2RigXC/TBj49SGy+gC3AvDbQm5jQGcKapIxAO+grv
hlNSQmJ7DIesEpaTYyOUxjagEHVKTovFotCUKXkJRZPDwqH7yKtzwOgSFBlkjBG/
1prdT57fSgenW7WcnM/XjImSDhg6IvePdvoC5g5UsIj5l2z0G29t0G84zjqbWbu4
T5njkjnHRS00SDW3sLHOnr4OE2ZMJ5/Y1Qo3jAT2QG0+2fKQeKEocVVmx0FQ+NBn
q9H4QumrU6Z2mY29Dazqq6GIs0NV7Wc6+3hyn5URuqxZ1V22ZFuSdzGJZbDr0C+K
wNE7UVJ0cqdkyh+HLdyfhqyDA5mv146c7NqQHcRsvDJJNCDUNb//wn4AnOAbs0eo
nEZMzRPDejV1B1mbmJT6UIl8cwwJOyh/DLb5/7E5u/Jx7xCV7X+9/NlMQHj75DXa
11xOzVahaGsQBSQsDoQ8j6sLsnn+btQiBpY8deJCO8kojLdKADciGCYCzr+3IxP1
2xSaaj4kdbUyMQkn3FuEl0gXvXgw8PbpOFHDImrwjCcqHFcIzRNnndszDNj5iKbA
SriPUs4hV591Q6TKyx04ZfUggilC9uqnsTugi1kqTgPf8Tu6e1UuMUTuYPuZ+58j
a48Tg7OfSLJKzbUqnRo5LMuxnU9BwSp6GGC97y45vXLNYpaXSMCJzKhQneXkn+u/
X0Bbi4iEG8hyEO/dWhb3/9ahntNZ21Fo7Bcw/zgPxGGyQEpMW9JqQOj+j9ZFrbhz
CdM8pCzdcGLvAOnJNNG3MuSd7KiKxdFtVW//qmIdbzGoGkDlnd+1PhGZq//XyAJu
XRvgtCEhV3j1tCNYIT7Ie7SJXtAhgPPPGQU6ED/Po/X3n3loFfZXUSFj9goTshOX
Z/LB1UeSqI2nedqz5+Vkb45snUrWe4lVGUKTOV1srmuzePr15/PcaqKND8kqfZm5
c1Sa50Hr0AUZwIW8no18OJSURncGzFZhouH/DBmkQDgajVfMB+j7xz/F33YwTPre
zds0EG+wiSXCzgRXOllItKssweu7lgWF5bF8XUZ5d2Z6fUrnPXrhL32ZmC1o4ABP
mtSeHEmXoP2H63VQflysL9mtbNnIdlXJ4xEtmlhioak2ttCTO4pHeQFDjdYiXtug
7TFWWBGHHQMGxVMQOzXdaulFYTpUzhZPdnvR4mrbus4IIcUiSlr2DmmVLQtbAuJA
gG8MgG6cGwbRTof+SwN6zUomq23rZ8iubMYw23hgABOkJNymh9QfzMRU93eM2cu/
agH33pCnPU2SZ6qIr49xO60IEOghMQBPBdewkMbEr2kB7YjWqXuTv5R2mDtQlL1C
JylTKkSlz18Lf0V1kBugVBu8FsQ4dbWI9baOMJc7lIEhl4nPbu64SNeAWMMWygPw
AAA8NhOCaaV8lGzY5gEeLpT+AxMS66LzlJbloCd9TkH6z5j1JSLSpgavmKGzeIeF
H9FUj57EPLrP6EtuZsJ3fQSDv8XyyKM4SaFLsLXwoMBBDWViuriLTCYT2d6hE2DI
y99SLr0zHKjzMb+AIUbKYvN69zY95FCZzAQGqmTVdtdwVAspG/QKVecslTC05cEF
xh2N97w/T5bW156HGASwO5uraio6s5gH9tjiyjxi9ZoqjURW/oEQ+vU3b1F5QqS9
JeyVqBRW+o0oet4nVYUjGZc/gd4Qvmg2Bbflj8wX4HV8Cp27AiHgap9xtfTzF098
EejFWycQsGflmS7rmonfXkgIMwRzpif/0VC5vZITvg05bRboEfK73tMODjRK4GTK
dp06NcupGr/+0YXWGtDvtZu9Uic9WiiVs96tCfQIsyegvLoonQfU9vjgGiPZz/P9
z1JT4KEPGTWrLdvA95mA3S1p3Kn+tWlKMTIxymFiQNMc2lYchCmsGaqvqOm2Jm9U
NrZkHmRxnnT2+Af8O1HZJ1y5BHyz8/Lj7mj9tGlSqPSHSj+kjmGHpvyZAm0awkg6
alta18zDoIsd4EiKfXtsCG+JgojXHbWvFD9T5u1RlS5CzlJZp756ef5cWhbCQsTK
WX+Rozkl+a14/9XuVyYa40rOJwNQ4MSThWQaHaNStm7qFInJwoGlN/T/Plc2+DPg
SoJ3nGYR6c3DY6RhxnYZ6YzGHytnntEWLB8HW1NzozM/2vjf81YbxtjDqs2voSOI
BuTJY1RLHqk1kDG9d7c9b2Ke5GXBJTu2B0l/PCqp++6LvU3rvmf84qNg6negB0jl
ysrM607vx/ZzIaza08YtjEcAlNsyX0WXbO5+gDFtMRF4iWef+DAPBEJqXGoSBByT
ikZxTTLAXZjs1ZofOyTe2juH8M86MnBkmiwPal1KZDdybSoxnqKNID3NDPGohtUy
iG3ktYD2Ch4WIMaglkFdmT1xAbfPrQ26fFnUy9sYDPNW0c0PVQRUi/M239Hdv3hO
J8lnZRsZCYnWiwlYt7Ov6ZrSKGex1hF6dkBR8ZKGEpbc7FwYOunKl2jbysb3D3El
kaIHj/EKMtjJtieVul2ZtQAbcfFTJHkoUuK2kx0Wh4xZ7W6tDkvJEzF3mLfKet5j
uZAiuX/bNKdH7cMIGitPimE1plN5lz+PnX01VxH3MzxCB12n2N/QvdJ6iNsC1EX8
oI3AbcDVNEi4P1VU6MVvxQZAu6FRWFKVrgFVOlbYAJChfHBx/Xl47TGiWiT4U+OH
YM5zZr2preZ0TqffAc1jYlYYqZlHF/acDOw8JBWbluT0xTXKHMeDMDCHeSAerp9d
zvNfqk6HYa4fPH4So/bY9ytmPEYW9DU51w9YdzPv3BfjW7I8teAwiIFqyFuInyD6
HXVWVuJBv98WiqZXc2FdBsxbopExQ4VSImcBjJP/qoYemUdGSlONzvcZ5z6cjpTd
PwUCOBdKnihD0hDtRhLVci7TRaG20OS7UsuoeYDJbICU2vGATsFh2/f//N4tbcj6
b6kQkyK/QXCz0LXGNYY/HwPmqrSTuXSZqp80P4YXCk8yTpoX2mmwfcCVbFndXtpt
g4GLOjaRYpl0Y7PKnXPAMORIVGUDp9IYEkQNXIdxY5oeEfXPvfNrYJSW9VsRVAly
ie4GyTURSk7ZIeDfdgStyZ9xZ7Q61CVvCFxiWSIqHumx5SOYl3URiYFq+uvMebjN
2Fm3GmXXDjvIpHm0iObL1lsil3n3cfdni84THFQwvU8h2kADGGkGtLIblA8By+PW
tEUz1mWdIoWkH3N6PyPAPmXt88TATmBFxsFxfqtnjbMSTC4OK95B6cKS2s3g0w0O
1k9H3WzWsMQrGnpZRwZ39zDt/ZuTfaTguegyymtn6CQsPJKf7+PyLeKDgqHD+o/K
pnaVe0C/zXjiuoyyi5AZ1wrmqyinibKDn11dB8JTHl51oKJgXEWT0q+U/wo1HiPQ
01VRdcDWB/gqK61UEtKZFMe4vJ07tOaHzBR/GPvZoAobq6PhdX9tS+baB3c8Wb1Y
zfwT8vag01qCXNRrVvMTwW9giEc9jXtAtBp5a5VbsVELgb3mHlNMA6QoR8g4/gQY
/I32Daofn7aeJ7A1FxN2Z3UOIpLp4JE2HLvinN1VMIYXCQh37lVGqKMMqjuUR772
49F0WDR+xabJbkr7vX0TAjB8iFGC2e2wd/v7agFsjc/ymkKL63nanefHrVZaPY5Q
Z58foEgPxZLCue/PSa1FwAumhDREnbALN9WD7QjrWGrMIMX/XnjnveE3BhjPeQGX
9lI0FFCvtJUS5KZ22E/JyUOIk58JRzLdyoKwk8vjC9ta2sklrDAyUFLQSxYIugZp
TXJv7RB3efbQ1C3/XMHIhYHdnQbWHIM0GO5x2SQSGypkFnmuyvXTVJHyvAxh+jL5
kuqifYx2KC896WtpieW4CM6+et7JO35PJlyzNpWbuUfp8x46EzIFtqjgnRL86OGL
VHH5dA/oZhoChZT83wvVLICqABNMEvlkLOUH+ZifjHsZKy+QKxFamJ5wxnxlFJYL
0sXyQhTM3ndUqrI/ErWNb1k+M2UsR7S1h/e9Z1YGoGgjmkwojGu1sV4SGDae3PTG
lCF3sZfgRIaeFpPLk34vMMCXJyyKBvB07mTUfqlsRgLY438Yb3pG4bj2aMh/UJ+A
nVDOI98cODhulhTRXelsOV7tQr7x3+ZT/6unz9bb8PjiGVs9vmYttBRbfmk3N7CO
ahKvwhYZGKLqlIoUKZZUV02lQqTak9RXnLLMz8v7I7lQk/98cTgRbV2r4VEcMLI7
kQblAVFBxrW68od7vLlsD2tQC/b/JPGIUjR107FOFu7SBoRWNQ63AWS52h9IGB+Q
RtY0o+/DR3pD3Zcz5gyBL9Xb5KyF0k1tKntOkAyt4bvuGgLios1axt3oqA4RR5vG
lJ/gFVXej7Ng0AaGJlOw0dxhAmzyLgy0amqzlGMCz/FJFzl8ltZ3YRt7fDGWin/6
TIisAXNVDhfogB7JwGY8rBOZjd5jB4Z4PDsBiJBWtkxr8etlXXglthqkbQ8LYBy3
ON5ngVCbKRU5m4CUCGEPN3GDeYQXLu0G0BcVsroeS5X98AsiCbZgXkXJhxfaPsyY
XwhS8jVLQu590NA+7CbjcgAsqTCy8WN50PTeNpTz3uWULczgCLsMyCaZb6qgSz56
c1BYbRq1nwqBo8XllvnF/R0DHQvWNrEL4EjCTeDa86a5VTtRmIlSHeOrG3Opl7YB
X1+UAssqV4MrNKZ0ExXCpreLAZIg3Lm6z1Ww+yLpfx5iK/Sb8CB1szycBEnrJ3xr
UcnPzPFG8P7qpeHTznNC1i7ijZcKZVcE4uSpL0HbAr7zo68R7VvnLBF3lqsnSNo/
3OK3boKvGXiS7LuyHVYXg+l2qu9xiNAOiv8cQhU6/7/+nfcdECSdGh4+V3xW99Pb
iI4AUIzuyMYJKMcYPudsiSgljob44ELHiVNSW4aNC1xZ9xcaezE3uK/YV7otLIVM
2mNELLvFgT1dmZMPdVi/yFUHw+k+jbbaQ4GZAMZqpjwWcWCRP4kZpHihmjG01eTb
QpMUhH8UdHKShB/0AjoBuprzYgUC0fgGjW+O/XhxfzClSF8xBZvT94pIfhwOMLIy
breYCvjejXW3qiDXgCuM3VkCdeTHzmdiEAunMhc4YopC7Y1QQd2nlfGMpBmb/Mbz
LM8s7e9krumoQoNBBrnXtmmwc5zpOnTdINiRzclO+AiQ9ESfQA1RNvhmSuV2Ws+q
dQWz/ne7I5JW9vXCw/z3YMPCy2Xnbgayg2+ztJ6GdSWUpdaP4CDV77mo7pYygZkU
50vzg7p5gK41bU17j2c+5zl9IXqot5mUzbWWYiI+wL1P0l8cQKF1mWrObHqYisRK
3H6O/sSF4fPue+078xUhCIJcHMhHk3l1Y+Oz+srScGYtfdLl7u6B67oY9UOftbLT
JXvTzyUPYEPNdgkD0JVIG6mGHiR6SiaGOIbbbvnHvwRxG21NnKYFh7jM848Zog9U
FRsU3CaP30do4sx954SDkQWJDz724pPQ2YxakkuacZNym5xSHOcycPu6QH5ouyoy
EpmKypPVGRKUDO5ntUcCfLv1La9MSY5SlHFIw1ibGf1SWXTJ2URxcQkuH3kJVmex
ewwFHhUFw2p1Eij29SrvhbPk/NvOvCUV5R5CAKMwd+2FLrVKaPgjfVMqgoewi90Q
q6eeKJ9af2JXXpFh1F44XRrsksAqXAiEVlk/6KzOeipmm/srDNEbcDq4f0R8sIja
zLHSuk3xCED17jofRqdnyXhcNj84OXaOszff18N0JObD+aWd7FbrGs4uJKXCsgvt
/vTwJ8ypSJyje2BOW5KX4ofz+gzBcRB5tDtGTFGpg+7A3BAsPLQDHWIsVX4Krfmd
oLpwJTOXYEonS0hheK7BZ+0MeIWaEh2hJE/IYM7TLcBC/nhxKk2RVGjINkGPQf+z
g4dddkBy4lKJIb9FdAMlt0IypaFgPrN1uxOByjgDrrN0ACilQqYL4oMLv/JTuqiy
aJOAb0XdiKLGJVyqVNbpyXDsZvoSEvDGOFioj4FhH/IAooRgOnqmJh4N0dejwQP4
f3/tpjs756w679nA2rLWQC9hOOMqoKia8Byicm7ldxobJYnE3ylH6AYWRR+K784F
1mYbZrRBBJkQhkm0Y59Bwg1usrCIe5yIv4hWppEvwlFy/QXR27bM4CA77HDguqFw
OuqF/Rs6I8udzvcpiK1TlJ+EwVVpWdiKjUWMyLh7nYff6k7iQq3M3qPSyzs0P9mA
dSmwUNSmE68nCmo9cNPijsUDWy9Q4JZu7gNb+Dsb9W9rbKpy9uI+l020pxKoTg1m
1m+BLtGxGan6QsWx9jEUIVTahdovOian3El5+wT+nemn3LL4xbYfosaReQV6Ij3g
lwZWVcgSmsr0H1jz+OGSSTC613TwRED8pfrs65kp5hyXz9Y/LNCFIx4FwNpKSeZY
xugDHfqYUBS857paFZRPaMFECZomWfIGvx5jHYlChcmCsuLwJdnwTH9xocP3M+QW
zo/UtwZ6oe0m+VeZQqyg1I1GXCsPmARZWmIO3yhi0zJINBSm3i+8mJ7ngxS20ZtV
JsCXEe0AE9a5B97aNBJ66Zvi212NgzK0XfTMgkZCLpa2cE9FI9cI71ykdHs3xb4+
TAfSAg1oKKyLkK+i9Qe9+dIfDdZv2pIH8tzNIPxISMbagpOiH5beuuRjzMRbxmtS
AE+rzXLUEBJxQfRile2nzhu53q6+6gVYTFVipMm8ZZNuNxkcN41mlloyViFliAl+
/mTVUlcxIY9DTWvtfY4zbfc0u2nm1rulE3MwKv4b1yYfjtKttAI2MLr5iGzoZJCJ
3VsYqX/7VPYGhtdH7HCZ6mtEjCeO9mRGjjTuc/T3OhmvhZI1lFD3OzLHEgyjRB0t
nHFknNaAHO4bXe27EdnpwLavj7nY98a5ovknfFHAif7XtTlr8WBvk9oVF9XeK8uY
bA9PSdXK09vqCS4S5/ZiG16eEnr22n6Q9nznF++UBMrA1oQ7AYTjuzP/GWfPLQF5
bPxITW0hXTJNW/iuX+P7Pp/LHQbwthd1uOyOYc+xtMknOjsgeDIvnjBYWOv2ST1h
dNP7SqL+BYffVV5xdDiiZHNmolMbw5jp7I4jr7+7V0K84sIAQAWKcQPzKdHd6JWI
u0pyzV8n5TzHcOaF0DN7ro3vTdDGiEzM4UykjaTjSawMzHvMaHHTS6TFx0smmFuG
/VO05HzE3DgNGY9w23R12aZfKQya0PTCoqgT0NbhfkPPZvpIPXp1C0wDXcZDieUp
C0LQktyPlT+ZbT2Ctuu9CPnH9K4sBvzBLe67N8/tLZSY39yzgiWc4EYFndRx+1uQ
ju+/wfe9KO7uhIQW9CWsL47ND8khpvAg6gONNoyUi2iGdJh8s9mKuvg5d7HNUSHY
7I6oN9MqfhjDRQE3PbxsCOG1luls3rFVEqoYQgVAnp9/p3VGAFkVpCQMZ/VI6sgV
C8L9HBLtz1d5/WoXhg1lfSC/OtLInSc7dPPWJ8MxT9hTNW1v7whNsNvGuO/RNbuJ
iM7gUoG4if2IJcU/GJFlydbu40DpZVhxyhRthCEkDC6T0z0r+jTtZBaO4zWyFUbC
WLLv/u3lpiacvWqen4beJH2hcm9fMpl1HgExZDcRsaE6hdIA9ek3gqpY0mckcov2
NjXE/10v3rcLMPyJXKeN6HaVI6f2DHQ5EKtEJmlvRxqzVsAv8uS0pGt3UDM/2urv
pZMdv8L/HmmwGByneVh9U4Gc+APGTKYY5iE9uvCxZfAD/Fzvi/RQfhn28u3mFJop
rPSslMlHMDO/uj/Fh9DpUsaR+6RVbTY3r2xANLafs6lqIK9kdBIT+KetqS9et0D2
aAZivKtMjbl8FT4ipHakN9Y8zPU7w6ClRoThQyj6gd1E6rjeXA7azuP/16/UIkxw
EcHTHkU+xL9Pk5MhcVfLQsA08KIirVsQ7OnA3zQ1SQxsoQ83T7eH1baYiJ0F5adM
SqRUpTaM0er5P+wybOSpKpL6sG6rd4GcuXtr9y4/3e/+0yBbQSH832EoEEFbpzTx
Pfn7dXT2Jl6jiQDamIOnkLLNXGb0IZNRiYfJihAs12PZXH/ombr5vu9So2tJTRU0
O5eHqRUY81qPUWEpdJkAK0a6w640roxduh3FRJjEE0aYNbGEltZnpZuCv58q+6oa
gt6n3akQkNCe18kYG3aSPc/e8tlehZ5YycHDeQEcHYw79uZEG4vas0+CS0w+xgKM
QZLGmnSW3J6BSJ3b+KN+PvundtntWhuO7ZfvyBIV03BXWgcENLXTFcf5A5KdQuIE
LhqVtZgZ71xpQMlZKAgwwTVv9MqZRsrA9HBup19MY8iiVkGj82RGh6MEqgaUzTBK
2pqRLScy6r4oQwyB51BziX+2MV3qbassDe310TBAtqx8EMFULz+t2206GR9QF8Ti
fHRExtl42JB5vt4uSaTca7iuik92uH4bUdLvEGqA1PI8eC7cxMp28XwaNfrrxyGR
VlEvmcwlE5w0Q7nh+96rjXvOdq5ekfcdTi1XfIG/c5qcl1tANFnKUcDiDk4Xym2q
iug47+0dcRRRmfZ+hiA6CXjLwO4CVtPMCfaUMenhGoksorAvzp7KWxh1fHXRrUTj
4xZL9gSz0RwpZzzuzOvQHSv11qZHPQ3yHZMM+Ozt/Urbp6TR9sakYr0axFRL0tdN
Uv9HsgvHdm/fdrmVa0oTQ494V7XNQXeqnLkjJm97mmVG3SIOrwF2v5yyq/BfAzZT
9MHsh2OGxRJ/7M69QBc9o6J0TZsLJExM1mpzCJnRZ3AwArRhuKkSDKLoN9DvBt1I
KytJ6JVtj5no20kh2UcBsytxeAE8WRRSSE6wWIyGnkIYExKd1HJ4zunckbSlMlNF
TZ+N6vyzwjeRsuwINyftQNMzjxkB7SgubFikSjHeqLFghmy0MQoE52fCyMGuXcds
g4vX2OX7xmPaqzLA5/FOVnhKiv3/y9jHaybL6OgqgwAipk2xMcLdOXWBR/B3at9D
cjZdCDCfDbSe3RU2vtgeDcrH6NWI7ZifSCddnv1e9gWJM6KJsOlCoLEP67S57vAt
ZD2l1IdXwO0Ot/IDk8xxfZ1716yF2xlu9Ie9HCnMs//B8tAB77IOGYWLApd15FHV
YeFhnzBSjV9n2th/r70PnPCIOFYufQWA+reuj2XxQPToFuqTSS0PhUqIviiZ2Y2O
0louIzbDFYcUo1acJNj0IBi5eDuCgFgIdgRNAPZWfPfVv7ptrpXgqkWJo29Izh3O
MCzNxeznoeKRcIKY/whNkTPNlAR7gp7vQok6sVV05sOZWebnQv6VaYk5O9G097By
mN9N1tGy5iRBkBcYttwLtlf1EoHGMoUOK9dte5vHxLZIpWPViBaFrQK/epbTQ3uS
gl60Sa7DWcX2QQ2tIJK31iEICM6+ZO6YLHM9usIx/tTIYYUyynf1exTZPt8FCRcI
zgUSqBMiCe4+uV6Pq+L/WiNz02Pp43co8ZA9/zgfhvWps6YauKja+iuxg0FPHl7o
vP84mdXeRtidxorO4jynQglf+4lEGsPrGfXiwdQ41RpXWws+IiN2hGrDyIIPwgw4
5V6n4VGOkwZqwQSFbQp5UrsQ5Uk4aZz24hsh0FNTsMtrNGyyo8jRQJoT214LzMuk
ocjcsbrh1ER8tTtZFlLUgZYo7hhqV2RGgLxcoqrpSKn1yFay669U0d16UmSOknyx
C55PFdASjJAuzah+Dg/30I9WwFo9vLieUXqhqaR937MyfVB2FAkfFPHmtfQyZ0xX
TcitplaxmRNnLTnLErFR+XJsS4FFKf9ZHtIUW8Uff1Bw4GET74PXGBV5CiaBdGE4
b64uY07erMi8Fp9HDpnMaQMqptLdOx+MlBC6bOzGA3HTD+2ZNcEcGmHbHX531F99
3yfLzgU1mYoDpu8ck4/ccRecUYJid3P596P7EGJXn4A9Y9c2ZGPIS2tnbm385X/q
JK03+WgGe4BnLCvUFrOocqQ8StcOCdGj8LiGM9jOwvEgT49FTfcYSRgy8EF9Ouv8
TTsZZgEts4cgufrIRCXTZQutrwhLtSUCrr6MXMXkEJQ2zggvgftt+5O2JlSX2O5G
96XvPLJCOaTGO56AwHU0GtPDh8OrC0/nQaAX0VP4BAcfviaAXQ+C/9AEzZXu60ym
G0xnZlMWI21jonPezYE+oTV809UK8m7l4E8e2B+2TsTj8GlRvwAFxex/y4rsPAiB
lVdNlnRXvjAGk2ar2QpZSNQpi570/3t6d5kpBSxrWFrI8/7esUoUAIyITfSWORYv
AfSM7f9+9YwT+6xZficYt+RnlizKvODAAlBk6/yCi0FNm4opwZ5HOuJ6thOnrPpk
Ph4iPXX6Wgk63j9NW9AEE8bWo1sDH4B4cnfs7H/SNdBaKRDOEHlkVOkltgXkQETn
gR4YGx4DhRQS0Y2tDaUDQ2kaLTExBsEwoJee+qwEOfrhhMi2OPgM+ts1fGgdsTgk
1ai4eqAa5jWlet4c1ju9LLLvtCupE121VCWPjzJ4Qq3xAj4fe6fHcC91zjBjTtdV
w3OGtQGmjUWvR4i7acw4jXBmB7l3/nLmjKTgY9EJvHdaz3V5gsqiF/VSQmtOme/j
WRYaxBeUP83Stfb/EG6di4ND4RzwFRsriaD8suEAgxnK1S+b8zTfP8mJwsBzJHOH
XAPQoluGOiTiuOtQ+tSUPx+vMPonAas5e4apU6KhmwKQp64s2mrpsqfQkAEjHyon
mmCRFw06Hkr6QUTimrW6hhQLYFbv0guby1/i/YnR+uCDFTW+39XoZqpa4dtOc8X7
6rvQNxdqkPs5cFxw+ROEkYDOAkWNGPO7vDlKsH7rMyrl4hPuMOfcgYPJrnzxU619
uKexMbdnSup/o/0nbSNv5iXxk+qones973RWXb+JDIDVvmOpnz5V5oJR1q3VA8m2
hS6SCLzcInJwqYdUkpqJlKipTnvw/3Rt7YkuT/T+2dM4VJcPa/8gFbWGEp+iBKbH
WjybeOGZ/LzSy+GDcoIXblKu+ywbnhu/ZmIchqH7iZE9viInbKN+Z7eZDvBgR0k1
UeK5nCTxeBBbihSviM2YKi5zQLVeaazOrZ2KrQzGFsK6zDw/lt4+x2NR5l9aexA2
r+qZzb63Wd0GTFsdT8z9X05FpSx4hxeySFBdpV/2FxjC/aPopB25L0UqYR/zLwg1
/DKD1Z8Xny3r7ZVVmjHz2edvHuwYv6TYbaja8IA9mSYQKTDzddxH2IORc+DydOEz
WAxYwc0BeEip/OEcfQO0gwjoGvdfkIop/opqTD/zgO33bAvc5zqkSOAYs0yuQQBU
qNl/gjglnxHDTyScnJ50svZdC6RXcyHnNl3ZMbTgCi7g+WlujsqK4v6zJBvtsTrG
31v2+v/i6i3U1hvtdUlslPG7ejOVVgeDyuxOf6G/lG9d1wN5uZfgzWDrm+Eac2Ga
aOxTy+OATL4yBGsBCqnBHwcyyNZ1629dZxBUpO1mJ8C6KSMNQ7O65DtzxcRRZa2m
ixDAvVzTR9Ku3caoaev/no7QhM2VwiSDinuCLdcs0rBmyNAD80LH/aPv6DyZz+7y
+c6sFPNtyjXRiOUArGnMwrfzaotbL1scH7TPNq9jK5WzsZoBGPfeDjfjpSsxw7JC
rgdG3EMMFPXuo/74gT/pJ4R4F6hQs6fKbMX7r8X6j4qpt6Anr9OogyNzRby8RN8W
PxRejVhioFuwB23Bp2VvF0fZhAdvXB/FxPZtgwDL0sr7dLtSXVCSXj1a5l43/59K
Xk8MAr8hhPnnbdEhEy3Bcvc7hNNt91e3reuxcEJmM63yvx4AsKkjRSpMV8a5KopC
ZzxWhcOXrylPNli3fowIiRqcQfRo5V6o+gFfUGofXVWeFftJ7aZe8ZClztyqH5fd
m79KAT5+p6NL1iNhtb5K0EQ/8JU8eue3uSbKdCXY7VJCpqUXOmyuy2DB5QYF1uKc
PcCC3Mefg3S5UBm0TmbX/VcnPE2YXQMT3/kilXcu0pQkxuHfldvzTG/Q24ten8PZ
bGKCzeKoWXO4JuLSzce+SfKHQ57qag1zeSNFcC4yKXaOUa9qPvfvxdqydrbVCnMO
gdP6RqnWfZm4accsM71blPWmsstbIsm4QfhajFxnNLR+m/lWq1DluMa8EcZoPADs
faS/hc2FK8ruVAs43n0lbl+YxGkt7K0tfxYiWJG8G1U3Z6CpIIwrNBWWHywmnMZn
a3Mn3O31jR51B+BTHPxEro/Wgnx7q5Sq0RiEry8wEGKLC9lOzNwsb19bxhu0USgf
bc3b/znXLpipUTXpmDkmNAI0B7T7W2ojN+aZZ3ZLocwBFG1ycLMpjYUm3U/6h4b8
AYFBJxW9Ag3eeioGYlXIq1ez0hlR/eNRGv2TePMMz0uQzL6WDTZCQUNYntCINnpN
xksLFN9dIDwq93TjgHkTegRHbWm25Uz3Dgu0iMpdDYfQhwr7ncCs4TEn63C7IUon
fdSZWbDaac5PNLDPfB7tF+WL18r0d/cgTYjd6gxy1ZbLycbKcDn8nXOZkVyyQAX4
d4WWc0k7US8xe3TJDtqLn/Zqy5OWe3GHC7oDZe5EXJwpO9zxtq3AVueZHOZERpHZ
DbrMqxjhrAgwUYuumrFJZocWGClO5rXDmAZNAfX4KXHuIoUd7WIdUECrhQ2r4Xip
HTq2Q8C25XDjYWmaFFOTOyWGN7Kl/BvF89fCJ917QtJD70J1yS1YOA57zLQMSwj8
PulbDvUKH82+wOc1F7QjuZAwgKXWldTG7j+ZGFBcygxXH3LSlJy+YkdxeyBsPx1K
eaW90RIma/D6hl8OvxIa7Dxyjsq+ERs+NDlcumforM7WIpaIiT2mP3umJvNdIqEs
nKOnQWo/+MYPztA10ueDduOBTQ2PmEVROUz1keOveatJi16JemyeLskP3d4u+PH9
PGz35cJ6kVV17hsPma30y6cYDyCXdOeNxaKvSE5P1MS/VZzrUldIujrqDJULGspx
BAW8dcUfZf2FmAAKeVuQvNn/3IjofRW734Z6sNa9xDllW9l5BBi219FBTh6sYMIx
ao3gaKQ6TwCbe9lJ9lo5K8mHw2mltay2PPjVQoZP/95C2Ut34wewG24LwFt0MnOC
UWZwIOpX6T042kW4XRen26CKPi/brONVkVsGpm2GNWJdWeZmaS3TdLuj9EYZ+fHd
QR8mRmwtANVsrGCqguSf5tOyy/t2i324ASGtyHbbqwTeNkmDjXfI0g7RUReggBYV
oD/KTf9heMgG09Ofa18tQd9SFGC5u4b3ZsfDJT00VSIC3HLI3m/msRgsZKvYNwzy
V0dDQfQV7NtFkWCq/gaAiwKhpk92nCE1qNlsp7ZNL2U2tCkyL3CI/UPD+lyIiwdE
qVGSjg3CdUb9fGXCJER3dn/U6y52Ppynqtjv4IQFpIKKu7/9VsIE3cMTxzCmrXb7
Nq0m4F0ZFp4Vok3ZshHOIq2p8G3nZ33xWvGSR5VD+oJHDbiVLc3QCZiXtAWAsaTM
x42hlXLpLIZQ5HvuhzYxeeq7iJ1Tia92Q060f1GDvYAfsZj7CAhtSsUkIf9jen/f
GDag7Bqhx601myLoNm9VMTrVqCyKWHSBSgdBMVpe3eTz4eZ8+owL7weSbhoY/CJ/
FT/ayaGP0AoeNoZh/BhFv2CN9V1rBpnQ7x483W/cp9XmoXYHuyXfrJ/jw1XHNoGc
+EhpPhGNo1KlkrDoHUzK95ldptP05MoA45ooYRfpD6Ac+Rf8HBgIC65mvczvLx/1
ogGH5abmUOw74gYcf+7+AsVpCcAMTdBs8J0oz01p8H+bhS1SI27ogmnWaMnRi/jb
VjT8svJ7wilI+LP0L4mqLpWJB3LfC2Y+OMnoLt+DTRjspspMUFt781U1HOL1Pgiu
qZGVW63h/cXYH/cUrQpivv7aHc/KLZ6XHwHkmmDiHTJfPjZVZbI51j9Yhilt6wBy
6LwKvVtCHpbU2vLBQ/skwaXV+7MNU4DNN0wJMxGcF3Nms4yLxi50Tb3qd1KzPPk7
MVghfaQxxcwIlyl5fXTKWoHf603I56HI0KnV1ZQomB4N353tbhYkbJRu7m4ZRCRg
jNTRi42kWmysaOQnWsIlv7A2RSIxU7PeGBqYTII7Ph71Dw9rogEM52qNX6LfG+kn
UIBwJ5POPwwBRzN9L6sLx7X8ZJWib8ZQxGTEQ4U0qebc0SIHq7tWV0u1yF2gNmwp
EtGEJNQvBpw8FjyS4nPemyj1jF8cgGbRJkP4PNjH9jOdo+wmwN+TCRj6skI/P038
9dRiayBz91jr0vkc6pPpkwxeih3P0KIX7zCaZLzD2y+KRbm/l0/lO1PX+IecOk9K
iSeDAx3/T11QtkaNbWv7+IKfepPb6hjoXwDuYWFn7xqtOOLAMfXl9FooFVceaDjx
Yrh3HrLkIyHXpBwu3XN7DXFM4sJIr1RAo6CHpXvHFmIRFDUQMHSGfqVb/yUME77l
hWx+d2VeIEoWwNEcrw/wlmz9VasyXAHNu5fcx8ynvmLxiv7KsbYk1BH9YZwemeU0
ShFlyIQoU0HRsH6YKSaLL1TkjvJhOpY43mGsZQesyBeIArCSyW33S8EHdhUizi8O
Kea9G7hgwWPwLV5guWOWLaq9pSSxo+OHQ7SgvyqwBns20PBvaaq+qVzOoNJNE8N/
1NQWiXSHfMq9bdKLVyK2op7tpWfZ+PSa1O61Cnj8poWfw/6ud+/P/dGC/okFktbV
NwcB90C+TAHBFXq6g7HlLNUHtWp00U9DJpo7R2AOE45XbLuyID0kJNs1VBaRv1Jx
YNz3dUgN03oew6U9BA8YtHM3MI1GdOC68gcPGYBpRODh7JN3VxODvMU4KunDckaW
BaXsNP9pXDoUw1L9X8QPKevR1NQb2e2RgIQV0ciL5rm5Da0FOpFjtZ/GRfmiLDCR
qv4w6dy6VY8aC4z0hvbW40KPf3Zc4Dz56EkA4JbB/M9DIzovyRFIja28ZdrHHTC7
YpZxGU+JJs4uJMxuty+U1Zc/Aa327wAhpO+vh4ScDaGz7TyRLj5dfcwLyWW02TjY
ZgBjS4rjDWIJA6y5JDhbed0X0TZP+32hT9mq/ubPEFBiESmTi7yz0tVy5o81JvE/
u5EMoG+fQ8X02i/re3+QlF9edz2Dcnh+mqYdQ3MK7py9aj+mj2mIkyNwPAWad0vE
b+FmNCl6QMIGnCLKNniJnLwPnzimgw3GYjiu178PLvdGmQMRoCad9U5W+6m1vRC1
T9KUlWGXOiLlCdyxLJskLkbc9oHLPTu/82IfRQYtJEbAeIPxbJgieyPIti6qv+xw
9yCji6TSiFgHSvTPnCXizyoO5aFeXKwkxpUNaqEhKhBFqqe7yKYBjp3mjosu3poS
x/u+UGY6Jvz0cIUCSy7lH6shQVjk+DpUwTP8vGSKRwVcOGe+VRHYoTPQNa1IMKfW
RnePoFMVK8xExTiUihDfFocbGFd3lctQXrLvhZMJoydPKrCufeNgALJLVxd+vIcp
kgZQt6gst92FmRsK0hrng8TES8WR+2kLrGrGRLMp9pxhvGBwL3Zbg9tTi6kcJ/1R
ulEIjHYsrjPvAdxeLCH/unufGLlnEe7O/zlOtXBBnSv18c2iBBd9PTyceAycEsRI
88AwpfNOONHHjTamP7hVO7N6pOjZq/b4BLGWR0MI6JKkcfFKcmQNrZ9eWjF1qqRN
zpX0vOAboXYfjKoXYB2m88PeKR+BMdxbNg6Gs8jBCcLRNWBYKdV0NNbamiO6tXrE
SWCecIY28odFw1lqRxZ7YJuqSZeuSALokdyC84JHap4JgRkkozgGcl75zu10B7Ro
h1EO0xg4VNoRwZuSfixw3SizgdYeLxKvociRuqFHNLYyGmd2dXunf9BpDcucePrZ
n4G3xsmmMFhy1j9jwLqynS3j+a/6EFlyv/71DLogLe8hantCCZeCqXqEuTameXMc
1njiXFQiP++cuGCLaZYyRq1DQIDHEaZQrv9F130yKpS0YwlcYI6+zXKTXw0+9N6s
+hxdYghYqOjdSZXgoTGssENFhOAE4PU4kQx4892aK7TSNDWRZtQ7DuzWp2fLeqzL
aV9b3yOzWa2Sjs3pq+0WAvNckCMk1xe4UqIFhO7SZdJCR7HACx0pIjo6zWEIjT+t
iU6xftJxvQElCuPjRXcehog0FG1HsASzfrizdIF5a++BBe+meD48z7IiSaQuWuno
HR6+61zLV5CnKK4y1MgDUHQeI4/IQsHcCB1G5LmuAplqbfzCl+edgWgmlJp8mZXH
kD48AR1yPZ5MKeEePf/D7HucjXd9A+pIoblxIzA0oc8T4chKkNdM7F/bp8ZzJ9Wf
7RCyAdwUOcz1+C9zyzXY2qMc3OKnQ7fxp4mqWe1265qapOzKQndxvnY/VrPo5+HG
wawm7xAyaOnHemz+3NwN4c8Uk8WY9NHM/MX3xh83nIkJze6QgUAWBZfmtSe5lg1L
YcjJyqt3tV4fNeIWnzb76Kzu9EVzyfKmBePrSJziqGostWnkWLP9ZPFoa1wCp8Gd
1muD7cAns0sBpzFljPMUP5+A6ibm0PTD8XnMkym4WrZrwbTBOKJggX82D1u1ETm8
vg3y2oImNhBgfquMEuzqydEbYoUGOJVV1KGLPmOF8byx6XT8SNJPlzY2S/+FPniM
NOEiuFIU2fpdgmQDm8h9GWTMnq3PfgIfN1cGbeSWPj8RoJ20HsjfomnYl13PIIvu
TkObGMJnMgUdPljHTEqFOutVNT0xosu+aqsf8uKcgL0sI7j/8tucooqgUir+Fy9g
OkvOTkE3OAHvxzkjz4tvrMRuXITKsDZQbi80YCFDJSXgVaFM7xFYXxryCCkZWKeh
tDxyDxkuLU1nNiYi50xY5Zd1A+3wbnTz4cOM6YN42XYWaMAvf+AGP75a+yJcz3fd
nn11jCesFKW5XotOVwlk9ZuCvVot4/50lib38JfR1WBggvI5pCh2/QzGp3ggbYwb
UvLiq7IaJ0pKCdoea42EEiSyDFNC1NkXS/54B7CcXDzSQ2YHxr2B6cVcza8AuBqb
TuB1Ps4cttckpKxSsSjGNHC2my8qF7pPb4IAUtWyh5fjLRue/WJGmZSpTkQlj9tt
9J0QpNy6kB2HAV/YHvUdO87IE5iLFQ4Qaf+ASH+IGNLCLSoYpKE6KeCe6m24Qro3
yIQ8s8Rp8ta8AyYbXTaTbDuyuehcvvlHBFUlf+CRCSy8B3wt5bENVm4ClsT2Nyhh
uWolhwBFs2wuZYl9q1lWznufx9ghDsBjPI0eMPpU3Txrq+UMx4uZji7qR6uExllZ
xtyURpMRgA6Wd3CjQrJmrrTKUTEqTFuPFxfgvL6km8vRDXhoSEdPteWf28dSjDPi
Ps3+25PzJ5FaCYxvnUSYZqxMv/w4Hsp9OpzvyI03ymLiOmGb4Voi+gA6ZZAQe8Q+
A7rB3Fvl3R+mvbdPOYKkrGqCaRcNd7ONE9xT6cad3khI9qBjvCHZavlsJiPtWG5z
Z5Kn9RLYdzf3uXzd0/OxY9IflfcTsa3eAq6T17zTPi8hc0iPZsnp6CQ7QTi9iFtk
iOADY8pIfcoGKdQSKpqurmrxeWfM3GtZbGC3BumDYPyUKbMQZLhQJyyZCsFr3KHb
fTxnAduBjJKzjpZpEE7AjKa36+XelZud5xoWOQIcc2IS/oRnQKyGq3RuGjJ4GMyA
nBkfmoCyB+KR7tVAXApEU/SzkFX7XK0IQhkSHiB8VtWz8jfSR1eq9x7qvgRnoqpg
4DwhMujnAW1OlrimaczVJHQFGgoBAJHY0lV1Lbaf7TQ4X+Lk6+gOBUX4L3vcczVj
jQCbwLzDTrObJ99mJgzuPeubElQAaoxRO0+LAoxGgY2ycEOLRQKGuu1uU/TP78Xc
+Q4gT629g702Rq1qAQfPZjINyWKCIe+QqQqTzVB3Q8hs5MNM5Y10tl5ZWdpd+sQK
JlUF6KPUIgigHjWfoIANsF7OfLsa3uI4glT9qtQopsENon05p5cfzKrUWzLUIwqo
LOtkwKF/zBVU12Rjl53sg017OhyOtPF6x0tQgg44brjKBhxEi9Ug/vUBPBmANk9u
b1Efa4UqNhuU9rqQH/Xu+LdQlYKQ3PCYBsAbo3sTGkUUdBoH/15KtT5aNY1VG+dN
a5QTpcj5Nq5UtZsLIMf4VrIGbLLgiZVvqk0xOW4dhRBcSCwV6RA4CylYcnupqjP7
Mm6T32Vdt7+sPZ9/1oTKeTX8vXnGKEGmcI+Z54hbXL3HK3YhjrMmpk9aazb/C9kA
xdQpwkl/fD2u8pMUSpZFPxM98BrwnbGctV5d2XLNL7rtNd4/bAm6zuaJ/DBfEwiM
b8QCLpH7sJ+qFH3qjf/tyTTqaCl85/vncr0WOx0ENA66sk87B4IISxNmdPPinq6S
nWafjoxQemptFKyqtkfJB7xulG84AF1E55azHrZEZlotNNH0YHBHbMCtSGZLLjyj
nZsDVNEw1WdcvUhgPhRIWMHdUpJYwst9JFP5wvViLXwrR0AYOFcFWRFrtnr5Gm8R
bcAyOR2GdaXcKFydkYGLxhcK4kVZTTmh6iKDGDzcglm6cI2WfjJh2tlI97ihjmPV
2tAVSvJkGFbTkW8Ajfagd7zljtKNjFA8GX/IDyFm4KgW8G8Cc6UPBWhz08ayAwuT
XcoaiTKA/EdYzL+1rVhw9uEJ45R3VOlzeGDnzd7JDN8zCEBFzELBlHUdt99tCQgD
wgk0NQ7ly+9k37sfICfvqBoGHPNusbYfkC2qlg2BeSzipJK6Cr8J0EePscFcGaTt
lzbXmR/TfmLzV3gIzqlT8dLaVf4afJF1uGzLsZhwVHjzNu3kQPVY0OWkgqFh2noP
zbpiISGS5Vn1yCVCyuDBe0tzt1S04ahUGVR0iYocjbetMH0iYR8DrvXjq48V68ch
5H0EX5GSdQiEgJ8QJJW5A2aTAQsKpRvyWOqISNuzUshrBBPIQoaZmENI0FLvD92j
b/Y7TKA5NXPh56JTrprxzOCNSpCKG60CzcNZaam34peNfCAJWqyEJyKxHRU8uUzd
9S6FXG4bwEytW1M8vA9YxRYG32fy6HYyPc4i7KqW7cN+DG/yh3X2SPnIa41QaN0e
rGv3DgA5UK5aXTcsHI/is0XtSmR0nj3dSOu7524xXHj1zydLentu2bis0ZDXui8b
g7pd/IMigK5Z3/BHh3k/s+Ymqrx/9XvhI2QcfXi9TfFanyRQ31Zof/Qe49097IhP
o21EirfscB2ZiOc6DRXTpLM5Lt8nebfjcfb1+2fT6s1zdPQqhYBF8U/6+DseB5Qm
XUqi/VW0qvQcK62ks3NKyqo/mJs0ic/pOA+wrHTTymjJKanxZzHuGy5KVffghrJ6
eT4Uz2fhYJIdR8cupoarMv9u4CREH90ycyQUHmGT2vSMRzV5FaNYU288LurKwZEt
70xWkgmaC19XUK+Q13x9ZNwxsiSkVp/ZxC1km5HNvYgukBqsZ4X9U4GSSJt1NqYr
MZh+irV30ur0zIcuYCjPTZ5Ug3MITooQmkjWQr1Q/+D/2MJfN9yDnQUZ8ddSz01T
4BsuyvrF5H0NGqUU0DSQxwEX9k2QQiEZPUwa7vfZ8eMQbFkFgWCw/6YdfD6nH8Bb
4LqHciaOfFoqlsBAUHYpej9Zl+tmYduSdWaBx/oCKKCS6SFf5LkysjMOH1UuSl5J
lVtQvzpEQggzuJ2D8/vlE/HsHgqK5DRclYVkMrwQHiFMHdxZCkwylacreeKWOezV
0J3aWXXXYqQER07A++ufSmMls2Y4YjRmdwTidXA/xVSfIF0/eseGdzvBUg/NxQOe
ORUU9WkYbVSMHekxUxpJY+8sq89OspoqLARqPVPTq857H7pnTPyBICBTc7S8DtNZ
32mceMNr3fM1TGhAN5GCE9iQDdZUZ2N8E1+hmcEZAs7U8qosSu3KiiqK3Av+5qk3
k/1ctmkDMY16SMahBXXyOi8oJyTrLBcpdkBofRSRKh3aKaEHhn3iOds+Z7dkTQVF
Ejn6ZwWh/+XbHN7q37JGwt72x6L9/nHiwgHhpP5cebcUPFlEtysPBgHlNfW5GwUM
USAQVrUxtNUZOQsx/UUlJnJF7/Q/gJI1rV/+uhXmEgOcldbBZKv7rD3BK+lULy0w
6tVephEulCpQ9BL5vi6LcUNkjFlaQalaDI+MvurDbi/5rTikO/TePeaCdnfNen1q
66aqgG6MXg/TSvAy+B48Zj+XXUblr2T9TGY2WFHO2zfYFj5lJ67R0RgNRvrmopvC
TCVSgiuabiF/JWLBUGMhjfI2pFctkUxR+gFJelmrEQpGp3v4AdblJs0ir01AHArp
C4B+HrDyKZg957hvMJOQRB2ayziUJUR6sMFKJhwIyDYREhs0GdJMtZ5s8R3l+Tr/
TW/25fJqyW2NLw5rmzeho8eseZ0/wACJ9znY2ihZEP7+pWz+yaboP9w2V10NNxv4
tt/VCS8DSxYw2Yc7V/JpGVfDnzHb9hfEDjZ0Vgp7z0ukh8u8QzyCC7QkOdLaA736
Wec3aUdzIJv+9bADqSSbWD9z6jIEj6rOHehFexkXXT8UDe2f8dPJKvruOfh5Fxwo
VeHt0xLEkRYF/c5/Kl1r3rbz4+Ibgvv4CkwGKSgjpNwXT7FT136xqBbF8HQuAtEC
SYeXHknrIyjjWljYGwLMLsKoh9oiuHhh4FYXuhckn+tht1zZ3Yax02K8Q48F0drZ
d0sEGKKCSJ69AbcIYI+cBFxbq1qOPhT2K26X0rf8VZ7uJ56NUTIbZCD4yNhZK1/7
hpJ06qvBOwW+gC+cUX4XUNecuGI9nWFGj4M+yrmVQ5eYq/FigLosdvNc3PR3/t/7
hG36mHaltZ8eqzi62ZONK3xde3aebSUHTpTMIlrmIt+tVGQ6PO1BPUDKBT6LaGG2
qGnQ54VKlME/32lZVdl09Aj9ckRg2o7x+HUKrjIDPv9IxpSjM7Hatmpf9gCZAFiF
c7UgRKaAazGW5Zdr0Vm9G+BNKBK1snP1JaN6VlhrvXv9dri3PPGqiJTQxS9Am/p4
FHxwRTpv3JVK1e59N4cW/N4NjVJFYRKC+MF5U7VjHXzGG3ni/Z9kTJAheR2Jt+0P
yvngVIGqEFQ8TlhXxyhQnzyKsOjcVAYNoxxFGNvvfux3n0pUDqcLe5vKbkmG0Km4
+HSQp+2Gk/khF2b7zZ4QCN6EYwkohXj7zMUnCPZjRW11uoW6AQwAli+7asLdAYhR
+EEmh0HOqWAh6nl9F53Hl2g3aW6Xw6iLBZEcrmkIIBdbYxDqcbxaBeBuzFvpDyhf
dhFgGcAE0btsE1q22YMteKiEVACJrcjqKxwQ5vc6/h67smRC3ZnIjGuciN6VI2uL
xottl5Lm75EnOa5q1vRP7bm/hYDbyFMcAey2XP5tUO5w8+S8jznTNjrtX4q1gHx7
gsgvA6QB5GLjsc++gh1OiJiY4Z/BmrYSXXUSTtWySMsp5TthdAv/Xsbc7pPLa1Pn
4nvc5oDU4zyxkkxkNpcQfeG6/wT5S5FSSAbF5yHuSAHG50VMjRWpY2wvyvouii0Q
e7cmFw/4ynO5t5VxpO7gpvJZuqH2gIatuVlLJQpZ33oJrRIYclFQEgWSn/L/eP8F
FOUoH4aYu+4ZO4f5f/UltVhQsAjKhpypjX1i/ybMXPMYTMLsAZl1jvLn51JA55ea
DE3NYxe2CBTX6mFR91MJcjxK8TB+elSGo6QX8jUtm7uMYjZcVy0WoxyXO7amVN22
gN2ea6NC91LZt2BXpj7bc7jXfmPZxEUv4GE5GTsz5rm2mNv2KYC8qXZK+DNZxAqp
Hk9/dkkon8+MMPr0CtmFEFiK0S2R0NfxjNE0q96TQlCDxOeH0aL48v/0nPXx63Hp
HBEnvZSZ1+grwmmvSdKIRFGaWfWiqLZRuqoeVDGVt3KxAPGAq4MTX19Xtfx6JFTR
oeTJbsYmenM939B0ZOL4yN3YObgbfsBWb9X+Il54UPKyASgQkmgrKD1Ia5lJyu4A
p6HI/ZLYmQBGHijyd4qtmLMc+V9/7jXZ/9KnCtMQHIfXn0JT8a6Fkq+91BiqOGd1
GLxgZLTgwI1r6ceFKfchoYQzvxEbuNHynIO3tKQwKi9TA+QVR6UCmKXTC47MwCM6
d+Y/3Hj0PsY+usCU28zkC4cUKC8Z3YkfnD9TOT8GyYQYp27MXN/vXzldCYuPW87A
sL6J0xXzCqI5cCJC52eiSq4/hQEvCAkewZebyPVd3O2RSnjtHSJ9LVGHIzlErTa6
VWj8vAJ3JBNza1sPBJYiGaDw3RLLsvNestKE+X8ZL7lstexn39v7NM0nuulMzOwj
HNGc5jbTNMC9oo5dqxOhg6UTm8/Vn7BIP+tcmKBtETRx6pA+BcZR5nUMHYpiweEP
bnmG4pfBU1oXcQqzhteaOHnSwSqiHAodufivtWZVisAyxRuyisqLsSTC+JL398Yw
GVzZdwSd+1KjeVAoOb9fIS3lvlHhLBKnnjomW0+FDt548cdeZC2Qhms3uDtBv90Y
Ev4nypwztM/BbgoWHCSIsVmqG2rXGOivfaCzEuRxUvaqOJVVuqDeqS5Ci2V725rf
aIa0fnFYoeg79DucMm20F8KxuSw2DvMeJztWUoAqtIgcWXAaC0KjjCwXT2NmIk2p
oIQ4kMAQgkXuOvAdev7dIdBlNQTBeZ5BK9tH/vGbk+djpNfz6fKBbcduDz+8V/u0
bzun+i5CStDiyHooLhsOnyTV5yQTQSFbhgLFC9eAwf64tkGftdUeJ/P4z99d2IeP
T6AIm+eZ59oJp/KWvlsjDk6S231Kqzazt/LkeLvSRBye5LvoQzItP0mQspqlePAU
sfW9z7TH5e65QFRrIK+I/NfQviVFEeMrpsQrQeu5YsxHvD1AZQGyC1tdiAF//XnI
7oWNaX7UWJ6wAWv42TACkkBWb0waUGulVRCUG3OQJW5SuwzL9eLt6yg3bt4B43qp
2QY8K62krgLXSchSD4B/IUXGjrufuhnRzYSrSmKVXQhCRr2ypABL3fpBmGVPJ2Sr
4LyhXCwZNn6LnKyEnyvDtimWybCy5OQDiDPUOjDKC44d0Ckdyt2Fvzjl74UjGTZp
2n0jkPTW2EsEvNN8plJ1AEJ0pv7X0pdyjRN67m4yMNXVSzmRjHIs9f3BHlNfqvqq
LUtkzo0Kr0QoKfhphPRhOF8sECQNgzy/Lci3eAcvWAMdYsH8SHts0weAlBDsaQeF
JTMK7ojCd4Il2E4YAZI/DL0h8tSNfxoMXNjaeVvFfOtXAH4wSw3aEymHsWlMewuY
Ty6MwovGdHXrRhMwNQy1Dv29GcEUt+sGvLPnDOVHdb+vS3MneF3796RWBLui+mDC
X6wQTqMzyEL+Vva+tPncMMEyhtjlP8uOAI6zKCejfNFpR0E+6o88J4vMkknygDUr
81fmH1x7Rot8KDN5lhOPhBmu1300eOvTAKltR7LFETk7kC9f+eHxRIniRktCb+08
AnnoiAYfvXKoEtk0Eg1kMBNzPHh/fe9MeSreJUkbN9j6kVDHIwMFuLz7yVwToyV8
9iWkYlSnbkhW0bz6C+aY1KMf5U15WVS32GcNpLbIbwGORQOfjUAd2ijZfRIJTff7
9QLHhaFo/GTDtt56DFYgTT0/gOLwDl0xnNASSePYOVrHdp4SeV5/ppm2XZhXNlN6
njTDde901vd/8fZ6Hp0FH1VDWwXE6A29OeGYHhwaVz5MwlXmNlRQBRCJe16BgTuP
xuGunwMcx0KiPX4xj1aOJli3o7IlDyma1xQnSiDL8bmTlqJkH2JK7YyHIMLPloq3
pG9Vwh/ZLv+RuYquePCYWeBwFburYdWNjQ0vjPXPsNIeit0ae3Z0gUR+5Dt2AzfN
fSfurJgIESrfEB757nwDte2oj5Hy0Na/qRXaMV8Nv6eKv5JFXqM4FnZTCqQRpvGa
SRk9YJaFCoAUc8Ef7ruxililCOvlAXMA4UyU8MlHPLbdCdNA3q/LwXRZ31VOBN/t
zirICU0l7EXctfMQzqCxT1OPblfA4esxjKymaneflMUFKEYyOJYNRqpmDct7L1MS
haS8J/IqUAZew7aPPMTtCx0QPnKWivRvOjvRRiMjvywcyIQTasde9GqkFbicXF7s
iEFKmvVOGywVFQa6oL8HpIhOxtLSXbWHFom1ALS2HH4Jye9JYnaQxHc/r6MJMldy
VsO8etqN2vSDsSEHQtGFDk0bFOm5USLrcFFIMj18XddWiJRZIRR+1fRm9ZHHHrh+
z5BRO0OU6DXmcskC3byU9F3PqtgB4cq8/40dIbKmjfwlcejLNdWCo8saz3UD0wrb
lmHJ3jIkhrXYwJ8mLUKtgd50WTq4yoPYwjnj+OlcwAHxGWkAlRL1ZMJxpzYvm1xR
FuQq5RCj2OCLVG1+DGtUOc0XElwXMaNULhS+S8ZYvfb8UUJcDQXnevShFRa7LgV+
Xb/FTkTFXfm3w9twp4jGdjYZiJnFLcULiGwb+CmVAanHJPUN7jrdh/+cjXFAMW/G
KWEQ2pBFeiLYvzhrWv2nnJ/Hn+u1wtQ4aZ8W5V20/RK0tbcdOOaUp87sLeyyouYT
3ZcUUMSy3svlnFlxcf81F4JPWGM0B0KuYtADrDlS/S1yEQb0f11RSadJgP8X/ro/
OgFDjVYPGRx2vZITZ+0p7W5aINS0SqZVmfAv9I8Znr5r/HGXVsspEIuinGbVcJD4
2uxtBxBSSDnGweVNWHzoNzyyXt54hguLePoTTE+vqLjtZZXPByFOvTlVHpflL/tr
hVgKxgtDQqu7OFiL/nZHbclXhPy+cdUXY8aJ8fipFt9rDrZbuucTeKJYC1SHgEvF
r/yDTAlU11NopV4NN+WK54h6y02JBYvlhr1rrbwovvMinzz3j5peCdn75ozlEcSC
d1K32HOuvQOW9E7WO01zhCHTdgsS8QDelYnTA5KNwUw20Mvnob0GtzHLgvax26pT
FUQPnwLuUdM6xsE1xoRCkeWC9Z6YXnz3J85SF3VzX0Jddliu4MqRt38998+jOcz6
CJQ42DVfZQ+r1Xl639Q3++SeiU/8GB+dTEufhA3dL2Kt5VD6pmMmnksWQUoQ+U+g
drT70GiZaZKrmS/v9rtVzOvnqmsvErl2XuqyQThSXO4aULf6yvJqej6UsL64yAGd
rcck3yPeYKyTka9ptm0J05OV2+QoSIpcbr5CMOMoXy6yh7CPCObYKA+Qthb9VTsc
ywo9aGbunfi7TaYOchNju9Lnq43uGwOMF9WcMgYqqkZO+/5MCVMtIkPI5kdAGKaX
yaOHpOx59FVekbnKyuKskIgvFDatjZ6YY3eu9cDdXUzR5N6BJQA2k3laEHagzT9e
gUdkQUbSiUiFvGZvIawVFALv5/OMEWgMpW1Y/IiXF5hW0kjfw9j5LgCqcCM8HBc3
+LuHeMneYcxpGEqfiUDX2LCQRhT3pCNicyGiZZ/8WSIR+fFNP11FQWYQIFAkt53p
bOfF4fN2CQodKgDsMpKRyQk1z+pclgJaJG39Emq76D+XizsDnESkfQcU+x3dA1qA
kLsFve1uwB1y+Kobati2P1V172LYIhJ/7yRAb7vV5/oA0R5ZvFkIFthDNOLI3VBf
87OGQw7Pxql4a9MeO9e5iA==
`protect end_protected