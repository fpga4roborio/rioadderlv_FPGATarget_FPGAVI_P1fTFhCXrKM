`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
ddtXksX2+yylW5zu6QL2Lhnb2d1sD00763mmSITNX595NcHTEkwn0zB1Dry37fOW
FufOhVzEJp80NC5qZ/+F0Vk7Ik02dIR0elf3clrjeJRK85K4e3Hoo4xn7YbFUIms
l/8VZSb14+JVGURjfswrIyCUotIzlzVYZ6gzoZwDXIi5gQIBf/gI+KxNXPaKV+PQ
Ufys/12rjO6aI/pPlqSm0hCvftmBcnezN2hk1UeXgOIuKZnogjOsf0iJVX2aOOWE
6pD/psybjbnsNB6kH5uFTA5frkzIzkzl5d9+YDm9OyC+k84E83I/7/j+rk4L2dah
QJOvksSIzN867/4Qt8qYTQ==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="MvBXkzurAa5VTw+1JJ70nePUfoQXBvZOku/SMmg4TwQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
oRtzZL4VJ4iwysPsC8SXYCzXS8Fw2gtZTOskLcDV+1B9Nzn1zTyNtlo6lNICRmmK
ZRVu2BmCc2G+fmzynYlNTnSa7C0Cuel6FYpxCBlOuk3OF2tzAmLAuDyOH3Z1Yjzk
a0aHuoCdIRKv7BrZCdALt03JeUmXKPdOmIlkVGFl8yw=
`protect rights_digest_method = "sha256"
`protect end_toolblock="Jn9CQpRhJt4rnzZPRk+dOpzAubz7omckX1MrFd4p81o="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 14976 )
`protect data_block
gD6l00tciPUa6pDNTk/+t0OO0nC/UTtBwLB41d4inuAUA3i/ALrNyoJVcBnAmEQW
ptbcNp5fxEUJjnOxnedyZEuEBxWRieZFQnkRdF269oPASLtWezOm1bQB/9nP14Sd
UDPOFBozsxi9Tc0ULeCFLNJFIGPxNKJO+ELzBF+94ByZHmbx9tGVo1WTkEssSJQG
GRmF5h7weW7JggCiAcz0lw2nIna1mBkq+wD3486io0byq06B7HW/LWdx44QDBYmt
OOBx3Gc8IAft7ZoidF/vQUnZRv1gIFevyZVXQuR8t3ZeJ+xMyoOyXNVsscrpj1PW
uRd1qymMr9Mm8BcR1adNxpDBQYWi6DJ9xx4OTkPZaPQ7Swe5RIu0AD7bwm6AUmvn
mGaPUfGJw4YBiFiLoNWm0iTOjgliKcKxJsZTuVAsufcCei/Vb6l/tNpTZRAL4Hbq
E8hA7kBFGDFk17IcGZqxPkHU5Ha/sbjqpi0mf19lKOcoa/wzCR5uOe26+Tl0xOlZ
H/isClInTc54hrtE8s07SUYU1D8k2lrlgFyuaDYAoIpyq1bhEgk/a1rhC/Ehp69p
4nNmX3UWXavR9bgZv1PhGF/Higs893Y8yQKEhIsTf9hZfabSaEGvJ87Fl+3QpL3K
uU3dfn9TqFDk1JP4QV3gfAt6pglK2xcbe5+3/LXyzHIYNn4BQN0N9ZI7+QeMuwsq
8/3gfYRyWUI/qLiAGRJ3Flqkrr4YPEQViUiXmoR5ZNXTPYcEOly/W1QdCoFHUBTh
XLRT182BKqZM+QVB6O2CAIW9zB4VKp9mkkionftGUMPsYoo07hdoHffLqeajlm3N
mnA5N28OOqWD1eq4g6PVhsbY6FzZVXFUFid3ZOq3YNXW01hyOTfXa7QHX/ue7SuF
v10ZzYzgDgO879g2v9hu9HI0VCHnj/SQ4TrFXGXZ9CVkeXgARoaKb4kBQN/FtwDJ
4TRSEaUGEeEUtqoPo1DMsFmtbxDGMzr+Nf9qsaebue38xA3WbvVdHQCB9fEebgf5
4OfdMQVzw3qmEVidyCFJN1Q1+k7CoZhMHdX6PsI3jwJJEeiGIVi+pqBZ6c5hjQY1
GbZUA34mpBNa2wA6+NLDdIQx8s2Mxc9DRWQA6Mx8FUSVoUH+oEsFGhp3zcPAA4B7
4pznXF84Mg0a/+nP4rkE+Yt7/mR1U1FomkC+3lJj5pOSVEYoNeJTlcub81JpctmC
fZ4GiqLeOt9/gG61ISz2pyIFhrwQN/qtTVYK1gcN1To+l5PmIjeHKI6B/xzx0a2i
/sywhthAfpGf5a8T8gmBjjiltyRMGaxDboLWyxmYQ8yoVu+T0eMjmS6FioeD8ZmZ
ydGcLMaF5m+E70lEAYkpo/cmIpA5w+XaW23DdECezAunW11jUYLE9Ao0Irz9tNVh
mwrn5tpofxe7Dv51dG++JQuCZh+JPZc5x8ldBFQ49R+kxGkjLAtcOKvKhOShZAL+
vZXaRz23No8Dhk9RZTyv083XpzOSSlr2X0Wg4P1DGn5wKVzTEUhrioujKgR1kJTz
7qdwLkWqwqign+pr0ApYVsHJK7soEYozGWsH/JfGgeMwP9c5Coa6bsYf/ggS63p1
wl6wMBPGxtLN4qeQqQR76cHIy7zUWl44iMGyiCjW0cNwBg9Gv+SlhaigerTAr8jv
xam376Dh0+mxkVu1zw0f0Eqp9yFe12YKYQ36whmVwFibaUMdasp6nTNtVST/d/YW
mPbzFKUfLrCHIkC1JvuGi9ncUpN5glAfjfaVM+Fl9Z+YMLkbHfWKApu7fEShGFkx
fxC89OaAHdNYOKNAPeaTIWHalWlj8EtHA0iQzHtSHPorV2bQB5xtBuYUTGLkOHSN
pFlMUNkc+HEhoCaOAbdPGnBJyApMkmShz34TI0OEtektaoKzCZMz5siXU1+MXefl
Z1KBcPCWB/n4xU3+sgwPmKmB8sU8spcG+C/iQdnIvbDfPe7ULiOOulbKKRrqDnvL
52j/Nd6dahRDljsmNVnqy2uW5NOCVX4YX6iJWKFHQeK3wbnMfrE9kUKc/8T/3Fks
Czp9EapxyhUFBfaKhcPiKr9X+360o0cHTlOwMbUzdtJX4UAen15GQNb/vJrpbTwF
mse3QN337mF7ADm5GSGrMP+g7dX2mtSQnlT5tdNUmKkyV2dNgZEtH7as1xJOhcFk
ijpEpGvdIq4lf/Hu05qHrofb+DAtcOg8YMPZmqJhIdPqH0s17s+Tn9GP/CDhx1XK
sPTf1zdi4iIeQ/65LGrfHacpxiOCA4XmC6fGVVIkVkH3D9bCt41WZDfVMiW61q7Y
NtXl8vRHGBStpT2TUR6+2nUvG6eDTIuPtpZaeQGRZqSh9IgaEhmngiJa6vozhaNW
1HE6GJ9de61GcZmoRu7E4Ci5pMPqHCafclKVHKpWjk/FHC9mkljFaLaz51K9vDk0
J65eyOQ2PXXnJG5dBdXwRrePVi5yyhlg1vZoRb9pDp42WXDeij9MJX1iit0B3tGY
eJBvLeeKKWCpNOqe+o6F9ZnYK+B09xabE4bB2QGg/XWBZsVcwWtItnkL7MIVKz53
iSE5kQqziIylVkcTiHaTw7UBBYc5AMPYVYGPBz5S1dgXBvMl38monduiuPYYKsBi
9sq2ZFYxwi/xbityRul02zb18ZfwfbZYbXrk14hIMLLnOoVBtEQiD5xhnwS8ijhX
TFBXM5+Xe70q5MPVw/m3m4v89Vq5/YGgusXEjxxr9ohynoygerZxOxr/Lip2Nl4t
Fxy4/6St0m1z7LNywiHzkB8Lz7sYJoNmeQJqnslhZadsRwOIANduNV59L6wUujXm
MHf7GpXEOrIMoAg94JnVGk+M8Ju2tafN6WWX5F/kLcvEJjFSXcYDFoYniD0Oo9tt
niedzdn2cZhOo0hhfxvQedh3cavQUZom6ZCUJvarVeo5Qr5wgvphW+oKtVqaSMK7
GjjSCnAhYfg+Gvje9AjA9z0gcciiQL7UH6PNMQRxTimRnQSwwMYcOiO5lJlOY9hM
rH9nZdtOSFzeHF4amPcgDdoASWzdBzFNIcYly5qsXghNHPtNSQBumfd17k6G4yMn
jhQGMoASFsWefW8UdfXsX72BP/nCF46XVTncjvE9nfZ0KFCi585dXTdBmD2tCpr3
qFwzmwqrl9oV4e+/Ychj5eU6qDPtONaiiK4wk60ZljbcBgBda38AP4hqGeyI//gk
S0KyEQR/OpAujn3LnJ/lV+yQbrgkZ66MTWPVAGrfaRD0Q8rZiq7VjD9xXfd93hnu
xvGXiXB9Xnjt/gTk+CV74d9NtFd8IjtdcIjBaOD1XOKV9r8Jkfy1vRcJ5q4yGEcF
s1J8yAYrZKTjaeKEMhzPBU6Zgw41GzspvwyPMvrZ59WqrTOg+Wgd9fV3hbF/foR4
iBZndbK85tErcEGXXB5GNWeMsYWefXG+gU1zrN9JBDjMpfE3WQSiNDoIClCm7w6m
UET/wlX8AeZiTmcReJ8u3dkbmyTXB8ZqdSXtroXdWQsnBJuPczMdPE0me7U9YGzi
l8vBoZGYlTFrUXkI+qc2ZejDjByoGcLzuk2aPEuvjqqaBbgqx/r/MbGlRZKxZ9FT
ALr3aFTgkEQ9V9hAEmjwQNA+Hzbc45WiZ+xkdtCkh84MfXoDgWzBjtCs9xOhaiSH
eazCA5BT7dW200+8QvwyDksG4K9tXivb/NtY/foj+tNRkNEIbkIQq4KOF21mYf0c
36b+e1Ig3SWFu3RLQhjf9bWc0+cIugtc/8aL09LBnBQAcYklp3S2W2+yCepClFS6
OJSzLzH2Ed92eky0erqGk9M6ut1DemSUiZLW+G6ZvZpmoDbJdu1MlT0/kkTdymEh
+bU7Lc9PSvV+rAMpLIFNxAi8Fbrovk5GN+1sYAOdRHDkd/dGqZVhvFiuoZxw40I6
FEpGznyI9fjCUtQq/Uw8riKnlDssn6VVsCZyCYXQ+hqDY07DWe4UFtbLDoPHzYuU
cpAiRIGbtZwPVjbFzm2pVxOrzGgZx6/qPwF9Kpn4jouObqc4NSrXcuburJ4NFs1Z
za5vdDxYCpLCtGYHMdp543VyPZ3ZoLp8s+zEVKrs70LU1fOIc4CqlaiAvgLxURSN
kV9/5tvKqrmprVAxt7KgFcYgO0SYZ0rp9K4WlcFiq51+GnGvzTrQl0c7HvWzxGDU
lUlhvrFYMYx5IKYe7s8T66y2htlfyz0YoPGIoan74pIGHbCiF75jc+5X/SMOS2S0
EOG9h5joy9H/TtD/f2G+4HAbKHvBRNEsSUvXPwYgEmioorjzf0ib1/DujtERZvIV
UbJl4kfrtYBbpl+YfatyYWwEe43MifL1Tq5nrmmm9w2QOKzGw31Q15nBVlqhvfy2
MIA9/oDjBGnEEuvNDXHY1HA2KxkOkTnE86PoAQgAIP726xXGVRT4HHeut+d6rWUA
m677xLouc+MyzmT3DAlsw834fgj2FGf+SfwAtJ92zXcdZ0U+Hjak2EPKxtOSqLR8
p05KDtry/ElS2Gp8oB4suL2EXRxg3QYUtBcaytCP+lt/ZU0T5bEW8R7NQOL+YO7/
8i8UIz9BCZRGwpm7d0CPZAu8pmQHVxsValm5G3mVWr4kH0r0dPV6PSA34YDluTmo
Cc7K78AEDq7rUKCDrQrZQhWfajqCi83OZ/6PYd/97zgEiZ0N2jv4zGZEGhpsaoft
pOX5F9jbyWP4dQP529EQWK+Vm63ck1c2ETRkdLKQQfk4Eqi5NCAjtvcL1tAJZkun
vc23NSplVO/cyzJJETAnbUY0iyElvYUBzWfnHLxhs2jgYNYkGi/lSx4G82mWp+gJ
ed5X+2876/W3qNDzjXVPkh5m1W0lY0OUGjfNeZxYVlRffjtEUFie5LRQXw9t/Jut
HpPKO6d8OXR24TVz+OuDYQFwA/0nfHlGkDdnB+lf8yFAmq7wA2eYeTBcJfECgbaG
dXqISX6rbOhamJDxxi4Qf7g0q5+bHOujKN0ILSChjDIoToE2u/1SOuool11kMOWp
vQZQaHN27Q5tB2NQZ00JRc0jA5POkYvgq7zOXVkjsFfVZgcJmfOQ5vf0/ldDJbJ9
KsCKC+jHcmjYsAy7jBLBKCeEh6SIvFTo/0NCaIJbFM59cy/6C3cPbrNohGshth6C
rLd3+uvVzSSF/BUGOJtoFwjLBQ5HzXDicLT6T+Yq7wpnmuCcp64LqpuWnXdI+/L5
CXUBEXMQwfxxkFxXDFS4lefl2+kMkMM4SKxWdv/Lkf/Bb05woQ+E7ZfdKS0s6Ud7
aGJ2yOoTZDjDA9EChazrS3kLFUXpZJ+Bnw/VitPSxBvJNS96pJx+RWQ1XihfswOg
FIat7s4vcjP6yZD1D5sj5Dm1pqEMlGsy9IFnZ4/XjmpX9P9JSxX4xtr+LdqjZonx
XIajk1VgKRAOITnllgU2YkfIJ4E/JRf2kHeWvuNmX3UJnz8Tt2qHDktAtAz5/7xd
Me5OlJ2X91VAMO1EYJMR3ol6vUq4Y/V7kEU59NQQvqL7ZTd51Ksn7HFdCZpL50ui
hzXbHINlfIcyfhCszEiVIaLt0q/x0s3EvWDOyaSnYg8ZPsxvZpecSjPQd4ginob+
zgQXKh0dGtH7UMhzxrbmxai8vdc4ZLau+AwVPQldnZkWBE434jxSj1tZTsWSIpAH
qB45G7PMywdjcnFgs/su9X/P+hztpQKpjVerR3kligViOsAxUBRWz5t6zBCyR1qf
TFrd8GcTzwUXTn5EuoY1+CsG/UVIhQ/eDl7J8VgjitBDoE0zFZBGNINFRcay4Hrc
psXmSxLpPybyZNEEuT8bfytyE8I1J6AZidC6Tc50hJ05hq3skNzPef0I9oFekY6S
iFZLqSeWAAVsLIRyN2IPmoIhnvP/C0aWY0yWX7vWErkps7qo/bJsTEKMzJcEntGu
YmyDk+YQ+MPX7qSYlVhg28B/DTqISJYC/x4sSJDgA78P2SXHU5XL9YilUiAmLeQk
EILSwtGrKqk2MBMQ8RjDMhX9mJk8ZibOvr1Z02x7Xa6QAtzMzn3L8l0eEjgFIA5o
oGfLfKxuj7Heiw3YWfbJOJ0iWdTuRt1Zg1HuB0WqFO0nEkIgmxtO2w8uMyLLQHc4
AH4/GDw4/hWY5/oV5CcE3V/Qxfs7XhwkRDWWPjG+VudRP1rQNZfwajKmBGglTz/v
Onhl1z+O4/TIJfHpRQ05Q3J1B/Uq6MpFYdTsdGUuQeuz1fGdgsv+2jr0GzZ6IBDs
Or+5kLH4oivMMuzy+3N3klETWRFT1tktADJEbkKxsbtORjEfBucIfGNSqH4vvAps
N7inhnn6zqrR/CFK2+VRHCv27qGbgXz1eQ3kB8EuB6g+Be27+MB/JHjPmra53V7G
+wS8rmDHDq3E8YxwdPvDsRpbGFTqJJZE6ssnK+S6bejVir1W0+iU2NX8d1ngdr8V
Q1WS45DO8FxxTpZ8CYfUhtnLiL5pd+uX2Qp4bgJdNlbgTpEGCmFIn2qxu3Egb0Jp
Or+Y2VLK/BoETiXMOA/kU3GNNNjhc/0e7Qphc8HfHL/uhgbD5KINJJ7O86Q3EI08
bvWa5r8T4MV0WCbut41RiKhyphJHGvStqfvVV5JpQ8+Zf1Ewu07zUWvJdCefiDY7
Q79E6JQ9d1sbBy/X7IkXfk9oFnXxMN54cFKPD7WzLciQ9PZrR4yRfi0/aaqWzyUv
2mU2F/uhPIYa6/E5XvlH3LCY+V++UM54XKpeE9fG0x9v83bIwo/S0YXq9NP/88d7
/eIEdNtUvRsfMXaVNge8YuieQGNpjvcRU1mmsqzfzgu4TnTt5caNLghnuwQ8TfC4
b4LI9OJS6QO+B4ReVSl3tQPSdNacWOXzOOPfR9T//58qmgj0WpssOFDeODA47mgg
d6mgrd26uWvdSUsp+gf0oL8gCwQJ3dqgxdAO72f67OGHMxL8QmNpBngbU2+9QlGU
yYhkP+P65Vg+nHG1Tcn9ur67pELVIlilQvzJ0bGZ4w5AwBgh0dSiz0URjRYn1hSV
ou2wA0RAHGVgdW0dKLjEHlObkxXZMcVsBoYq0fa6q6mDWFP7hFCYy3xJwNpjNRvP
JVn+ke36fMso22U2VMOBCF/eiod+QNlUTV4eh+Eotqz1wbZdOr7F6CNu7XActpoI
Vpbz3C2kk85OgucQMoUtiTPBaQs+nIpZiIBlsqrYwcZkR71Ig9OPENjGwrzrgood
5xcDvJevdGEr44N+pYcKaWqzS9vSCjk0mganGQemKAVZb1OIVLsEnp/godESXsXg
CCXKWpXbhrPom42n4CFl4C7+j2/eNNEHGU2pTlv9CVXyWgnYFaEZ5RlNx8V9FrTA
pcOZMp9ui65y/37RXPe6W/6/lgzxYjEF7nBm9qqkY6CIZj1AGy7BZl9TlXBNaTyy
vVCwtbmXgtoibo1Nvfht8YWYY9vIukMOQJsVnIlMD3lrfTWnKAA47SldtgXz3b++
XclLQRngHd0ytYkVt0NN7h2E9A6KOyftaWFXy7NpZBzlYfzcSHsT3qsvj7DfvScO
F01mS3zcMuyOc/pRrVVzHlU25I0EeN/MmCIcpBdB1NTMcDqlHlcu/BiBifYW87m1
vn8KabB644KtWvmbHSRjihecrjJOhPYQ6lLWQqr7xrFePZUpZNCAn4Bu6DcHDJmu
d2FkAK4S/TDyD8aC+ZKuaHRZ541LLF8xY3Bk5fVRN8gHl6wUdGATM8VbjuTmxCF+
GF11ZEhWSfLeTBSCTA4dm8Vn+9RZ82gn9lFBu6n7ngWkuFtXDXk5yv0RYcyEaEnI
j9JKkTcIjEEgldVbJBkebgabbDpRSIAjHDTbktycShmr7fVSH0g5IV+3pg2MdSQF
Hp71yUG4MAXJiLPjs+bT35KwA+UUaeaeS7RLWnQbBUm4vdr4s2jReOjOk2PXN8ze
wA74orjhAGDwnp7eCYyycIpzT2CuDmIA1nLjj/hfKDtnFFs4VR81sYpfL5rBOfRW
fV8GHcztBVN7kLwTh8Afaakw34Mzg5VKZ2mWFUfJte3WF4nfW3fiQIOUfGcq5q9y
jHMqvdL8q44MHwnqkqsM4IKB7MDnL3I3CEFpGtIMhVPvh+N7Bf8P/lPRAoewZSKR
IGe0PrsmoPYxu4dOtI4hmwP5eOW2MwKi/Da0SxiU3rJ5sYuYZBJR3JfdjAWDTKqj
sWMP3E6yeyGUnVvQ2I6j45WHN5jiuQ+Mt1raSy+6k49g01vcmwQ3p4ldijrIizde
HvM04GAmqt1znErmn5jeaJwcxdASu3NEPk46Tks7uv4lrDeCPo1yJj/clxENtgQQ
M63OgvzgbYHdMqapq1UmBLbNUK0+IIBhhRpspFSFqhIciISLL+M25bANMsVbH9bf
xR3euwhsdffUA/yVJdM4UjiBCBSrZbvtujG+V4Km/KaMgcv8xD2+9u8CIRQ50UOl
2yWj/2wDNnh2+PDP9s4y23ZVPPoYAYHXcAXaaEzXTyONN2rPODDRFgAtIM+gZ1r4
ivpRNSd2dabvVQYD6JvmMnUXStitQWdwn2gY+0p3gSFbxp/3dg3R6qwTU6IfUGfS
mIX4yeGsPAX8wvNwMO1fdX6jgFDPpStsk9seiO5cXsTIOEVtqKgMs0ZBRglA3YNG
gNIwegxuPgxJDkO42m2ovHchMV6nI+lYJV5WGp55Ct0tne/nVrUlRzQhtMQsqd/L
HAGZZ8iVIcjptWUl0jUZuI4BiaUTo6txEHDkOIwk59VZEplXJo8m9kdzjzX214I2
y57L0KbLbmA6IE6g7sd+OI9LtwmQM2gjU1q4KSknGpV4N6g3B5ArrS+SOV2y72L4
Tvadot1uPcd1BCo55ZqisNsTLW8AuG6P/+UfvISe6mFTPc/9B0iAKT6ORETn2x14
F/tj91195O6TMmfQ9PQU/GWgae049lY+OXsmmEuJBTq08Gt9gsT5YFIpKBe9rGFU
h32pKXxT/Tu1kM7kJYb6mz7zkvAuOqQeDpjzhQdY76WfHNbpCF2Fhp/YEcZqf6tw
2cxcHQXOcJgH0z7r0p+Mbynt3IM0lr89BaMQoaRyDyz0WuXLIjDBJeKOTaJx6bTK
r4nZnuqhfiBKTeUa02MJbmx+rlhb5ZRbX0zEWcZ8pVpAAaFtDYQTfkRTOp4DbRKo
wYLBkfZ7iapzAHQkygbgKcmmgr1VlAmXJkbr2nkGnd0iyyjiz2EgcDn/yyYv4vZj
7NuwfTYMgtMzIvMPDNbq5DMz7eF70/9HVKMblL5HpPPgC5V9T09wUfbCzmKiYufH
8t9gaAqmbhBxkPzMokFJAYXeWvcRsJAGhHEzf2uVhKVgE+nx8bJhTBXFY3ksqMOA
0DAA/BGFmvPsD3bK6iuneaj7DNA4iiEo0E39rhmy79POTlUrT6Z1oAm0Q4JAeS/a
1pd3sEiNMMz75HYo/IOaDsaDoTdjI6CxUQcF/XoJG0vFiUySdpn7pWm3ymID3Ryw
i4FlWPghNnw26+tU8hc597mZqruaRNczN0h4YYYY9kKJvT2pHi3J2Da88jmbRVcv
3321p1jCsAfDq1HgnezttYl+Ry3Uqz/NIH/Inp09eBi6soIAkZ0fd5Zfxh+B7qTl
zwH+RhEI3q6lxBaUphgWSOqEnl3/dPI2YZSfWQglQeFZNql89jM3V1M2HNbq3M2Q
+cmd5AgZ8ks8s45spM6C7A9uoap3K5xtU6rghcUI5VRxmV0tXZmguyp87rEYJL/i
JcYUODJzKFSPcabXnAQ+EYB6BYC7hT7z/QeSqOicU6Ujo+R5Kjkf55J9FdImVXvT
tgTcTKqvYLmCDnyIlOA5s6T6Q50bKEeAyrTilZEaZaA0l7LKgKIFWHAic0bruJT3
IC3jfzMPoBWFskIc2MqOr/DFEOFGBG5jMNOwep3+DqyPK6jleDt3HTxOAMDVLOkP
td2c8wqxZNO0GEenXomzBFUGRaXOGJkoDK+P+MYgfYfUQRXCf38onXkOuMqegqzV
YGHPYAYWlT+OaMQ52CWPXKcsyDUyz6dGQi8r31Gw6uB2oO4CdR8eKdD/JVADNdL/
/5q27M4B/UigIRfoao5OzZEK1H6vvmfzYqW/UabDJN1/wo1v8vA5Y93k5JEosNaE
TMg8lc+DiE4kzNZC3FVv+JgHQT/dyb5JGg3I7y1adZuhLEgWIaVnLMSEoSKrUvtX
p730nLsHqCZbdCeKMGZyCXxPFxZHvarpzCmtGHdyquUkXge0BpO3sOuO96phAcLI
VqsutLLPjmpwlM7p6DqkTDNWF44YjarPXXee0hGB8NJMpL37WlRR/LaVG+keN53C
XpL3oRbpfBiwDOD7Mw5lrbpUVFwxuPRnlxcKnOg1evqaeb1gQYTSLzJOyyLXLID+
+cIEd7DvTLgFdsZRXojCgFroQUXFv4IozuWwWvcjMXcGe+ehE0EqfpuOvErCbImV
SGjrZdCD5QFq2Jp4otDwm7GZWH0pr8AVcZ5GVjD8w4ioz/7AXDZu2wK13gn8p2EJ
Fi5rCGQQjwi+LKNtFbn/YBcAKpaxdpweTn0TeOt81Kbks4eUOrHaYnVMhngRWyog
DyefeWrR73ZCrVU2+PRUsY2H5qpFbppxq5mGI/8NaPolTTWKj2uva6TZyv73yfTS
wA4z7Qw/fJw6Hg6hHJXxDSW2X5Au2hUOyrSexvt/NDkN5fkBLQfHUCEhFEBMS4OM
lxNzhcLQa0b1ds8LYuJCWCWZC/aLkRmGBL/b+I3rHpBRhIYNdDnWwbZtmVQMSM1X
0VdcG28nwHHR8Oahcf80fkjRPcq2E84js+P6DvNQNOW5HN/MBrnxFqVLKOO4KXZW
i7/huKUfxWacNTV5vu5XeDxkhsgb4Ckrw1oqrIhZlI0jp6WTupjswW3jQObOFL6F
3qtL6WYIfFbhrauSK8FdSp07mdyl107bOjblElJXz7x22oLXH8NZ9XF2sC0QT2in
gUGZ2dqfaa4SLU/VfWIrYVuC2djZogW5JUEA2UkLGy+e5Dq0XQc6NHjhUW3Ig96j
kx8GLKg5+sNgto9s30djk3uHxYBGwUGzHCMI+ZPg8RmghwJTYwu5NBjmeQXk8KZp
lLGWMMDlcgAE91nCFBqWKAXbbpdsvdsklyBVPgH5syx7oKfJ+tk7JitdfXBk5s+A
vF7vsBWxSUUraZ1zN5Fx9czzEBbX0AKCL8VZ/eUTJkWnyO8BU+FezRVM5pMeZq2r
+SRzaXlLVrcVl/Y02EEmM/7HsvCFfyZrtFtTa/yjzMd4Twea/GxX34E8+yisGll9
OivQoNI6B9ukB1LMH4Rh4Q6IHGfyDxH20/boKMXEetgm+dSJsTBK7BC0JL4cFiSM
c1YSqScYhxebUgmO7tlUGRTCyLWpclBWslRNaQ1f9Z2779xH/JwlGMvjM1JIlm8A
wLfuhG4WXiDlksAMY7SiVOOX4KdtFr/YsMgk29SIKKyJUCqxbXxtfMXHCTX62Irq
GJAN+FqrALFgcPAGKaQ6cSIwM2WYa8vFZYYyHkiF6LSdcF0V03y4QSdfootMPQcr
ocVtxLeadV7G0uiLn4BYbiaLomrTy6Eol9VF1k3mftyZnZ8gF40VXqkvSZ6/0g56
S3Dbaw74+mws+ycIOCOPiLF8lPrN44nexT5UpPLZTs9MFBmDj6z5oUQ6vIarmhuY
aQtgj5QxlY+YXBibL/keKggNZRYJTM2WzQpyi68gu9o9iJ3tRQL8vOBbiMxCe0Yt
/rWf60TR0ETcAPwIrIRwJ3j6Y5+RSmyE03zKpv+QDVXYjRD8qNXelnZ/csB07Q8r
1ZSSjoo/fPuKlI5OE46W/rdq2+ZN0NRGoHyrEgTADRXljV5gaezCty55oUkRX65r
v+3CN3AYAuAQoBQCHJov9aaoigrsl7uC2/g4sqXV9xxBHJnIGFQAapGUjw+gpajV
9jyFdyxfws0e8upxu1C2H39VxBSmt1Fy3nO8CFoWsXrpqvbBQjTe6GZpt5DLlJ3d
6w+BNgXBA4Hb0//B98TjfG34cUz9dqTnkK+2915eE6Vx7ebigc73SoQGLnB1VvCU
8mps2vi3HntKn2HjPu7fF3z8zcW1CWXDL/tGHKYqXpWp0eYhAbtKwFvAAnqDENHl
E6ddr2HPj9j/vOMi5t6XbQnyOzS1uHR3kh+y3s6PdLsU0XPMhjk3GqrgR//yV53N
2M0hGSiALU6F71YtgFXA0+PXVDLM9OdArqFw7pB05440mvENdAqT0xFE/bE0FtB5
p16NJaVqNSyaunvfwTO/jaIpWpm9G57PL/sOQxEV91I3rWd2EMyGnXHsPU477yBC
skyQeMqk8pnMU7Gvv4vp0Ek+2R5J6jgk5O/2Rp6MDTeSGbpns4nzENJWlKSMWaco
h6TX2JNsEMObKtgd16nUnokmLtljPptR14cF4PrKJFhNsBbm1cfTz0NLsQuoHQ7t
iQ1V4ylkY5SAwhL6mjE1sKsaYtB0rPP5BW6o7mkoRQ8twT30C5bNZ8u3XglIDOeA
oS94K9umcgPi/F95ydwGVpE1/UeNoJbF/tRfXcbTjHMbnDovbHCvNMESwVD79sOq
3kZ7CGRGCdZzIoNIQxzaB6E4yFg13hFtKlH/3ClwpgAzAJWC7QQoIlxffnAjvZ8Z
DSgQoZ25JznrEfomCxm9Mmm4lWWINsQZ/x1A2scd1zXb22djSyVk12PtVNpRZvUY
MN6CrMul8a0zCLqRQbXASQNMweX/XgT1k8mdg2k/vNbnFv2yNh6ygaAvcrLFdicU
PfGTL7sMWX51RB+xMrfFpOpWvjc9Qz0Jh8SQvXUX6ROb7H4wjcs3eM2lhw9isS2B
3yCAtpE6sYti2OEcQwWElxOLKOCOcvjpFxkXf7vNitm5x7lVTKgHGm5sf3bM65YA
o1dIMPCVdHZuCvjSYe1E/RFxhlUCdO0uByHIEm4PoQGUSpCJIjd0XjfElu45lKex
qQnfs9T+p7q5mm5ZP9wWuBHELq68Vw8BEX0jnZGc6F2Mh0ZfDkUnN7iNuN1ihQvB
jjusA1Br2nR9p/blcp481ghhB6qYNjwndzac42NTiVkko+INrkokUcdRwRmJHuRR
VayuOxaXS8b4uA7uHSaU/Mn8JpcvUQzfAZ803Ak8Ypo/aTllURAHInRQm6EsebqW
ooltvnrolJEfprPf5d6BCmbub9V4qIN4c1ouShT6UAWYuzqwRSRNOBJnLPQ7SvgL
NAjz2d/zcOYgKswZHawYel9vhjb4f0+vgFVc9ikVjBgNxKpVx8AUmHzG/k2UXl+n
b3uFy7PUBaXPZuU1I38cqmc2cRI7KJu3eq5rNKmO7Krxt8NcNO97LyViGWdEyWuO
21L/m/0dDSWW+tXIhwSGS0iUGBJmkPf6af8575eJHGEQcRgL3ZVOjjeEAKXyIJ9h
995kpuksBxlEig9GZta3Pvid4LiCYRa8XEn/GqKBTfHtJZlDjxTR3Ryg/Nyu6FAs
uxlxmSrm6zcBGnwRlAQz6kOWytqPJqlGq0qanzSqSjtck85KZt3sf9mhiWwqVUY1
CIM6phG3Nfk0f3AfMVzXY1yw2xJaQkIoKt9kDdvzrkP1U5jEYdypHLHbm+LPASs2
sS4xWoLr0sHwXGKlE7txXrRpFv/d6tYk00sKTET5qJ6yvBIN5Yi1jH+q32bk956/
xaFIfh/jJ8GjEUJWyMxiUgjWWz2Au0gNsEpKJjfmdtsYkWAIQO0ok2w8SXLF9rkN
6yqPrHjDz+n2OmFlLvOy0ekbzrRJVpQ4JSk0TBkgjuKxQ/E5GzSKUC2avUr14LWa
p8ykrRTKPxs5xyho+Uw2akrPQrD8lUKhjS3UinQZRkaM1rOFWzE0mvh5T9nT/36c
s36N8zGASZP2REFzOT0X3FwILgyR3iHmmMX0Gkr+xzP3nlVkpfDyg4K6+W1jgNt/
CpkgIj1Z6oSxvS5LTddKO1JEpK3eiVyVonLrVpGofEq2Vq949aT9MdxskCfH0PWe
1N9Vbm8XLGwTV98NoP5xVwYcjnBtT0wVoosEFeqqZrX1rh8p52XYJ1QsADtg4mQV
doIO9hvL6ZCsr+X0jb8UUwaN6nvCRJQ4Fw+CmLQIfvckR/y/wIngmBDZPcx57Ozj
9FabOFap+AgNTAF/bHwjYJJvFF4G1z9iPGQr3FfFCmfaDhVF9/qGfxIt9hWPJoAz
JWzSGhujBiSxeyTkFs0hFe2ureOdRQQVkcdlpxLINzu2ZpBrTiReHfrVboTkvD6E
tBAwkTJItdkoUsv4PFDUa2CPVCFvwhMJj5EKbw16pEuYJAzb9QY4tdXwEpEIMSv3
fXnQbkB8eZgKFF1/fGgOv/BqN4JVyKGm8LmsuHUHB+vrDe5QBLHsUdpCyCUtlPvS
RT9wl+n0cN8cTyE/xasqTc2ENAOMCyLBn72YlBckT2qPrRc4eFrsgjRcSoxGEV9s
OzHK6CzCmhNBPr27r8A28CkSJXL07O733EwoPT1uk7yijtMTykK9St7TH3zf1No+
n8cBGQ7nKJRatmgzFICTdtK89UIV5Ynq/NxV2j+YJS5JVF7y9ZeS/0enW8Db6LI8
iAUJKj9bKQG35cTZ47PC6rDrjvh6Ht6hmMK0otDrzkuugiwVWunhF980iz9NHuEK
1FIRcvZBxnTRbRRlWySL5JydSYV5UalL16oulLCP3gf+OzMAFI2khIgBdybxu28v
bORQz0oIgOqeObNMr8Nfz1vvz3ePzODAs225XhiaCYpRqori+rvAPJaXwPDZKB5T
SfopaaIY9lQ46g9ZUwdMId+2OEs7JzTA3yZr8Qvi9Z8wMlSkXN13stak6zMUk3nr
jL6p8zpR+lIUuXSc26fFr2/BznI/iISETAR48NuljYR6yQm9Y796AGjSmhhMPNH4
rmiQ7fEFRLi9FyQLPmDSWSOMOcDbJvI2oE0vqNEyZxt33My9b42eVR+DPETapUwg
N+VxLZ1EhBFPyASN8g7+nvWDYtgspeXOudUAq93jpUY8Nd2ZrDU4kgiURmiatvls
UUtwaJGw2yPy4Kto9YRXX1acfbvPqIsiJUxxWPChZgExwyTYb6xJW5juaUM68zhd
8AYLV7TzxpshXnhCUU61oMuvtC4Jh3MstF4jSq/nASsiY4ki6a5TY1n9+tZJoXyu
OVgPKS1YKOc22MPNS/Fmk9m2vMvFVfH103zva6mm6iBlU+jyJ/GZSMF4bXTHBCCa
XOUA7go49hK3vGadhPRc8ZwUkaZwoeGKP7XgoKSH4e/Xf9LUPuF9GhbQJKNl88NS
2lxsuWK170h9ve55Caj2ih4GwiCEyUhT4YhgIMabin9+nIRNVpifL+j2V0oSxUVZ
UHMtJ1001OzbHRCJz0GtxPKhansJoHZs52xeiJRYcJqd0LIKpLAgEPUxOc2yGi8V
aEwoZ1NK2/dYjo0Xb4uphcyl3KOWRRa8j+2HqRzajHndd0qkOp0ybDy3snri6oS4
VRfnBBsc9XT65CiudIv7xzKVCkby8hALdO4LTZsDWBUmnI1bftomDd/qJTbwUQ6N
eooBXZOKmgo73MntLhz9vS172wYJwMDCLPliLZX4GdfwGX7TP2KvbhlG6Syc+Q2W
KM9wZyNF5ALX57iHH2MxZmCQPWnlM0ayxBFHKgIWOXzwqmeGTTZKkJ8GpZavmueX
J2WQY8kBrjg3H/OYSa+kGOQ+7Wze5HojkGsMHrS+GO5upaje5GVOeACexTpPUkKi
NEjzWzqe6nBJgdtxxs5X5e+u2xae78WkCB0TOYl83SZzAndkv9bS1aKSlbb5iBwF
NulAZPjZFVGhUru5+01FGG/kr4sDZ0lTzbPuy/J05BJpL8H/8rFf1/9pucXCKA41
i6B8tQAIbr/951dt1YqKvxJkijc+LeOtVvpCBIknleSsgIvaXaVkT4QdcPOomg8F
tJS/InSdwQ3xEerQLvKZB4HEEypbv0nNFbvSOjdiDK050+2waVty0YxAyO8nPvHL
/9AgwqHVSyrGR2Hk5n+CiNjwzBGTvMDPexAAY4BFixD28A70JN0BDlCr2wlGvh6+
vD3eVQ+/Plo9d1r8rTEgYa0NGJXOrn3/AqPAaqO/9tXJ8jKNlVLsI2iNtDKZM11f
iijT8397GQKfAja164PGHi/V1UxYBleeGmlLxfNUQmnyTJVz/FnyOfi0In8mcezN
lVZ1VI60DFy2D6jhGxNxA757apUNIn77hd0R46MPDPhCTx2QP0XFeYLdCd7bhQag
+QHS9VjXG70As1Sb0iSJ+Dv3rouqHs70dply5akycqKSIpz3TDPMYQFfvPN0lSCR
AP98pVxyLCxIVkO2QGM2y60JQrbxqEtk91f+xDkQskx+gSfGyPtjssq2I+2S8Df9
2iyNesm/SOohTYamxZ5VOaCBqEzg3t/3qnuZKkilY/vEaw7mzk93bqtiu+6kZzfe
iR4JMUdHHPkKmemYeRuvqoH0en4/OOfqGyKJvJ3yQQGwoYw3tTfclOSQHr0XYMmP
ElMm8z66wPg99WpFJcM/WFsIvkhGIXWV9OkZQ9SLVADhleCHMNZqgVmapVKVhiTC
nZnLGoZ7a+Iw96GI8VVkGV5f4akEt7ejFiJzeUHagfevYsKKvf/FWIw7HZWyxcaK
rEXOgNK+NXTGiV73L4RjY6peRMPp/o8p9t1U7BfqhvNXbuEwQIq6HZpgNwmdUjlt
+ztfu44RDZpv671f1HYTurMIGfs4uhxzmcHi5h2r7tuSf4emaJns4QuUtcACvZUx
L0dKVyTYtV6+HhEYlT1Hu7ZzSlzpykw8DlMeMMBoysPBIk7Oeu8hhvjOH4lRuoRe
ugt5f0zbXYn9YzHzo8P4euHXICQ7T16bndrhP1ZTCZwvqce4uKpApslR7uUL7x9i
P/YEZJjkPfiqe92Cl+NMoWkgvl5KJhqfd4BXrRR6YA0WmwyI/5ZccbcZZ+2sUqLR
8mQ7urCTCvHOwQITcfQ/YCZ8YclsmdaD7mAKcy1nA4MQltp945W7yYBh/1dfnpnP
g4dJnx9OoaJjh96JMHolz+p3/IHae1co7C3/AEyW+eKZd0F/VwSZ0K5XtgqjY0MD
7Pk9YhUyFTo+wg3Bky0F2J9OHlcqoj8SVRb4OD2Ki7FpJcaGN9RVHsIMVYkIVvB1
uFAcf3fWe0zv+TSrV/njjmd8OPivJHDzW1oTHcVDG6TsCbLxQ0eibqJKORGVRRyR
SFnqr7i7wN/ZXmbnB6YTJp1Y+PmF/JlDyuUqrE20+Hewg2LIs2q7Qe3DShm2rzL2
nhxS7Uu/a1+L6tisIBNvZMrcG2Vz3E6zDhnILLCd97DIJQr1VFatr6EAqJemTOD5
AXQqWxACOYJZ7mYQ4XaGtSM6HyMgnrqAjJKcBA2RMY3tD8ga97SyqEET9wibK87H
i7stjEM1oVaF+caewsv5s3mq8bLhwJS9Z1Dn1IHnmB1jnyA5kEyGZySdaa2Ag8Pj
f2DM1d8DdtqSbPQJYxoBI7oDoykhmlL5e6FGnV92Jv00sQvxDojDPpb///M9d7uH
JGZKVcTNxOjMDYGU7ZZk2y3DUGiYzQOmKYgQbLPmIRT728yU+iluLCccZ90LNvrB
volbLx8YbwlfaoxcWR6fRK8VXrFAlpkS4k/dapPzD7XN2ErFlcFnmepDgH7B6sVy
yfF55RVS2ojhP50l0XGvM0xVEOk9yarI13IRdhYmw/Sio/nzmJTeuWuV0O/OhaYU
M0M6sDSya58EBuG+OfNXD1GA6/ZSgOsK7ZmHHl58M4tTiwaj3DWVqh0aVYXZmXdh
x3HQPLZr4l7Zezsb+tpTqybkfpQyvKcHOr+IgzzYz5IqAUMmdDsSjZd11FsEJfL/
dXAbmLmJst8A8eoD3KE1DiNAhQU9nvlUvJhUFUvp2oC8sbky2J9PkY87hHSBYynB
yeWo8bnQkrcx8Gxs1LbBcZBrfjPhEqDypxZzpXmrezc41vlmGL818yeUuSD97A8t
XaOptMNt92ny6k2fQIy9eUgg3j8twUpUXGc3K1jAV4cjOCCwaddYTSjnMZ2rt+Th
+TYscbOcEtssqxkq1IKixHtoQ2d1eKjWiAoPrAS7SLMMz0VF+gyuhZez8ZadGUhw
704xnqNMkE/6FzGlofheOSL6dnOUrvPO+5ZDLKinl5q5meqsEb/dnlnYNIn4Eu0k
syksSG6WguzhL8OHxB0aOeaJKAYaIfnZ+lWEeD+Xgvl6P132P4iae2zpa+vqPlW0
eNZ+eTLyV1yZXiamaDfSwXmNKxRR0fBcTWrRtDNfFp8DKW+EwUfsbdnZlS+6TbNv
ufOwAyp0EO0swivaO2TbznT7giVBgX3XvcwQMsrECUozsl7LfnKX3/8wSU/T//dC
DPRgxnRlYI2k1F+x3Rj5Rst0+dCHGy4lqM53/lARVlj730lbJxaGEwC5ioLRpiuH
KqIncfR3S07bEcDUaw5kZELaZAIqdTJuieVIRobLtJxZXfGyCO0BvmN4q8tABY97
7H8KLnqaHxiIHc3PhSUz37F3CuFWk4StQE6SX8Xs+2C0n7F1pkgYpRTneNaYHrAu
XjPSel7AA0xtd+QTzGRkJbGsI1j/+xK/aj5jNIDJ6atyGZagFDg/F+6Qm7/kX4hF
z6DnkZ1IRRnfqUBQNZngsbSE9qyuiTteIXSKc+vUv/eQZ11lHTqOufrrTm6/Hv6+
va9kZZ6Z65MXZGIHZtP8ctAeOQsNM/biWM/RqHotKptFmnJSlkDFhEZtgQFu4mpm
r+KbIE/DNmbzf4NogcWhA5XwYdk+zKGO05TlWwQthU3iNa0zeAeHTukMAYDQ6Xa0
veCSkygISQcVQMsk0dwEjLSUrInJDejZGNSsgCeQuxEbYLaKVL0MEQMu8rlIy2F9
sqqDaFW6kI18Dfk37timZ8VMKtIWKU5V9nPjF3ySRvXlN+BuJUf9UU91AAUZYoDC
eZ3ot1NWXoB8mlxI6DeRJrL13HHfBbMK+VJwrKbavvQamer7GVLwRzdr2ACMFtty
sdYDXBG3DPDsLstT278eD9J4hSoWevQM1EWJilALFq0oTaFB4XlG32gneWiDtSue
iOuLA1SNELkIltBY8S3lojHXb32q7tn8yAQmS/NDwur+n2l20YR/jKtMnaXvxETE
lki61j9aaFaS9VC0oZs1QzHjhj1UsD4BOATP4plHr/ORmDf4ZcvEdOvber3ho0gC
KVouPklmBFOpUdPidCxWQoTXTztMQaOFXsjyzb/aWJpKRsUlzJTXcFLTbo5R0dD7
IBo574ZMuu3Ws+KV8Em6tNoelsyRHtIpbJIJh3Gi8FqjkkgnFdxgTCH75MCGEyQX
R0/qwgIXjkjzMqd72NTdTYW7OXBi7A7eKLucbm9yZZ/gOUZ0SpeU0Owm3ILGHwNn
YiS7YQZsk7qJUc4fRBEdNbpTDoI/og7JxJrtMUhZr2v86EAu5kAIRonty7RxCneW
yYvT8eq8vaYBa58Vt4uAVQwuiK5r1qxNgy0luYV2Bk52EtWfDEL8zFp2k93m7iHb
Q8Z9/cizgmG0cUs4c2NtB1QCR+QBxDQqOzjnW4Almwr5LDo58aLqxoI5RaQRaZSy
ulNo14h1Js4p6yVQ0lZXXvq4AC4oF6MW9obc0G8DMZu9QygMFdyGwP1NESexXjWY
ymhv/elLtU4T2W+bMtKzwPpFHmyL4uw7GGxaHkqxoXnplZmklf6d/fag0wDoNuzh
yeb8NOFOSMYp7qVJ++tiSnPUaVJ53GaWX1Dqk8tIvdcGROVlxRa5lpzn/rKPGhC2
3+kMpUmipSDa+EQUpgz13/qbyZzfxHiMg0SPnXYyp6k6Vw+zzUu7DcZt0adjE6xp
nKm2aRNpXpFKfKnGjnyUFZFwplFuguhO3A0OEcMKp7qalc4sjYRf5Xnm3Nnqajhc
UmCIM2lALaHFVrPpEGCaqMTbZ4dt9MQ6FHgEm4j8rfDV/OiF6zsfyEKXsDBmZWXI
t3b5pxInlm6YALGuG1Tu6Of5Xs2Pjdz92eBeW7xZ7IxmsgQiXhPPOWjX+i3+tMlh
AfZnw9/DhMMoj1GIYpzNjt1LByq7kQ2iqa51NtUcwGtCAeW8bq5J8rsSFpfOVLto
`protect end_protected