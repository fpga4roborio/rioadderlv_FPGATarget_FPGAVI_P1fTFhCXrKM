`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
ddtXksX2+yylW5zu6QL2Lhnb2d1sD00763mmSITNX595NcHTEkwn0zB1Dry37fOW
FufOhVzEJp80NC5qZ/+F0Vk7Ik02dIR0elf3clrjeJRK85K4e3Hoo4xn7YbFUIms
l/8VZSb14+JVGURjfswrIyCUotIzlzVYZ6gzoZwDXIi5gQIBf/gI+KxNXPaKV+PQ
Ufys/12rjO6aI/pPlqSm0hCvftmBcnezN2hk1UeXgOIuKZnogjOsf0iJVX2aOOWE
6pD/psybjbnsNB6kH5uFTA5frkzIzkzl5d9+YDm9OyC+k84E83I/7/j+rk4L2dah
QJOvksSIzN867/4Qt8qYTQ==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="MvBXkzurAa5VTw+1JJ70nePUfoQXBvZOku/SMmg4TwQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
oRtzZL4VJ4iwysPsC8SXYCzXS8Fw2gtZTOskLcDV+1B9Nzn1zTyNtlo6lNICRmmK
ZRVu2BmCc2G+fmzynYlNTnSa7C0Cuel6FYpxCBlOuk3OF2tzAmLAuDyOH3Z1Yjzk
a0aHuoCdIRKv7BrZCdALt03JeUmXKPdOmIlkVGFl8yw=
`protect rights_digest_method = "sha256"
`protect end_toolblock="Jn9CQpRhJt4rnzZPRk+dOpzAubz7omckX1MrFd4p81o="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 1280 )
`protect data_block
gD6l00tciPUa6pDNTk/+txp9YJ6lFS7W7YO7BrMYAvj6x5dueVnllZWesGWXkK4/
dR7lrgJAmoiN6kmqMp1E6aEVmrJicH8bcGscpAs8Z1+fv0Hk4cMZH2GJ2LLS2yHY
Dxza0e9G9MWBuShKGpqp803YIpREhnHfDgoC6+cG34Qm2NKyW/K+wsz74TSlj6C6
DOkhXCpEgFK4nQ4j4bu21UV2gZmyrKo704iHz+8t+S6HHg2Heg6EnRZTc/s+qd8l
KEyaYQ2eSfjnuAuNCferGMM2mdBKe09/E9xpkqaHy7/hAqUuRT1QN+3HCzR9wMOQ
HGao2YzsjgKx7IHH9oKheWQ2HMXh1z2DgwECnBVHDQ2wnGn/DYaltyfiL3tnzmhV
2R9qjUe6P0Py2JRGlugklKauqhV8jROH9NUM3sTrXiR3mnWi1ZyD2G9OK6i+hoCE
5rFvKh+OVg2RzslrDkFSaf6I8r2wyz+z+sQvcbdGQ0zuJqN1zbUq6YDAo318pGSN
1/qesiLNcw3D2n+KnYi8vwEeWnLZnXC4WH1qMNoF8o8lzvSonY5gr8HC7rB/jxRm
56PXy98egZ+mj4rkLKgzZk54+Hpw/tGddDjqTv7yUxOfn09JKJg2p+SBq6Mvfsaz
l0h5yAUJgy6rxKM5qIQqz718PzrOiXLtvKjCiixb/hpP9B4AYbJ7Q9SvNE7R8cQW
0kTHbsxav92GEorMRKLm9k8kVlmNf93ytkwkIn1q9+dc5mMD8OCdvPx00+VwoU4y
vi3lu9/7TWR3gbW+dKF+4ys5h3SHZ0B4PGUn4/REuxrMHRNrl4m0fE8Mz6U0I1a1
smaMAMQt1df9PnPf3vCQJxk08KVV6M31J/rb9aW6SuoVHazX9NTpq7VDzJ+lml3I
iH+x0N40Kjt45e1Uzl9uMw3Lb2Jfzy5hnGLCBXQ4TUDoIJuC9vgMtZdmzarUOkeZ
HFyyLluTBpAohq2AuFCSjCNZQUGL6OcfvxJKjOSmZJKFgdPy/ln9DFfM3c6AA09E
HGzZPPO4s6zdUtHa4IVUQCIUzlFJ7H4m2p3DqUgQypFB7jw8A9es3VonbbKS8SkO
bd8ZL9471iRDBnfDyeMzOlqbPfZFMIKkDLgXv3MD6kG//GDd9sJYWsErR2mslouZ
gFJT5nSrq2Lu4HYzzy3sguFvGzaKc4z8mOyKLqFhhod3a0L6q0JmbVJ0PYXnu5gZ
GGWs0iKB9SPGWVOS27tIBEWGSwTppOtIhzxiYegGnruNggsxi7HbTJ8w9EiNLlOK
8wMxqW+BnT/YFUBjg0RAdhOizHEJ1r/HOlaIg+E7hbun8W+3GCNwOEYMXCxi5eRN
dX6kc0Om0ZWF1AUhWMoMXcNXg25Ul8HXYp3o+7r5vgQXSKetXkQGImi1ooYJBqil
AYRuPchccYQdimX5WtQRgJBCKJeIpbUJ6luukyrSvPCLyHqiQrM9yTfkNg45rs4J
ZhNF4vjd/6n5aX5Clx8R/IKjBurgzS9skCmqXMxZGNYzSlug+naEo357qyJEL5oC
ba++uU2TDQlae2ilWoZ4pUYoLoavxrtbjfVE3AOLsc8+VJKGQlrhvYpaaprsFRvs
x7PLocVfkh4HQEtjdeGXupGEOovlpfBTdPeaa0sB3L/BaM62y+H+OS8iDApx/SC1
+SiQPEP8yBvFLS014mLGI2qTZKF+QOljuRLi2JVnfwg=
`protect end_protected