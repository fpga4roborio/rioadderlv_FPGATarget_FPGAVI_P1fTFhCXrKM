`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
ddtXksX2+yylW5zu6QL2Lhnb2d1sD00763mmSITNX595NcHTEkwn0zB1Dry37fOW
FufOhVzEJp80NC5qZ/+F0Vk7Ik02dIR0elf3clrjeJRK85K4e3Hoo4xn7YbFUIms
l/8VZSb14+JVGURjfswrIyCUotIzlzVYZ6gzoZwDXIi5gQIBf/gI+KxNXPaKV+PQ
Ufys/12rjO6aI/pPlqSm0hCvftmBcnezN2hk1UeXgOIuKZnogjOsf0iJVX2aOOWE
6pD/psybjbnsNB6kH5uFTA5frkzIzkzl5d9+YDm9OyC+k84E83I/7/j+rk4L2dah
QJOvksSIzN867/4Qt8qYTQ==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="MvBXkzurAa5VTw+1JJ70nePUfoQXBvZOku/SMmg4TwQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
oRtzZL4VJ4iwysPsC8SXYCzXS8Fw2gtZTOskLcDV+1B9Nzn1zTyNtlo6lNICRmmK
ZRVu2BmCc2G+fmzynYlNTnSa7C0Cuel6FYpxCBlOuk3OF2tzAmLAuDyOH3Z1Yjzk
a0aHuoCdIRKv7BrZCdALt03JeUmXKPdOmIlkVGFl8yw=
`protect rights_digest_method = "sha256"
`protect end_toolblock="Jn9CQpRhJt4rnzZPRk+dOpzAubz7omckX1MrFd4p81o="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 10496 )
`protect data_block
gD6l00tciPUa6pDNTk/+t0OO0nC/UTtBwLB41d4inuAUA3i/ALrNyoJVcBnAmEQW
ptbcNp5fxEUJjnOxnedyZEuEBxWRieZFQnkRdF269oM7mNxgLZtjdTN/sjYJ35DR
q0D+xJRoe7Cyaor8a+2kBLgkEx7Im99sWYdQ9+nrCiAgM2l17+8i9kQc8C0r0Mrf
DL9JqzULkr3ac15O8i+9Y8ieHlmTVw0+/Rtc5bA5GecmBIRRYkoP65c5xnlW8Cho
Y3lLPuyzSQpyhWVfgWFOgye4C41NiPLt2Kodn/nv2GMkN1ovBVfupEwEOfBaQTuD
Wi1MlI1eVQzcN5QUmny2hxBSvENP6ci5zUAIefj1BIsq1K43HpBLxaPR+CDE07pM
znYJE5vVe3D/8pI03xp3Lu4MkxXPGZyEr1MjKRzq0VivqkawXHcehMRbuiMuW4k4
s9IBrfow9QXTSmStg/G0ijcOPAm+oECn1lHwnm8yjTR9BnVd2FuC71vHnTeb1Hfe
OuMJUB/zZrAoNFVRIDuqz/y4lyyPB+Wl6aKro7PCOWu4h4MbVkyX0oqk0GrN5aUr
S8L5b+BVCTY7O+KanzCVIOfZsnVizUgNjPpOrAUZlQVd9WkvjsBjswLj3PcANqAo
Z3Pm3FevNI2+cWYW60dMeDit9qCNhBvf6v0qMLO7S3WRpRaoN/9+xAYfa27N0Tpb
IK/dQefHG5oHGNBuSIQyWL+Rwk0UQF4IbHH+yV9B8lkqQdSQWlKi+1Z+9IzI6Vp0
6eYoTM8JIm20qRO9Jdp/XVppxXfOwMm5iQuF7LazsPyCSEeF+eQdF0YyW3R6ZXDk
D3DNnXagNitsT40m08JVQ8dfMhl2bQWXKUA6pucf3la6LO3O/lsiTJwVCZaRkXqI
GWj16/GoU9foWF5vpySG2BHYkpBlR1NqVFjNPYTFeOBEhSriNnstoDxeL7AHVWDM
R3UVNNJFfaYYRnHK8zkiwO1AS8e4a5rvVQYegeX2dtLydIGstn+eySqXb7saESWN
zjatZlEDEYEgyYKP4DOXQ1mEGR/p9xWf0IgGPCxSB+vtNzAs93h2ppxvpqbcst1N
i18VFKvyzkcD3UeY+v3rt7swxVBODFY6ECrgKh1TbhMC+4iQrF++GOUOqB+mNvZz
oft0D2LKglh5peB22BvObzWseISJn1zX+v5nROB6rb+C2C0TPHtsnHXyd5TwSsoE
Vd/Y4uGoCD6WarWhFw9Uz/gwxF4Q9LZL1vMuqfZ1Sorj5DnO0cPpwOVe8Xu06u1z
TKJ94gcjGCKQ2Qd1OBIBiEHTfpqWXixKkwkkCzVjjLy65QNKCwN/meQ40oSdOAxs
TyWwwbLSzJJhS6qOIJO69Vj8T0H2W5RtBnXGxEFWugxx6ur23WNtZmtHxZADLhs+
GY6WeIIbcn9/U1jhvMuZj9hedtw1XX47nWBlD6bcurl50wPcfOt1RBALhTpA6agM
ANvnw5i6eRdhyTvp3G0L9Bv7lY4ZfZ1O0aEkuTd/Rj6k9bWFMz+AfJ5gZM7cCedi
UE1yCnwQSBMxNySjMhr42xwzERuEZggRYfbpmgxfAuZEdyrYD63O6Wx6bAJSxuCv
8BId3f7xaA5Ui51JBy0I/TRpCH4jyeV6LbWezKSSln23QFHd4fDC0vti6uH70YdV
TCLTFUbZIRAvkFYGWRY66HP4IdE6EP3sD0XvF/oNGPRLr3RS1D1Om4nr6KZz5XYR
/CdI1l+WO7KJMhgbqQl5v5Ukqil1jHCv2UFuwyujwaLvpVzxsEGuHgv2xoWGevkg
y9nPUn5AG7X4it3ZPeFUSlc1PYoBfsVCtY0sRUVU5R9kZC5kxNyz9dy96VfExx40
TtfxlmSauHDfRdru7ny7SWYM0lkrgXgbW2raA3T7Uf70PJ8YniYOEuu8+yE7p8KB
5mChS2zlWT8SzkKw9J7eRr4Deo3t5gs8rftoO4FxnVv33GjJs8qe6iPDVCh6pVqp
etloOJsb7m9LyVe3todJ2ExJDhA54nGkE6FFf7eqEOQ8HCCV84IPVgy8P/j4xzu+
7xzul0rRiMzg5/NibMuUQOzoWI4QzMAwEaurUHFMRd70FADJDT+WL21H4yul3lOU
L0gTRBbpj9C5p8mdJ/Vlr/V+Z8oSt8aV6iESBfu8DVLP2J4uKijg8KjZeEQt5uyx
d4B+7S+9Jjto1ql4t7stTfz92pHnN/052W0G2428eXQjMM+A7tdv1o4FyuNDe4cw
JrzqanFhnTry2pQJe8qi0m06eqD0TmDCIYmT+ycWMhIndTKLrZtOZcu0HzqVXp3a
P43aqhqMaSDlJ+0QvLW2gFVG/pGt6vLZg29Aew6IM0/v8XzmvbqRTq9Wtr6/ZU3q
6Cp7Ojh1h4Pc2w+UAyeE6bqo1yvLBx6mTCkJcGe1z3a8oLvANfPVZCdnVWkhbRyy
PTmCz2Blfj7mutmtwcL351SkzVafutnkQYSoXqkXvjSBwod84XpQeNjDsBos5iNR
5uieO+nipxh4QD85vlyofvSX8Ot4gYF7T87sU5Ey9nCCSBCVPasvMk+CweL4yS5u
0VIQmlBhQUU0AzSrefnDCxKpZ5RBHe5CoP29qEb917Jo+uiYcUoJcIkhVrs6DyJx
Won8U3TYTKylMUa+wAXxR0au2laI6BVWIdCZGw2knzoUd1QTVPznPfrW2/olDGIu
aVfr8/wM5h42fn5AWoDgZzLMUVK77AEcPrbFk0ycwUJM4WH12fm+og/dD49mU7vP
QpVAYcndx13SrlVOPfKQuK2VNHQcIGuL9eF0o6tQwvhJhyyTO4GSOzZ0FxiyL22K
IQGhkaaYjm3yx4u2KPNlUdu/+mIDEqVlI1HQzpAT+uY/SBbUiEo5fKCAncApEuVK
abaJHeAcmaVzl7lAqhT2nkAyzDgSskjNkbw9x1SQHnuoVSLaiRSGC1rV7aa67RTu
y8+c2ItgIqR4ugUhxAQAC8j9KOkmqbJU/BBN8e1qmF/iIRA7/6XPyJWPFl1Jnv7q
tWYNbo2IzWaJL1lM6yz2Hk+MTpwRJCYEVcXWUyAgz7obgVGZowrhjchGXXBrYg7d
ctdq8DTBOfolWaqosakS5wmoDlUC7+MeDBTULoNHXji4Mm7D1dHqZjjSJGMZ4969
h6CXzJDzPLRG4MA5rP+wGhO1id9xqzdSrFn1V+/OJaAVQn5Nx7IiK93z0PGZ0AgB
MSZnTaF+/rcl8K1q2WhykR+eSy4mJ+3yS44Oa4qE6fAWwBnYr0YInyo4h+MCoToh
ZHrSQtT9kTQflpGETmSop1IdJS0QYJtWosPNUpMyMByMyS6dh9LhVGkEM8eeZkNG
CqIPogsQ2jt1KfrjdfjRRrejm1bnnrygvKFfg10cVMW6IF1CocejXJsxZoi0ozwW
gRuZOxvpvKPHYR/r6bMXygS8tOAoWr5vYo7gD/WFA7oO58tOi4qZmlxzv/QzCHmd
3XAWGhGpI2f43RiYKtY2XE2kOXqEpOB4LwtE/zwXsQrkMV4Wl+IFkKobJH6xkPh0
alXmwbM/FVb+kGIPAUwSLVE+2GtDLgrE4e1TQikPhcuXUxYRd2+9LmhePvLmR0Pj
BJDwaWFEClzTI2Md21/x81DJHOeAGan1/9bi2YK5Gro813ejOEkOjybKBdQRg9yy
MlB7kH9HGrUSBHStHF66PFGBwGUSWU8Au2FUz1eOw7krRF+S/5dS8IikPU4SKFoL
OYzchnc0b1abfmCbK11lYP5TcqYnyHkm7jsCHHN4UmjnQ2x6imQhAf9grMWU5j5E
M4cy8BfBsd2BD0OLAXYey83tWQR7yqED4ykkU+k8sKxgqoFqLCCBzWWkSX/aWaWA
PeOQ815xL83hhOyB6HkM3QIF+qqawJ3TCQreQcbHEgq+7eLA9j5oTU/tphrXC7UF
666DbEbadWsOXWstlGS6Q9sl/o5ld2aOIIqoQCC5zocgVkhvyAD9wNlyl78ftZ5H
0eEBfIRTQJxsifYoFpQzS/MispKVSid7hUlVeha4Goh5SbNrxRc04dlEYlWGxhrB
4mhDPxFOdA0Ig6kXSEcune8uzo23vcWmBDmTYW6P5NUPDWP5iwHldVM9sUXmIzG5
hTBL93CrvHFbZpv/CJFYKsL7aUp/i/3MxqYvp4HghJdbH1UqmZGu9k6NqnkRRHKf
xYVnSDVyY297NeCuBjd+X4UENmYKnPfF+8QLXMm0Fs7G/UuiTcFflQnKCybFYvfq
P56D1ikZ3WsE2R/voxlwJU7QICZSvwVw6X6TerbovFMVOkw4yspExaG36sEh/qGx
XWHQiFlmmPo2x0UzER+qUvvToSOvkXF837H5bYMxbWrU00R0FwVDyBjRJmdOQ6Ah
8h+ytGO4rYEl5CDIPNsKWN4rnHxe1z/C8bP0Yc/Z7pRdMcYKbu78TAiR78a+9hFi
He+OSyR29wm/ARZdPtpZFeXS4OtnrXvtR+hNYtkMhY9GXXGEJxYa6iEiNkSj4fDu
kxEuqqqNihtpCVj//cuXZf/8uFlSo5tzaIJ8tJ/ctjIj0Iq4GAdsWyWQ/gGYYyS6
JGG/hwMAfmetT3w5Z2vUN3nw64P96uzEL2exkWCeSwPArwrQWR2IAqNxuNFcmN11
vpnP0BvzBZyVDDZasUsHizfVs5tFCtp5YXU7qrs3SU1UuJlacIEoBP4G9cFf9kB4
iFhmtcKVWbIOG4xfVEny7xnjvrCWDvcvS0aRrWyp7Rs5VcMpjMIDlFEd9oDIBc+2
FqpszN746mZRFwDq8ad5Bait9KVbpYjvwGG+hyhDDFJnOg2KzfuYmmWhHcOogfCj
65Hx+TGEqhDQBZg9RDcSbkkCH4g17xk11uQR7mNvhMxdKSYnlHdaKurEW3xPUIGh
0pqjHCupF1ROAr5JhYO0HAa86evQtP92wCDqgttojAkEzK5FnVxyTCOwScH/105n
KAB+spQviBKnvjNhh3+AFgcpKTtL8Aaa3MC13fot0YoYC2QdV+n0lCzQPLndO25K
cil4u0WCjMkk8QddCbW7Ucf8yRtGaxNt/RRbQmkgzUW5iW6SyiU4d8Cnr05II0Rx
gqTYENUbt8epfQB6o7JguuVe8KD/3rT8nA9dTi6efP0s3Ehfo35quHYO9yCLGfew
NyBIU5ww/VVoJqCutZGZ0m8Q/GLHt1jYK6adHAetP4Yp4NN5fVD5mKEw//aIoGzM
2JkM8OFOPZ9Tdzl7k2UAXk+uQdddaRef7BtWYkLNWorIIaeO7XnVrRNYVRloojPk
jvi4WDlmymf6UJithBmXX4t2wLw6fzA1f1yqImwy0QbhfkH6vYvF2e3mzIgYJSnK
UxMejUdKSHlkRrr+x9gHv+/o0raIss45wTyugCZ9sCtKmR2nUOzYRW4wND51hDCs
TizIc7sZuc4SaWUlntFduHnbKy9boiU2HH3YW637MXAYbW0f5/2BI9efl6llibJG
G+K1/PpQNyGPryPmWLNkMbd9p9pFr3npx0eigOvf4LTLCdBgcBQxeXpo5Wq97yD8
0NUPbtiR6PenQga1AnU3xadHFr9jOfK/0q+P8mF8cEhbKYMyDuZOr6cAszcb7ueA
WQq4EGpk6v8lu3jvCaweWpI5CEpGZBmhnrfzLCHBqWWKVyPEc5/OEvr1HHffjCJp
lqMjy3OdA6ZxxGwb3h2En5WCuD3GCv0TQRc39R5UNnpKRmpdhY9RjfgdLQDsOvF2
3eMjptU+UKJ36Pmf2gMdK5CSkABN+5/Md4PURAPaLqci+BgTmGM4Fomk35Lbk3yI
90W6DdgjR4SBh3NDcQVzBCI9MErXPJcuEKVOgo+EbMzOJ8I0oO8PmISLB2E3U8L8
5kVKrnrtxW6Qf6vAvpLi6n3Tqo34N++RNU4e5DDRxo9+cjAiAHVP6zxvqQ4f0SO1
F/+sju3zfFV87wRL4xq7Jg/uKJncootw9qvW5gLnayGWopV+kEgZgP1c33okSgfu
asg6Imuv7VJ5rGVtXM21fpsCph5QnzNg3KTS+cwWz18xVEZlXXyJCM5wDJuN4pkQ
wOoWu52rLdOZLNX9pnBqmLFvgaV6FdsuhDNPtVYxX0cAMe7pnHXyQnTXQiEW2VKw
pOQ3tF9VAqPGj9oetSTFOlglH1NMtRepevAmEmUaQXPOnf6KRzZGK+C4nPH5ZMpG
cb9G6qLbtUVm2LCh08oMr5dR5Ik9ydBaHHqPVFCXT5BgxuQN7kOV1bTKLzUWMzk1
2GNTxmymBMBGueRLpjpMe2PbhZHWxKCuBtHaMN5JoD1Ve7/BdUDb2hSOHCxvpWBT
XRCXb/frDG3AhNxrlSHgwqkU5cHQM17EAAuzpxKfMdIa5yXgLQimUJOsPaD/c4Pt
AmK5jP76MlUcX/4ITL8KvKyH1TKYR00/OqoIiv1rAAQt2UDgkGmQ694rjSK+Td8O
YmZq78O/ZtTH9/Bsz3zx4mX7NV5DmCApOQNOPW0KeRrMVSq9JKSXRQxZD5bnFq/T
OAwUoxzrcs6BwfJ5iMQgUO+i6Jgs0/3LaiB16zxwSyPGRAUeU9+B9ZzUspHq4ZJq
qs+KfbTBXTI95xzgsutHKYymXphuSn+B2c5tyv9FxLcOgkffxvsfnf/QPwFeS0VS
bBrVQozLZIEnM7atZIltv6uDHTKJxS6JHbi3IlNSp4Fz9IA3Qbe82pTswivNW1Vb
Nw+VTEg4AIxTqp06eDYWbTnkm9/KlBqxyc7oVhyKQtDwncKJi557OfcSK/8Npni/
ojrJOXyhJ7DvUDbizYgWaeFXVMjXi9tJ8hDyP4UBwu/0fHyy1BnSRBd45OTo8pZE
zXjycks4c56CmHoihJ232O3PJCMktaXsbaiwdYDJaX0OMtRAY3QVNK8UxcRjm1nL
/Dn6ULTzCSZgvDguVzXb6nYmbU7Sn1oPTsq0gajHBinqYvcvIE/vAkT/23+KSD06
9wk0/aHW5+Ck9c3zJSXvK/J82UlZ9XG3yNyW3xWRZKEQD2p2H6oSj43JMmbw/w/9
kiyk2JGiADE6fHFmnsLm7K85FSDMUywTZdn+0FASUB665eKM7qubE2nG8ns2bBNn
rNOmmfZWHNqqStXVmwERMhktBaGdHp3WeCCe2vge64KEvI43aNTEJBKaZta+rvOl
fTAkcqsOHXd1c2DfwMTSp5QCnU6HeqcLglLYgQR5As4Gtm1IjwrgmCKMoxs8fLx4
NDU9NOZXi2LMklMz87V3NZj/X/BsKGMcM0nTazWAH+ZPSXn/uAcsqD2+VcAZqG/a
gdUqML4gkVdgQ0QlP5A9Hlqz9ABtw0X7w4tLP2M0wrXkAoUb9BfUsFLRLyqnEa5Z
pFKC1eVSL0mjc/nDMgdQ1u+aJ3vPwh5k1dR4nf7aLKnYgXmy2/NwYW9j8IQgrSNh
0GHZn2thd7JjnGEBlY2hjV4VOxUEjo3w5/2Vu24gZrVuhdIZeHHP5G5ia6ps4UI5
5XiVFxqvpX9IO5Bm/KFYpWE5KbMm+x2wG3EuH/76d37TfuMmX5V3Cg3M4wRjs6Sj
+JTPfCmwhsTH7VbOBQtv+kAKL1BsGsoD2LO7sjTouA7GFMrAe3MLN678v709VP9M
BgZG3FLTJT4eh2QfDJPkmPQCxgUDHi4yKC3crt4zSG+X8MVgx+lEfkzILEDlgWdw
d68TGXdO13uY6gbYEtRx0O0m+UQjTwuUzziXpBZ0B1fMLMgwGF9UoFeBFA7flDds
S2HHop3ftwHsa6+/RhDFcu3CYqsi9cOlHwnZXLf6Xerxs0TbZ+HVEekEoodAIeHN
kGkFM90ch+z4E0sj6ZKdSu6glqHb7K51Vs8h8e6nxFf7K41juhLqhSe3CzsGwLuM
JHNfCNvXBsNE1ksTsfuewcN2mpNqHT6oyg0aR7/YZGgiSzZjgrT6RnJ852NkawAL
aS4oyaKdYis2u+kjZuY/3IHHtcpkmvUiXEGDvOVvV34OPFcHk/0tXkOx6yqBTQj0
k3hUMVhuepN+sJeeG8hR/iIf/hC4DB2APNlCAbiP4A929s/UUoeFwRqQOIHiej4r
iA4ZZoti2T8wXbLB37xqc/vvU/48tAWcMI3J/PUTx4kJxkeG/Rq43eurd7x8m29U
kqVe5gmEApI9qxMTV2guTtmbs2DDGKG4vh9UlkWdjtIIHtbtbdgPDOuaMdHuqMWQ
ME/0Hy5hlrFiQ2+jD6Un8PyOtrty+mhky6U3kKzINxj4ytioDHr+6CRuQ9CdV3U+
3Qzp2JfaGUzm+h6tzGcSpQulczUtOrP2zrjiL+CEZyFfvIuiFPlaWUD8++5nDFdP
A0SPVmDH9VxbpjG4Iv96l3QDkYXEJ0f37J/O688GuxO+YLxthJhsHjZhIgi2EzJu
4E+4/+yCOuRqGcqzzDA5gCPqUzd3HSBRfNaKFw5m30Z3GffLQ+Sy95V/94aYQRad
w6IwytTj/+lP+pig/F+ot8w3IFDon7W/kC4ALUM7zY4gqg38pbsTrKRpikLWQYRn
G6QAuRdswv/slq+xxNgZ30Zg1dwChn8Sjt9M9ZccSSZm+UJNnZx6lskBUEiIltoh
xH9gAIWCN4K5QvAWB/uQzJBi7+VpThHnePzcfsLKRxKJnQFhrRQrN8eCZirkyBeR
nbxO+ljrtDIyFEvmhkJs5aq7hmCCqKk33Aze+kbr4OUn0YZpBFuWUAHT7z8MVQL0
SOzhX5yychsVfFEyAI6VErJ07YuFKYn9IiN4Vv/51tNvrZrUWuTTIXD18pRCBuKQ
RWbLA3NmGh15VQHTRN+Qfor8Jza2DI+qRqjJqs/uP6LdT60rmQyyHNrpvueLNscE
KRANUgtzPgFs+ChZMe5L3elfkD2yix8+YwK9IS4dUQKUld1bvW4n5t3lDNkO/tNL
MyD7DwU5I8zm8H4V2u2kWCSqNXHgYbSooPGemkhANX1SWVL76Hxc2hAtr6ieOinD
V/Aw3XepsrL0btw+tHBls+xH0LABxeyTb/nWbnO29zq90YcI34y24QPNuUxK/f3c
L88H3BiF9QMzrLNmmacyz1BNqCmQEXu6ojCTnZYqyxE/WZsSUa3jeAfMnLlRwey5
1Q4iEUE0/ubV6BFdFbvY4giJMSAfTi/Qo0ZeTnyXvVd2eJRTyTSrDjtPxpfxhUwA
82EX330Iz7V4QQH0HJsLL+MQN4vXnbFtIBMN0nXljf0oaW/ZrJEapT0cC8rSIFgj
2r8V1iWQ1C1nQjOus/FZ+Yl7fVA5Ne86HadMi56KIdCgYILTBdBCIFUq3+I/ajP5
9/4zDGgu6wE1U5fqdR5sppWbMxC165V01oW+rfwWw3ww9dzp9OclvpK8GJZg8xD7
TNzNVxJ5erQd2C8QoieOU9lJ2RLMTlDhZ5xz9wyFT2hdIIwflMnzdWCAS2KwHkMo
pTlYxyAiiNWDchKYtZJVr9/ho5+QA6Z80cQFVLkqu1CO2rYRoltsDG3eAJ2pJweS
WYVMAhuGhTsTs8BOa0p47P7gQahvXvcXz0jGCjhx+kZcQx9/BlNvPUjddCPwIKhj
VpyjCbexf6dtvC4X4Atyp8GViR6o7aAfYnGQRaGSL/lBCm10qW1KA4i23fEeDfdH
DN5CBvwth/OdB34zj5TY8uLW64Y2BVE7ZYcmLWL/a4ODSyhuI33Crzxr3L0kLjHN
sKDf+s53aTS1Kg23odiHqZuLyl9KRMpO8SjF0xMRIzVNyou7p9zD7fU8qIStb8hG
/isVmO4OrDyeMTE5FXwWKiXfdxepCG8aHWtY9Wf9cqPMDDKKG5VYqAN3rCcQbY1I
pyUFptBwIvpBFpAaWa/poTW9gpsYb2PNGE3PCKtTObey8tICW0VjTYEe8f9VQUKo
DKSof6EUo4D596UQ0hM+v7hmugAw1mZUnQ2XUKTBzrbDmabFZ5FkhclSSrKWr4k0
ZWbmcU6PbeGNoTW9Dq0mZ6fofq/CWucgRMsOi+qVCs3eC6K7/aKQVjKJbW2YA9Wu
G+8CPB/Pg5Dsvl7Sklp4oGQwJdaonU27Fksj/Gdt2LUg2XzglUls0p+svvuneh+1
N/2xdNOwpxZhR2E2Ll9ZnA/6Ro9tJ0NwePYoSOH3ltYsvz6AUBXqZoDcRmpFvjj2
9ZjjUD9mbeGDkW7T3K4UIl5UiLnD1XZvHuqQsmvGCVxZtgD0yTZF3CyXJTyU+yOz
2o+nwjM3dpPzC1SVqPGhM/WoOjCMXjQUaierf7yeAOnF0fF8qwRIowFWq77WLR7x
fgjc/yi4gUvOboOsNneODlnXiG7ARrNDR/W5ztFEOikvmCMyb5Nph/WtP2YibeKf
MDPAi+EP8K1f9qzExxRiVe+wohT9Mo76unMfYEkt6EpmuvjCxl5HwkAMOdAwUgaR
0EGFRXgGLjoPqaml8gK3JW6Mz69e9Q68LfCmS59grRvxMzEOR5wTUQsVltIfZMBj
JHfZEqBEAhgFM3y7Rjxmv0h9/WhE0+Rn9JaURYBJdbTKdd+IhLyZqvFgszV4rhKS
GG0h8yEYbOrC4NuqiImWKl+kDwaKfhGSw23isMTd2EjYA7sRyk8OmUA9/pvRfRn5
/RTpLYjYPGyQm+oUdLVEsKjYAtDpqXaTZAMHv3XQGziNAm/ANJzBAyLoeo+T4H0/
6AjlRBZMnza7VQ1Jc7KvMe1BUFY3vI4XIAAqUhOU2XbLEhPlFX7l/VUuhPEEFSH+
hhUIcv3MpnnWEduDs0I2ekL2iyPqoCSpSiCdYfpr0/Mfcrl9raNdy/sr938jRBzi
00QNEDoRd/WFrx1SRIP1B21NWW044s2Cl7bNk5BbWz6V69NdyPoHX7RYJE4n184x
Uv6uo6KAHh5RrWAADY6+rNDAEsdZAu7T4rK8ZwchKSImtOqW2TwKkqgJonKcC/Ul
E4byE0JSUtgYwCCB5R3+eb2FbOmhxPbD5Qk+A5Hh6T5QSzEK0Pe9niMb10kvNO8b
TIq/I5490eIKwsBg5Bx0fUYTnDpxnVhJlEEN9Br+irhBtJK8RcJ6iVvF/lNNpRnS
fOCE9BAZ8TtTOmCYD8u9WlU1TvWnP2fnl74t5a/2bvaGrACLDkk6yGAX3rOZCO3e
JSB2sLAjFlObHl3dkUt1tfUoeLGj/HFKzb4f9PMEyxKgOSI7gSF0GgR5YqhjehMf
wuh5ckhPcffmUmXkT9vn7nHoF1+M7njRH6sVdPOamY3r4ONqBrErWZ3GD4ndR3xk
LX9sPq3zQie78kO2ap1gVi3b3mbDnCIpzpA54wyZtiFz6FmB16hjv4jG+HgEv1aA
pbiax5wjkhos5YOzzwQNvFtPNUmMcANv6Q5pAsuvpFGxSw1cTd0iEfF+T1z1lcbj
gdAccj8w503QAqpKxTyha/3ivipkZj0AmR823tGjn0GTV7BYK86/xYQCtWKJCDE/
ogEY7mgbc2V/jq0Y1iOl22iv7GTz5Lmnty3L7r0FyzT/srYlJUUy0lHY9lkFSiAd
Z9+hY5i1XWUKpaekBKcdENpUDt3TX+1K8pGE9PdxuZSr+Dj3xrIiOLrtvcwatFD8
6U/7BaKUOzZZW3dv6Q/YRQDuoAmw+p8tZvuUD4qS1lBl94Z+pb2yf7KIHPUd3SlA
BSceYnfuruRb65iR6rBNo6HujWLyb0/ZitWrIaUIgnBTOu9ujGa4yXsqH4WOhz7Y
/cayz8PhR7y4SaD7kE6zG91QQWRh/VyvfKGu5fgWR2RfCYqN1HA5RuHA9E2qCO5s
4bjXWr6sARdNieS6XBr9NKZhzpk2+y4eoY7QPFEcolaHv6My2gtYZeQdWgXJmog9
vkgv/AjlwoO61dmnONdcZSBsJGwd8vx8X8AoaRdjupDDtAzP1N/VAYcJrI6pqQHx
s70l0wB8jltz+J1nDH4aQBAsBMYQeuAHrHuncm6HDKoV+Zn9CPIrcuw3bMn7ZFjG
HyHqUCmK5zujb0Ay7ovmdRFlMAwfUHDMmZauO+torkLpkg7AQZejBYsAPR2lFKaM
XbQ67BqecUxdvB9G4azK4pxcfJj0veubZNucuctngEISd6gzpB2mI6jSP3YlRDza
Qdla4EdvCa9xFkh/85XD8srUeqUw3IZXLkRYnyqAsrxg1kfQz3FpLbfQRly8iTUg
cIHcqIToRF9chcnY6En4N4CzKZBBI6cd7Q0ONdZGccVLF+E+NHX88GRI57P0aU9t
O4UOp2S/oyUfoB+kOfkyN7P5J3k1hnDQrt4BfAFLiX3yv20K52loyn4tFczm9ElG
UFdwuAqBIssK64iiHTI5Bmm3wEkE62sHUkJd/8X3LFLFXfEWqZC9D4AcTKT+WBMm
NgxJmfWeIxj/ae9aHHF9kMQQFJlMHOYv6Yp1bZXa0Ds2GZ+07CbsdJGYt2mQmOo6
D7XdMH+y7iDL1OkCIasCjjJa0E7gLMTQsGYm7lOOQhg1x1B5fvkrMdbaXr0yG1vU
NBnpW+8xRpKXu4zcAY0gO9k1jJH4DMFmIcPx3mr+MGrNfg+UkLqjM7y31zdaVLo9
Zlp4Tws8jtXXLtZ4uPenOTms1cSi25GZUDVhOB0Ow0wsEfS6P3oMhuddG6A+FaZx
nLPDQkrfQUeCKpIRbTJV6KXxA7+7G46VRaVkA5WcimvIFqXAXfWCFTUQlq7m9P1o
SWUhHTvr1R/E5gKe2vlw9eyQIz/ZpbGcFbviZADVYsF26h6gIwju69Vt9cj1IWMq
d48mlbfIOy7nkBcruG9XV7E21X+Cjr9pG+85NJVq5xe02nB+whzoYH5YHzvSIoTf
PF5SuIjg0vMtviT2DeKxK/grw5Wzb1NGM2izsuctFn8pE9IHXhjrm+FKIYTIcINe
5GrsaN3IV+Ic5Gd/mAMmVPCtqL5b++8sn9QPpoSk16M6vjZyhIw7sQA/Px+szhh1
27tpZiXbOy4zJoxuBgqgJmxECjrBqZE6x1s8sbpLn10flqOtckCp6q2pTuuXI7p6
JgtsCUhgzLG+mvXUOYZ1ho04+2ylI+nmFyy+xnYHL5IkKouYu8Ieg4+3KApMgoBa
yfMvkwxukTX6tiJviRFVTd6+PYM9I+nOT/mscTQRjQ5psWQdatKmug2j2JTs5bXQ
lGIqnZWYHAgbNKsy5x/3TbmyR3cht4skGSFJybh2P6371glt7M800UgiS886Es0W
a2Q+1OGzJdw9MTSWvZ1+NJKmKdlrd3oCdyrEQJ5kLB38v0tE/7KpvuHBZFPkSy4t
hgVEcGvFiEN/Hu98HvHUm5HrYIXdDD8SExoORTwNeUXWCwL37c5WxL+1aUyC69B7
IHV4Bx4fb2Q/vRCk6sHtzbdgf2C1nrEsJhcRohkWSK1+3dYO02qbKxPO39aVkgdX
2eSNTV1dMCvnSqZK9oLTbLsy7xVV+iVm5nZNmKDjCQyfsI/fOivVYpMyiiCMyUxr
OwK/sFiLEpZYea6LlZWg9ff4ng9DA0w66odatvMqoY7+FoOOczi0sjz3ZzDHyftx
Q6YteqAWgJ9prG13Mi5n11z8xsT+iE6EEOyE53PiZ1lCRIYlu9T59iG2n5YFvn1j
BzMIwjP+URC5GpYft88r7dMhIEJ7XHUpnlMf8AKq3J2Oh5loRBUoVH1Dss1PMsU0
FpG3OBT+LSROWMMuo/yRfRV/VKE0ImpIrRogoQhAFzu9fu0ugV9BmLaisQltdqXB
OqDIaXKKrVtb5+8Q7YcLJDx0OwYsOmckWO5YFQcDOyeY57AS3RZD0uRfJ4jaZgsy
/KsmABTkaDGfQ8RlExqcFlAk02NG5tCbFU83z/01t/C76IRinexVQ36zc3otJAep
HnGoaEC4tKNAQAb0iPV8kqa2sh+I8LkT6EAyShpWxiXzu+4hsHQpIhJZ6XQS7BqK
i+beGl3BvpI0ozLO85VqXp4+QPBzhXZFOm4KWaD+jNcJ8wcQNbYVX1hoWEVtop3Z
BJmaqx2RcbQc2NsxCs8GVpIvkzfA9fkjJdzxQUnWgtAzXs+n4Psi/RhI18+kCNWf
/fReH3nAOIgZZF0vNOSvG/4HCgd+A00QTqNrjQ3bsUN8EbG+qsX2T2nN1PsvMfVM
wNn33oBLEmSxzTmbIuJkIuOC3mGWyiUz104+NaULkgY=
`protect end_protected