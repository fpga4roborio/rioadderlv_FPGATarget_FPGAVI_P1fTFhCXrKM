`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
ddtXksX2+yylW5zu6QL2Lhnb2d1sD00763mmSITNX595NcHTEkwn0zB1Dry37fOW
FufOhVzEJp80NC5qZ/+F0Vk7Ik02dIR0elf3clrjeJRK85K4e3Hoo4xn7YbFUIms
l/8VZSb14+JVGURjfswrIyCUotIzlzVYZ6gzoZwDXIi5gQIBf/gI+KxNXPaKV+PQ
Ufys/12rjO6aI/pPlqSm0hCvftmBcnezN2hk1UeXgOIuKZnogjOsf0iJVX2aOOWE
6pD/psybjbnsNB6kH5uFTA5frkzIzkzl5d9+YDm9OyC+k84E83I/7/j+rk4L2dah
QJOvksSIzN867/4Qt8qYTQ==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="MvBXkzurAa5VTw+1JJ70nePUfoQXBvZOku/SMmg4TwQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
oRtzZL4VJ4iwysPsC8SXYCzXS8Fw2gtZTOskLcDV+1B9Nzn1zTyNtlo6lNICRmmK
ZRVu2BmCc2G+fmzynYlNTnSa7C0Cuel6FYpxCBlOuk3OF2tzAmLAuDyOH3Z1Yjzk
a0aHuoCdIRKv7BrZCdALt03JeUmXKPdOmIlkVGFl8yw=
`protect rights_digest_method = "sha256"
`protect end_toolblock="Jn9CQpRhJt4rnzZPRk+dOpzAubz7omckX1MrFd4p81o="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 5408 )
`protect data_block
gD6l00tciPUa6pDNTk/+t0OO0nC/UTtBwLB41d4inuAUA3i/ALrNyoJVcBnAmEQW
ptbcNp5fxEUJjnOxnedyZEuEBxWRieZFQnkRdF269oObfnLK4wyrdgiGqQi5kG/p
xZtbOk6GQBlohRtNxGj+lQApCBTGUBtPF2xKh7bt38afR9xi1c2Mc4UAWwmDwdL9
Tfe+FbXxRB0hzZ+heXx78Gfd7DhM1oYP7/ff5gYc8soqdYM+wJTMF+GclKUtVdmj
SsLvbPfChjPAVmhG2rR5kd5I7L2rGW2IjpHjQJJQZFqUGsKDaqH/6Ty7xF3RnxeN
WtkVJ5tJJAsgG4UBUBm4jA09eaaEwy7HiEQ1JIyvICcimBoap8S32QBJ1STt2IDb
fCQ9kgGLISDxkZkDd1M7KXA3HD7Zo85ezv/eJLMdqBVOgaMRhNIx3wQz+rJeP6V4
VzzYJpeW8j1Mu+WK5gS6MKGnu3RCxbdY6O9iOyymmJ0sOuvvA/Et8u3rmF5Dlu7y
2ooW0aKu4dFIp1BezaOpqpY2XYT5jmWqlSL08EC9cpV8t6cJgOKgwziVl+roosxT
n6cE0gJMhrFuIHDqhptjMGaerLcTRSgqiDEA9fQUtr60QEEgERGNr6jjr+Ye3cev
Q50k5ukXAS1I96PE4Lr0YNgdy8avWkRH0X7Cir5UB1K7X9Pa/Mlw5n9ZKsm+Ityn
+iUXdtDBdiRm2oIdJXpDncgsU2i8Ak9RHtVD0KKpFVPCrWFzQjqat1aHSj3Lv+da
rF6unyfVDkdhEVNAuIeWbFNE9HslCY1M0KPap50vWUFZvm/cucJfJiNJyOUEhabZ
0oJGj0D3ofuO5VOtbbQK6ImIY3muh2Cb+CkfPHIyo7O2ph55p53yaWFqBzyRppjr
HeW+nNK19ROx+yd0RxJsvCP+/IWR34zZ3HXRRGr5T8RUYCpbEI77hwBihCqcLais
J4/XA8n+b7uzVBYybJ/FIUq7fQIvPiPerJ6AlHdcBKmCF3pByN355vn4dZ8wcTw+
vZ6uyi9By0kSVxsIca2HiC7+dGpcC6iSShGPjfYekYo8b8wKqMXraV0fZ4Mx8sdj
pmcqeGFS8akopDA5l4FMg6ovVYJlWYMpLL4jckfZQeean4dOrMu40Yl96s/8jQOY
CHQVXOq/JbifN3dWm5t2ZmviZDLvN5rZ/wwJ3BnDn0MBf3Yjou5u4j1CPK8CEo/Y
7mir8fGwcH3zgvXKLxieR6otLGEH9ZCRjwnqFNb5AIIci8uMu/ywRDwA3Wji/JLC
BzDeGr0/iv6+RlVyp2n+tsT8QzNCuIhcxieFpBhpF1/lFF0m01sNXoiuUmEEUnch
CLAFXqn16VwcoS5dJkjNtUuHtWiIzwurVM2Mpx2/HV4bgV+aDnmpN9JZN4jrtNa5
8qiObDi/lp8hFvlPKsqzqByJBAbOj2LMqHgvqeSXSq0GUDTCzdPoHUDIAEW+2joh
MtfdqIwAP7VuZJpkph0wyUAkqUZUBOrLmBNWUQtkpnbrZc2hAc3f70z4EIeNpfz6
xKZHGlFGR4AWUr/2/mJSdFvcuwHtQzcTT5OSITQhvrq4LlKesB0YQIu/O0qRNBWc
y7oY4nizmxaX37uOG92pJOi7g/CR0ipyK84Iv0SrOn09zQOo3YAxOPuWEeJptowZ
5iHcpNyi4eug8tMh47afgmwQAu6IvtWWxE6cOkDQ5xWLHPdafl/Ys4Qqzy2B74fA
iBrr4CG5rR8YRAgalBy5wTw2iURsqD4UlLFk+t369URKF2DhQDi04uLYzNndb4ae
403g8IWob/hvbbvrmMOwzu9HX1F8Ivn26MBl2Hk5bnEvsKC1jSMIIxw3qD6AKiBO
mWaLTxJQZ1MfmzhHOrQStM1zZNEW0j5upUNF9TXcsTrOUnaSkxBlK3c21R/5loew
bBKk88Y+NF/nDq1Kkg9fDxSNSUTjEVd/WEfJSGZZsd7B+luC2Du08tFmE0EIuIZG
sDxCV3IyfxQ8UAS0IjC/XZblELVeEGtPTSh1sbRYHIy7yaiC2EGLuk4E9nMchjkr
K64LftuSgl2PrtK9vw2xFXfdEvccjvNxHdricoIarsh9/nQDEGqGAT+gpI57S9fl
PY7+u+Bb58U5ib5wArKF4k5Ya7aywEali+hqfq8Mfwhkdg33RuWL5S4T8B9Z5KXG
gzhCFQHEbce1LsnujQZANgjGm/rwZPHZeQvh+BvE2PIjOpR6sxmBNBxPbDzuT54H
uucUUWgI9ogM2hoZ2TkwaX+N1e+Jma3Pv9p2sHvjNbP1O60QepzdmBX+KR9o00+4
i2CpAWcQSy7Bqgec0hVxfaaSCgI9AmjBfNCDT0IiMMMEPTb/+ZkXrk+Z1v1H5/B8
45FJHkItTOJTiA/q3fKhy57MqOSHpk2tBAQGLEQiclt9yuFZmsG8xbcJ6Ta13+AM
OhzWFFbs2a2BBjFI1y6r3rkJSKL3cAgaVDmQSVo57aWh+RUMrj9r5WIDzEYowQCP
YejjAdxruH70g6bS7PhNiyoVoIzeMzg1yBMAqaXWkCEyyrSXXqi2vwm50vIVtcoJ
lGoQx+u1m1XrddJ7Bkdv3EGJkWJ59KcNCMUmil4HqUz6TbDWk+mqJk8ugxsjvctk
VK9n8Cl50sbl4kYg6obztzS6azbsTalNJ3iI8ta5p21CtZPaMbft0fYi+7sZKGYL
MS2mRcwC7xIrTmn5ix3bqbVEHI4ENiJF2bJyBI2Vui3YIOdBijLviMVVT0f6lLu5
3NpuAYVN00eTK//tAwT9cy/oyT0gNe+85PUvIq2ql3LCQlXFBQsObrC17p2FjCG4
MKc45VvlXTBl+PONhxcqnj+OysLubdoVUMV3qo1mDm1Z4OHvtkVjnJXgJgbT10IH
WWOqkAMvLycHszt4wCsCiaKql/35xJkHKLh6JUlc+FuTWl/a5+Hf6ymIRGsb/beX
GrqkmGprbcb5ghksJnsTPU4pvj+4nDGSOJLiG/c+J3Oqst/TyM6RfffOPdn1V6xh
myh5rDhX8J1pChMUByAdjVS3mRulaqygyC5UtnPIjFnkKTSWNwihHXHEBsVxB+iU
etI/1cHXwfHrGgTFOxeEE8CASNhdSWxn1HmJ9kPilzyaIbDXb+EKCk64sldIJQds
rRa30d5K2DsCUu3jOqA7y2EawovJ6DGx/R+f0SS0VXwadokAlRVCN8kkUQIjX7VB
ImpogXM2K4NBMKxIgAqp4xACvwORSIuQfRUZ4oDl0lh3X6iPKq716sfOrhKzcE+X
o3JmNu29diOQeHy0tslcXjWaPjOIWHxjmadNh5rshjgRMsDSsSvT7OToHy4c8+lv
im3Ig8ctGGiwhHr9Bpq+9kJqljsnSlllTxSErmwil6n6bLR+iaVYXwfJjL+dJThz
O3SjF4dZMZBhcFsxyXgZoqJY8bFx0Ldzcdi1muX4gGBxapNkupEMnm6TUSTB+omd
DGha88C6jw3Ilu3wIjI/DnjVT6uQxF1kwn4Sj7tXS5uKQxz0ScIL3P2gwO4rjfvr
oywU4UKD6OV1zLjXAynAWY0schP0yRBo3uBY6Qj93rWDrUPgCjKTUbxUAXYiOVzN
S7EmjRkvWHbhTWWTjm/tJqj8sbIq9luPmwuDlx5GsxsoIZN4Evd7gYbm0uktaI8b
zimiOKtDXmlxzL94S/TW5cbJ35LHHD44l+1PP7HOHNQwGxJjlHecCXXs2zMoy9SC
eJnTHPVJzkEvCbc4VhudiuZimCsdCwf76zlV+ZM2jXUU06DxomkB9NBa7tsNR1X/
JaSY1ux0YuDqW/Y8E2EPYqZ4a6wpG8JJdzLid+nG3iwaQtyVVU0enUDwMz9MoSlb
zUAa5xih8Zsjr2yQ2zFvwMN2BFGt1h6MRc4ytZUZm+gCC4QgAAkyJqt2wuMaccNd
M1Ce/wNTwx7DWSlbKhQCwr/iUvSD1exrlis1XdgpSvpcTZ12RP/GeMOmWHWmYpKk
IVkv/rrcXi3HOhjMvSTyE2t1zMMBJPc3rSZfFhI1PdMiuhTgkSeu4M/Wzjq1Dv7K
6AI3bnjdV1Qk9AqbbkbgIOmRN7gCbCuSd2kpYrfFSK9BRJ6SslkFvJL8U85jbmpE
gZC8QIW92vB45iEyDLktbkcIPLHvtlj//3bwZeBhFdqSjK5gXYMa8YFJRuDShZU+
KoBKg/3pLkPUr53/m8577mgpgXrXAMtyJOMs8SrXbntfis/whX9weppfXkKqh8j1
2bFh1ml/vc8LrtJyNcNjxtz9m/MYa/422GRMDCzXHXmoIxC4yNxDogBAicaD0iBL
JhM0Vllsyzeiw14ETFFuVyxCmZCEWJ5MgX3N43nd6xdLtDcRATYrbfDHUOseP538
W/CnpJKISfrwmQgSnOrBT/MQ9tAaP7y+WcClGv/TKRZ2dASGZUtvg5rutIKz7mW0
BjLkxQW3XqvBWTATXcfzbMR9zRfvyrwuA0sDr35gGpd0w4ugJw+bGiDrC5JyxLvg
gIs4lr4cQuBMuhiMkmMM+YBehbhjTHq48Fkl6VWwyoD3eFluN/o9l4pGAliKlljP
2PabvOj3HoOVW7wAdzHq/GHNEp6FIiNCO1qqE8JHqmyj30rzU7lG9NfT+dNaNB79
ySujP+KMVIFCgdkU2Ep3isfZDYtPQGAWY1jL5jCEl+YSOFBKvQdVZWn+n81hv1OU
nQLTxowZ5ig9/rZLLTf82D9mPgdCAztAqyA+bUC57955YesxlQaIcnmhk7fFI8FQ
zsoiGLjvr/et5C0uCE1rKaR782aN/mHmASXToEq2GWFkBXzRBzVbrf2YOcF3IwTO
PDS6YKCezaOoXjYmBqVPUg+/ZN8FaFI7wrzqwTAjZI7LWSW3nWzmh1kOY/NSiRG5
UDJEQkuL/npQDpu1AqzMC5ITI0My/PgwWEyYoVzyjAIImrHXsGEXkbd1MKTffwkj
qWqPuMJ8KjNVzfxcuXBpV2nnpkqX/By2u6/Ne+Z3Qa9M78v1V4yF1nL9PM6kCEGR
UuIXQ8yl5D48r5Ff4F17TiFcCDpM1gbyu5wq2n4fhZGAWqZWfWwmCfZc2S6h4WoS
qFqvmLfV3MDGZxseGiO7xEzgjWDfLh+SFu3jXJjo6yTlyv0JRPGfpaNJgi+zGiUL
UMLbMlJkmeAmr4PdyqiiaKnwGJJy359GbalsLiyE2GdaWAYAQnc4DH9oj8KoLBDR
NCJHqTr2A/BPh+hPszsZ9bv9JU7pmTvMSjCWRK1K27NTjlgT3IaPJi73iZDLzh2t
SfBXcfj8X86vBNBwDDryNUJB2HQywmFVeyVaoTnkQdPnKgujSFxiHu5RTGMmTAh9
7XZ8eRwoKbbX4Z3FxzNSnwL72qH3PDQ1Ioinn0t2DDOVjHLVByMU2WTrks1P9JS3
kYnhPZtj5mzOG/4xqQvWtpjljAT9h2sg3LDEoCd/rf+/ANWXO9VucNdTWJVABgXp
YfhZK7IUD0GDyq3Y6j74pHQp1q48pAUe2KkBCFoC8O37Qtmp2BSXNW3L2Z6niwIi
6PQ8Y6suDeoTsTw5ezVEWsp3qhfkfwvX/MAcFiB5s8usNtsJor7vQ2SeKx86yGWi
14wEWKBM+50Q891eNRZMTaPYA4pdbdb13kh8fFdOdWqXDL5lIqIb25b7VAYOha3h
f1TBjsuzY6sqlMa7asG2NefGRjyn9DXpZOQ+bFNqz53AKRwmOY6vW72qh7pWK5J5
7cd9+uklSPQka6mM7QAhY2h84iUfkPat//cUCdgMeC5fmRNu5ocnuPYzgucOIq0Q
dFZyZwlAujMqyP9SsAZfxVlNygwpu8ygyFgsbBrz/ca/xDrYziCR4dcSq2ZWeczD
uU7M1lllFADKFSuANgd8XA5FM8mJ2k57xwO/vftmwf25LwJcKqRTUzUksqdYhkLv
JYIb6ppauLTmcgIssih+FF2x2VaVUA6JQyQO32hqDFC1RNWhjPDwrAdpkjhrzevB
dYczWqnC/fvlnxD0ol+ZKawAJaXDt77MSNZM37GWcy/7rA1NOPG/h9pUKcZ1boCk
vBvM/bvvp45T07xetICZkj4wm0ZJFa885rKRTXlgWWao3/gzwp7r8vLB+/+KpU2S
yFufKirGZtQ7b/TqdoRZzUQXyYxhhxdMz5TFkHCMRkvzw+rE7w0eLY+3IyY/H6Qy
JR0+Qm5sxSxLfyCfjE53W/NYWbpHbR7fQ3COa/+7EBiHwKeQgR1NalZDVzKpossp
xnC7JY99lBl+/dDgusi3HpVbvawKHpukUTYolDXzT5+pusWHwKtDbcI3YTspfPp/
/RpuAC+qUjTR62vq+mj5mW/MwSUojxYeaEK+YcHAAGgtu1U44ZmuV+DTdg0CZXKx
6DuyItc4+Q3L5N2F1Fb437oKFB2OXfe1zud/aCF4O/bCLt3+MbuDh8aPdjI3PDON
DKdjiHUHOWFVApkrlA4u8YGFk6MjjERaMkghvGLBH1RvDFBqtRkxKQYlaFMSNKA3
MSZAelZAMxqXk+F+SxkADjbtUPBB3Yy6RA3gJI8IJYa5/NrU1FFVIEM9jqjbDyLG
QbV6hsoVMCbPEeIEx48C0KP1ijPNYNQ1kHvTwRE+BLIjZ/AJWW4Ore8xvhzn17kG
kzBGNnMT4kp+6mnv6fuG+YR1K1j651uHiwYX+4Z9QnapPEnk3BMyrOtGi0Fcw7FN
Tk38OI70upUaJSSy1meTSmgLBEKNXwVOjyCtPgKK5h44C8edcfRXls0YObgQMsRy
VD0Y8H8q5rifkOTu93yAxN3GZ+eHf1Mvp+70svibB6TSo+ivRuFruwx/YNS/tuIf
zvEZR/VQCL0M4f6+yhtuCVkJLFHbkDvHN/inGcVqoWlyltb2AX7iAdg10HCnm4s1
IXAT/HOqfjhVbDLmuM6ALEeDcPnNA/E3X2Phx686nYnXAgVuf3Z+HJE+NEkAXxRM
oHxOReIJnq7xEjx2qm1G+0B5SKF+g+s0vqJOIk6K0AAqmB2JDypf2U1EuBkP4eG9
YDhLWpe6HfbkWfMngj1DtXKzkE83XchrukQhFxlkpvp2qkJsxkabdSHTnFRavZ9I
R2spBmDKkZPugm0LpffqOzh3s6vW+/T32yE+izgLa4u+h3SW3dlJ17YN7s15Epcr
+k6f2tT5k9swsfi4JkIq9OWkCOU1TMMee/OV5lJogSmvqk7ps+D4usWaU1w+niin
Eb4HxsRypLcIQFN2lA6zYA+S9fvUW8g0p3YMc6LreGA=
`protect end_protected