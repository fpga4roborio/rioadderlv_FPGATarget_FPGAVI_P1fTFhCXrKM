`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
ddtXksX2+yylW5zu6QL2Lhnb2d1sD00763mmSITNX595NcHTEkwn0zB1Dry37fOW
FufOhVzEJp80NC5qZ/+F0Vk7Ik02dIR0elf3clrjeJRK85K4e3Hoo4xn7YbFUIms
l/8VZSb14+JVGURjfswrIyCUotIzlzVYZ6gzoZwDXIi5gQIBf/gI+KxNXPaKV+PQ
Ufys/12rjO6aI/pPlqSm0hCvftmBcnezN2hk1UeXgOIuKZnogjOsf0iJVX2aOOWE
6pD/psybjbnsNB6kH5uFTA5frkzIzkzl5d9+YDm9OyC+k84E83I/7/j+rk4L2dah
QJOvksSIzN867/4Qt8qYTQ==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="MvBXkzurAa5VTw+1JJ70nePUfoQXBvZOku/SMmg4TwQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
oRtzZL4VJ4iwysPsC8SXYCzXS8Fw2gtZTOskLcDV+1B9Nzn1zTyNtlo6lNICRmmK
ZRVu2BmCc2G+fmzynYlNTnSa7C0Cuel6FYpxCBlOuk3OF2tzAmLAuDyOH3Z1Yjzk
a0aHuoCdIRKv7BrZCdALt03JeUmXKPdOmIlkVGFl8yw=
`protect rights_digest_method = "sha256"
`protect end_toolblock="Jn9CQpRhJt4rnzZPRk+dOpzAubz7omckX1MrFd4p81o="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 3488 )
`protect data_block
gD6l00tciPUa6pDNTk/+t0OO0nC/UTtBwLB41d4inuAUA3i/ALrNyoJVcBnAmEQW
ptbcNp5fxEUJjnOxnedyZEuEBxWRieZFQnkRdF269oOfwVvfNFWKZx38b0V+Uxog
4dOf6PUeE9gsUxBzRc7tLuhEdqZvB/U6iXlNqZl3P3Dn4kWPmJST4q6tAk9gP4dj
TJ2gNws/0AdDrhR3xE9lnZ/H03uhorAj7oe3GxGUlVdpcXq+AHt3whorxokS+xAo
sMZQk2ZzXCrbzCex/e7jV+GHouLcIuXqSVRXEfNmszCbyn/w7XzPOL/+R4VrlIsj
VfpysEvTTzqdz1jb7eYrRAtWF8pTLMdAJ42p+egQFcUf7/S4tIzVSYaJPAsRzbTW
ssk+dO5SBFUUVAuBgWdmuOYXQJUi6hhKI4lgMPdmvKpfYn74UQkxCTL6p7J8jDMT
U/5WrYTl72SqQ2ZlresBWf8ckGf3lP18t+i4oeE3sDk4LZumlc3BAL7IZDuc9esZ
5vWxX1HbkUTQsL5Sosg2JNwqpiQGMgnZPhwzwRJGaZt7EdgQuG8QNznoZpSIPPPp
KluVaaFHHAC6/GcPebw5mqS9A9gZXBZQDuBXMMqfWESFWl8tld1Z1PTfkdHq/GWF
aeuQkKRd+bIS318I0f6OpSlz9kc9AcT6Kw3Kq0EiTshXTDfQB8bplbVfg5zXynLu
UBsXmaIqn1s8xHWzCUVHuTZdXVD/Enmi2PKOvlY5oGJP6V+4kGfDwpIfjfcWtYDu
Db9kQdYokMv++LGGCPT2LBzq83qSjTaZCZeFXd7WLP/vVQ3nVctvZ1jzTJoW4Pzi
sCV9jGACgRD0qKHIweXm0G+h66sBdseyozAamRWp/M3GmLGdCUGYQsUSPRayUL5f
a2exSxJYgInDMk94ETACuyg+S/OT2uwyNCJgEHy0YoAsM817IVqXUGqAOf5tqffc
dSr7KNxukGiR42VrCFIZOrWQ7qFswmKeUL1M/NRQzw4HN4iPWE1KdjL6iHDkLxRm
fb+9HayqxO7Mo83RDtmZSfDZ2Y4FXPo58OwSa0/69RQTNraktwiZmZaBq4RxpfnK
xT1aQfkt4YLDqANfWSfjMXtlEThe5p1lsBQ5tNwraSjz7664rgqzZw0pTBFx6gj3
dRjFbkf2+SDkHFRk4XjlLtP92wQ470Y4npraBoiFRIkrLAVneZmLzJ+QkKU5ZqnV
n+U5s/VAMCRV8VUIoVSIbjN9DY6dPY1ehx2hfMfvy7VjmqaWRqvnYg0zJUNTAwZH
euaLRVKM3DpKmZF9SIu5OU9NkaP3lQlt9QlRMQyFdz+x1Y1Jg3DVxOJyI4qAkGXy
fiSU2OOzmBGYhyt9c7QwcdB7M8Tp16o/rBthYotDKGc3dS54sD7MMurAFva/6sGD
khiVPWHpoa5suhjuuZbsmP5vExB7aj6kZO3DXDLS84TlDR4PWkk1ahQv0ZmlK6jI
KYuG/jx6fq5C9pJN2uQ0vvJvuatax4OrVkxGZtIiE5WEv9Ee4Nx6olkPIQSxT5vg
749tATBT386TnFwkDHXhK9hnI9ww9Vd/M5NUNPkz0u3grAnw0o+rWwak0rnYlsy4
ytRQJ4LzKvGQZ5xl+WKoqHA04NGG4uf5BwoVbT7iKfNoczjoduQPMECqao/raE4Y
RFfuR8+7G9WsuFF09RVQ1NcwRH+3S0hu0ZCo2i4GuQRIMCpbQzJP8FmQgOFcz1x4
hPY/8WS5kfwoWFxsv2Y9MKjiO11Qe4EXrE9sTgF+pJ2YQb6TYCT8sMwmRH2QInQ8
KQG5hjs0LnCXewTbT3sWxQkw1ebPUIZKTJKMRt6v3OmR0wgwUbb9GQXoPgZXpTEf
eqGyGjxX0bo3XzWjW/ZphmVyg5682Vx1IbDPjWqZmGnOCiIHjR+3TN5ntIU6KEXF
iHxZx6bFp0nuKCkf112HAfx4ZGfvfuQxJJrC4KnPXa/0jxTxXvZvB4s9luiXh1an
KofrKyZPQHeSEgWiAPHBksPsvSbsF846w2+W571UgL7aA0xRcyxkOaAG84Mu+Q2P
iagN6ZfV04hyHQtklJuVEcpQfl0yDRBJbXl+RfyP0t18XtFn+g3HoawYs1RPD/tF
kEQ6gJr0eqHRicpULkiVjWAHJMM3AVCGalRkc2UfR9CDODVldPQBajHk5YVas0h9
UcVW0Pk0x5hcNLuEg+KfEF2yHKTp3lYleKwPleDzmpAo3xeLeTSXPITivjdjGOtk
yyAvqeA+2l8CWhr2JCgLDgwdIdXQ8Hq8bsfiUO27S3SkYb9lt1a+JWhk/CuMv6em
E7qUi0xJ08pAvqgYMcPQ9N0BcJVhIl/bOx07vosuSwwRnaCULX6RHxy2tFLJxaPw
gSVSI1xnzRzoOLsALUhq3ig443mfkURckY83k7Q7M1kfYSFpxvgPPTtn3c0xpihr
wCOCWNrDLbZNsgdXL2y1UKLK7H7TTHOBiFq3BnOxx95o5L7uUSJm7mwBrudanMRt
40VdvSuLr69I61EDcvDz0OOvNG/zNJuQDlu3nqUtq8BlMPJoDF+DorClQb32ZbNN
SA/P0SKPdt7BOKM1Y8Zc0J6KfTFgx6C6jAfCUpHmLbrSfpGgy+jF1VWAJFDPDSqd
2nOKengReTIqvxQYNjpnkoxro68LmUn4b4v9owuhYHYpQcfFZLBpHV89hp4sPlgq
Q1PStFR5tSB+7kuEYUCoOlc617O+RLZsdi2JrP1g5PlNedbAMl2eFt4QFQCadWQI
UZ7C7rlnjwE5YCgeTmLAe8KUPqN9ggMsyyZPMI6GfD/z6c6MX2ziP7KlNaSCm83y
6EMFKLahQVZdx4WMFQY6z8znzygVZ5e5eB7Ue6N/D/aCz+4WTsk4QYrvCxKH6zlh
qj3Tu3+9Ai0GqVIq9ZXwhTGk1nsJVWrKY8qNPHhmHr6ndDEgUFjCkCuDUKdfTs+j
C5OZRKjAY0A1j9M5WE71+/rBIoxIW1j8lsjptMCt+URhuQRz1D4Hh/x3Lj4SJT0I
jT3IXBxJTSn9KMdVC1tLw/ajKtwK+4/6ZRh28wA+JMCB68/Jz894FiD1rvywWLDt
0TeZjRr/I+SfU1kjVyz9kubugFl7On+VF7pfTu6GysCP5JvD+JHBy7fR/zpTZxI9
cLiVMnBZDbIgMHvVqfI8lZQTgqrBtNmyHROgz72Qd+rNv4rcmfqPAwPmooOzWHKC
joj7acGvpT5jxI80VtuLL9pqrL/VD9sSesevs8igvGDL5sY7rKLWw0/ewgmxv6+Y
zNtmyYzZS2lu+c+KuGY+k7P7blNzJVrElCPywsF9e4xhegm9uIrjaTPkfdMkbo+E
+tzTf9eM7ldAHv2kcVGDvNu10nczinz94ZUKTVsnf/YUMp80/6PUC0xt9Cn57cVo
zF8oWl0apNKG40XWk4h940p+EYX1kcoxk7Cw30RH62wUb8AH/3qH7kMddC/ryOO7
f4rJfGx5AP7ME9oacoQCM3pcwZeLj0CihtzWkK5QXjCNGlMfQ8DGt6rbCh0c6gmS
6pk7Vt2NxrHmS+nXRagiWg1crgeLcYz05JlfL8hTDb8FWBzk8tlMu8Pw5eUALX6e
c+d6+mjpXtBNL0/T7XR6Bi2vskT/tq2OtY6PG909C9DDcsKYZuwQZOMSix92vGgY
fuQ1OfxhnLiOjIQSPZPS4r3dWdtWJHta9YC/x5KaIaVoMI1Npie5ssfImHqMtKSR
lCz1zRXps+zKfFmr4Sjp6qHWpmRmq7CjZZoUG/SwSPMqRbTVp+uj7gGbDFlhlhac
NXvwkto26WhGlmKPebu6PGLFL7pv5FLrmIeDRucUAwNeGvidVLAJfOCHADgoSD8o
UY3hhzsgOYA399raCwcgN9ShAxolGA+x10ZRKadBpZSv+JDs8EDBJI6ljezy/KeB
/TX29HgjYvKKZEBOtHoA/7ZD9CXAfeLK1fs0Fmi1XUnBFJENhb0By3sZgRcBqxOf
Gsn7EdmO0LM6PhT9ulzEy28A5tk7tc/V33Ixiy67EurAMJe9B0zZWyWiHZmob8c5
W9LDLKwBlPAAIiuuxZ4zJE3k220ezOrzbiyqNCQRRMEY46HKem4KDUrviI6UUyEB
o0yC+6CNBnwRL2+6OwWsPTx3UFl+wU93JRfY7ekXou+siToogU5xP+ebLt5FjkIo
zJDnRWnYsbtp0kKUlX6Kb8ITN/iQ57V8qXWMkiDpmIPNFRCZb4P4nOr9IYbRxF+H
L0AdAenjFG2GZZcEPKWzVi/Y+KkeL3yvJ+EuVT9bXbEuFDaLKRzgEyb1tx5pGlO+
Hfg5dULH0mH2EvzlKYD9TgHv+JAYw4FfUQasucKh+Vg/KdPGXfHARqQdeBwBzDVW
fIlmjcuQP2rSGICm2pm2WlfsGFZ/0V8+gehgjNcm1ecWbB4GzAmN6PUqMKnFzrQP
bIShHIE3ivVYLo1L91/beucszOuVl8WCI2dkHcu528BnxrUP6p/eGUSmC+PYFkge
Eu25cgzRuIdVCMg+JY6c3rvJ6SR4hXm7Sm6N9+F6/+E9YSSCWnUsQAPHBiDpxLJc
NqsQCxWGZJJ1TEmfnLhXFvL6XNyvE1jCU9lVwSB5eJhXlPZw7ZcLLEdO5Cv7aiGw
dTLSHWtDAA3u9hx47mtc3HWf+8Ivfa7axOI/owL3+Qg=
`protect end_protected