`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
ddtXksX2+yylW5zu6QL2Lhnb2d1sD00763mmSITNX595NcHTEkwn0zB1Dry37fOW
FufOhVzEJp80NC5qZ/+F0Vk7Ik02dIR0elf3clrjeJRK85K4e3Hoo4xn7YbFUIms
l/8VZSb14+JVGURjfswrIyCUotIzlzVYZ6gzoZwDXIi5gQIBf/gI+KxNXPaKV+PQ
Ufys/12rjO6aI/pPlqSm0hCvftmBcnezN2hk1UeXgOIuKZnogjOsf0iJVX2aOOWE
6pD/psybjbnsNB6kH5uFTA5frkzIzkzl5d9+YDm9OyC+k84E83I/7/j+rk4L2dah
QJOvksSIzN867/4Qt8qYTQ==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="MvBXkzurAa5VTw+1JJ70nePUfoQXBvZOku/SMmg4TwQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
oRtzZL4VJ4iwysPsC8SXYCzXS8Fw2gtZTOskLcDV+1B9Nzn1zTyNtlo6lNICRmmK
ZRVu2BmCc2G+fmzynYlNTnSa7C0Cuel6FYpxCBlOuk3OF2tzAmLAuDyOH3Z1Yjzk
a0aHuoCdIRKv7BrZCdALt03JeUmXKPdOmIlkVGFl8yw=
`protect rights_digest_method = "sha256"
`protect end_toolblock="Jn9CQpRhJt4rnzZPRk+dOpzAubz7omckX1MrFd4p81o="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 3664 )
`protect data_block
gD6l00tciPUa6pDNTk/+t0OO0nC/UTtBwLB41d4inuAUA3i/ALrNyoJVcBnAmEQW
ptbcNp5fxEUJjnOxnedyZEuEBxWRieZFQnkRdF269oPsI5UaPdpHiya5z/5ZYLMN
UUXlRnfRWE7kwZ2vfSnwJFW5Y+gxeHSw7Wb5GCzaVHZhvkyLgBNym/MN2ZRklWXz
VOU0sDdkODofi95nu4hyx6YXwx8oBeLNXgnIqZHumqsNv0XsY/zj5D/ovD8SGEIm
Ne/01myeSFfRU7yn7j2psKhHHgV5eyxUtF8C5yuu65bcsnh8RplDkGWrwwxTnVo7
snPmK5r8l8Ef2rpkf1TMNnWH/GKcbC8GxXRVyaGvxc6PMUoxDgso171G+pxcbAQX
/yC/UXPxiY2sOYt+U70o9vOQ13bOdzKA8/WHSkpu8EM5pYwv/jHG/DExh5+NO75u
R9f7+JemnTVMqEnmH9PBarrqXLLYM2PIwD57AI+Vpggo27V2HDeRzIsV5OkfwjlH
JsXAcF7ccNJdyc4zS8zcweRbusUodwlgQyoT01/igF4Up6cHkl5us2s6iK45MSh+
fx4Pc/+hXsWhZw25mC+oaGrrE5obHxXJrDer4KZIijnbV/cMx0qkMz+lqNH1bgdy
7jvbfFa0oBWBQACYIni3H1fVwlFV1HOh7zOwBH/Bt7MmmiH4Ru2ihSVVOrfiwat9
t22oaSAyVOpQ8p6sf+FL/QptJ0mGQjQeamUudYSm7c7qGMyipn2KTSivFZDYXhzE
BbY8n9L9u1E5DCb0SEUdTdSVCFR1rnKA2bSjgQIVE9FjByZ23d5GNxEWoHyBvM8U
BMVPFyx50M0D/kkGgCJuTAAYR6olATdXOc3PtIogT+Ibis3yVCzP7gvnJu6pXHD8
BcfelwEGIVIuWaX1eKuwDqUBDQ5alejTGTXiPK4jlSXkpqS8+tXKjN1HKz4smoh5
Lt39CloZ6ZLEbiuoiLEosdIa0a8h2vA35MBFJDDKngSylVy/eNGyo3rnUiWU2QzW
0Dw/1HeEH4mTFvYAbGJax90A535gY3Kh0aPUfwjb6PKioh+2DO6ZRC5Jrq+E0VyN
fxHgf/df/MWeCkSw6AwBJGYcbsV0qQAhk9ulK9u09ccCoP+Zjm1BQkEjxzW7uHk+
lJpzHB+LfiQ0ZjxSgrHPYjqM1hBQtW/jPiSUD8vLx2M1iSCRunSOmpTmpdod16De
Vf0sAR29T/ZE62eTi5aHnBRc1XWnjG7ywVbDbZXDYLLk/MJyOoI86mwVzxju/7ZA
U+2ueTYvsMxGezrbRRrD48BVSK1Xc+SI8d9SrZw1G4FL+LyBQ6m8tJyAdRxERnpM
cR4PPnj1LXMEu6gj9yH0l1Es8yL7O0s1PD9iXJqrD/LwEdVAcrlfpm++eQptjaQh
xTIJ2jfZ5ChbFAmm6pju7VovLjO16cgfi8NfhDjlFDz6cf3FdIHaRVJfumEb4is2
YgvDlUiJjpG/i8UElcD4d0J7HRrKJRGFrZwa5wcg+Eog5QrqbOvFaxy3uaSfMUZ/
0xED3VAwxZ/Y0fl1fI6U9dWaTIiADzFFVcG7hJg6IgomsjxmQjwoC4KtnkpBceH2
uvf6ozWCZzso2xlzaWMubDrBGjs0WEu9MpZz4zomINGf7KIab38mk2JbX6JRiPln
U2y/Hhd1WS8CDRrcMQLJByYNQY+Njw/7gWLkyYHKJWlR3+4E0p0ZYzz0mY38BNKu
d4XZ+Tq61bU/PNBb8pz9G284izYXzTbGxEkeDqaQT/OUDLXDCbgLuPFF3Br3/kVg
zKmyQurUIHlOXR9WiXYQp5vgE6GpqmJcL0qJMX+OPhjKSYFPdYcUqIp5l6IQL4D0
G46eYhX3SIK0UhH02i+XJOSelxn59j3uZ05yhSmRU7NnvfhBj3No3DbMLs5O/KU4
c+Z3Ley514LQP4jkUa9NOZxDaAzEgrgb6a1M+6jkhz9qY82+o3Lhd3Bc1Hwmvof2
rbZEjgplDg7DK5I+qXgmzn5TceEZDQsj19aPKO8sto/PzLUWCPiCdTN1vSNaoHPg
4y2T04hrZsrkvrTS0I03Jz11Zx3cQIn1XEbC6Gjo7V2vZx0a0eaWEc/fPnBsL+QR
UrpC3JRcYz8vIyPsLv+kjTAl+AbSLMGU7hkWOskZPtHXzCQdoHX+aCkBTScPAp8G
QrmDypu7gpsN6NgcLw1kNhaxD7r4zHJhBKtffDABLhMCSh9bT4+4Xp4D16vwmLzq
USsVW7XzkGPk8HaWJkG5x9j7QBsvWG2vFUBLri/sOs5lAiBXL0GjCQ9Wi5g4nsaF
xxUkP1KorGnrMKRf68Np2ADe74EBq6KBcQ8snMMBR6LAtdzp7bD8XZNmIRA6EFZh
l33CFUh7EO6NQrd+m8tD45CDoMWxHGQLYxSNoAuQyVoHUlEFDKj1jSU8xpGXTl3c
8axyjJOfrUFP+TTXHUN8GUn7CcW4ROvj5J613La+2gBBmBmdwVafPISqsbMJBIC2
pNrmeLBlvqr7EZ28i/ctFxYaiJcZHcmEjp1CIGCssr+XCWeZkC0Y+B8QZB9An87D
/cBVCSH3zE3mmQuXx3jSeRYayT4+D8uCkVOBHa5IRN+xSNg0T2UIhP3gnPf27fvt
tvOa7HzF6c0u0jZix5hRdEJkul7JWlMyF7jW3ZMGzkHAsHFLBWgoFhfYbviza7bX
IuodVEvOb6LDE28rLEHNSHuv2H487P6zGIpWhFztXPlFtlQsVfbs4wU1/4bbMUjw
RkhJvCWZKurpaTdmlv7ZQY2GUvumFlBRF4dzbY59zDG/stMD3JL4X214uwaVJJVX
5EyJq//y6DTSWRZlUyrpNPQZr7grYYPOJ9ozXNrv/Whj2FA+mjnClgCzmYBiCUaJ
kmoekBPiJDCcJh9m6GW5m51lwQYkscaswkhwBlqOKWpZrc6PYrIcCemlL2Wupleo
DsNTRlAcOMU8ATzsG+UK7osz+QP683bBzdAx7iiWOQ1yPIEhuOi0+IfTpVg3p2Xp
LqNbK4Gd0LtuA7YQZXXCazvxdAsDcrpZ7zfxWyV2n10+lLOKkiMPSo7oPI1DCpTI
HOE4y3ZOyXAibfMsvzKq/LCLFmdto0n4AzU7Nl4JHxkmEwHpp1fzOSscYTmzWabR
S7I/edQEAguG7CEwjUkH15hHCcSqv5fBewfvYd7zcaChj+7OOjJpf2PJgIeOxMvR
mxwGGVyn+IzGQXK2QYd9FiAoJF8AfZkf5nVRCtIilB7HQ5+Hl+AwwPFii4PKIXij
XNbWe7k1UVmhwtkw/xSQLOMmus5rjxibO+2XBF1UgOgNiz7FtLdTTL9k9DJ0RI1e
krkqMOh/prIy99YXgJlkqLhtTPYMioatBaKCSW14o5Q1sX1kLTWtWI0d3IKPw52G
PHIlfX37fam/rVgRXPV0bZFkzI2LpBaFZJiB96LhlGelPG6DeC3VrQSx+AWC5i/3
uKIzedoqUWBkseDf21PnXxaofupfALd7xczIDxlqFeFxaUOrFmWppHKR7ZOBdS8I
q2pgflKWCVWETWJG0lzBMkAFIkTK7iO3vgyD4/+JpMOxoJk4Wv2Nk3mLZ/rflA2i
NmyJfIYRmGylabV25JxwHIxlCvAyH4qKui+qUL0C0uRnPVl3VEYP+InZMu2IMJ2J
YOmuURZs4kJKywd4kaBVsc2Zxg7b0C3v3rA1qmzBlGdWy0AzSronypJfQrjhUeyt
e+BG0fSfVN5TJE1H2o4m7kClfIZ6aj3XpuLWP3KhbP0v1vEPZH9vqo5Esuui1GpY
wRflyPTAnakoRLPzGDB+0EtY4T0eBxldx7B0Yziy+0mwrPsJOkXpWpUQzTLDYhlN
tz8PJEN4GDwMM3Y2ZS98Qffu+5Ko77FpHcQpvLO/KrZD1QzA4QisKrv5MrgCtbo7
CIrzKL7ruh0dur4ekWQygBkyrnihBXYb3mt1kSzPPL7KcoanLhv0tihLdit0Lgmo
KDKV7tGobCipOdLuS3zM/1m0Kl9dNSAVUyBgnQ8QPKFyfT7nbo32L6MnX18we/1Y
Ot1GYBcRoWOyV/06XdkFHrsCPth05J4zEs5jhsFQ+Hc+n6aeLwL2LACITLBP8EqR
5fNLn6B4/b+Owzp0d/MaHK9wIxdg4lDiTMnPkDf6UqRq7SNzNBZU2lMCKVrhEsX7
/+frtB2akevjuLTc3/mmJ6VLktoUiESvnINRyFZYr2wKocRUG0+7QoghguYQqhqq
zwVPjEaDjeMpwEFk/IPA9gHCsSHbBdMMnFhMlm3z0k0Ktd2euzBqIYdpBQhgxiTC
ebSzmworl5r5j3JGDsB/5r6rNkOyvcM91oglI3k7z7JwLZfbX92dDsnj+5a2eRA2
M67Yw54KV7t4QByKgSQ1/e9r9zGj+bcAP5TbzVspnD7slyyYfmXK44pVXQAOlA/K
kBRZ9pqcpZlFrvKZOAj2sUaKJV3j2PBNG4uXTB1M84EhWcqpfhSkBT+RF7re7ian
QMvTuYxk0EbbxIevhOsaQJ3Cv2wuH3LHw7HCFXhefG2+gCFwvQE+JGTHbYBSLfGe
dbh6tETvsDEV/ExN2DRw8sUJA+WXimp9IQO+mCWGX32HYOwHSUFBF7FxajTcbZHL
JO/AfORg+ExdWmoiH4W9GaRuyv8gLtmzM3aqUCslz08jWw9gTTQirkyPduLvGIRX
+wQ/RxxxtynjvsWOxUIRnWXL0QjcQxIiqIZoh7a76ju2EeWA+qvp8q39zSsypCGS
fZMZcXlhX/XAcfBA9Vf6YWIUG+TRSdrtXPle9Dd900Rujjhlov+tZzBmzG4Y4O+E
Yv1aAPNSqYYl55RDLd3kZGiw18hZq34iCgo9qj20FdOorrzHCwXkmpLGCC57g9S+
Gz4Ohz8NHeAWTwsdszGpcQ==
`protect end_protected