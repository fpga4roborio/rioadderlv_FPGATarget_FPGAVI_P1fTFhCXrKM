`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
ddtXksX2+yylW5zu6QL2Lhnb2d1sD00763mmSITNX595NcHTEkwn0zB1Dry37fOW
FufOhVzEJp80NC5qZ/+F0Vk7Ik02dIR0elf3clrjeJRK85K4e3Hoo4xn7YbFUIms
l/8VZSb14+JVGURjfswrIyCUotIzlzVYZ6gzoZwDXIi5gQIBf/gI+KxNXPaKV+PQ
Ufys/12rjO6aI/pPlqSm0hCvftmBcnezN2hk1UeXgOIuKZnogjOsf0iJVX2aOOWE
6pD/psybjbnsNB6kH5uFTA5frkzIzkzl5d9+YDm9OyC+k84E83I/7/j+rk4L2dah
QJOvksSIzN867/4Qt8qYTQ==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="MvBXkzurAa5VTw+1JJ70nePUfoQXBvZOku/SMmg4TwQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
oRtzZL4VJ4iwysPsC8SXYCzXS8Fw2gtZTOskLcDV+1B9Nzn1zTyNtlo6lNICRmmK
ZRVu2BmCc2G+fmzynYlNTnSa7C0Cuel6FYpxCBlOuk3OF2tzAmLAuDyOH3Z1Yjzk
a0aHuoCdIRKv7BrZCdALt03JeUmXKPdOmIlkVGFl8yw=
`protect rights_digest_method = "sha256"
`protect end_toolblock="Jn9CQpRhJt4rnzZPRk+dOpzAubz7omckX1MrFd4p81o="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 27104 )
`protect data_block
gD6l00tciPUa6pDNTk/+t0OO0nC/UTtBwLB41d4inuAUA3i/ALrNyoJVcBnAmEQW
ptbcNp5fxEUJjnOxnedyZEuEBxWRieZFQnkRdF269oPM/dJLjVQfa2HF719sJBwd
Npecl7CEHEQ8y0mI/p5uGS59h6iorBX6rurC6s5jqyo0C6fu636DWUlpejA7aBJr
LszXLBalMsY8wcav8v5dmk9X5v06l1VabIuCkfDkWH6413cK62zXDbj/l0FdPwaW
dGYvxmnlVkn4op5grL0Z9/nSG5S4SSBYs8XRhLFhkMLSbI19IKIbKqcWbovbjJnN
uGY2rbKfKFnz/Rn0fpy1Ni7qSIqLaPVt9YCI1sZLjnjBIGOIsOEoD1OAp7c1DVS3
fHIdCgfUdEwcZ3n1digWmOCAIJ0kNLEYRjgRqRJdZNV555tQ3vlhOl7BCfCb0PFx
1QwvEev7q9/e69PGtM9m+h6glQ23ZYXhnA+HQkH8FNSoMRrszbxgXcrkBgwN8xXS
g6tY2jdGtGudRTdO8ouUXbOjw997qWg87t1Hpp6bZv6X9Ssfd+7pvfIp/D4Y5At7
/QJzTdYbouv/U8jEyyBh2MiNX1HF2J82/t+YS+rT4C3HHplJyfdMfs8RCYA+rgs8
D2vOnhHiYO6jJzPVuD4d2F2qmZ/TDD7eAfUTeufjKzOvBnH6BMH5bzEDXGHdHYVy
FPUyP4o3z+MR3G6hJEX1e1jKmsj8zJHz0hgnZTeH4gS3D3wdpI7deFDKcqpKLkMX
GqQVOtgZJEGd3U/lpuc0f2kORtOj0OqPqwRg4zhWeyVhTrbf6sICahJGki54bDxw
WJsYLKnNu4z3fS7LJ2g4S8NDOIxSnBzqrhWOUWae3xgUAaNGwebndqp/IKMc/1Xb
DHAXtZ6cbZb+ziwBbIHEGyqFKnviMxFBDOLgSe2D0CeDlJiKjUq/92Tvz0NGpjbl
lDlHoI9OpJPFTIu+jwzwektqW6v15ojfj3jZ/BlplQ9HWdoBKu5Jr4WN5k1bS1yv
+8yjyTtBXnTeNCTFvNYJUWWc+O7m/+1+nacpynm9UJlfVBhVTOznRglaoFU8nn0N
V2XpI8cTluiVRXcqmzic7gbmLq4xj4XztdvVdhONjqDaIx5gtONFjioVQU616sIa
tNAeDScne3Zu7KxZwO0FuZth5l3lGOgT9ByTF/Qe6e/19Iv6S2lVc3qd2u0NJ/R4
R8Wbui1jvqk+57uSkWPwEgR1ezGgtOC5t56ye49AqKmDwOTye3vGnZvA7YUkagPk
aAS5T/I9dzhaK2jusI6H1mqe6UiMylGT0ddqbML0OAlf6s0GGzJCyTpAe5P7znC8
8/2iPzdNo18+gtF8P2oYhNj3Uk1aLFrpj52GRLIjcbGx9BOw1BHlZNup+0jiZzjG
wh55hR/h8vq3Ysz8n3o81obNWj8DYgkDfvrAojrDtEOfdEO40Z37xgJ1rSwnQClE
XViiBCr8sXYcQ/suTTvjoC9uPcnQwXDNC0wblXP8vlo5SIZw1PHFqLu1E/vEuquT
5nO92e6phuVZPn87TXvBrFHOi5dvsOPx968Yi7i6tvoM+a90It/l1rTMnu0MTiU5
ZUaElAMvbz0AOmb+L7/rcz0dTB4FQO25Z7g2Tgb+KhTPqYmYA5Ne54hQbSxhu7eA
dWraXxviN5U7KxYLO6GfWaxteBFdzPsypcIRdk2cs/XRBYLYIqruUjVWPn/j3F7Z
tjH1fJ7lzgL7zwaLVOrK42flk36IdyQAg6r9PmgMZOSn6vqoH0dclDvzpAnr0Spc
cS0GxP3DdkzqcSd9R5sYbqIs1ivtxazZswhYsauI1UODpTRFInFhIKuTwQbKv/F2
5iCvlIXpNhHNpUutvRX2cGE+p1P1Qhq/TnxfQLpNFTML5lrznB/e9HN0HWKaFIUF
xCyDQDlOrAHJbkRDk5s4SmcfKgB63a4+zs91fZWoSSRhEG7CoZgCLxKzqja/I8Iz
fszJfDP2JaacZM9Inv+sVQ9f+2byNy5s60a0l/wvUXyCtP0g0XDDn9+sxjCaJfO6
TYnL9IWKB3yxWbho36UBxlnJntYV1CCXzktkoAiuXzm9V61998/wZDnLVekWTTJg
frXq2na6KmC1BzhvU0TsPshdGHegqS5FP9A3aya1ljI3N8HSMbuABbcVgiiIEktP
2gyGQdfsfQnvdepTYeiwIf6epNGyeabtn0hinCADWNNGwAllqm7kGVUT0UZ55VtZ
GZBp6422LAyk38y9GS2jBh4VUwLMKtBeOeWFlaS3jrHPhCn2e+M6ClolEiA9AW4j
PeiJoZm6Q2O3aXiF0gNh1tHVHKjzNaMhY33XK1KENgyz+wg9/wHJEBPc2AWP+HxK
381vblYMKXLi5FhxM5YxoeuU/qLkiqpb27T3Cy45V6gSKEZjhYhhnLPHrkJYvq+w
lCgW3ggQs2q9n1HZ4gJdP6/J6dJku6Ll4h2QBDekCl3MxUF3Dn+LMIRE+EugZrfk
zVkY0HcRjLf2TsSmfBw+hPF9OaZhsI5Sc4iQKsdgxdNSUMBNag6mop0/nwCNlUqb
xBT2r+94VIhP1aVMh4+SZaCdIySr09mRcBrWzAEO2ECxB2icL70cONHhE3Ugwr5Q
GuTL4cN1DGqL9eJ2R9xjPWOQ6gGSt6/9YHFuuTecpCyy10rRlqgP/wCtUkZEch0a
6GYLoQ5yE4X+e5jmDjNiGIhJwA3kkWieznPzpU8QxoWojD9eQDv3/lOURFKmHKox
mwThfoG+lTnjXObsyEAcc3Gb8E37F0hv5MPgeq7Q4NuMPSIlLG+LZGxZlo1uspU7
rydO283eSXC1einV/9aG9+mgLi4RabxVK1Bkh2b9S04Wg+RzTacQrSpzjToVpKk9
v0ZmZ7rUVwPA2RTI5SQupmzAqc4BhD0Qua+zlOe6sUkyN+NvSey068n5gSWjL/kw
NqOPYWEUBPrccW+SAEImf3vPJ8LovI+ryNVLzFDtCbKZ8FTEHYgmk+StJyxJWbmf
8Ws+6MMhuEHVBwPRf8qUHOzItXQyZWnOQO2LZWxI7d2VavWTJ2/JnvgNEfZzmFwJ
OiqmP9XsVtg3P769uLUQLxEl1e4Q2FHLTU3KXIT5woBj0kHznnKIhU5uW1LMDa2V
r8zxLdEXzpqYMQUxlmWA7iwVkiJWRApFIVaVXy8B9ZFVerpvzibX8H4qJKJ1OemG
s0j1TLV3TKo8KIahKsm161QjHnYLf9ATMoRkpl2IDALqmc+hIJNKDP9NFCEiiha+
UuEWqsa4jt8RQReSUbHkJmYDAPoldGWMPNfKgh+r2TNjhpcdghDAqE8Pq645z46z
6SQ1fpgcpRiB2VL3vVya+8emOdR/WGrdlo2lv7aIZkodxbr9nwQDTEOOpJxi1/GY
/vv2NsnSz/VbVi+ssgiJOkgCYIRJ6dam8XY/5JvEElUkI6QWI1W2sWdF0MuruKWW
GbakJTppNJiNyMIdQpr4TnA4b9HhkAlaU5sXRsmiGyOnWo3VHfhqQAvrClEXQMDk
aEBDR3Zyt+9lmur7b1geYz2CkG5ypvQx9c9Rc0E+BOXTLiD65oz9QHuSKMoBSyvr
CrqsczMsKIYnNTpDjSotulRCcu4DfNwfYltW7uI70YbWApJfJJG/qHfujmLW1tGR
xoyzepqYJlfmf3GwcYfueYKLlw7ROHNPmkdu7BG8DRV5TpoOufZ+BRLQg23g41I9
wOEkX9eJ4LCjd6MH8RkdH9jevdNzHtNaF5vt7L1Mq4ZdYfZiatrzeUFMhZUsUYOz
tV4bEtIpwwmdWDjhFIfPWkcNWXzB6nQhkezcFt4MUKK8o9fgTminFqIaBEIGetcB
1nPv+qE0xBqfFEe8lPXVHB1Bd9vWL56E3pxZSEbiwNZmJQ4wgBI0mU+azPCPFVM/
OEdUyp5KGpsdGalphQr2PXFfs1pLbL+jhRvyaAuLfrKZh3CFQ5weth3LSg3Al/Er
EGm4KRyBeF3oMaXzmbzun/TFCqtTfsXgoEFm9/fDlzF2BLSiDekLARVTcfV7smx7
xMMiWWcQ717BG6faHwDWdFelkLWO+07Xm9+V+riA557q8ZVRio5MB+Oj/w35VGu9
0/vnJd4DEYwaK+m2VA2aSoBG29qccsQ/Z4yALETB1ik/ujVjqmhaUvvb0KFWIUBm
KvKtPPoeyhwcy8KixKxRQgoOqSpkCLQeZL7Yv77EteJb7qHKUWZNqCeCMmnw2uZP
s/kXEHvxeRgfZcAiBTXq7znzSI4CW8BJWCjmpdORaNfzJ2EHZwn/i/66ITxKcA8B
fsTztivqImnhBkMSQsHABCNfzM+kkdLkP4GrEfzDZNlHow6mKAwupjVmL31iugnv
NmS+VEHjDz8zK7PQPgK9q0jOkHeuxHAnAi4iBQUvIDaZuzwu7HIERMzSv/eQMdE8
KiyK5ns71/sfb0D721X6XnqVmkK1gnVJsV1CKT4msLXVepRHJDcTCADODdgy69Er
N3ix6EtYHDE2CMgQ7QCE3+/WF7Uz6AIilz0WCdblAC8Fy1WINwPgD3E/zpp5plih
A8uODVXV+lq7CxGF5yTxLsX1AkGyvansVG7EZZe0sfj2apGDdIwed552q3FzwYdk
wFJSC4hd/MgCGifjb9T2HV6KRUtqTltCiJWy7yWTiPmYZCTufu87qpoBgngJTpwA
URoKed6YPilKeeyJHgT6mz114kUk/Hxq9Qaim7AP0I/89Sbq/TvTE6KVqI8ffZ00
6PJ4OZSmKNPERY2C7k04fm4U9/1eI49cp0A6bj/VL4oyhG5ZJ+LSmTV8nTzVZWV1
KzBozEYsQKLyRYrs1JbTDT+MYGIqPHcJzfm7Se3UmW9+b39HrXyRld29KsV3CTUk
pFCMODfTEhBnV1VfgIh5YtzqycGmHlVmVvPXlnQwTEcAL0kK/qxsbi8NH2teAXLU
cPBvq/Es+8OT8yNcqDrSJVsWfBI8ZZha9tvRbDI71m0KDjGDII153EgL5uq/6mfg
oZMyuBFe+cxlc3kI9gTrYjMitQXChiUNnwIh0MHQoNY54z1La2zeuQ0jy67aA4ji
k395fEGOvLpi9TxxnfCfuT/N2dINBdiQlZ+VSS/CR99avQzWeH06TL7pOiCcboyk
uQlcttw5ej7f3wRRrlQ4gxgsVPG4QvfyYrCFRBz+0aoaoAYBT3e/46o9t4CESET2
k+d2Sj5G9B/V9pgMxj30WubNw9dQatPQC9pBJE8TiGC7mMyYtR+rnRkJfs1rugih
skmT41qMVPJzavfBwov/n3sXKE5mKie2qpC/8as6yQZDedK9erON4fo1gQ07ic/1
RB/YKlj5I3pHaag8TjJsPwvZlH4UGjEmjX8+0bg4k50XuUQBiobbRg6xSa1SU5Pc
HBJIwV5LalWuxo+pZupT4JyZAIwIgVNx7BdXfPw22NgqvpOVge9e+2EaxDTfNokJ
/pf0tQSzqN/fe42pfY/QhMJg7+n7v+uC+nwFfy3t2IEeva+cwUlrlGPmcgYi5bH6
bobbGLd8sdJWL5WrrYZSvupEBOTbSCvXpGODBSHIMNWdFNv/G2R0X4AbX4pJ44o5
GG4kznNS72iKtI8VItyD7YjI9SgQrP12nZYNNXoxahvnRgxwQdJ9moWV0+jIEv+P
kZMMLSlDqoUeVP0hrAVWGnAQIC7uDkMDSkIh4ic4y6Tc8+nGhV/lKWma9TP0DnbR
VqSpX3VbLDBR1wqqvYZU05Tig6/iyx/amqjgLUiq0fybj5W740OMWxrUsRRMiMgT
B42YCFQ7h3vTbPNCcO4aatHbvQVgd6NuMucuAISMjg+SvNcJlOoetTPBEZnEG99M
Gtm6OiqkrMbWu4tatMI13dlC86Y1q4jnylkWwcLz995RonO++qqCALg72wuFLrQp
+3VDBWbdaRvHrVHZlohNP+VmgmtYxB74dMWEWuoA2Vjh9wGamItHjfxuXdOhiDNE
iBhrQgon85YuRv6qasBldQ+KBnBwctZALSkTJfYTUw7Ia0zhV8C2Z4rpeoHDLsU1
LqrAODdnW6Fu8RXTg7YcgdJM+vpUJRk0SwIDip86rwKuoNW6HwQdS3BH43qb5GmI
Cgc2C0CyCWAjccrFv4qcpqpyom9BtQboGUN30whAXRNTgIJNWN9qYH98RMyacwkT
tb7H4l6ywYtqkiKUtIktmesmGcxwyUaF3vfLQlpptzduUHUuPlV8DhtYvjx0kEpU
cixtPaD2NV9+hXjhbJx9WBn+/KqBrx474dNypxnc5qi4Nwe4BKVMBNHmOndAJBsi
JkNg1dJ1gh/rvqD2Tb7TRA+VNanyj8uAhaje2PGpf97O4msneKuwDkuH9CNi5zqZ
dhunjA93WPaL7+pNWIFNg2qr93+/9PaMmecKGLeqaP4186ItuF7jxebdkx7UWB6U
u0pZGxcN1CxcQM0S+rgH8hIMHMSobfpq6CcHxk7zWVNu/ld+oKe0tcj6dmGMP63s
7zOjykjWWt2NWIteGenQLjCRK2Of7R+L8y4VLLyGPEx9g3nWaB7Km6xPujq20qBR
wGPFP6lEf07MYF+F+fUPoJSp7qPXox/SYY3FUqvWEcndyVKclVNYZRRcldA0IIRi
dT/BTrdq5agixAQ8dOp4VV2n2fDoEIL32Unpn7D4+6v5PZ4Qatm/zAj9TncKCtna
XdsLg4H/0MYPvVB39osayWAzz0QgRbLSjchyF52gKvkmCJx7Hf7ejI0mwjH/95uJ
CXoV3qFWUW8a2WVfgRFYjrS7eeVxXOifrM12OYmP+OXxu4dgKb5P4oigmDP7WYLP
807Gb1zgwi0m/gkdPibXyQU31WlL6/wdQr1FrKM/hlkP1/2vP+ED0iOrP4O+WAXe
a2IBG6rsKDZjNoNiMv4SXb7fnD+9TopEp+uCXyrP5j19n4UB7iB5BiDCuRvUkjfl
7Y6JmnHNJNespU1xgeMgWk7QRXtPAJcvtXlFQFjWgEmfuNaq88PgG9sqDCX+WiPS
wz2J+/ceuM0U/DxmuP4MGb+FJBQuwhsci9Jw4Eesyz6GBbSkg/JSbkv/rwe02DRW
BpF9R4RDLLxkjuUME9LvXNHOkE0WV3lj8Vg2Kc40q8m4kdYODxy9iNesbgISM3L3
n/YSQwshmqiq99OE/kZiCqXFVpVOBA5azJv7/FWBxKnnGqS3Fzim0b2TlKZC2WNU
mi9XaHMBPocIbqDMhjSQ2aIYuyefaKaowrMv+dB9lk2in9hqpyPa6e+WeEpJHpeP
j2+QB5LzlGndD/nbZr8sLB/xntSUPOj9jOkaX2+l0LKRBSoblwRDbyuY7uc1kip2
hA8bkvBINhUQTTYlu1gJSSjjWDecablbwdigyNsIhgZLd1KN+9DU4N5F/0mNMfuR
alW/IH+3M68z1P9REPRKLNd7jiEFMTvIAlU42G5NeefDW6wgvwn5xMRVMn6fnFDE
d7NbCGVY01vQoN3AE5aNBXc7hyG4PiHdUQ6/Lznw6FBYVKpzL0t10JD6Ob+1RJJt
/BzlV4tEbTbFDowHWdjFjFWKOR92r3cA72d4qF42QwWvTYOIJ9YIJIKtH25cu3wY
ZAymR0ZBorMDzxOqbOFKdr8hLWYmNgicac3tUg+ZhzE44lKoCqKvyKA4V6ewesGa
b+pkY17yg/18DkSenaeOPfBd8quZe/JUkg8YEhCoLAiu5zJIZ6fQ4F5g0dRzbSG+
lliWFp5hFOFd0G2/byrIxrEvtpT0xaOKl5hBT5f1Hs+rw/xbF0YxCP28/cp2Ded0
vAXLRqCxGnWXhKP/OKt+Xrk9UeKLskvfBFeA4WpAZwCJ4Mp81n4/LSsgnF3ZodMh
4yHXbvP3iZr+FH4FamHY7cUNmnIuDXVs2dcgeVkGAM7Dcrhcuxw8oz01H7ub9jO0
h5HijUxdDhLHHe8FBSIW1NouyhNWOZ1YvV56UtEh/IkxJ/dTZhanHm8Mp6eicNqP
LCqM7GV8rGeReJnJfujKColbhiVcMltgbnYHlwTuBxrOMScdCLgU/pJ/XsrXRDe6
WgXK3R2L4wzkqSH0GoesSfRQujDvC+TLRCUmnhJ8t5vzYRpsOeei4NjsEq0JVBGl
4ak0PvU+5k2MKv41rBAzaNnx5P3dymQMDdnMuqCFsH9vrWUJU3erX/d/LYGiDyt9
pZ6Bg19q1BRunROaeLRJpmWCRt1Kvzl2knsc2vHgQMU3NvATA648zx5uvm26YxDa
ErRg1HK0gic+DolaQVpepZlm20PQwp4Gtd5MFp4zsXN5s51yvlrqt2RORJq0J0cJ
E6XzQuKnnyHUPsDwjRrfU7Q87NW9B4i1+n80zSUOSQkDGwx9l10imjVrXx8YVuN4
546D2+hnJOh5TZjfS73n4OqP9kCR5FzOXtWeJr05YY9kcu6ByoOImzGSK48vySsS
/Cd7YcgnXCdXJ22d0uWoIuxTKD+lY7MvovWUBkb4cNCkpQ4kClbMUx20QPB3Omp3
tS1FXYbWuScdlQhjkcMtSviVnwxavO8y/gdjzqi/r+dCzqhsJDlMVyw29NRUqowM
8Q5Oofj29HyD9SuNjsbPabAVBHFXaA1SjNBprP/MFkffX5W3Ymo+uJsR8Pb1vj9H
rgra/DMM27rs/MeA2pYBWJCZ7x1PCAcpzvnbNbghKlPlqUhrfc8OXFXZ4oa7NRHh
npFP5xVk3lTgUwzzHkYuMSydmIAhkPS8PB1r/NVb3/IvPgIm5Sra3FSDCegiF9Ic
Ki18bPyyAEsg3rH75j5230Qg/FUgiMIlvqkJlSGudreBhNJp7AiOVMIGqQ7wzmeo
g5ikt05RCgXB2eaSoF2WN5ncAbjkH5q6xwb+uO05eRUc1T5hf53XvGLzSKInueai
+C5U7gQ6G3jcwaoipEH+cGcMYjOx1bezoE24F5drtuI8iYRwZT6NbV+uHXP5kEVf
4fSxA+QUAJNzmU1a39xoIM8yUeNyVHEAhqx+HgTWifhnu6u7l8VsE2Cub3IKonj9
/LVhUcv6X155Gw0QeURx+B3maYpkRTQz/ZjKnQqz9A7ENH3P85TMfD3XgnkB9ELz
xsuX5H4J/ZJtBqrb/gYSeRbUEPMnKVC6eNytSwceYmlNBGU8pGwyjRGu4aI3PorD
QlulwP5KPuHztj46BIj4dhYwDMvSey652hipCaSOAJwZLzqg7DJPu1MMH+OpCyFp
lRnImvTSKU2hm5XkBbtbFpin7QkZs1lNjrgnxoj7aRtkQZUzWnJ0AF2blvlBKi91
ibKjwNKVxP5SK9yNtn/75ZXcJ46xc39nfo3Gtpf+UGpnuMGMMP71TuQsy7LnR6ou
6Y78TST2sPOBbccm+bYuHDgECpdypt3MJavYblwY769QHCQFOV9rOMNWbz46yegq
vB9iMFKDFaLcJnvcfKPVQX942iDNuJd29O3J0m50hZ524JfZ42ifHXqHLn21lYcI
8j8m1wDnOWbGOXAR8bcKT6ExZsFH4CMP7iYgn+1QizpDtxv3TZoEDGVEmPfIbPiv
UIeETiQdcthIi8dHZRZYNUKaGxE2V/aYhf6t1fDsR1ysBXvwkmAWIA2gcyfsR9sL
oDlDrkXQY+9fS6/NMPoteS2anhnuAzfLXzKHO86HJXkskP5oigHiWBmXIU37zo0T
Z89sb9IZYYX7T0ZQAdJLTMx5uAuHarRKjm16OSMeoW9unw9xmWxNlnurE/OobXpk
2XoCa5h6X4dBaJcV1QS4fBQ0IUGfquIvatShANcOSJs2xRNwtjLrfcnnKOIHMU5Q
VJzfKgL/Xmq4/gZNMFY+MDDjRYHaF6l2MMsOJ+KaPZcG2cHyGFlgCH8/93IXrNj2
YOTEA3pV7VXRTV+7CeFD7IwPBioNqzS4cUSW0cQPbMAMN+PznWTp1TaBSd21Xz6f
xgl2onG6JwKAFjjsmZE+Zv/dp/rM24x3dmVsZWiUqDgvqb1AQR13pvDO1Rq1AUID
vMC+lCL8G66qjJSwcxDh2yNFYmKQ6BymPJ+dY+XQFdT+6laTJvV6etHQCo0Sen7j
qTXx/36lU2XYVgAM44X6nssfQDIrbEeOLgJQqMrRTOqhHd171WL/26n4kbTWQzUI
IyYC8ozWQVPs5a5ihRZ2DuTf9aTiApSyFSv8hX8x3DU+cuaf/0xNqO/OcEUekyWd
IINKtSbg377pKf9rFSLBx6f/9ZPR5YQkSuZYNMux/WC1ext3XgH/fFz2CUnphh0X
q50Ip5GhBB3lqpF5rr6Gfb7rG6t8G3s2/mH5wd7UCZMksNXC+ERJy418oLTnBAaG
J2tzMrbeRa8fUhqB63iTcL6s0J0/bSaItdO5qWqpd8M9hr2dvoFkysoO+Qt5IpLm
jnB8g5jSgi9RSBxTeMC+G16vxhN/6z8/30nUmHB6cvmfXUWPU6XUJW0AJWsa4W4+
IQQvUF+qyp2QcUz3cb6manH5aW7TXB6Ycp7foDkGrRt0wXArMe01VQ5CQUyAkFi8
3Z2bCC/PnfSfL676RXhzpmLWjCOObFjmeN26wuFB1838FCbcVdtlZPe8GNoaS2ut
GDRMsHOgajnEnBKr8NqjznuaYdsPJSlgX6el2btkMKstEl9JGOt+4+ghBYelZudC
VcKoSGRyql/c6NIz850WhM62RJMV/cZ85j7FuTjTQNLje9GMYlU//mR7lg3eDdv0
hNZ8IaTlE0ZdvcCpSRwmgritrrjkBPtDmzTJdPgLmlFFtzigmbDQIOquyihTB9ug
rfzWo6up1z8elq0buaaKU/S1qNEjFop7p2Z2ni6GqUFk999bV5xeMp9GWqu6mf5B
QPdeE2HiMuegzkckBU4ByPVqJuDvlig5Qx3+c+StgdmNOlITqQ83go2CCMEq0M3L
mdfXpfUePpPx2QykkWAazq+SbrGvirDev/S97W1syyszKErYhQ0N6//g06sT4HUH
QNTVZUg4ZmvsTeoU1z1b9LzJh7VuYuPD0nN+djkzLr1mTjDPSR8c/ZTsb0vj3W7q
10QHlfsFOcVld6/wanY+5LQ+qcTEGEdt92nZ706ZZH2Fw+b3nomFgyeEzBax9dne
nq5noUArxdjS+31GT/VRvuHDhA0b/zb/dgxUmHqJ2fkPcqfwIBpp5E70bE5Ylr1H
6beSZnqbNGFjN7nnC71BLzCEdZCcJ5DCYeP5KzLpFy7mec9uzYusmKMJ1ftJYeIW
4hzQw69MM4pIPT139XIuXF7b3ldzuQwZiWWJPfQ/YH2pdqyAeUoNXnMbqJzbwXnM
86POY1KxD0hniQ0rxYCeGejI70DibLigfPZTmc+oaSrfqiEf95HuYkEggQNMO5Fm
KWh7khoiiMtdZzZhGFrDLAnZJO0irQ12BXKMctJCKDcfSvzK9i0VIXMHU9yV9RR9
YCVVwcvF7m0JX5P1QU/oYWFzNitBiARgDtv3HTpOw92Tg7ZxOBfRWH6ZvnLZqMde
wDxaJ13JhxmZlkXOYMWEJ1CRaqFNPjcdXub+jaeo1Zugw/bd4Jd+/N47yKKuIsPl
GeFXyIbemmxQmuBE1oG11o9lvOiIC+VA6Xy+CgLsny2hp9RXdim83BdPC7ad1PU1
IBmfmoYhTdArxzz0CFhj/BYwv9RxlNjoNXNIy2rnlFnJ8hH5f6FVGhZUvkxfE48e
wrn/it6NW3XKoSLOk8nUHVhwYDe8FNYPO3q8C4102tOCVQEo9pX0zWWY2Byr0JpV
8OFpf5evz/IL2fyJXwMsaok+hhsHvwqLug685YMXbu610X7ybA60V/ZfjoUwT+QP
O6XPMaWnPBB2RBgd/UAoLElVWI5RoOUQYDwACDSwxg4Z5/54CBsbS87WZxHbIC8p
9xh2S3LAPaRcgbIOKhex0UiWPGk/T9BiI5GZ3A7Bf08hKhjXgxH0Na+DEwnPSAJk
aEErxN3kUC5dlNcbJej5afWE4H0U8u0zzQOO2wnJ2KnMLJRXVjYs0Ny7ebjNHAP0
PvWS+0ZP1iMJQmvn7LFMQAkG7imBs2kRnrd2mjxZvDRMkba60eZeqaFWqMK4Nbof
gI3QHkpCcw4sjU1b2WJgQ7NH2d2W2Ibd6a+SElHd4Yz2lGzu54evE2Yjxp+fVK2+
2qNOsCp6ODRJuH1AVVHMtKZOOQxHzheY0Dwge8DEG2OmD4PHiH4AjZoMWkoTmgmV
BLbhucxq1slQ4RrvTLLKTCmhKUmIuvUN1gxHstV8KXyGNoxZJzySobfNZ3NKuWpo
wFcJ3uolIOrddgKx3SBAVHhKAZKwd+uLEpYtQ8kREcH+ZPyVUqelbxl0sZ1FWJD2
03HO1hsdL8VWfI4l6qccwzr8Rqxc4JOc49bMD7Dd9VsFCbOu4oj2Z3PhXwF33W5D
fDuH+l3Ue6NGizBVkMZ0Xlo/JYXkDRwwPRkhsledhjgI0k1zYzBgNW22/yK/9ETN
cZOUhSh+UO0cOINEb7k47AG7FW7ADRIRnOD8ewl7DucYfnOURMuBHBvG6pIU0Uze
gUvZAtmg5lTDUObskT/zR0BRTpXpVoUDoCpFQ8Xj5DO/5i9EHJXmUlsYwSVI6tVi
SX2KIZKeVGKm34mg0OhThwVl+rKIZcqinuGoppbrHsC4e8eEfiQbPghIeomdxtD+
lHNTbcTIY/XcBFS9OuISg8wkxvSHkHciuYlgWoBT6jdlUltRiudfN/NKXBwQ0BoM
en0t5fF5PfuDyfFe/OQ4B56cfxTHwrtbk5OwLCpjsNMHJ0xsjrOPFP1cqEo3dB6t
m3gNs6KhBgnf8uH30pX7iPk0TTj8qg9tAkrSxMYF3W19IPHQRegRv7lRCANifMFI
/c8ySAiGGDfPIgtkQJGWps2zco7ch7p7uetdCruE/2ZjtkM9pk4I6yU3fAnfG76d
bolZv2+Mfw+H4+pdNU6fnwLBdMVVDNr26HWLimPCrp5dVChsq11rMeBXRm9uVFvl
XCKOltpqe2rpOyO6bSS8nqqTdzEuNEbah2l2IPPtg/7ZzvVRbQUX/bEvlpR1wyjj
5lVVKWUuWmfWjosJxpn/yhEzqCeHLAtUphPqvNllSKpjaEn7utPH4j0umP77waz0
/KC2S8E6Exlb8ptitSAvdvefoVdeZpPwNQL7JyCAoYvE+kg0NyhhephxbHvWJFCX
QLjEVgbXGjAJft1sipHBDVKnqsfLlCF7KWS/xtgUamZiXOuu3m3Vp8SKM5MqU0x6
Tr1U9CkkhE68z6y3fOsmqPdaX5XCtBRNmUoWvZn5wRUo7mlNLB5f2wJ74MuoIY2H
6jOnVjAJDEDIx6qpDGHdgh/13b4raXru1L1DkUbSmN7RFxFsmlfYjKm28yyIndXn
FjWdFyuFOix6cleiwu/c9cnsltzjnhJGNnOFIh8o5X59MP1k063KP6zRMjH6daSR
0ptRX8U7CjLlphrB2IAsvyYFb+b37gGve9FPh2oWfEZmRvOBtlhxHM5gKJA7Owan
eCNnEtrwmO8Co0xI2eGVz9ysxLJZrMYOO4RfME88chphv4w/YLFuk31CO+M/7zuw
RA3/eDk4zly0Uig0q7Igb+B4obUtlvhTTyCf/aIAbAwBlDtdS7REcXbY6LN4IRQo
gsOMxZDbeV6QwqvAzMm/xPkmoto/zZBaLvOEdcLehgK8MDbPXMoqc+TSdCG7ClWb
Rdyx5RKnVKu7VhGGX+tqkKAAG+frDG1hdCcLQ3MkEe4ecyLn0w/N/SIc50GufPBU
MVe+srocTuwnbq3ps1qqHxrLqQv+tOoZVZtrRbAHyp+8z5tD6DKwm2IM08uYfsxQ
iQGvZBls1tOHO7E1mpx4ISTmS9QDBPaTbsEhV1zn1GjD4mgGo3GDyyDS7MOUSZ9G
vb1yGuAXTRQ84dGXxuc6WMPfPH+ucWIOpI6UdonP6TNUtEX+I9JKmMsVZngX0Qo0
/A8cKZpKqeh45H6ScV7Rd5smJbdbbPQ5Bu3oLvEN4kmoIztbgsANkPMr3nCKL2t/
J9xNzoqxFVtiMfiF7Oo/73vfSaUYaIXBahbAvI7ROBmctvS3LUsuzVriuq+V/daC
tSr3VRSAPVLdp64ZDCDqenuFfNrOjlX6Ne7+i/sL+ptIgXpVtQCmYNxCXV7YIa1i
fMgdkj6uXGHx71KlZaKoU/d8LQUloy1ig/Bzbmy/iiYnGfMCeIVaHF5ELplkJAcj
kZ7OGmtAY/KdJ3TqrRnuaeyoL3OZXlG+m6scUZ8SgAzTZ+hyMxOSiXjuMse8tTLc
PNxBvEaY6aKfSttddcxim7Uoy5pSKOMEjKMDgBpwwXNOnI2jhfn3jrhLCJ6IRhm8
m3BkIq3c7ynHZVwRmQqrvXB/+4ypNL12wn77Mk7Tngomfa3NTusGoAq3nqm0angI
XR450i15Y/pO0hoNB/Hdz4YnGQsODYhdS+7yD0PBlc40b71/C+BSn7FUDbMYiNQg
TJvfP4+Wcx0qR1YPl4bxVCEd0+D2Uv4iebWHNOZhZBWho2kR7nlkgVyc/IZD95fh
U9NoaqoalvPdO5BPQEsHIanrmzdB8SauDvljqIUpSdVd1zbYTKoi1VUl1Apghky5
H0BJIZKvAFJQp7S+Ea1NVFGRnxQeAEJKqes79PctyJKGWF7DOG6c5Ci7gVyj/sXe
S7pH2CfyIYeTEAmMTxtG4dY6xYFp/pFYycdCUrwvMdcC4MqmkfOGjKBMaoQjwERS
aWUWCukjL61vZpr78IvDdou+euiNg2W0azf1HC64XgN6qDQjzoRfCLCc1FZqwZR3
LERP55BN7rlEJCX0m5a0hcWHPSC4rEokYDc7YAGijej4FKPyNZeK8ttUrkvmIaO7
RUfOFsHU5Mb1VE8QQIt0/jVUjtx1Fvjmwr/lhaGyWmN407qsuuW+Twef5K1QRg4e
suUxhB9CLb8Tr585HxvYvC6m4FBdeSzvJaffqPek0opLdhfrMr52ACIljf0+9yH3
ZT0+Eh0pA79cvz+RmdTTtIov2KvuWH931FswKzV+/iJwMAfg5ZJ3CDNJSDXHQcYF
umeUCzcpSXPrN31BciCz5s9+JdO1tqs8c0/7EN7w7sHP+N5UyiehN5+GB16hu6Qy
Jj1umlQK6pJo5nrrqYxKjGQ7eVeo+PgbB0ofBMnho7nzNs5mToDP/n7FqpdtwdiU
PnFdx+pXIS1y7vOgBQ5iXzQE1CArgB3Kzc3zd3VHVd1s1OpoVZ++b3vFWseLNDBR
pUwdpM2u4io66BEClntPrRdyXHDfUo5Y1pRRsCtCpg76kByrCCPdQ7PyM0qT2/VC
zUHJXV1yjLeV2WbF31kd7z3L0cgYpIwU+UpOEhwoRbSR7xvw46rhnC4qenw9OGdI
Vo01zZGLkfFvIWCpGV86Fw5PRwgPWMVwNZvOOwsEhzl3d7skm29ck+pfBwyMwPJB
GQNiRTb3Ec7yNHa38hzCtGBwF2ral8hPhUnpZb76FHc0AtZZGLN7tWjoTt8KGclt
6Yl4ZShxI0m14gU9edOLT34OpNEsal6wUANWNMKQp+IC/7AiAUVlSWSB3bq+gBx/
BEH8f6BnmjabvhJXywph2YEEwJSecdoKHXykrS226HAqT2CtUcl87yWlQov0LXYF
ducROYKlvVUS5vfzv5KeNk8RBdAgAZx+rRuU7jowfdIpigfB3u3GPwYTswBfrWAW
ZNb2koY3P5Za2FNkuLuiRUOLyVfyoF9Y+7jWime4LZya4HOcmqOyYaEGjYmqUeoP
eYHrombmhiNQq1Ryp2HXMaq41PWnQi2aD6y/XQcZYCz+XfnPflXrtStl4coLgADJ
l6++NWk/5+9AEbek85PN/VwJmnMjIrqdlV43NDrV9Du4oq4L80ZFcCAfwcO18d7X
JYFTrnasbwaD0DdTqU7B0GpuB0D1TjpCTP8R4OKpHWpvh2vziD6nMwxxdo6IyMPv
3euRFjMDJMuB5+0ykGUpcMJrVsP06ZWMcld8izF5IP67YT846jBIGnr9B+oX+zPR
kTbciErWJ46SuMNqqr08W9CCtN7L/g5LaSnxOE6caTDjNzxOLfuPnicNxyg7f74G
Pfc8HgPIoaG8lRsY0mdWjDwWDWI2J//7KlIVk+3z8nYTWOPMydiKzRLrgc5fer6R
HKZ4FOHw1kDghzAz5IdfatxS7cTWwsugkwAmtWB7ltL0fPKscP5JpiWS5vmN/IJS
kLlx4Y9RhONXd6Qh6ER3GauGbrAAdYjTKmJDBokuDp4WPXwbWyxjsud6V/ztl9PS
5ta5z1n4YgVONUSH0xDWfhAzqyQTa6K7h88igTI5WlT7x1SQe/n/1RZjMeDWNYeR
6sZ7XKTjO5xaZFt7zcSQbrHHLrNQvgC6l4yNcmeOMvzvqW4Bc3tQIJYHo3jBsYQQ
qG+e2F1RAq5C9PJO44LP4fg5EmtLqOZGNBELpM75oImnXBeHNluNeuy29yrZoK/M
mXjWUpygSubKC68oDd4DUlp10IAKPZ4r56O4CjAHyL9pYht3atunofoearuBeToM
ZHBh800ZHsrPGvVbEcDsTtjWtom+djAIV9HbqjkvasLLvmi+qq69PfxvUJlXLqlf
5MslcQLCdeqv/i+RUZD9kCYa7LWHh4qO+0ONaTnA054TZWu4qOXuojC5Zjr/RLXw
ueSwKiY1+ZbB2ueiDg3DKuC+aXWfLU85oDm6xrSrOQPHxhfLfnwSRqk5nxHIamEq
TyyEsAj4450EJ7BxPdilW8vkx/Zs5vAikF/dGNr1R32kzYMojx/DRLD3aPYWjPS4
gNi8NL4OzhqxD8kEgRUPz291MoUF2u0RmW6OH8EJop5eCpZcBNDFUwFPNv/Zk6hM
0UH6MZcEdP+7RzyuVAO6RvXla26xO7nH1vZs+/U/aRJc+Yo9SyAY0mMiPgkur/hF
QtgP0ZudzogdQuLC9KWQsQXimIbByLbRfx9Yw5GRo0aprIlPEiQ/P+yR38JAudpz
1NlOLJ9NJZP2v3gEXeCVOFGflWYABWV1goygm6wnhVl9FRciV1DtM/1ndSfTTkIy
SfnNOQuUZPEPLQvupJvCCnXx0BSTNlKsT2ymedEVtERV3pAizTXsIr9SEpVa5/hZ
CMtnRkwcIZIsWJ42I1Npm3tAT9GY9OBcQ9AtQZbUiVsk7vaq3wgLC+5YB6dfmafb
NzAJ17iDdjIbEnYBBa7ke69V+UFdgAbu4b3940DoCLhHdycHlNQ3C8/pYQJkwK/T
nCyX0vo4PFqYiIQbK7jpqhXy5LnChk3oBMB73GdfBGSfY5Bez10a3RX+SE2No8gs
1ul0JP4DW/XkCEsYvWtSO8VIdg49mcr4i4T3ZNnAXgAUnm2ZOT8qGypkzg470FAI
Ys/vLqq7ladMmp3n6fHvVnOs2rpkc5mhbsmax/ZVYAcat6So/OYhylhTmq0xsmeb
8WJcTfA5iCesR/+LGJ+0XNDJKUAb8A5gDzVCwE4kXkJbWGqh1r8x/IB+XGMO1e7c
gSLn3FsGukpiDmov6FtIQuMX5UjS0/OaH7hhUN384wBnMgicPh4+qnTiHu5ICe5f
+ma3pMxjQofL7/fDeijTsSimHuoPZN9VvIrfkDaLmymGtlhteYsLANd3SsSZZDlT
2olkHrxp4PLG6tUWvXssQWv7OGTUD+l+Z4pf6YYEOgI2v15y9hfaWUhC0JQ9YNEI
BMKMziK/jB48Y9u0rg4L0SK4JVIVWmsXReWbR6jlPeImfa6RNGvPAwcC8oR7iqQ1
/8SuJDZodwK9dPa+KZM3CpsyGp9AJFgoh1kwkS8HuyvUdgivZTpZqDyKXGpamkZg
KOHsLO1fsuK5cTQM6CwmUhkvQFOIqpRc/xqouhwQHFJSlQgCVjsVVBUhze7+5AgF
smMGAEeWm1JqvySuDp0iW3RFZdY1c93D9xuJkZ0MCo6dK96/ZaWHuv18WINwlZzn
az9E2qhI//jVA2o5I9dOglja/Bf2K3etxnja59fZwkGdzhP07YhySvKaeSLVMtbW
eoX3t5B+xik3ULL8odkI1iJ++h6CbjtL/GxR1irNbyPZSaOINCYBGD2RZ+HPT2uj
y1eDjt/jE/Hh47seiPPyEIPtKI8ZAWswHIC0SO9BICWxAkd19eSMATh1EUUMg1NX
RQPfAwYBqnz6SFyrc8Q38QWFCfQJNxjnaqKCGbvx56lVyb6j9EPcG7cd+x9sujrV
en8u7xtp7YfDRhIS26G8+qBEvq55rDvuUZmRbtynTPDWpKyY2WhtKFU5DG9vX8qn
GQ3eoOF0vwhYQV2hrd1AgapYtZpnlIHaUz9ptObgPwOZN6fk9xic7eYcv0wkXws7
exv4iEet95v9w7Vr023e/89PAG6AmlB57MG760NoHtT55XpySWeTV28cNWO9zdvP
Ne5GBkIxCxsNlJgjl/0t2f7G3+YIUyNLjytS3AuyX+ZGnAHYRPF6speRYgQN5/bt
nCJE6SHkuNT79kGE8r4BolbjEGztNztFT3630aadtjbi/jBcjj9AQKe4qazW1AoG
ywOVIOD/BZ8AHbU7+h+4BPA383/ZdHFTMoz9UVns3MRurzZtxcKcx3OziQNZWENK
t5vEAIRm4ZG5WgX4hv/xUQpGxKhyfdBE9zTFGJJLnZR7bg/Zdoz3+CYOfFZ2BAXd
j3amig1vOYBD1+nLeE6AusN6anv+obM9Vmep3d9cpJI0lnfxlpipgmPrOIR2j38h
UcZXcX2YAGZRivhJNY988feeQTy0I4lSJGm2HPYgQ46HMUta5IgBjOHmM2aRbPrQ
LKU2Zq0PZb9jdLYDNtXuUTMzS+AOLoTHaB+5SCrJio3BWrMkZA2jdhP248//10sR
OxOFgR+twWD1RG4PQ323vFQxiaz6Wa0ssBqo+sABUZReQ9c0kuX8UImY/0c6700G
WkVYx3YYq8Pkwjh/Qn32xMcMvzX5L6Tj5CTO+JJgJgIIVikhSFMZ+whoDat9spRy
PHBNkz7BSoUKvbA5DA7xZ8LTnAiwLoI4LyaVXoxn8ahMUkAl9KqXs5HPGBlI1NK7
5JtBtFz26MEokyISVZ3fU8Q/zmElu7UzdLeAMPLhd0e9wDq7+mDoNKNghGL8r8Xe
KGomWjzKawm77/mWWMjA0xuwHAQusGCQScVQL9bzqKXlefOxxQ7QJXUm1+i9mK9Y
O5g3EOnW4QR6POzV0/J4D2TTNtoSl71Ycvt+fZBWeRvh+Iep0751H8Dn/3RQBpW6
L9yhlyebm8gB0CeSP2jznrQAFIQLrNBKSW5+lMOGsUaY6W/JMiEvvbnpTDSAtWl9
2tF+eyPMxKTrihVuQUduYOJbkSFj1Y6R7/fWpeknxX+VWuYv9HavYO6HaIoIFSH1
CZZPjDYZ/VAW03sqi9EubTrhcTPlTN6hOEUQH1YO/duElY4vXvx1rqzSI05OBgsW
QeoOaLInUgoJl6NUPKDspicHseRx0RDdP55DZslrzZpZdOjYpvI58yUSdTvQYTAG
dM2aBlLldO2uqCZJakfxOBetjM1PSNp9WGY9ub+OBBJOu0zf4RLFCU0jjtv8dGSL
sTJcvkimcO17crzINYdbYspcob91V2lbOEuLfUUt53hzFyDZe9cwQwgYkCgO8Cjt
HMuB0a8W6pecBebuDhWLOULOwZEccsxOhoAHOgwVzOCnhpgwOFmFRMXGkS7yrG4y
JRWVBAywTPSO6iZzjscTpyY/ATrGHy9BPyJ1iyin6WGbiY2ilpbQJvQBJYhLOyGn
S8MemWUtoStaUAPTDK0Fj/ak+dlfPJgX6kJfsVYBhKbtepY+3fgagJ5GDm9yU8HP
AbR3ghtW8QAjQARndH5Njj2NykPZGO5WZT8JtFE2Eta+hsKCc5QnRSfyWO0D+pAh
BEf9A4N0vdKHRdxf0IwreJRxg1YafNuio+/o8w7ipGrjLmze+VZxLghIg/v+/XrW
BfOmHmzQ51185xLKukBJoyGyLa9SZtej67D1XAfdwn5Ff7G3atbucL9HbsGZi4tR
EMxbgTRXx1/m+l8ceOGCni2jj9GyXHlYhjCt1ay2Gigr9n1O3zOwR4rrFtHAyU6a
OCud9HTTazLD/fqnUxA2gcTnBSdmNQomHId3Ipk6fH095v0RtwlZ6lv0PImuRjfd
U/uWKEtu1Wc3vh3gN6HOAYHtdulRJAsrsgac8lV7L+9rfgVPhduhiLbH+CpqP/zR
vshE0qLlK+kJm13TXbtdoEcK3nEtC6Hi09xFER3deGji/61dGs702xY2qH8p6fEA
L+2Rm8idFB0sL4MCvWugv0kpHP5TLKeEzVOhiVS0/CuofCuA5g/xCMN7PDKVWdaM
Q7PUl7OIIXPaj+i5VbVMPDQfZSqyYRgs9YviXJExPeHOZVgBMYgGEIi1PMO6C1bW
7Q+Ha0ssH2VGFUgYD/3qATmDhMfprfojeaIW2feYw9BVlFcneJ2lCn4cWFC5YNqM
5eym5X3lNX9mhaQGHln6ZzaCLjvyI0GP6ovgWIUKOwMvcqzrdxHKsKT4yoJTIMrm
ct2kmCWNaTr9vm1Wxz0aCoJYuu3R5IDfT+BF/qzzFCaAY/mJs0Ec/hh33nF6YyJx
pCT0E2B21OlXmlmJFEhHmEXNNZdttjFyMNKdYBxeVV7PPU1t53rWYzVWKlZiQRR0
O1WbgHczwv6Ox6KqrpiN8d7cEh6IGCjuz0Ue5Dy0tjJk1hjHuge88D09VBOh/r4Y
Yntw8cpTvPFhQCsJmKrLh9CKuMK2KjICB/F2CJVNAkiVo8gF+wJZNtpQ14+FhQCp
3I7/eAi+6UIwEWVKN+xHfrPcjz9LBO9sIE+Of2U7XPSI80TCJLXIkFoZR/TD4uAi
KoV97881/jqwxdqt3EDljchkmAWGSKWOWrTdFMMLdqcOsrZ9G2PXhr9B1r5tvCCB
0x3kUXdz130Hsx/26Xywr34hfhk8gF6F7PKAdzJo121wTegs56ij/br6XL35UJYo
4aXLnT4G5V8t83UHQeicVZt12P586FaugrINmW76J354+WoNFHuWmOhQhIXyZq21
+txTkK+hGD/gWbh9wW5OcFkPifTEvGzA9p5DkVNsvElTtEF4SHaUXoxRbeWMJLct
R2IopkuTKVDtBEl5IEKTzBet9p4n3agdgdJa3s4tUl5CTfy0ueJuVlDAbX69CPI8
5YBUKNLRQy0ZdzjN6klW2MsqkCI/qkSIkcNTSyLvWQvE5JD3wyecGBO0ZZN0pqzV
qRB7YYcBLaqL8WURbr9U4hs9MZX8WOHf1LXy1FpmrZQvfCjrb6jqrO/9t/sapf4m
jS+RitoQO+xEkwOyodRZjhVon8eqXrzYrsTcyOkjvzHZ2u3624hEqFbdISK1tb/M
jlySkQsHbC7Sixmdz+3L9NRQaugI281pNOv2XSh6xDnsPvOHAu09ukaUoDPOT8gY
euoyjlqq1cVHhy3wTA4veKu+5h2RBXTEES1Sv8GKi9Jl8MLRPU29XUGQAs0zK/WK
K8w+3J3erh9I0GrmNY4+T3w4BZDcCypRvyhWwa5ocwOhENLWuhLs5FpQZiTuHU6O
lkVaOq79+tNdwpnv7hU2p9Xv06J5wxRub+ag2vYz0JxyvF7BognlpvCFsVGTMIo7
vAy/BUcC/LJET3fUER0wD6QpF2AXtikvsBmuBKoDVvtRM+BHWkrtMRpV9UZVe7e6
459/AubPMjrKFRixT34Uc+A3tYm1sOUwnnPLxvDZA2h90f/60ENuEnO7A5J0jRNo
+1ULknnjPzHrrT4tQSxWPQzxpglm4vGVbvuxXmXq2lAJ1uToJeSN74MHxnzXbBV+
HGgD1+TnjKtnOfdX0pF6QfJGK0YRfjJVwQeOzTuQbKUP50iTFFG5tH54W/Xbx48P
oUOpp/EZccvdz6lEGuvb7dzwwUdjeR3LjnwRyvdGct5Bol2h9n5YVEa531w27BIF
saXBz1zA+OnAjyQGkMni/cYYHsC569etXkeEikUTYASnFXVWkA1yedHCTk5gJXtI
K05fHOYQbwNReT1bP+mITlI7/4CwhYBArKw9xObuoAyhnfY5MWna4iaPTq9+ifDz
MOmow9ypn30vxbJDnkRmteZPko6EOadPDl9dnPY1SUxvR85RiKIn2j8ZqlM8EvzY
FMoeEzKMa7ipXqLvSZsV/4QpyaguyuiAV/iJDqNx16LgfflJRz8IsHUd5Dn6Adxq
m3uj82vKmroBuyOD0DpQge9Zi+G2PS/HwkRCCaILJNfYQUs4JYEJ8yvHe9T9rHPy
JkZVFNWNOjJIG/25hccVAt4Ox6dZiMjzsQo4p6sr3BSK5dpC7Nds5qiLUIzJehhX
8wLEOe6r0s0wgl6jdIJ1VgS/bfqh+K+TFyyFY2VEKK60bk62ovC3dq1fpI35sGOa
X9lsTG2pWrtEr638frRpkq2Eu7ZnGarDQco3BVMHC218ProeI5vJJreXgTSWlSzm
QsNy4x5VlSQIIFKCPGEXSQWcPhhLLB26O9KG3nn9ezUhpqHoNK1mcVLjcXPrYLWy
cGwf/KytGdKgPECoqFCMhvz1Ya+h12sTmp1Vpcvj+cF6Au8BWxrlsLrHX1kyH/tc
4a4vdIhjdrnZ/xLy2vLGXT0kqmxX65nphf8OMGQqmcYN4R0VW6X5ERprKJhSZiUM
Jg1V6BtgE71IqHWMktz9+bRUPaPAljPMWEo04PmQC858tP4kDu02M3Q8VbfWxZ0a
qKXaKJ/6ARVXlM0kH6W3mS2YHEcSRZPdlGbTjPapK/u817HGPZNQpRw8LTv0mT1/
O8P8ZyfO7Mmwxm7lUocSucbijkGu+NbG9NXM8CknWKob8mh1In6QzO6fMGPAvR62
JhuFrLn9zLGpR41DCp7Gt85ymShhTr2Kdxqt+ydDl323Bu69UTh6bzMEd9XIs7k+
tQxfnaXAlrEMZphyWjAQG28jtQFwFyK76rQ3HEsQatJbZ0nRb3SmonYbcFdlUjhW
KEHKMSYD5z0lKpgxFtqHZ+l0P+XNuxq9ub5/FdeiCrSrIs9LQ8dIG5f5vVIswlkQ
8JDkC6pEa5nU3oEYBnBoY6OEOWSpODQaDv/cpOwbYr60FiOQZ7KhQfdaMMwb5b+z
HdxQEvrcNwnN0Z/V/wyr87MyM97h6FbwCg9LA1lfoWYSMfsY6iXCCOJWSE/YjPwj
X0mZTRgQARsA7IvrmWdbf8fX7QpTf9LXJJehcBiy4iJ8u4IVSPhYfZr3hak7yh18
2YXOejAwfEcRa6FnOTF91W20BcSyiQkWcvP9QGWyYk6ketVBzDRwnj7l6h3QYVW2
0pyeiPvvQkWAchlPiv5bOCNnWlxJJXTyiG0lZbmG7+T82v4VtEFxoVK0iTy2jqMF
bpfWMa9nHe2XGY5XWPkYtcmt1VT02miITjLrNpOxIdT0zL4SeoJ8yhCFlg8Fgxdd
7DL+63GuK0L2bQ3k3ERFdHCSzsVTPmy5pBAEHlh3z2dzUwVLqFCQn0WlafP3Kpjt
Qg3Vu69h2z3+jNyAcy6MwosedahRERxwLCdmj1MyvQtRaDs2MLaKtvHOPZpS6Woq
GOM+YgchKyZX4JknU605pczv8n1v/GvlHkeO9F57OrK0W0JphRzkgjJGs9z3iPzS
BJhgvniQJk5bNP0z5vql/85sRitqb+kdt0HkvF54GeMJH8pJsTbqyV02HTZHiapd
fMwnjwaBMhEBnOPuw57vYlGnjepe6tlWjwuj8aApx4fMET8xSrguxGpkH3aSTlt8
yBJzIRlnApksT1wLOROoCpTeYy50EDYJxhKgkTAyNcktNCdhsktBr1bEKeD7AE78
LEFFqa5ENyI3BFb5/xzxXxp2pTUjBW5bWTRsMNOtv+pBEiwwW+PPqIrRTsuE0D+h
ZErK4h+v6cgNlyxL3MPzsfCLK7Mldyuno9u/9FgO4G5zmVOFBvlLpmfvytwPrsf2
p/T0QqMzq+X2eIovGstz+pR61OuTvyCP+5a6tW0FsUQ51PJYeDip40ayL6YsywDw
a5A28hHyhlkYudXTP8TjrEryK0jIRqrHaut7o73gytDCEGEcGsupL3Rng+HVYhKf
7UYXyo6t0UjYJsPLwCRmbIWAA7HokWe281mdKTEI/5jrwDK2QBO+r1xiqdAVKqAn
VYJ6BtyRJ6Um4xGepscJ/iojmdwHgTiUv+C6pbgh/krJE/w7p8QdYJJaBoTnK6hE
XxzAVyYczglS0EuohWdR45Ei7Hf/Bd9XkccyfE/WjSJASSXWR4adkh5+c6B5BOwO
bbMui7aH+Sm7sjjQGi/I2PDMMm2Z7IOgVZmYq9UDhB/wjXxdSP9J3GzPm39dCVtz
42WN8mFZDWyJt2NjXQVax+VHdvKzSI9y6antMxx4OaRfQTphx4ZZMlQMDGB9Bo/C
uKRBUP42DBLwgGoDQhrD9Xd16uarNjdkfVKdyUEPmCAPAp+fqqbawlZJg9qkb7QT
ggTqu8OZNr6eVIctK7JRmdKjcuazYHH7sePk+6W6GKUN8Fbrs2/vybBRgVGNIC1I
ZGJ+WidwYrJs9jGy0ELksFZnvt29/zQfArwYO5eQ+LZYyms1VzkwoiJ13tPesfkw
fC72ANxM12mqPQmOzgEqNhzCg8YBTthqepPTG0f2vgYdQJd9icRsy/Nkpx59vcCu
kFgsq6+k8MByHLNcaFr9r5m9VE/3GKCQn1h/P2FFIP0mDSbobcFj5h8rr512oTE6
F00/aHlYCwixG8aRl4K8vnEjr7tecTdn9xH6nZiu+gQ7tWuFuRYiOxzsWT1ehpzM
wz+NlLULSnxZIGB82E+4uLsVlDUx19MaZsz/lzLaqs5lFpcO8dbfeQdUBkF50TMf
BgKxDFgagDDPfVGBc89ApKebFpc0G/tqzRRz+D/XHSvrcFshm/cRupinsXH4X/v5
8+STyDvtMUJx8sRbdloCwjWaopWLsF05swDrsGTkZcrBWv0Z0LwmY61WDCHaUI5V
nMw+HcC655dbedswDH0TnVLG2Y5U6kK94IC5P11TdGqX/jI7vwdbOq8VOBwuRUen
YDSy+HVzY/mSfho4M9CdDxVHE0zNoYNp7vXUqk716ybi/9nbtcdqS6J8tbp9cCSL
8YbZTxVR8A7UG4zPjMZEoNGB+IUqZIwt8nXjYRjRvE+6IDMSkh8z7JgELIcWMR3o
X1zdFXA+jqz9dVriow1W3hbc1mPHSqng6Xr5EsH+KkFI6ySIlBbu9zexmzMCyim7
kctxL85GmSEPbpbkYskcMOWwdWKeeamg+8dp2ByDFLMctaeTEqGlGzpHdDt3Rn4I
MbC0eq8CKE4dHjxqxlfdTDzsvDIUTLduYv2hrzfik7g7SsY7y6BJoKw4G/ndeWfW
ZC+E+Mx2QBJBEni+SKVyqlUnkyitZFK9nlorPV5NnR/cUGKjW9TueErtWTpOFt/L
Hxwa6PAvkOekibi7ctiBbcknquuTWah0JHcN4a5Mx5H6uOQp+M4yKGIaBHNCdlY4
cHkMSjAB3fMRZkeHun//m41nZiWq/uPCYZvzT5MndBzsj95MqbvPRFZrmv3Cyh8n
H19AiRKV3w/OQpTnJDreELKdTDwRBFd7LUzl8ImEVmY42AL19UX6snkDnpGxz0KR
7Rxr9EU9rgD+Ma9POFzkmupIuEgTfdzxdcM1VDrICvPyQluE1Cfwp64lCX38Yjbf
klj44Cuy7Z8ImMjpIs9WoEgWWPIGveVIN5b1/tVMbJA/XX4aj2ZtwH4ojlhExWj2
nDBxvs3rUEgQvpmV3pMuXT90GyVgWWu8ltpZr2zmIj3+lCNpLljNg5P+TzofQcOv
ubBBNI/mu15xsq2o8ME8q4a6OK7rvyXBgGFtZXjd33oDEi3E+khPsMOKWr1lRhqS
Y1TmgidxErDRhm0E5banN7jSQDHmlAmsX9gcrzbxdmIUlYo03IRvA05Mqcx5xE/N
p/CVkXFoeETVYr9Mex6JFjg+tEn1bu8f9ovDmZz1wTEbxA3oTbGqApi/eFSQT5uH
Ld0OvFmHGtxi8DHtog0UlTFVpKUfksns3F/prHBZGMG4CeAhMFzHYCNZIrF/0X1c
P7q3+R5uyLxBqoMytw2KHiapQJRXCGMtvH0PBn57J7JjVVXDPeUu6yR/mLPaaudZ
T+aMsPj1uOT1zPcb0ymoY4OwSjtVWBoFUlH6GA8Il3dHdFKxms6BWP09udOF2I/d
w74SmNkwC8q6dhPCtd0quTXwEjhmFOxuRFqFSwEXMAfp8C2qUJl3B+sYbFYWga0t
sCCZwfwzXnhf0wAadiXO6No1yKbNp6PZl3kRNCouKNhbbma7seCowp1a3M7ER48r
QbDUuRYrC8EqEneiacEzsJro8XKpFZlV8lkT5JL7IifHZrzqYVodYwAy01atncXH
eqXp6zxuWSwOmf4nPMMqCvzV1qXbcyq1u9SwkRhLyWplBPjoAEmSAxHOrhw6iHQ0
pO2uKzoSXAABsx3GTen/Bc68z/1GoQxPp+VSA7rHW44mrqBo6Oa3GUQtmGe9BxCq
5oy83QJAJ3nGUhjAClKYvy3gzlCSGudWQbc9g5oTofS08MpVJX61z12+ykY1F1h0
F4DMyC2uOABjQYd9e/ZgF+/I5GKiE65moZPQaguGA1smDTYM26LZcznzwctBIKp0
PnkXM4z7K5ngL3nidYEAXHI9JVdVfUUgqlbRt484hTk+p5Z7nV5FjSRB6Cwr6vCV
2qGkKqYqpkzgt74V3Y8iV6b/eN5YVzJyJaNSzSifyjIehScJRpkYmCmcakTSQVlQ
qOK31V7hRlqy2HmdzY/OdGHcfe0sUMMgEWxOJLu/HsGNjIlD+rMDvbfEwPUJePpe
TyTYRprn5zbgD+8GWCZb7xWlBgWb7U7WZ7n4nAbMmSaKbGrUkuKS8qYYihDC1D5V
Bsu3ylML9UYxw7Olnp4lhSG7KjtjrngHbkLjE2nOLS+9itlkH6M+FNCK6RZiHsEq
aH1uRNQJuuncHTsS46NTNrHqWsQjt1D5ySo8+MTgV/uGb8YIwQIjh1JANoZRYlz7
1pR+K3ask1EMZkVilmn+ltc3G+KPhQxKWCcDIH0FUDTw8fYWHnfmqV51y2uCr3IH
6HhsghIfQExPWGaGiH/utb85cquAy6ntK8PxBuOSH+Z/UUXOEDlfvH/3Sx+4sbJi
diJbFEb7BAbiykaS7SFWKX/XTuCdAGAzKu9OvC3GrhBU6MqR1YeDfuZP9KIFOHBy
R8QkCa4+H/6g/9R4+aZV8R2PPpOTLnPkiLJTl4wwdHWi2XkCX0WVCXSaAocPGi/5
GCWkkNMdRdcyDwcfIwnNApPRGHkcroaljvILo2S2mKeZALS9DsRgvL3fNdKzp6HR
TmOtqKrOSbfWVVy6o+e/w5VoF7Gtpzd34LoReV4+SQaI90bQNhhw8v/bVskj1yFO
OVmwsrGN4EPGKs13mJeva0RfCK4f6VyLi3PqGwfufEQU/exydTIMjYB0C4ajnihk
BOgem8EV/LpdslYlcbsWoqT/WCGrFOwoXd1uKLFgZXdsa5eCUG3FHrQo7CLYHPv4
LC5+RQAzQHs45Jqfqjb2kyvhwVBTmdElXGEprO7O72jQCfQKypaF4WlLfNagGBH/
NoR2ji3hZt9IQylf54figBImJ9/oSh7jjvJ29k/mbvn1Ub7L8195mm0U3vmIAH7t
MJ1QO/p27dKSp75HUk+KdhmEs+VwIq1+q8KTyYuQFPDlkM2ozA4faxKt3m8NMH1i
EN7q4LOI3XTcRHDDXn4PfBJH26FaMvw12fQ1RgIV69fPk3WuA4Iw7kAh6Bo4r0ns
AnwNShNpUYbQZW2p5RHnqguJlH0Qg++c9MzGjVxJ9iJ3MRBXC2Npd8zK01NLaaP2
eYCaaijRi4bT3hmInQetTTFUG/f0WMJqn6olaLhM9u8xUs2hKS8dSNcapBfDu8f7
J+MVd6qiAA0jF3atfKe0yXq7UjMSDeoverYxWAzKg4u5g7WHGZ1ifcJrlokOUBbm
bkqeZw/FR3EoPaMNbKiqxtQLH1qeXxzCLgQIpsXwDToqEcYYaR80ZLijFfw1ZOEP
wIrhagEkXw6ZPfjYojmqRsE4Fz71BmR7FUMqG786U9xdXbBd0AgbwLGtYzzHIvxk
sQAMBvLI8D6FmYvm2NXdjYACx3Z9VfM0OE1t2F1J8qqJWYyH0yiWVFbokkk9Bldu
vRDSTTq8ZQ4b2u7ueGPjj2d81BUYfy2P3QsOjenY7aX4AAOc0TD9cvdPa5Vx+EI9
wCkKGFw3GFVNBTB3DYt3p5at1yhwRw/vo650s//i8UjAQ7qnPJp6ghVwYCOjD1Ay
ggl5fYcqQwbnb7fpy+49JLoohB6KYA4kmZ4VX/5YNVC4f5RTV+ersj8i8kfmlptJ
3OORv2I1rsfDx6OxwAIqM8L3k6SkODH8sCoFiFWQJgkdZuXEF0RfjpmLU59A7yzj
2BimmPmgUM1yzcWsUTmWJ4WZWWt7MQOxJUiuqdwKsaGsM1Dmn79az0F6Z1iRUsm+
k93cS1DMbNC6pDiAon5+j+HqJ48vfWyTzN00LET+a3lt/xaeEeP1TysZeUFLXLmW
46w8o1AsFedxtr2SgYJ85VblzlhzU/jHmUOrtIdQe2yN/eCNjAmbUbMzBGxKyhmv
exbWjqWAnYvZmHKpJ97BL4DLT8zfjSH2MI75rZzkOczkIHQBp2b7/bdbcmmk51IS
QDlU3lJWOc1SqEIIpR1+8bd3C/jkoLWT4vzrv+PlYP/1Dsz+tFjZkJO/Fr8fhG2+
gr45DDrNCp2NDUkKGhLaSduNg5JPZj0OIQH3HuVef+qXnAMJUcionNjWiMRiq2HN
9HWu+5f+v5f+z/qLIc5S+8R2NpEc8snMk4KvjmUT7vqCo2O5w+YLgWs6nGGjQD/a
2WDpgJY7QS2xhkd4NnfLDWQZwzEBkb56teJ5616UeJ+rBRd/QLM81YUjZEjcpnBk
RL7woGbfa4PH6B6MSoM3btrxvXC0px9w2f1Q633Bj9yYZLz52IIgMnQGZqEEEcYA
Y9turIE7Pegd/b9elBPL3wnG+Cka5W3R7MAcOcZ1d/l7W4f+Fa7Itq50aEpjNGbO
LvwZwPuCurvzHYlSuDQbRXCdQg95XzW3+MvtoQDrVWlaD8kW2FQOPG1ifCLaOHa6
sqLrSRCKi7h/BpulvXQ1LHY2biwXQyv+UB8vvYjczAn+sL9BzHcQ0SRCNCka9ZNy
TdV+3XDBMBjLq/1NxtsANWtBEYb/OM4+z0ZnI9MrbQxcDF1C5bpO3QtUcFGc0QvO
zJgRkDf5yN8nF0ggvw2OV7Bhvb9nXiOkAdnBKRiwcs0KC5CY4fwbak7GLf+JzNVb
jOqGwisIF2MJ6lsP06gIKLwSjrbrm+KhWjwR112UtibHTYQmo6uPXuJNyk60ozxH
boPhxR+gXfcj/hIZ7pjbcxSWZECDUoUtUIYJryVjc7Nkcgbda8m90qqR/+j9xvWh
CAj5ODJhHva1JD7y6Wzp/Fd/jZQVRNI6Sb38USRjjh4Og7GOTibs+ocA8aJH7Ibu
auu1A0eRIyvu+FgdPVJy8vc78tttQW/1+DovdJOmgePGKN1RiwPSjHGJZNjED5Wx
47vYeGBf8dYs1h4daV2d/c4C5iwI/RMNTBC165qONoKQ4WXegNw/HZ7NWZ53FY1d
okLtwixzuBrssr0V7zyHK612FHkgDePwcjniJQnbB+CmmcagBTwi4YS30IM9MZ13
a+K2UJfVrDVEDktoaXjub+wx9mITpeza3kfMf/O65Op3KNjL2lqCbsUGd5tnQ95D
DvxLkzpt7koYO6yW4yGsrjSPZnTdnzpjaAVAVHVqqYyR3z6dGURJo4lpP4SiIHCU
h+qckAKBag3dykOPRYRq9IjQ+6DgkMd/EaW7axdK6B0OiBwk97+sVgirv0gAALlC
W18tdxsqpcUYCofrOq183ksmh7ay8a9bwOuAWTgr9dANaZwaRcOBwZE6/j2Luz1q
pJaj477skKg0KrBUdDFlRoKFJCN/s5nDleXaGebEG/AGTtmz1Qdvv5Rk2Pmk9/Eb
Ts3otZlZX2Fb9GmkiD39DfeWo7E4hWXmGGqOPkw2Vurc8Sh+d4bsPNN+pHP7mw8t
DNlCOlFQYwktZuR8Y5Vd71R1pzE6KUsqhjuNJzosx6EA99tzi9G1Oq7GSlGB5bS4
LIIeQYURH2cNAqvApjH9wORfOpOT9S+N9mKSFCrZhO1m+Q1M5m4qi61j8B11H+oY
t+CYIoAZtNWUUVrT/dSceVvqDF089q4xLyZS+55Na910U434Y58t9GbKk6bEkK2M
a1h/n+AlPQTMCYr9i78s8fVYSpqbbcfipytLAI1ZVv8osxm31DqboBM4Byb5dMTU
5liWwesNRSJBP+5jnPn0u6HUE650AXa0SVtTdn9RPFkaf5pvwvW1aVtwmo9KZbLP
YfV1PosjBZC/GUWd85du99XgPXLwmfGyyF7mnLVwd24msOldOZylSu83w1V+SAhF
5YIKqFv5xCp9fRQviCNOgMoNa7O/3Ghiq1Gwo9x2LmGOIwFS1aDTWCz7wGeGU5Ou
Ry4jcKjyMNx1DkwKP5aRwYOOvx8E3f8e8T/Bgk2YdWAhRMpC2IzQ4qnes0sxbCoL
Q2MdBdOAX6hlhyux43BsIMtvusEi0oeQRCr6vTLg+0leuWNvCfkpueeBH7VXhvlR
b17FM6v9ZmVuIVcym3lkz/F5RoEEvNvC/g8qanzt+rd8KWhGKxZAfaBvE5LY+qQO
P7tf7lxNOr+5xuzVRTI+8lU0BwJeHccQeotYMrHozx3wfKiW3N32RojnWfq7Wber
e/c4qWZYM56svyrF3TIk0cZwgcg6SizafnVbhV/aKOUAdlh+8iWHkkeQrbkEc3vi
CHO77DzmhPneJNoCyZ9vW9J9E0J86AsIvb17GibT1m4Iav9hdQopUjKZBDI7poXG
SrXTANDSFRMsOKeQHwVELto6sqEaf4UJUw+Bqh+Zb9f1J0AhxiwPfQ2Coo5CKxg5
GyxIR8f6xblh6ZvdnVWB2Zc5QTKJVn04cRh6XOB/OHjF5n5/2fM+d31mgaNZhnD3
4Zuhysxz7bc0VUojPN3XYl6xvcYz/2HaozNGZEsX9asPjyQnOsdYD0Bst2hj/MJv
jty9tLYpJUMd/2jyo6sFSKbH54pQvdUUi5qpGkkiDd/gzvUX59fOULsuRuSVjSt7
ee8dAC+Y9GViuyZGAQxbGBjoE0anhwpvZINdFiY15Z5xukvYVJiHYPaB5m6E5NEl
mXTUIk4pB8Zc0w+VO0eVkxS/Vq+1oF6ABgzRO57+VCV+QvnAA+cHVA/5YPkkRe7/
rB38f30y1clV8PRBXs8q1a/+cOlgDoaAbU22iEfyZIZTDKUJVUA9JZKZaLnIT9Gk
k1yID2HUQ7mx/j3X6faBleCnx9qyqSCWFX0Lw2BKHolmV9bN4Xeu5Jsfi0NZiFD3
PuFSHuroKp4D5dGhxxji+NpiuM10WMWuSD0HS4rmN4nuIOH5WC7p6cgXZEvXCLt+
rVYEFmoDt19PZDKd7CeszCifw+dEqsCAknIEKJmuyIW342U8zgmmFs0bW1Rn2tgU
H9+8CWT0YhkYyYgtkmw6K9K36H2LpVX4P5Nb9HCAhsVwEYyEIbUkVoJqv86dBxOj
AGQ63zqiy/SUEIogjpMBly+pFXbMp3aKfL5382tPTzmzfCFiouRzoVyBVKlt0cwh
FyA38ZZCQEzMSouRyCTWZ31oTL9xTD6owR5rMcGiC0tyR+2AJlM/6ZUpl1JCcdKq
aHIJ7CDPSdpbENG968URXCEPxpOCXNBANYSX7ZvoW4AuMU+VUG6HuJfs9dkPZuDC
T8zdYSiTB+s4kog5zazdQmOLeWRvKV+z8ssShcJlDdNjjNHVKQB0bijucV00V8Av
AquegoKFBemyZ1i0xPcXu3iwBgT3aw3ZpkohtRtp/mwb5ghh0VKLSGfchko4Gt7x
Rzh/nIIqNdSVy2kj7QVEoko2lhPsd+PHI5OiK0e4+aYevTX5lk8YqcEpeyboOcYc
xYdTwL+GEOyOIkYpiSprHzkWPOvUYEWV04e3HonXvZJ4HMrElDYa+I2G3gh23EnD
ECmwv+YwRXdKEg0pliWBfv6XbX86fQbPf31xSv3Rs7drujc+51nCld5wkxYbgzI6
F3ABiwQhnSznGxVBInbGsur/9RxSPg5rYLyGfWpG+Q/VCBre4Eb2braHmXR+yMg4
Pcx2Ani0H5nA0RZ32aTKI4lD9wh7xWI7UyCF3TyqZWqMgOpdN8FJ9hghKEFFUS3m
C1JbPotfCbfMiI55SqY2psL0e6ZE1BSBYMcOhnsEY5znBKSbl7PN9I0ITQH3DnYy
g9E9v3lxeNupHxufKw5ZjOm5JaRo3FsL4CFb8diSgzlH0qnBSw2m+Bz9KrZsY+4C
hm0ZRhqrtdjzoaGW7P1TpI9qebVOeyPSr2nlvmx8RGBVjChNUojHKViX2ry0+qma
n3fXEhI2B0cKxUTJdqumrcLmmYHaFGNtS3TThaMy9SyXM+i4jL705xTi4aBkOXIF
YhQT4fdqXpquNzW39Mmy9Xu9S4WDOFThoxIklqf/+0B+jERn5rQNcP0ZCTltPyki
O17H9azQow0yWWY9BXbz2ezj59xUs7Du+zRIMFK5IMKezOO1lKTrWMCKNWWPqUpr
A9ym221P0z0qxYaDm4j4OgLXYfViCOYdcU/y+ndjE5p915wkiZ3DwEidXnHyuOG+
BV4SGNTJMBHbIjHX1YTk/Ws4P+B9jm1EUSRAyWlw6ul1BCfd0f0PTukdslfKXQgk
5r9qc3AXtAbndw2iQcfbj7YUpimFmFoeBH9qmz5SR1FDXujzTrnSCzSm2le6MBkJ
QtxPN/5gQ+/IsMzDGbMyrKjGE8Tx21WyQck4vZK1lZGC4Uw4psyC34pLVsbv68rD
VRCjl0F4WmNudBeys24jteNmI7maxsNC/QnJN1P+qXiBd3ddOeFLlb0j9DO4W7xK
godJewSYu32kr02Y+kzMOr2wpHut7qXFEl1CSL/5i+spxQyUA8E/tF4H9/P/gr9x
lMnaLfMHU9WK9oEcH4j0IUV8LbCUjZJoIOf8zBMbOzQzVKNBGJZov4WpFgHQVnFD
l/FQ4pMv/Le6AkvcDypJlu9X/nJ9BAZgQMLKJZTNCx/l18ZIdADFiiQcfowugOtW
5D3ejehYTUtUZqqkoZAakCE5MSX/OBfJuRS202zDXWzhs1vKGXCQrNPdYCk9ouVM
/phxH0clRXXPk9rhOMXHAN+2yHUEinUyj+LgHDNHN1OA5L18CaMqu5FYGEs0djW9
lm/jb0Rzx2bcDxPw7pIXVKr4xteaedjrP3qHePkT9g0cYlzxxlPVT4EM8x1u+de0
4YxUof6ZnaWDQQICNUpC/jLOtjKQTbY+nm8R8+f2L9OOgRjuimDGwgHhzzqK/Sfd
xJYKintovn0LIp6DsXD5A0tVuUl1DMt7wSVi6R+XgZ/bfBd/VUG1ap8v1bYcNP5R
RsRHFK58hX49jXM4M+kFy+Hjfi+1w7Cq2Ra/279nHDC0LxUlc/FDfSQdetsyr6kz
rtdSA9uNqHh1BjK1ByISSzIVjsO7xvDxSvgyYpCcyAvIs5OPgIat9QWBtUMHIfIW
f4X9bk0URSIiTsngEc2o4eT6sxC2Y7s/vIPF7mAmXvsUzX6Tt8HRwF5K65qmQU/j
W1qWfK1o46zVLrj/F3uzAh/Fmqc7VTHe+gMw/jXNYe9HzpiSv4prbGxPXUgrs/Jj
4h386HQED96Esz2eEwfv/ceB6KU4ib8GK2K+j7CAyAJad179/ZBNREZKGSEVdwMg
x2sU3R9z5OapseLgghI1ZFENZiEs2sWpERBxxIIadSAQhxHKMuooTgJ+5wj9uJ2F
M3L7a9bDnvszr5zte+gA1/F43ereWn5d085MdO91UGNbM2ye512oKLBByflM0GQ+
tjKDqPgnmW116KOUG4odkwzyrPvPbVs3OmAEI3rlOyvvoRZVtBpMUoS4ABZ1hYVx
YDbyKu9MpXSIzsjzggCQV0r4ud0qvM54e5IAQAJ66HTM46a1m1Cvj31G1tDyfaLk
g+7J/6nBdqq/514yQz8llmqytMaeEXmi1AtQcJWsk7nBIqVgd28VtczRhqIuRWAn
t9fPFL8fs3PWLj9+OuoaI7Poj6fjXfd59tzR/hsM0tO04MyIMFe9m+8ZLuzXgcvk
mrvFju5mexASqC7cM4Bs8Pb+yimNFcKDlZ/bLWqETVXiSUsah1hcdk6yYCDP1tjx
EuXGczekz4hXCtzj7HAeu0tPodRjBk2VvkuXtDTmAT7BI/q7dSmNopR84xrgyZZ2
PQ1/PZ5TU+xJP7q2WNLWvxmZF7x3/pydaMD5k1DW+IhJWFdoAoNZpLmdLuBUuqST
1dmiuOZqUP3fn1n8o/1o3sczE9SkVYKL6afHeJPFy461XTt7K0zI4M/nxSJdm3NX
vJjvbkoBpvatRjQGAvWUY4Hme8Mm6wbn/O0h+VTh81N2I1DV4J6DfEx//Jl/7ISO
ojbMiXFR1oIZpm8ETBkUYnD7Aade6Qk4Bh+VvfVnDLfdeFOageHdFZO3qqTU76H/
dDvhxvqDW+qpiUi368qjQO50AiYehV0cqxFF8e/v1iml/vwUGodqB/hDIkKt5M+M
rpM7rdQPUosGYt7kHFtogXDZ9IvmLaqbJ1y2RWIR7S8jM1lkdf7M7fu7JEExNMWo
FEgnCbTsUCQF5doBmezXk8E80ZHBxE5ioBWY3x7TrXOI/9Ku/nLLYaaN6Am8nV1P
EePDeNKjBXTV/d5PDmGDfhf1W4hBxfgTK+BTyIlsJFszutZtZ+0VEOp7RqO5xn6b
wfb//tu8cY3jb8rTPYW+4zu1R8Dtka/AL4Om7iZGpBrhYsRyu+d50ON86t18rMvK
CR5PL6HfbfBgUuMa5w+GPJjQRMSFCiljZ/GHyq2ta1H24P9G3Efd1gFq5rLyAc1G
4KdhphR1QApht9gvIJf989r6izXAjHPsurMEgGUo12AnIcta59owQhasOIR4uehm
DlEytQa3obXwBfNxOGxEHMxNgvJ9M4oOJqDNpDqgnAAQrXnFpQ9aHinIt1EyiFDK
2GtAp1CB6nhxKQkTHtERrr6pf94FdSln1WJW0n5YWwH9PYbPv2KCLzJRExtKMqjA
a9wL7Twps9O4JMB72ixNoRc2F2Q+SAkz/X/zfyG6Wny8m4pClxMXDP0GkqCr8rDz
LzuFCYgX6inU/YnAFDxd4EEb+J5Uw5BhnnqnB+YOUgZvrHngxUujPcT+NtB/JT+B
h67PqNGg7pS1fpKAPJyglyutI/4HdNrOa/lgYcUEDIBsWe5/ywNVcOY/Y9MuXtBW
nKK46skfBQ9dMgs1HNHYmzu9jc8POf/weCHpzgb5CCsHAaFJJkt1zEIK4VfAp5Ke
ciri67twhAH1DuYjc+9WQgh7oAfhHWJ9QpwPZfG8y/9jgKX28l9kWdLUvZAWRq2/
WRRZw/snIImxiTMA9wIYybh4JPwnrwWNmpdWgmN7siWHqlhlPX/IJ6zhxIc2vyrR
F+WXXeYjL3VurzSMRVDvuC+azlxJAb3q8P61K1swXODKyrquP5PARX58U0Co+zqd
pMG+XCJGhWLRaBabxattxeEU5Y7MiHlehCm4+Iq4nth6acjgjeri2BAWIWDyj5xf
SQH27IPT4KKIZAILOhDJbq0LnCpq6HUru5ygn/nBR6hlNAJCq4OidHsCNjKAI/15
TvCR7MMgZ2fC4td4i7MOtT42GhFvhFBLGSrDl+de/TQE3mEpX+fWtYdavWuk0GtT
X3K1HfrKVGetA7PRUs5NmD5Q9OfMAeQ2CJ0YvvDsOt9HSWfnl6KxrmDdlknzbALO
VhhapsoHoYe0vajBqRoe96vLZgw0+EgDYEagXqGqe0aUzt71s0SX0rGd3B03tno/
merqYB28t5IDW1RrjsbtH4UFICG/AMkA6ox4ZkHWoOaev4L3GKPD0rw+S9NBzVP7
BleDE0373V2/vufqzvJ/j5gzIvUhXisNmBrjM60LQbjQHmbC7xHeC2lwlxnDLtFW
DY8wyAM7/+fnvuRE737vdPxYGfjP8tIGaaxc5qOuHIwfpLLPM1F0CJQ3Tflvg7/T
fIcbFzRqjUujXEVOx/2zhcwOfti20aI5dkm5LhzJHP11oH/YKYSdufmGRZD/h33V
pxa1dnke0epAQusLlMfTKwYcXnyMKIPKNpIhuoDp0TllPYfQnhWeruWQUUYKPpMR
ELyj+uE/Y9zKdNQ4dAgzTI9I6qHqcXrZHcbMT4PxfAnwSUJsJ/Nc4+FKDXlhJ6Qw
0EfzzRNVRI+U50wNliwv4KtmH8uhZqSj434uFe1SPuw=
`protect end_protected