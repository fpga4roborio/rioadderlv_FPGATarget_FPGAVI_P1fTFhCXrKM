`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
ddtXksX2+yylW5zu6QL2Lhnb2d1sD00763mmSITNX595NcHTEkwn0zB1Dry37fOW
FufOhVzEJp80NC5qZ/+F0Vk7Ik02dIR0elf3clrjeJRK85K4e3Hoo4xn7YbFUIms
l/8VZSb14+JVGURjfswrIyCUotIzlzVYZ6gzoZwDXIi5gQIBf/gI+KxNXPaKV+PQ
Ufys/12rjO6aI/pPlqSm0hCvftmBcnezN2hk1UeXgOIuKZnogjOsf0iJVX2aOOWE
6pD/psybjbnsNB6kH5uFTA5frkzIzkzl5d9+YDm9OyC+k84E83I/7/j+rk4L2dah
QJOvksSIzN867/4Qt8qYTQ==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="MvBXkzurAa5VTw+1JJ70nePUfoQXBvZOku/SMmg4TwQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
oRtzZL4VJ4iwysPsC8SXYCzXS8Fw2gtZTOskLcDV+1B9Nzn1zTyNtlo6lNICRmmK
ZRVu2BmCc2G+fmzynYlNTnSa7C0Cuel6FYpxCBlOuk3OF2tzAmLAuDyOH3Z1Yjzk
a0aHuoCdIRKv7BrZCdALt03JeUmXKPdOmIlkVGFl8yw=
`protect rights_digest_method = "sha256"
`protect end_toolblock="Jn9CQpRhJt4rnzZPRk+dOpzAubz7omckX1MrFd4p81o="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 15184 )
`protect data_block
gD6l00tciPUa6pDNTk/+t1gcgy1iCdpjTkA/bOvU9JA+cpFEv5u/7dp25hHk7lLT
6tYtR8HgwcLXTcx68BnPlzdPHkVIv0lwXo6yhFVkYlDWBcqD9ubowgKij0UjlXmV
p4anbpVt/gKvAYRDYe8Q5F2CQ8AIsxOuOcJ2vhCPchS4QF3n7+oG0MKU5ZyzxTu6
z91WugsQ7cx0Td6ysKI33WkLDtnLus7kpoyW2jwUFaJM/8k0THa3cuHPg4BND0cq
JmI8xpfVm9BoVCwGXTqNWemklg4h/zUHvcUrdnzyivAPM1IMKQn5ltPvY9C1wLmf
UEt9T94ZNzzUeMWQgLK6tLJI3qqFhFKEUtEmMI8bd5ksXf68kBzJ21ELCW8HJ/KF
8UMjke31st+n5XNAvcyrkYTqu8dvppPTjsISG5Ex/clev6IrRHkMjfTtzLGVnDck
wlshFd3s7nXPwMVSLFmIjKhHLIpsmS/wA1NXLc5CL888xRrbzVGJZsoRMGy1gCQ9
aMo7pPCX/uDVr2MUvFmzRxEvD/Ne6SH9UX1irdEPxJZmOXWl7FqIsEd4LOB8oT/j
ebhjoZrpfMbxRSnR2qnt0zY20q6veoQprbddsLmGrdKdViTBjkZbfM2RJt4kTMC2
L2mgmpS6g6/8jsfWiU2bECKc6cD6sJ3g9QAzGBm0UJS8zjfuyf0TxQjrzxVNv+G3
pP9evS/5b/DdPw0Lnizwe60ad+dpq2T8JUIBFnDbzdW856+WzO40xVQcOTZE4zSt
z+9N/qh7qVs6BqzwGD8/VTvkFLH5xyy2l5BQEoMS9UlUxtGTUXO3ANkW4A43d/yj
i1ahX6Gp5oCYhM44L+c/NNTfwG7+T/hb9NzEwIc2NDf3AsHY3QtVADgX6614RzG+
fW6SALZdR1shdjSdQzNUHlW5GR26LWMVcquOV0ioCdNASPsOPkvNX2ix3WNf/HNc
J/A+Kv6hUfjszcygUrhL8r1lOYGWm7r4/QHyQTfkL9Ds6ZTytl6+hNlUyh8vDNnS
fCW5rgC7YeiusxI2Y/V79Lbfl2LZ5/SJvK12PNmlxXKB+fQsqlOAfJVhaEgfJeff
CoLlf0vBhzxgNSojq4Tpbn3Z4wqZ4tGgYJaIXpoMN3CW2TJlf55EhYOyb/0JBmAy
Hx/7aEepxCRx+szRUnwLA4Z2IxDBCSaKdYfQepZHOlZUS0T/YskK783jhZWgdjS5
BiG34ApoNVVf86ZlRCdtg1jQMWZrUfZS3LjDNNqDtqEEE1NZadnF84jdhmSzUtSF
LjUDgJA9NMtlfFqvbdz+aOZcfXlMeLUzs97LSYTP1bYzy1+nvZ1bbzXVw/h8gwHB
wxm1yG8WMV2Ykj8AILH590uW8SXnwKnaxhzvAYf9vr2+w+AxUfCsyW40x6cv1ebZ
ucFsdVQqY1lCjO2m8UvjgttAg4g1YV/zZW4p2lMYMegMFTTXwudBa9p/cv3tZkHX
I2b70mC2LdAVa/0Mp7LohQDuJNBVuomiifLDXnkvYsulPOTh5xdQ2WM6BF8Yz4Hx
qnRIlMwHWXb8+93fqejlOoxSB0K5p1KX5JlMZPEXltprRl7aETRn0YLOAY2YvzT/
YMQjiFYPt8oHeVae/GaJOtriJ10rrn/y1YuMEHA/J8vZ9ddJAEGwl32kNfMGRTsn
tw9/GeQ1CwvNsREDvu0FGndJLew9fC/1ViBm9OEOHAsxteqUNm7XPnc4m+Z+FFW5
kkO+DnyUz8T+UiTxBD2hiaKq1Nt5PHCGWZ/EwtmzIBH5zEUCC9hCyxbuiDduwDxh
obECeaqAnoF1/wTSlSd5T0SLlsedQOQ54fQWun34g3dVRRsd15Hma6hd95H14JJX
OSp52mqlHXvpHeIWTd9C7AwrjqvJN62BvSfX2MDBd+05dZ1ucAJ+3mhnlz1ZZMZq
Fsi8VgjLsggG7GVKHtcPuqCNr7qO96dL+VIXoB1rRu43ZHjH5LK1Bd59URrQFqXX
aLYx4TvvEP4EtEr4HjJactnJTk4f0Q96cgQCMV9G4kKE/NUdoUq5Fdl9eg4zcLRW
ZF+ICLXpDKJDtdNCPkUsevOi9vCoOe2dv4awx9aLGjKxN+2QvA+1uNxu9E73X9Nz
P9VvbxVqSj5w2P2SlDsznzOZPDE1aBFP1n8gJa6rIfXJ663K4gpzOtVKjJn9ejE/
ntrbOX7JX3+uz+6oPVsZVXa/PVyec3tBwI+2BsB8BR3JbQQgfxmssW+tfeIwaCHF
9LEgCyABYbGNGt+Xx/Kk9qy4ipv7JlZE4P5cwKEToX0NzXY3vo9eeHoUSXQ0phf1
2oJvvJdoUEup/t3kDb9aKufhC8hHBct2JC2dmwcjo3TCUu//UbyMlGfC4z8xvPPb
slNg3/tHLB1Vq3k/baXHuXMymmqkVTsSWP4TRSi239eoSbnF14AFEcg1WBpO1vvT
wx9tnpXR6NwhQE6lvjX0HpWOSDW7TliNWAdK7IkKA8by+2j5THeVXBeEZzfMAs2E
jT3KldUU/BNQlpyPvfR82NYIZbgw2X0KAcMAAQ2uWSXtvpBGurcSIRrqLoDfsjP4
77BHXVksS5ABMXGMGVKBihNS7OzSxhTNh9V42h0bNEWFjX29FEyyL1LfFA1eZvwW
sj3MqJiC9DegeQmshBG0aa79MDo/ZEX8QVS4Ooe8hyToKh7zY4cYh0aqkl7adpxC
EYmP6mmlmxgsiLvpLDeu85uLq/cRFPKyXSU+6VXLjoupUwsXSZNDUdlvHD7rQraV
Wg5H6OVNvfXWG4MXmFhtIpass/A5gXimvr1gGivb21qj2ZmL4mUSUgFBGUa7E37a
BBuahi2gmmpaDRdiLHTTNvGGaq8s4oCuXBYqs/JPeC4VQyZOJuIs7VpcbmkUYipJ
chq+GMSaBVpl2jrZh5QTBzTkVyYhqMSKJfGrM2oslKDflstXkrYq+F1TpT6DGY/C
W9X7DoV7IhMpVKJ0CH79elVbr+/N9FCJdxa7wZxMzNjSTeVfn/PDhAihktamoOS8
+qTho1pCTchINsvD9IKnicFOZafCtrGqQL3UE0emLwVtshysGMCxz5GdfirWgbnB
q43QItVoVKufZbDc6uP3jcGWj74gEHnzvcVzfcvmVKbAPzYcXMCZSHjdj4QHa64t
hVIn4aglSZclsWjxMBZOlqAJWveubUmz4Vlj5Vyk2YFFQljCZNsH+86wOH0fuNxm
mQgj2PBqpsZtcFXZTnzHtt4iVHwvYRSw0Wy7Nfd0Xb7dGgekGQ/LCfO6oqfHnFst
2Uo9MiXe+wkQSUfsEeM/6utsYH49qgyy/1S1LVl/xsEJUnZehVVrCKAXq+esUSuu
Vl3dhAcTAv4P8Do0fMs4IEKYGd0tR5La1WcxdRWHOJLVA0p4D6Hwz6lWWK7xnCuF
k+Tf3WE8x6drzb2CmJbT35KQIaHwoDx+mEHRB1jJEEKKjYo3k0xcHHAFtvQ7wq2f
oY/0cUXGZf+wTMdT+PdYROyoa17jSPef1RVi+Ob2w2aRN8h5jmekBFw6hQIF75Gd
TVHIIBg4RoMkS14hQ6DaffGg4K29STmAY2GcBggZVnBrmMKPIHb58kHIo9EZeg2y
cOoJeHfqXT/Bdz6APXva0yWedJRQMLrq6NEPnqaGEYyFM6K9dJG/Geb/rL8Db0a4
D7D8WBS4NMwAp7VDW35K+oUn/RoyC7/l3LlzSSbilP4t0pnE5SZN/dQNNB91hpE1
wfMvyNa2DSL/E42WEbnnC9NHZ/L/Uu94MNd2j6gfPhyTfdbAYJiF7DBNe9k9tpBc
hyHC+KNjp1O9RUT8C+Ev7DOAVlwFKHu52R472uY0X9epMz6o/a12XNw2hRX8Mg8S
DoQ/j78kk+CR9rPonyArO6a/euzkKD114R6YuZictosXsmd2y45uUzBVhFsJ5GOx
nWh3rz6N0xCDNjyO2vGoOaVkvDXKAyuOI1wPiPubTHkiaa3roEsIOfIGUWHXxqU4
nkcC5WIj78MdklkY0rjgTUDVVb6cs3wUx1x6Upld8J6912WNZbHbYu5itik4Ye2Z
9/4hflR3X0nEgPIWR/loS4nHdolOnFt10K0Vd+R5oQvez5wf8Tlj0VTemILp2JrR
/siXh1xExAd0WCKDKq0aDzI3XUywlobUUoVg8pG3cd2iSiOVlBR2lNcH7OT041xr
1W1TY4UZ1SbPytzN1/Sj+RKQUw4BuTSnnqZAGSrxkd407e2zHM2jI76k8WyY7Ptl
KF8p+O033ur06wr0l1Mx/6PRAfA/oVxkNdPKRmWbUvJCHcy7JLUS7cG84DwZqZyQ
cvERIbPYFxcLPgU8yGUOQ/5VC4CvdJZQiCIKsYh7isMQm8Tz9Bx3L43oyaHZ/uVQ
HaoJJh4Y0jm7IXWHvusxng30wqxXXpE8lH5LacA1hkNjBjRCqeSrdgUPjFJxWr5o
1oFOi8pLRHj4nC4l8rY4V0Pjgrgv8RKJHTbMcTAvulXStE5S3+vJsBaMWRygBXXt
+MIsR8naDG7AH0Kjif6Oi07FrceJKsSxs5fXikzuocmHe2kC6h7HxCiPdK0g3d1z
CXFAe0K1Xp+59hWtZIoMavhi8ufXHExsk8ajxX07uRq3GPsHFUCs7UPbr/EBjwEU
CmE9B54dyOLy72yyBnn6Hm6TAGWjtDQhz+CByAKk0iIemDgZWax0aIuFn3N15WUF
ZDe0ykEGGOr4Qb2Cst99aGJN6/f0Ysud5qEj25AaGkSkr4ZJCF+ZxTF/JDQYsihd
gdd7ptUtAPa2BXwQGF9FRJtxOSjO6DZEgGWzyzizSICU2Thb4V0KkRkjv7OAcNSD
Y7mC8D5eucs+YDar0tIgfz6mlL6iBrFhPPEM4crIbLLcCyJJ6CvyU20UtLqsLzGE
dIoAaGRi2URyC41rp96+xodeoZ2M8yjfSDR5I7S59EOEWj011UPKX4OZbXNC8bGY
FBxXOQOw9HMLAznR5UxpTSjHCS6G/MBKoH14YZt9b9YquqKzD2xsB4LLU/4RNrZC
8ZRYd5SHBuyA/New7ijfjRrIYK8uq0hYfqQXiU0K2jk2qcB6r0GykbsKTk4BEy0d
cczdjgChad9HBxqMY/Ws7ifon5d6p0AUrCLljNu2NOGxs+SGPsBLI5yGw8wjnT1j
k1VEoZXXZB/5t5omtQxFI9gex5yM2u3KVlvuxZOBFlIuDWeRRNzNkCVCDiOvv7Cw
9GVBllGd5xTSS4fL7ry+aKGNrynON9EmyMuUCNBJvXKu+qQsqVLBmhK4DVX09GmZ
hIRpC64GWF8gzKqptQbPwjRl6hPDhDOSDbw9nXTXIbP3JMZzlUoiDY9RbetjJ4sd
3toStBjvI/5ee7j7aE1AnpuEQNUWhd3vhgSVbReTTyRxK+CMgq0SXPFoOHV6xlCn
hTm+fGZQwgOIdfttJtt8aywQHNLPPea1s9PE+Qv4+lUrIfAGM3yvQS/ivq7lcV4g
0AwhL+nwZGDkzcyuo+in/i4pb0ZecIGsKTHIXwGDEUTQM6Rk4ONQbsNg9RhLkQpX
G/BQn7aYZemsqUYV3qs8O4w49DWQWXMtMxnWq+jN4FmixlCOmfI4VI6thBgS/Yi7
kddlj21WtayHUziSV9KKJEyc2qOTbHu/KBU1aqD+xCEj2TSvcGNjX7weE00xq3el
++2Ddx+nKZbc7dYFfmGzDJS2cWK+9DBLzRxSKQfu9tYIBKTmOirND35Iy0ZXo4//
JXq6zPI6bZFfUD3ZdiV/06oAZ4zALo3RrR7sjnm0erS9oDv/NVmGDDuxi2/ZVfxk
zt6Xawmr86JFBFDylvzNhKEkHuFtUhX4Mz2cvytk9gyGRQfWX59lRExMwBeDqwlk
gpxA1i8fNTrDN1W7Zt/RD2RrIuSpq4UgGadcYJdSRFZYL8Qbik/KlzV+xyfHZgiK
4Nnl9Ka2OxknxO8xLuhvZul1PM7h/YIK6jLkraHtfuu0qdPKrEjheRlCEBrIKogV
vzIv7PhaZ2ydk94aZagSfYfrrLxkIYYwIWwhgcwifwl9eCsP1KR8epu7aV/ToY28
WEri8v9JHh91flDbGgLA4ps1jTk/TyXTg1dT2H0NupJGpzfI527tfbYv7vDQw6re
tft0E5IZulQRa0vK9N5bteRzfHrwlrFVuDK1BndjxvNETaAnDGautXQvBbBuCSZO
8O7QbAeDxTShGZkRfuupW2GmvtoZgvwT8Z4IJPFMI82l0RbfVHTBPDs2S2p6Gquq
5fziAnWZX5Qbj+4Xxr9QPlBStZXB11gkVZuhkQQZICCCThta7uSBEw5NyYUuUp3A
U9Mhd8+IbFzpkQN/p8YMqdX9Nv3vZoQ5CwhzAY1kZK5WMQIQ1ryNe3njdGbKrw5G
Ps+d/ZWQncwT7yGBISOfjGFFx7QYpFWctZa0t/o6OtG3qxPCHc1FSXsc2wY/tr3Y
ig1Jl75cFW2xBwG+6KcQWLWi/iB2eX4bIDmXpqWYGJn2Jl7M9uGdjjk50Pi/SIYA
RwdUzBrr7AmCFSITUgB6ImLUiSd7YlSPTCloqyji9y3U7/+H6XvS13Ru/nJOTWDv
oq6TEVl0wc9GYyxNbw7ZPaqqXMXC9e9SriMOJ4olqQtMlXDaYx1ENA9VFJUj4fPU
LmIJ7t0+C8jfIrDYPB6ipB5Xl4lGacaba12dpLAAw1leWYA96Ye9Wrzgh1ZVAjpJ
1nm6lJ6DdganYYOdKkdwVyRLzMnw3uXnxu2OXXyFbcfHp+d5zJt7F3JIYjjsuKtQ
3x8Zv9vVU5/rPkGrpfWPVuGiEMOfUQZnx/mO4jxAv0D1oXwirMSRBWbh6V6IEEbV
2RmOcPrs/FWd0e/HtQxYxu9oRTdjGHUn2lU6+5xH0xGPH+VJUwuIcNHXLCCulyYP
Ap5OQnRwjJCy57v+iA54Ee7RhIwLhg3AZvv4WKvL8PltF5I/m+87xSGl2Snbtogh
dIGvY7AqD6Iz8GK5oG18PymIoUXLLsfAmqzWje9z2cPuQ8Pko3pR3dnXAzXKpaHR
XxQGEEJrXB30TMeO2gBb20VeoK3CxZToOJuqdOZDsJXKNn2WNPg/fS6CxZCIgMgJ
jeJaTZg3H7kC1PIQ4y0eKO0eX1cXzgodA45Bh+OVrj6L0Q3+b628yM5jO9wIOfRb
Vi+DdtyiRxck1baPWScw5ZGZes0VMEPaEGMUKXimFQ/LLtkB5KovvxXnMdqrgc+h
NoQPVTP0wuvQcogZvTTuk9eB0Di5wG1sXCwE9TEjxDLc/341Tgdc/+dtuBKQJB83
AXrip0nlzW+hKlFxTfNCmDsZYlAd/9VOvfy5og8wE7zgoRf0yF+TAvUtw3ijCMLm
vzEwvjpklslyjLkcUYsW4VkKqZ4h3KbbdU8gBlexy0cr8Ispk3zTZg3F4wJgYq+K
aDvwnHGSz3cS9hGWuTEXdpZwc0OW2zAaitFTxQBJfhfVt+xxuTx5iDsHrv2OMw+1
UqfExnWvRwWREMgKyYkRyeEmL5mx/N9BGgnmFkZQ/rO7VHgYlG3C7bx5yr4lbdvp
w/kHordij8gH6lC8eSaiJgBRpIr1TskaAyGFYn86/mJH/yBeJ7Qmq8nCxgBlNb8+
TA2dQwIN4rk+2KW45Kc58/32YcSXBXJPkCkEuUddW6PXlb+PD23AoQ7upEER4lmV
LlfJF379+eGLglgImHVmKlZYjs5TlpZp6pk0Fn4qc2ADH5c91HbB1/1L2ouEuMTU
AQV+8tkWMrVNTtVVTOl1Vz6/kj8dx9BduJnZhBGSSMS/Z+tUSIz/Nh0pArSLlpbA
9fC5MKRoPrT1nglptlGKgwUwwNRbq3prDFL6f2+kijn0AWHyfEHTa5pJSKVouuev
hfsC7CPXq+8XubjBuz2j+BOLgGV9Ok99bi2yphJ+bUUWdwhaX90rgW4mPR0hrR7o
h1t/sQTxKhb3Jz6arpUMk8gDCOLFja5Edj3VspUX/ks5NWT4Bwi9VubunGFCoQU8
IwDa9k1fjcfIjc0L4cWZoGTonStgWZXaZfCQSe8HtNK2DzlQ22TOyxftzhQjdZwl
t8emwbY5dAvEYJ+ySFBjtew9F66VkymoyjTIbHRK5Zk8P3S4LkjSQaC7zetfDmN5
xGFVv34XVrj1byaFyaHeXH0+8ZjT1LUDZQOrPZAWwZdmGgxqKe8rWCz+h/8u9I7E
gvET6ZAcRlKXNKXcYz0sNyg2Vsn3hdSesE66KhWT4GiT/mLSmE+SwoK/CbonduSG
mTpwcBGGxkmXtHlHS6Nwo1XT2BH9zCk4jxdPkCDbp7xNdKRekGl4w0UTZN/jHpJ3
/Hf9grtUOAO+P5K6XXFsYrPiPa8wcp7SascWIB6+AQfsH0BnuP7GLkealzhW8PpN
AbDfQnwdR374h9VlLHMU1pF5dFJrs06SYVDBkqT2iodm/r6+FN8vu+9WC+ldq+LB
pKhlEy+fx/joNedW65avFaGPB0W2Rd4z6r7yMbjHVtrxgoJTiJ3+SVRIbOPeUW9J
0nyRxUtNLFxaQ6lj92GNe3+YT4W+eUGeN417WDegyJy0kvBNhVftjrR4//Opty9h
+LKvA8KaPuW+WNgJYAy4/SmdWcUlwM7Q1qLGGZcczRfChSv8i5SlZYkCZsYQRWcH
WJT3W+yyqaY7J1Q+9Qz8VLdJbYEAliuoK48EVLMHdZdSg6QkEnDJg+d/eRrW2qim
HdROCraYYkvEgt4/cl3ls5rvypaLy25DeGqGr8VUTFaGzbftPSm8pzBIgh7YF03t
pcJnDcOHwnnyF1diTXnIfmSFPFOp3l7Vsf7I12zIu6EcHlHZuHmh2Uwv/Pk1mQZG
+2qX7Pnq4m3oiKAYJhab+HFO69zHAzmpxCEf5oAioiR9KhedNmAoKjoZZ6s8WrD5
DN/0k/Dth85tEx4Imk1fE+qh6mpdFVClBIGgwbEeVDw6y8QPBmVMGlmOhIIuaYoN
mmVxc9i1l3pQukV9KjLpBOorR3CNYYey2lwspuS+TtVFdfqvQIaUEcHUfauU334I
h4oqKpqOiUSoOgAVhc5jmEUwpNY+9zYqqSav8LYWK7lLpA/wEZviKA4Wfw/QzOPJ
VrtkXMCxpsiyn3nFOw5L3DwYT47IQUu/xI70XBOnPSIEzlPkc8XpotFoDDCju5EJ
kq9UuBTxGe4zHqAo/yPbng5ECTFnRlv859yf8Yf99Lv8NcPq/M8x+HbUSiprUjG4
1TmBXllUrsBbj63jsVT8uzwvuQAaJo9aY+59gYkCZS3kee6uAumfp1oJUw4gTqAs
lKvPGGGHR0/2vJfvZqQruDtIEGh10kwc4CoSKkPoZkNzSSdsUIVSPM5OUyw7qMz/
hAp+Ibwho0OBpx1/zt1pgm0/OHcmat31hlOC7tKohtHBO5RvDMKC2M6UGX1SXM+g
eEq/1CHM/sGNdsw7pARgP56iaFwbk4AcYOvaj2/BUgDVna3mQXqLo7UihDBMG7EG
pjJ9XIB6AcQy94EB+OblByj67Qu1cf1zG4BCmh9R2RC7zScZaZmdtEyS+cTN9kt9
MRrvzevCr5ZxiZixCV/9PZAhLT/H4WrZ4g2gYU0Esd9f6uG0YH1oRsgkyTuEgnOD
EcIA58yChaqnTQY9RfOVrx2hS6qy/0AdDhoRTi4yOBtK/rsREUbuJ+nfmzGidkBV
14I+pcpIYH9CFTNrR/a26ySveqz6VfSRI4bwC0DDWELsUl3KTGhjdESGedbsY82C
blZSUooSQ6hzt6Ty/YYJbxwms653IZ0+U/tWgKyX5Rj/RuZKSgi0jOCpZ1MkGD3C
2gaLCuWemHymzCSCX0vMh4TMocl3UUOUu/9eyrc0ERvYH5IfAo+rxrf/aAVGxBE1
QAoC90BNmuxpn1FQg5dR/OQ6kwwgHkwUNQHoLiVaNEmUXKWbc0jELhAgjQ990TEh
jbIx8HCsghAIBQTXTiPv5NOUbvf6CD/qRsiWjV6pzmJyr4cfqkKObTdyYWaVf6zi
2AlhhXxqCSaYps+Boa2AzR3V5TtRVhlqp8L/slfxQO6VtiGRAA2uYa93gJtnnvzg
D/VCXOyVqchrNu/WYYlmp8qOmdUyOyFTw/vui/F9VUcjOR1JhjI+rNOQN1Tm286G
GukuS8iJUHEUBWt3Tnpd3YgejNhgORKmRJGfq5tCf/3rMVk2bGigSDLt5XtcnYyA
iyr4uwFvygm+yiwq4YJNpNQb9t9/ZJ1NqirYjS7sanHds9DC5ENgzWfSJ/tL5cK5
oFNJw0dILbatXzPqg7et5dzWbFuWDVSIbK+PcvXwu3WVl5rll4KHC7mQrTlJa5Ck
ZJHRTX6+VQ2bVBy00dD/WBrh+kHqGLc8f6Whcx26oDxCjcdQyxn6eTW9E7p+76O4
q/bn4rXwKsT6mfc3uONGOoLev6smfTgJt97gWTuhQ/dtdrRZ1BPYP+T7LwgpnwId
e1bGoRuhU/cl7nWf/vZKRBkwzAhGC6m85hJkpjKASo8MkLGfuiNtVzg8c0mNh2ZC
fqyWpkM2T9HLkbS/j6/TplaDUEyzhh40vpecTNAzs/gU1OyLK/0vp++jwDyLesVX
5rVhEgVFKDK881dDhTgmYsrE4XLzsdhU1xRV/i2uMq5tB5dmKDoSZeUxZu69tgVA
nZgtcgnDgaahSqDVXrhRbuY0nEWLG/oS4HZSRSN9fPRc8CZ3siA7apfiUO6ObrZH
PHrZ4lOx2qZRWm6nDdxD/bB5NUUvttRUX7oydk0f305FCOEBZ7zJeTa4/EwRRG5k
b7UwLs3Of4tF7JMHhXRG9WXSFMy81Fwf1MTcO9PIAMDCNLH/5T016kAwYDyVtwHq
GM7GifsZXvKEtLJInKlCvryiNbbx9nagUS/xMvU6zuc4NTnfysQdhhZ2k6bMZGOe
IJuXIEuZ5aU2e2NmenW/SE1mEAEINfC7QzeFu2Y6Nvw+N2gi9a9AzwvlEDJIUfRZ
fTIGH3MhB8dGRNduTNUTfd5D1m2xWnJF+DSyYvDM3lCW3KCehd2CZsAegoecPCeS
QqfAIqcpaTEgKoGiVc4r7JTgsyzhBQQLCZQ5qFEmqOzVhvu3RLTS7nZif8vIUHxL
XXVXmM10FsFRy8msfMrFZ9EgBh8nJOuTncv+fzmth8t4GA84/X4vUi9GEG+Ci/qk
Rr8gPnOTx89dPaFFkwxO8v+nn3tSSR/VYLP4ZHCrrn9T9cAhF6x92cLVN9q5bvmX
OBDEpO4ZtXYIznxgSGCZhMnwzzbHozFmGegt0bCsK6ej8BbYFVUwshUWu06lo0KQ
HV6g4UxqukABQ7c4uiE/Vs1Mjva06vkAPnC4OfMCWwmNke57zHA0e8X6ID008tiu
7+KrVGtquXuXiGMmFeHACzppl1ei9eAsDceiqatgyljL/lF+i2+z0NMgG4B94dB7
jhBw8WbW5Jzq+gB5pMeix5t6i95fduEP0xllplukVz7YHHsaeIKXeJIekGfQ/hmu
5Z2lwzuuMx6mse7dRHr6oqLVy5mcguZO+EPQG9ydH3t+noorkv0MGEss78MWM9ML
blBOnwGhoKZo18ejP/arDISJMtTTpkLqatfUYkc5FMSrLhBkgLFphWdNYuCTWWmw
ypbDjc9zkzTKpAkUFZVW/tdAy/u/tdQbXli8jq/DOHGIVQqnZRZlBd1mPQZKASmf
ipFYUcjl1d0ZDvHhuU6X578ULr2CzNj1e0lL++0nLCEDdnbNpioAmoB8idLsQPNy
d8COM/xXocfqz5Tr/qRFpILbZwPske3zCWfpGrwW6nRRVy+xZh0mYhP+0NlJKPo3
W1YpzUmIQdXk6FI2ACAme3t/MOwbINGPRdKrfTv/57hwuY+pua3/z2iJUs36jus7
RiqwhWeuhKcFwvPQikVW1v5/LlzVMkLoHSLhFHfZeTGUflUHAfFlS5P4/bCp6yAk
a2S9StISq/NL7SNpDfQbIX1582mWw/BniAWxtI4VkeJGTPG2pwNQKEVafOqqbQZq
D4RiTejOgz45PGK+HFzJzJ0V93NdEPlH5wMnjQweRjWR80suVHC303s6a4VtQ66L
M9vSHB6dSPPY2aRS/42H8947sXIktiZ9wM9DPgDSKQX982uunIeLakMnee2N9Vj/
3/oFHd0KJbsYZTJhiINgjVst6aDKhHmHssBBiZA5tebGikdos0nF2vtjJDZNRHfO
eCSmEdBvsxG187AOcPkw5GYCDOxiFBzKCYUHLY0QkqFNi5VgK0lmSbx/ohyy5V7W
8QaZeZfgLJ/U4VHH7FshNR25d42YEWSfzBJPygxseOLT+qqa322GxCpm95EXM6+2
m6FFf9e2yWbne11RReaOsf2n6ScoQ5NiEt9qsPKV5ucXKKf8NMT1TM5MK2w+8+tZ
6s6KRmneYKGWlwX301zHjcVX/WyoaHKjj6hZlr5KZT9uVfchroHTM1k6jguCpD0E
dRM4fXUGCXNIkXrA4pMnufTSJRboPviMAFuFSk1Z1qPgtmiZekXstWrkvgqk3s0c
iZ+U1Y6WdbOw4qPU6ytpUbizvNhHAgRkhMRbF+hbtuwlKVE1jvFIg85r3rDl+P+c
hPr4uDpiXp0qpwUgQg2hC3tzTgaTao/noId6RV7aOSVK022D2II3NwA8YNpNZHkL
UKYbWeNAgBgT2v9Em0u01MGifq295q+ly/IFjVtK/I0W6alRuYXemjfKMoPGndyq
h9LMAMLjE0IdLky1EMRxQgPG6iaATSVY491iHgU39z9H7FWl8YBEb/13Ev9EZPnY
TwotI1uOAmHrfPT7pnAarpIPqd2r4e8qYds8w4iajLPb3F/Cfc8E8cBVOhQX09pA
53tVqefS/MuVFTdPFSZJ5x7rqAxWc8pl30ObhkvPyaHAuFXQMeHC6TcRl5F+/yfz
DFWBEV/1IyuZyaG4SjJK95ACrQvMdByGft75r1SK4uFDtp60whR+SKn5HTDU1gyW
HbTjO4cq8e+oKdKfUPwEAqpsTdnqbPRXIkPok6h6ou8zEM122B3MtdQRm1bdR5rJ
xxaFRBmLYNTfhsuvTrglkgeHFVLv9Yk9jFKHj/aLkA/XukthUweic7yfHmor7Hm6
i99PnuDY/DzGYBZTX+uUlaSDQp0ztHyTQ+Hbk04jLTSeaZQaFTvXjHCytdlmvV8q
RA7S26vN3IzMu5jNroES4p8ylxcMBXXSHneEWyWbYMX4RS7EqCKzry7WC+qqrxoS
gI45MQqSk3LRHu7XdPX9D/5MZZbl8mLRyDNDndtlDTTZCThc1b+gEiTy4eva6qvl
bIzqWKNxja/hNqQWqhnYbTjYWs95XXq4/0gol4cS7b3oNAYvweDPcDs+pHqXIq0n
WQbU0j6jEG/87Ym9Fvt6FBnj0YTJuTKxqKcWsxg7R8RkAkNockwIcMrPDMPOVDKB
7jl+gIa+FOR3RkWk5XsJ1yfdTI2Ap0mOoTOqX0c964mnmSIO6pbu+z04pvH6EDnv
J1cujmZyaRmdNi0QiY7c71xCFospwn3Hutqho7GdLc96GNCQ7y9cwf5mlsMMe6/s
UyjzvLEw9bOeB9ScBQrc8YiqiprI3/BjNwEHy2qBj0oUe7zyTR7w80ln8WsMjH7U
yroD8AA0+Hvm2y8CRQvFhiY3AQ+7bYs4M7Au4bAlU6SUotQwQ5wes+0CBHrKUmbE
T1LdkawYW/atuXusLmuj3mOwCKj6igktLuFQnP3bhDbHAvmayp2UZUe8tkv9tZxp
NKHK4frL8HEKpnUb05DmW/+R+20Hdown1uMKGuOSomUlF7190nfYpl5rHvytqjNI
Wc+5EfwZXW1mCdjGERbh0Rzx8JfNkmWNuBIz073q3wE+PoZCL2sgMmaC+i9nkG2F
j5N9D/r8wiNMSNMZQy6WNfENcuw+R/P6PMx3MHlPjdtoXtJpEqC/4Ej+jrYo9Vte
DlVnlB69h43jGILSx7HMLAkOYO25ceGKW+a1M5N7+DsdxykkB5ifKzo2Y913g5K+
cNSQlI811CSGFX1J0YaTWf+ZmVQFsdsKRHa7azrgRb8cH2GjEVXJY0tud+X4rt17
hgQ8rMFoMX+QaXVm2nTnRsmLoKovlKWtJTAI0PzSUP/S8fP5SQXiDM7vhVrivhr2
y6shBAHNLz3OOlA8TRN63o7TGch3NieJhSltjFEKaasL0Gclt+HI7NohCjjtJVqj
9uA7pEicJvHjZXyBMGjWuYUjsF2gbmTh+NpbKOqnbQK7s//XGxTIrOy87FRKKkpP
RZPWsYxB85Zodvhw05I2ecNPI8hHC0eNJTDU7bvY7ofdZLksOozo3wfYmGy+CUje
33398+6ZoTg3YphQc3dwOdKy+5D0wOh8fxGm7mrH25xT613hLk2AIKaF5nbUVAbK
ox3SuH9d6H8iRIKR4JPTVDN/AY6BUV9VcOaCYYbtwgbQmkLReVkzYOg7Zci9yL6i
kl/9dQehOlVg92e8iFo//fZAseP7XRBm2xVmjF0q91djeULebNoZIlMgrhpAoVln
3xT2FPqH1YcslUlIIxayQgKIS44TgvPOauzBsXL6gouqupNWh+buqIXTtkqmHiOJ
OzXKl8r+y0N9dlUQEH9U65rSQ3pX9irZCmoKPEcz/Si7DXFt8Tfydj1o2wOtOlZo
nD2f1tlsiI7cnaZY+YrWFR0Zq06sIEqmTR8MTQdwolunyn84z2BTR12jrH/Hpyox
YOVxCiO6AP/B910f/jqUDtOlVRhhwtqT0UbAYEdfsXy+mgwBJhy1GrMYjjW6M1ob
T6NaQJovngnuWFHIDAVjx2bL95ziMZ2T2EaxdCA1TlMdg544Ef/oriJquUZuxXmw
gO1NMom5vMBk0l6m16r1pPoCSoA4rAplvMHsHi2b5OMI+2POmAydtOGgNx0xuGC3
NWhQLGE7WuWbX3mBZ6DrGesM5kyRhoQ3YtcATV5XIutCqo4l7oaO4KIyaafA0jHV
85o9Gsw5N6z7avhm1pKaJ5ElIQemkKrJSTPGFQ4RwZ1y0kGqrc99MsO2ad23p9rR
dgcU6jPq0/0dp2ZtAqz7aQUiMthRVcxWQ8iB5W4Erf5nJslYcKe0Hlunx+9IDBL2
6pwIsSQkNX2XgR9gm5M7yuuVikgDltRdtNtWT1/IJKEnZn5Xg4gj0YDbh+IYG5Im
NVYpb+IlA4An6sRp/p2P/VH9a5DzHF1OvBJWv5vCDzsg0fdeymwqPjY8TC/xROp6
Ifc2gynuXJLlIhzF+6lPn8ny57pzQd1V4iM/MIy+241IZwRKVprLeE0C1s/+YSqH
2NkFnBBBdOEQ+5qMYLuHcmJU9WDD+vnMDDvxAdfHf/eu04N843c7wcie1EqeCZSi
LfoSsvE9zhs9XKzokuQUhb2CfLe5fca4sIhITS7cIXp8iFk5Tlb9r74aQ0H/DlML
FSGE/8JBVsuuAHllOfUXYy05CLA7rGLwIn51ub2Qpls6CtYIy4k9csEafCOf257C
ESnTex8ZZ/xTInXuQGMYpuShYJKfkQipzBa/jBn2c7ID7ZOYzfVhs7HKRAJUuFVT
5vmfrGKWFqy2PYyaMEaRNgydICXvjJeCIPP+EkBgOwAwlQm3JFSiY0aM7NKMLDmQ
fM1gpHPyDe867uFHfkRNWrpUui434DuaP0+WLiQhMW4mp8cB/rdzg0MZUgnUuB0o
K1y9Wp9FKxtsj57RA6JdK4y35HN9zFHYLgALCdoWOcV5R5zRIZX3AN8q0EzkdcBC
MK6amUj6xSokoedAK9Sqf08GE92uS5c+CXPgFkJxq06JDLvHnMAEKeIWsX4uIbNw
gYdmU5G0uPw62aKobp83SxAiOrYDxtSzWNNKl/r3FW8MenJGADz6OO5cuIhx6o41
VTSoPC3nFpimpzq7evJtYkld2GhO8IdIP7pJ4sQe6+Fxj5xVioA5mCCh3cV67BgX
SQgoFSUrXGAV9+GEao1mmQ8A03bTCLDe/aMpj71jDyub3r1q/IzkiutcpqN8ic1N
V1YREL02eUXELvK2vxEYCw5v7sbdGE90vuNEq63BhdGfjTfiduDg71RUoCW61wEU
djhynZUWLRBnDgClJzG6Ug6IZg80S140IxylWQgS1RZ7eCloXRvymGgK9gk1Csnp
DjIq+/3x8915USJMysvnMvFydSfpUIcWXSNq6Jth6VA6PgMGHOuIq4QejFm/Isxy
Ghm1Zr3ck6WfdHycQrOvq2FY2TWpdyUJ9NUEakdd3pb7XPCMUW4wzipgNxUG+dO5
Pn/5WWWHxPjI9tTpvDj4xQYWAH86/FZzo6QNb4spccbAlZ/89DiSXWgrCdD9lNl/
WD9r5EfbYsRWrKRKAHMdqFg8cBuCeYWAl0KHkQaKEWi2MZHBpw0vhD30cxit56FF
s1yPXJbO3CiryAfoVJ+wyrY5Iu8I9eeBAlJzUbODKO1nZzgSyJZLKFX0d2Oi5nJJ
dSZSt5wBpfBwMDjN/Tl4bXwFZ5aB4LJSsXY0S1HrptvpFOOvLPQL71yiWuC3vbI5
foaTK95jmDv2Sg/N1LdD1VoZt60fFU4+T8sLCz1WRZvXIOm49lav+D5Fx3ZBQd3q
RrfGQIdOIq3O6iO4TbfqbG7MJPtjubNf2CyEZceoQu2kLjtpy7hVJMS8HjbBoNAg
Qhd7EESe+iYzY7vrXd+CHtQPbiFkrrlnUL7vk2I15xIT7RpoZmOrqAbK1zygvKKT
CnOkpsRy/QOw98z0ro1w8lDkqpXlcZcRVMnHCoj88qOQ+djIsyMOuO9xVtyPsQ5W
CEzE9Jdgw8NWOaaO6HNVqA2MrBsqkTuzJLJub1y1wRF0/ruGrxGWlhw8cb8ZVE6j
KofKG5V8YLh/MLzeJDJjrWV7wmnbQ2h6FfBxT7o5ykAcjhEmgAef5Sy4it+TXh14
TsutvDIt67BTvfKa/kxJmYTCyqjycpANoLL6gwHS81t+uZSIUrJ/s81vHn10nUWj
I9gXPvpniqg6DIV2UIVXzpib0CCpSsKLJ14MPrQiZ8hYFKSrQZ6OM8qbwYK4NNm2
Kte4q6Wk2HBvuKttN/lhD2J0ahrfROrK23jcO7xO/O5iU47pfmkYBlfZu0jbFJYr
Mke6NTXLfcarU/P2xb+6iujIghbKWVs2aEkYqPghJaWTfpAn25n7SfL0f9ATQbf2
cuUcbDTylhBzeWE46XfFYAoAUeyiWiTQc8mLhhlriW+F7FrrjbUmK7p3UqEzD1m0
PYTyt+5vfy37ZLmy9wRLZ+LOyTb5oSWLkDDnVKjrLr0NBbp3iyr8k4y0ExShVlaq
xIxLAU0nmpC3ZJoCRZwMhYJu8zlUCA2BnhEBeE8i9wtkTROzYmOyt8UfR12bdlgo
a/g5f5cTBBce5caVlTwGzXUoeQvxYmw8serxc/nPYYzgXxec1tXc/zj4Z9mc34VT
pvGBemUxezIiplG8tqAQ8/HX0EytLgEbOChQsQ0dtxjiOmKT78VQsOy244iQ8W42
aSg4sHTLVHQR/1Fk/9uLTA2FDwkCI8ctJWrD62s2uARQrzCdeYyr+GRwd5ZGPy+A
UvnHSXpdqi5+MnQTNdj0gjxmSVZ2UOzmsCk4twdZgIsf6SR1BgeDrz1toEocaG+Q
uCZwbBdgq+gPPe2/Vn1BGkbDX9vYcEcqDOxuVd562LfSH97vyX8DFqmF23izcRDY
P8uki7uh5GpzkUcEGwEKRZX9Xn8CRN7Ce29F92AeJAXAqYJgDtiRspH0naWsVNYk
No/VrexnUd8jzWhYYc5RVMWQS96r2TrO/uvDQooF543bWkFNoaXiscLDzMkNWS34
mDSsxdtV0Qx8uEj91QvbDXRB1vi3zfDyQY0H8hKMiDSoX14xxe7dp99+nMJ3YrEe
8in40UUCewhqnGzFTLjUmKpqOxwX5zAl1UWAUxUhUQ/koDZpps5qkDeYp3cJTflX
nh/gIvrkbZh0QFjzcCaXml525DVP0rt+SHHsBb5lDMS6saA40LGgQqeykEzcuxpy
3FbNXG+JsaA0xf3lN+vIz2bFZawgvA7GT8xWr1BxHLYktnDJ5KPXrg7UH3fZwpWc
5oxzyrT0ekzlvape/zVMX4/O+rlYhefp24r8/20HOGUvyntEGkeqfiLSrjhcNER9
azGyddY+tXu0WBs2tN/6aF4viq41eGZDtRj+li5ViabGaNB4QXTvAo7BOxa/UQCu
Lg5/3hmFO4dU7Dnlrvzr4tHb81U8ePiNZ60Ub3pIsq6qwcjqCMxYoMs9PiHvDywn
M1uP5lIeibSCl9CNF+kfBkHlZah3f7UtutBDsNoHGdJKMIQ3pngG2ZRCi8P3WMMH
a4Erw73ocP0VgsrdhPFbKikb61QJa59uvPt5dZBjVHcc1+azz5qTaI5OMFcgNWQn
lwERB68lMENV6Nq6iuGSlelmTxHjG3pGvigElc65WPBM6zRWQ1dlzpskvpuzFg33
F1E27v9dJpDigbbK2b532OyrdZ1SBHyGrFDqQj3vIO1DeMBvb2HPZFijHuAWMzE2
SphPhMrtgMsJANicgI/PU5xjGmAeZhe2xS0/Iqw8DRRFx+hjO8uSI7ytVRt0MuFL
E600UKgZ4y8jAmZeMBMgtOxTDK/3i+AFC0FMZ/fB7UMw9qod/F7hfJov3zpZaqRn
J8rWFwwvck5IZ8OtekCwTbGb++0udwApbWUWiDPYxJLwIWSOgmUCUquVn9xEtjmj
vFpbl66n3DrLbIPJVUcUglohlV/lAmyAo7VoN4sdL4stUwtGMK+7yj0H5WF3XMNY
PdOKQjtkqcjKvUGe0ZcMyASo4bZBaE0QpKpWB4f+FwcoVMBFGK3YIX/Dy361aw8e
pYQVRE2fgZH/hJpg3Jq64QX3M6Z03Qaug7not5mwOKIvcvkdzFoZqFnB18wB9Q6B
BST4pBxbN2TMjZSDVo4+9ZRgv4lw8COxT6kVwBe2V/kJikk1ZySFzQRkeXyFaxno
aQxWAbxhHRf38VexdVLQdb12KNO7Xm6U/Ue1y3EGsWoCUgTQ8cvW/JEvoMxn0wU1
E813WELBPcP8DRmwzeeKCBua20gngi79fFTguwwb22zfnp9mZlsqJSmS1mGPgv/g
2dqZLYTxElJSLT9NDyRtwCcPH+xMIGNeKo76owgf6AgRYHy72Vit1iR9S9I9rr+4
jzTToYalnE69RMpirpHCH9Jr6fFQcE2RMTDqR5rM+13c1SK9KOUD5poFXqFTejYV
aDOQTi4tHe+usPgZtBMlSMe1CqC8bHh4MAfci7x3sSxLNKdVWdo6uU9XVHS8FZIV
pYcpd0Hyk8+l9YoRg5drQWe3HEEnwD07S6I/WNu7Es3cEcrvCOk6lUqtEhRlBe2K
vpEHHtVNrAdarLO0xu1FtjDYDtwF4qzZ3iOgpmHDLJvPsZynmd2MKwK2K22c6etU
6hh48mJ+qSon7VqVx7tZ45M59k6bna5d3C6A7G9bcX3sO3ta4W/Krqt3kl56t4XO
62YUkacI37jImDtfIMhKY9Mh6QcvZLg6EdvZc3kGkunWNJNG+pvvrMVyAWw5W7Jr
sdSwXOXiza2hUnWS+/SiLhTxdVkEXVK0RgWnoJ2ku44+4RuWRD3mleJu1p2uUVEp
qEW2/JsyAsP1YwcoN5jQNMkOU22w2vtVVBNd0t8xp3oVQtdZwGlTYkAAU1AtoxYd
lJPg4IVi0LoyS1Jc8Kjn70hrkurv2mM8g/Olly6RM3dmHMgXbMR/4+wjjAHCnjvd
xfuHSXJtkM3Qwwek9qd3sb07CQuWr+nzugVx8M3e4iI+enWqyt2ne/Ak0z2HTrmq
GR+4yJ+LFnziGGqaLXi9T4vIaI106lRGumqPhNeP6CHiWLbxk0NMy8zwJSTLQ8L8
eL8LrLvNM7qECcq6SAy0K+4YbHREl/9MrbDZ4jRbgXifzGotFpkWsTAWmzoBmsBh
UP1uhhWelG9cfnVoOCmGQU8irIqJyI1wpmtss9HkocjSOxzt8YYwn/YPXxYZJUUE
ABcXD1D3zTWC//hXA/nnrIzUVANgXsnNw8Ec/XkpobRHC8ld300xmJeuDxoKc6fP
d2Ff6CWI9CUuD0Pid3HDEITcVtGZ7Num38oy6Xr8s/z7OFxp8eI0/cAbdFsemC9m
GIg+Jq69B3AzV4HsnujU8BdLz1ufqCdATWDtA0dXK4DdiDT60MBkCdNv5QdIxmS8
9gESTktlyPk57WR3AfbGQxq+NHiu3DXHeYOiNaabL/8LdWqrNkYYuuC9OBwiEk5r
bVzoS6TDeIXdORmXtXAOwh4AeOIKzF+R/GDmJC/eVBFxcg+cD0cYYio2+SA5+pAR
FKM9jVgKdeotQxN+lbWXsrRQRHnhK7OYPbhVaSGv0A2kfpLPiIjMXI2rgeAM1pTF
Y/afapGMyh2jsHeVZsiUZg==
`protect end_protected