`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
ddtXksX2+yylW5zu6QL2Lhnb2d1sD00763mmSITNX595NcHTEkwn0zB1Dry37fOW
FufOhVzEJp80NC5qZ/+F0Vk7Ik02dIR0elf3clrjeJRK85K4e3Hoo4xn7YbFUIms
l/8VZSb14+JVGURjfswrIyCUotIzlzVYZ6gzoZwDXIi5gQIBf/gI+KxNXPaKV+PQ
Ufys/12rjO6aI/pPlqSm0hCvftmBcnezN2hk1UeXgOIuKZnogjOsf0iJVX2aOOWE
6pD/psybjbnsNB6kH5uFTA5frkzIzkzl5d9+YDm9OyC+k84E83I/7/j+rk4L2dah
QJOvksSIzN867/4Qt8qYTQ==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="MvBXkzurAa5VTw+1JJ70nePUfoQXBvZOku/SMmg4TwQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
oRtzZL4VJ4iwysPsC8SXYCzXS8Fw2gtZTOskLcDV+1B9Nzn1zTyNtlo6lNICRmmK
ZRVu2BmCc2G+fmzynYlNTnSa7C0Cuel6FYpxCBlOuk3OF2tzAmLAuDyOH3Z1Yjzk
a0aHuoCdIRKv7BrZCdALt03JeUmXKPdOmIlkVGFl8yw=
`protect rights_digest_method = "sha256"
`protect end_toolblock="Jn9CQpRhJt4rnzZPRk+dOpzAubz7omckX1MrFd4p81o="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 10416 )
`protect data_block
gD6l00tciPUa6pDNTk/+tzLxvdHE2s3DQL3/JqqujQBC/Ei+vcAB8wM3doqg5vTg
mdfn9XB1bLOis2CVSfu295W2DNwHfMSTc/8BhCDRnTlLIX0UCJs9Za0+LoM0rMrV
T7EjVWppbP+Em6PkVKCwlmIQ7JKaifJ+Y+kjw9HCGboYo5074hY+K/CBbfsBQY86
AyoN0MKhsIx+eViNgnWjAw/QlPdiPAswm27LDiDhPtMQIY44FEcHTxEUdh9j9Xq5
rnM5429uT/JnQ8KqS+aqHiJceOKpKM4gq4hZTzhikHWRJY9/9s79PEcxmWKesN6K
W3qEljsH2l2Q9dM+MKhcPcbt/1byzRvjKOg1sXekurEVHPeCLvwh+5Wye32YKpCm
N6/Hq+ZGuWf3dAWlEUxR/lCKPwW7OScjwjEKDd6xjXpNd2KhSaHt37fK8TlTwpNr
FVfDtF4T+x/klcKqBHEp5215VoHo06UZRR5xzzEfjYBm26RjGOrN+j0aVCKV0bUS
0ApK8p/BiYGem5YrQ7iwLhKDwLuhHHjP/n9gI2ksanS0uSUVa5N16T//al7R2Vwd
S2Wk2lsZffTmq7rqqI2T9G2ClUP2j0UcAml+PljsXQYBlmkBMyhOGk8voTvWnA98
twogYjpVW3zRqqdEn2xzYEY0wfMzivTvp//wWH3tK+o0Pz1IkQaV1kLNq/c8ybzX
3ijdFHbufGOvdV4iobDQHYjmQ35aX21WR1DAqrTGrradpM5kbS1xU6i/wfFsUKth
tl1BwC6lncxLdhcSaqUdBV39MvuoZNe2LKvvDEbodR6dKU83OwDFCcexv3usUWNL
4M1N8VnabCq/l0wEilTJDAlBirudB/aYrOwg38i4PCMZB094INAyuhIBnAKdeR8U
hQuATSDrWSiqiG0+TMLo2AIzoFsH5D9p4fh8rW1dmyKZuzAjBs8YxAzPyMOjqaxV
wM7zD7hRkGXcbrrceUaHq+w4ak4sthrL02Mne3BdF7LkymxT1I7J/KxXpu96XBx8
9Oz5MozZU88qhFPAJgyf0yCYq1GyVB12rJLhviftvKRYLuNLLELBdGyAlNP/n2lt
u9a36WIB1GtFfuFrlQtw+6BungEIeHS321hNU0roxV2v6LSNtDw8tPdANnjDq/DE
gjmcdfeGk4JzEeuh2g6kEby0CmLFMrWcaOg+fSFQM9hqCPtyvjiACfu3peYgdvLs
EwIuA8BjguF0Yn8CLAIjNHSWmkF3ExkswIKM51+i5rHIcT8nCwukuZU4iGeL+ylI
DHMyVmY27OkOPtQbW6Yk00nSnYOZBUydob+m/07FW1lOgCXptm3SuG91D/b3x/R+
jz2tIAXmhOD8oox4i6fQOvgL9s3LHLVq05qooqBQvBVTRJsGbzxsThPoACPJWmxT
CC38hLC+X/ckOGKdBzckxYV1HVx/pMxAXDFxhtCDs35xPlZHKGKalOmjPTdNzQPc
vzR+OumLOGLV61vugL/L7gURfKLy9ITwP0vHbP2c4Wdb+U625/8RFbW/7S8LzDPf
RhQPMXKX60ebOIk3qu75dvsHcwjayiqVrWM8KIIzMdimBZ/o4KrLgBOUZbp71T0w
xtAtMNQiamnCBhE1LledtDl1fO99FKEYpqK+LMOYSx4uzvDS6cVU1N1SvcQP1e2U
bc3/M+ifay5U4epMQGpcV/OLBRIg3yDRiAs0fzljX8doddfVHO9Zs2Gwadx1+N2G
CHdvxlzIsBcjjokiOKtJpVIwxevAKHssx+U577Dzz8NQ5XqftuIMbsU/cMLEH038
VR0zGWDMHmUCO/PnUcp7OSLsDs2FLKYcRJREs7Eq6059uTWgjQTM8/XcyPj3er5O
dEXSiXaiKWeiV8GBF2X2iIVqJVQBsoAWF4wqG4uiQemF6+Rc9nS2vluK1H3C8aTt
xP5LhYggslV4diGura6zn9XCzuXvm/kUWnKtNBn00Xfst+0aeMcVKLxHdD/YU72i
N4Xmju1LbYzKAq63axUATIW/TGxyGZ7LFdRxx42G0NMDIN6x2orcGi2y5fG0i8bb
rAvHIkbRMhnWuk4WnLLprINnuAQstm1u1XV6q4estg1DDUK21xZykEfpe4cXnKAO
UZ6EQnRnb+LEL9NcQ4FR7KMewfw8W+0VonJA4BB+93DoSYvusrOC3CTvsYl5Ktri
MlTZlEIeQxz6GTXayX7kkwYi8pZmSkR16vMm2Gc5EtNpsbDqYodnpmAPVFOUlZPv
nY4sJBthed2XF6fjNETopFW91OnfwwFU7VFx10aFKWOqWSFyfV8sMoxttqiqiQ8L
3wSWpeYBy6E20bY2fMOsn+LrwpYY0hhnGwaiLefFl4YIoaYexXCQ+H6TFPUHX+rG
UEpakGm5CNscJVeatSSPrjHUa5fxBAMqrPPbdEllEAa+04TkJQzfZB5/33NEprsO
+mUYJy62L0RZZSiW+5jd40nY6ygGikPeV6woN6VCIiBpbIOBTcThAz+Jcxp3dkE6
OS8x1xV64dQYp9pOw3H0WlcTwt9nxyz91Rf2xHOGueyuj7R324kLIMp1zJOo2kvg
OuohIYj85uTcUyYkvyBGH9fo/cJYjAtayoKLARR/gu6c1p+PfHeyUyaymYXNyX4W
UbFyK1EoYZpncEFj8hp2/UTOmun5rHewxBNG4MchLZOOVEKXCyN4O7h3K7FdskUA
WTH7eidS4KTgiYjqZ/U4GBVK8lV/v4ncHXuUlpWlxytbCPPca1fIPeRBzRzojTGn
MGnvaSYyIqXb77Cuuw8nOp4f4qyx12DgcNaVj5ycND4blC+RV1RMdpUJS+TJzs7j
JqjD13Ava/YSOWyAUSuMIHCrFg/axQpigGJX0mtevHUyJeMqBKlv/CUBsD0cInXo
W86qgD3MUWMuYhSV9XSta3c+H3rGC94DYYlx17nyRNBqyn/nRNMkPTPbQ0d1p6ES
cl1YQT8X7GxPqHKijwoFY10hI8Knl1cI0ob3VHQ2AKxH67cUXtVv/AmvA3a7AnZ0
bjp/TlfdJCINPXbuUvEbHc/cMfkVNOdGHeDZYdJbn3mk1HRSJ31B0OBFSuiZngy5
3SaIUTK6xu8B/2hAkwG/Km/DsV1XU5jncwsJNR9LGewJUfzPVjl1thoz35W7x459
EJ8gE31ceqNgpOfAuWlrnd/S9hbW26gktBw0GGlniGip1CnEsAxpLx5EA7WQntOD
/zs1NU7re3XeiVEo0JAt94Xhl5N69/UDY5xO0vA+lc6Hg2ILUDcgZRgQzZEsCedt
j3h7S4EOl9lMglIxWEAnfk6uvmFb6vJbjA5/eVdzQfcnj8uXj3VJbvIJAjoAlpkd
r7Z2lvOI0PIQkeIlZ8TaXCgI2umTQVtmuvkZ4u4RV3VA2gM7jV8bMweERKDikFaV
ariQwcl8IYDH+ED04PN6pzxrdx4Ozlwy+enLL1rxWDsZWTLfxeDVqhdB/WlrrFpJ
y6WcJzpWA+4+nQXbmoC4ShhO5Vb+tz6D5ttVz+fRiJrklWBpcmggLxVYE8nN+4uO
DzrjnyR3ToN0VlMYhQKesW3N8ApdDabb33v4futDOI1BcEsimRTVjaotWy4pKuKO
oYfCxTM/DIyovxPYbgVMOTORsY1OBaeugqd6/gOy9F+mI154sHbAFaCDgAOOCpDf
7xR0t/7/77LzR51rL6kU0peQJvhlMBHaM9QwB7ZgnXUkbkDseQaugS0mgvlleyuJ
guhYAvfmpViq6oah6vk8sxoFTG/4KwoJF5F+DVUdjw0iRp9SGoTsuwoPbn/zKG0U
56yg4xSQXyzauxqcJZkNSlDgap9mbX5XoNRGlaMnM2/1PapwVfoBxVV4+rI3xBlF
9PMS3TMZHr/zTLVbPqSI6NC6iA7uEVd9QXo3KDWlOQADCN+iCrLFXr8TIXbsLjvR
RVDF8BOtmyWmwcfpwF9XPbFxBbADWR9O/ad9iC0ewBc2z+c8pzMDSV0qZ6m4npVB
BxSh7gQbMYMjOozM78TE5wl7nwfKYCEVDTK2v7+p17zwdbaXMUD1cEp5AI85vdXz
f48Ad8Z+/ILRqbSf7kOYX5LviVwITFQ0tjjEEEWGdiUuyjrB7oPDz/Y0StAkruZW
Z7D4rRY0rKFp4rNY4qEghyu8MlFCW0ojP9HC4sM9jZnASsogqggJqpLAFZgUPVWK
IUzHiyWsgURKV8hgvVJQFRl5sx+zFP62+qjDQfR1tJPptT9l1LhDXxJkZ/fKYFY0
PoElfrprlCBe1lvnRXmiCcxJqBkjKYfcViOIOPzgupbKDEBI6YTk7FJ65r0UJsgh
fJyYiI276d3+eKWU1lxXEJiN1Tn+RcDe7Xb/gV2KauwonEs8WkikuV6LJugeKVPI
L5Hi9wAycPRNDFB+5RPQjOBEp60yIqkXHGR8idxKtvW9Mp+spebkFf3DRothc8og
kje9KoAyU5UBZ3xqiPYaAs+VjHnFc3itPO+g5UMNODLMe/8994YXGypuznpzjLr+
9oiCaM5oBDrXgC1J3SmEK2rGjGz+wlxacYYmsR9BBFfZhrzaqUrxMQG/r0clEsht
es3kFvEJSIBkozvXMG+QCamDDHzZlZtFOXlgXk0PsFSVaLL2/h6aOb7n2C5GJ34u
dYxoI/3ceTAuuCtpZIBOVJrGkRsUrE+ZYMQeu8m58n2z7jBQohsmpvBHwfzpudI6
rAkZ1mykUSLUzIE514L0lD/4fAGeeiWksbqgtDimvFtYMSYAs6lEv2fdSQhPAa1v
i787nxOLDrpsga9mfCskICyQYg746S/i0e4AEBzBgflzrx/JfiqcOYY5kaMtz9tG
cFV7vhCZXjOZ4T3q3Iht9lLw/7jnmGrP9IwTpPTvflE8I2vpK+xUKGFbFn7gV7QG
/myrHz1CvgPcCEPVbWxeNGwT6MWgf5SUhXVB+JO11fEy7RhKmPB6GcnMYYplpFJr
n09G2JVuXt3bGvil9AVqwDAbKk7ZCzgcUjy4zAHR1eUxs9uND8Rz9LOC4Azwn5O+
hTwUgscHTl4cG44YPxbdor2WFZaLLkBLjHqNtD39A4u2lRLncIrZ92Wz6AnVWTIs
qnvSf1S/rSkCYr+KqkYlvZFCVbDGAAhvGz1QMqNwItSlJcJ5f73cJaymyOOQxEKY
MMCOfuroUZqsxdqQkfME5jNGsIrgZJDIKKYKMC2rREZbfnJbEIUIJ+dmUUNQTr1p
9p5lM4exYBmfjz70WsTVOz2ZnBbGS0TU4ZDSVR+03HKxKGUuA+ibcZGdzrBBCNVp
iyKJSaQK9t84zFU6KwbXlxdu3vbA35vkQGc22YeG//U0wJBdZW82ZnSou+wIYAby
Fw9/f/uhv+lOw27QU7sWTyi5U0Pja1yuHNcrA6/BXE0hQRgpDCBpwV8lSU+bfdzZ
Y9l6C+VJ9qXfFXcTx5gS8XLEQqrD3g9nj7i2z5cNuz3eT6efmWNr9gs4DyDLnSNf
FNgRz4iSt6J8a3OvMciRpbjjnXBBx6M5pm3qiXfe3a51BD4pks8a2CWecy1ZVdfd
VLWQxf9e/VI+HTgs4fIL6lOiDmgpbhmh+S8GbNneO+2lIWn5IjS1Rtyzil/hxWEx
CQabGZRL1MUCyRm3RrUnlbhCfVfTOD0NUsM0223MReedFzgO6VAPxWzbJ3DE1hMX
07jAIuCarVR5XomLt7DVY2gexpb3PPm+n9GugVEQo0G8PzouJrobO0KAxZqwK3GT
YojKdY0b7dX6hfTUZNV8dwifQw6nAavqhuz+wl5vgS4i1iXFhSdCgSPUyxGOn8CW
HgaPt5cJ8YfS0Cq9DEuJH541APWr5HBg25YKxKIhUGS/tX9mjB7i73tjuH/KK2to
nLf6PBn+IqPUcis+bQtNZBB6n1Rs/pvrmEvPLFpTrQG9JwCHp9ZJ5t1Tbc+vJJqZ
ZRC2fj2r5qmrZCQzEyElgAnbfDp97zQ4AJBY/YoxZuJYeaJnvXs7AaWTiaaDf+33
+AGhEbgA8fwdeHiP8AS6coHB9tiG0+3KqR2mPM/CCxA0GRbA+OcIFlry3zybT4x6
XEDycJY4hb1keQlHAcf5yeSXdC0yey2iz0WUxk2gVPW6IeN5pBd2+/sAhRpdC/qT
GJJN/p+saRWLYd3oMkJDrOXiswgntSSV1lOO+9tBM5XFFrDwpZN1K42ZHqeSt14A
gBAq3EIA0tYYOTJYdO1Ni4M1avJPQP+rH0BMGxoqDvuw5Q43adzIVO9Rd3pv2xlp
1Nh2wt+Vqpj6+TN9mbpZLxbOWSG6Qlq442fAyG0+LjcwV9rXHmag4oy0d7KnMveb
8wIgHN5rZOpXDN8hi6jqHPKsH9n+2YC4J7aG7bp8qkltl2Vg1dUN0ulYDrmzFHIx
+wksOHFcD9JCK9oSMVGNgbLSWuQ/v+fQ2BKNKFhGkhIhtUIVl12eoKLB3j9aNizf
8mVt0w38tI2Il4oAt8RslPKXS7Tkah2CXBM5oisZEc8c+CkGFuvjesxLNp6jcrFN
VqBObIrd1TMuNrVf76YgisC5qE/aaKt4Hr+2e3Nf730J2f3QUOSoMbGKGc23In2r
vzoxfCV0jUA6rGQiszJIEZnZrYZchfA/Rflou/K2oav3tkOKn2fOlfOD7Ht2Z6y8
Qr+i4VLkou8n6ytvm4Yt+Dq8NeFyEvY80+UAJ3kLnlkFjwytn6tZvy38OpfBGC8c
hfyxSwGjioSHvSOq8Nk3o36jWmNZJdZFV4DfxCtxeJAShsxyRF6ms7lkLBTYr5CW
1kC9xpGzcNyaoCOUUIJpHOEbJFLmrK0DTWHoHtJRDuIhxpn9ozQf3kUXbGessuOg
lWEEoonB5/0VeCP7b5QOhLa5j8d69ywVPMqbtzaMicpF/uvkgXLlEtBwCcC1UOtU
HeZ/hk3VmN9bmMUTr2Xvz/lZQMNhI/BUyyEGR4OGRlnQWUJ+XL17sVTR5L02mMQ8
qNqkb+RwS+FvEQWAnkX1pU/i/QW4Vb5Rl2GZpSQDRYDsbnIlWk9pkcZYEQdqHigh
bI+htitoZl2yTLgzb4QRajZVS3VIE4lZJ4wLpj1Ap8CoGCjZf9IjOkp17k3TNVye
8RefDyxo/p3+hham9LuL8tRt6Z2+dfDbYQqCysv1DuXQG+9ZFNx1U1LXWYPu3oW+
DFRgwI4O47cgfnFD2s5BWm29g86bKr020jNEgwLa9uIR2FpOgWkuo0eH9njplEKn
6VkF/84hTzLR+DyZnZ58gPPkgNmk0vsM4+UDbsPkXPrCW5nQQIbEI+WDY46Ky/vv
QJcbkHmEkoU92eISwVRz7cBkKGchePZgqEc3SJ+QI8k1WkW+b6RyKUhcT8RD7nOd
bImdBxwqMSTsz80VsrdW9oFvqn2NfE75iZmJLoX6nO9EQXJeolfGiZ67LMuRllVV
kt8TR1PrLoKk6rR6NSXZfqQJqxW9rqK04g5eaJdfyLbMNF6+WnT7QmX8lAahS9XU
aUozf6jnc2KZb4PKWss4O0dNR9ldrZUGTGX6jsdC9WctH4gXS8nGNFUDjZmGrCM4
zvajk9ItQf8S2QgHJ0IPWUuaF13m9zZqKJ0l+/SYe513k4qfu7Z47626+l+8JfIR
wL1JBQ3IUyoAYFL2mm/3SoKYpAlQKrMe+gg1W3b0dnKjZFL4eIwwuQJKXg7YAhSW
oy+Og6SG5fjYKKMJyTD6TNEaPASdBTMAdZp0wLMP1s8H7jm7/QgDDya5HLqpTXZW
27aA+xCTAMxxbHLp3ZyuvV20AaakfVLHQUDiNIb3ZM+Nro+Q6FPwPxg5VLUCnLP+
N3jRWfNhVmX6L3TCv7XyvH7zaSiOm3F8RcCnSo/9IshiYnPs0OmO75gYcJY3orjK
xYYB8HwBaKZ3ruaWO2k1SJdLn03Ux1pMoJM6KnjWlfb2NOtjV3JIT0Klnn3qiy5z
rjpu0L7RTBkXPItt0OK8BydgpnDbsWGeWYoeBGXTLHFE+HtmpwwEoK4IOLZZJRp8
34Npjj6tXFv/DvsUELtd3706IfIGcupQ5zoGAONqc3z46T0q4mBMcSaVp1pL9wnf
27ufN3fVSeeZTie01e+VBnCbtg0EX3M8QBW9LZRLrHDRElyWvWlUQfdfXvAJKdPy
tyjyPDJcK2uP7oXgLy1jhmcUaXdKLY4uQVPE90aI25O4YTy+bmEXSHeVv0RSe9TG
Rjd54Gs5V2oo/xyPDaxD5l1gznsedsRKlk3QfvlxNdC8ArUG/0OwS71n4lSZY3gH
7C+AKHwsactb7RA8cDUB4lzrLIMolDLHEj7AILG0eWymO+yXKjAxkvKHVasZ7fJo
hvG9AQ1eNcn/z9QpcJY4ktpo5ICj8cV2WK97OXpZA9UTbVzsLgj3e5mIyuO8ducD
Xh1pxhr5tIKdNeBy9tw3CA4/HLbLQEWVgHVvzgBC9NQAaWGXlULL+x0GKEmx55/Y
xJ9+HZ//o0BmPmrb7J5JAP+CPhvIi683oT5T75P7CSTnvI6avbga3Fv9i/mNTZY6
ET1HHEc2m+rNwbryJapuCCGYua6t+eyHGC4fVyQOSA3SmaGD//qT9mDg2oaIpuBO
moCbFbMss5dOEAierYOFAV49Tfyat/gSoVSp+VRbZf+1Eibdo9oFjwnwh9EiRkdc
BQqyt0JZA1rHbqhBIZMtY0KdT/BImF8A+9yij4hKmkkEkY0/G7vERRSZqTK1L8Ch
c4kLuKTCzPPHrUVnHRZKbgLwlXDqy9VZ/ETHc54sgtwO03CWTvQG5fPNSu2ZpVUg
ydi2mXEXP3euEzrJIKzRSvGF6kkKC1pj6YvnZmeHuAWEz82QVLnwya/ZJFbXjlKa
H2ywRLCFaRQrK2uw80Fw5RA5OAfQHjo8PmNVvXWlJvsMuz7UY0n0b9i4XxNiwcZf
acmtQDc32FYArEk2QX6ha3Wce8hvrjbDxNHeUuLaRKjiSaa80pRophAYh3lVoQZU
zdqBvIm3uajK5XbGScWfJDhmvQhaLs/BUprSTwUAHDzGMqD/OtOujGuEKMrZiSrR
JW9H6WQFs55O6d/QsFBZSHlstcS4vkBOHiHOpiraxmhdMpQDMDmVUtkRIiy2shRi
8LTptLQAkjjs3DAHrzz1FVjQ2pMJBZ4qkHEiLsCkfNJAFAUeUoLw2np8DZ1IPCwZ
OJDy8Hit1dKZnOITCVvEjO3lw1Izh8L/+D2QZLclr1XcAMyBWK4DfzfB05BnQSxj
fzB9O9vDSOjSA8FekoLeOU/iW/cSbKt5s4/n1umc5b2/wCrZCpH1tOKvy/DinpHk
GA9ozPIWeiIh7RdLuPbem9bRztBDNcRFw3g02yuGHY4jhMm2YDpJtG6z7ypC/rlu
/o09Yn81JThL8u7sKprOEdvtbf9nyB+mfquaoh27Smpxbyt9rLhjSnZOEp1rlLc6
7BlZyopq8uMfFbO0VxEaPXMiQKq8FwEMncsAqlBEDET9WVArENgWKTQLlLNdP9SQ
Tb1bRzl7QQBFhZ6ty77R/D8dPdZzWPuEE/AFk8yf1t6T7aaUEkATFTFFPg1l3F8e
oAwAXkERIuIzSGSfH1P/qBX4JK789ROQgFsfNdFdlIMTXMnq663VNGLlo6C7mBhl
Eagjv/Q1vIJz8QfaJEnRRdcFze9OGjMYG+FiQoajpS9l67aVE4joBmtG7hzMhPTN
erK4HDwkRHesqbi/dxkU/b0pk2oU0hQLhKhv+o86N2UJVFeG8WA1jOqkE2niSbnc
45PJTpu6nTYu7PYWshRy3CoRdr8Beg1Q3hIljFCRBTEJfqQj3i7r6hq9hp82s6Ta
UnYaE0iI5B0Q2WSTmMhKoyB4jn58v+1tUmhC3GQeDAU3mw84IbMnMepBihZn3Ucc
p535la9mtIB/l8Oc1cQtAlQVxZmoHaB6Dy6PcpiMDUr0RNNeqgJl2Jl2+/eXx3jc
EFT2p56fKuqQNhH47nVLrJon/xIfRQpn4OAh20notqBtnql1KA0MRZToaBbr7fS8
nTVzSIEmNVs5JedFfkeEEzVAx4Y6tgM6/0cAO1VzVOEPvMnFUbd+5bH0KDV/VT6E
ZR+Qo4MLj0rerTzKeNgSCMfIaazG0h6ICHlNUymFUB3c/GriVrseF56G5cuq5hP0
iU5JdPt6mXtx9EIaG3hAX9SdwxLH6lo1j2XRHqjflvJinkXQuYqmOSZT+2Ao6CMG
zpItiPqvZMRNxX/qycKrRO9z67i0dTFu+fTejWpHNc5ZQw5aNuoYKVG76zqphecf
x/pZK4bKBHylhzbwxwy2ZrH1TSeAUsDK9hTksQ9hVsuUABavH37D6ka/yE9coEhC
G73t8tLEICGDeQ2M8ceBReqNfvnwmuauqMtw5Gx7ScMC/ZN0ZXsEc8E73/7eEdBN
D4Fk0M0+2if24XjVXzFuVygfDvoa2qLnm0OBfn1xQByRTskoAgzF+kuBn/7OLaec
tm8jBdPBDp1mmxq4chwTXG4maao0RHTPKNRc0QPX8tM74/FcdUW3dyS/rGh34Fdn
VeErMvf9+StLY4PdtfZg4H3EwfDHY+e8i3o+zlIo+5JYIlEIr5ILaYYLYuA1oXCt
S/7Y1LjFzR/qiyD1QM6DGSMrAVlOfZYoXu7nKRAfSYPWijEaMpH6x4XKNTiYwm5J
SeN0qhvKgBRvSLL1s0G8ny0MbjeEDW5yAoIMzF/IAzVmHVn4InIQpju7iiREfZde
19HZvV+1PWu0Vqs0vrvUvatAz22wH2K+OrTB7Ksi5C3a/A61IvT0RxNBVZKHAPZ8
bVxBfAM4f0s8d411uA9rwU3JqAkxMkSluqEkCP0kAyyULToCEjJ9T/UVTB+q593v
Uw/0Cvq09h+WVrYtEBt3agbyj1w0GxLOQN162LJPeF3wwU5D83zXPa7ifDnJ7xQd
Zmk+Mf+JPnpbO7Z0D5DK53sBHff07e8IysrUG0mJytQkkoPqF4GCiLrdpZLCI+uS
J1AYzx0FANZqvGvfunQ+Yz2JNxiz6z3+8hVVvfXrIHfcmJUhrmIEC3R4DVeGD06k
LsknzOuzdPs+u0ZTGJNtZja9qDvnMkWKI6aEW4WADBq72GjdURnGSjGzUs7GsuYl
QxR66dDISMIMpKGPWAnjVZE70arZ3DeOuYUnBA+R5DcGH97CxeyUFo+Np78YoFGI
c+pzYWOTYggWm1CHffAuJdu8be3V/eVXKxzNX5j0nU84HCe5rH6bmCHCE+KyasH7
vmZcltYp6EkpkzT6MdKI/UpdxuCUC5I+5U+ABemGlFCrmrnTfQJEAVRYCK93ngEs
kA0joz1IJ1uMrxSl61su3MgqSb4UIsXMLOrh4VuegR88tu8Dc9yz8BCWnc25f3op
mwGe6kydNQUulYjXDA7Ev+Rlp0BLcGethU4EUNcte383hLwdp2ToZM09t/WNIup/
gcx28K8OwJqlgO2G/oGtbXeLLZslUml1WScJOG+50VMOCyfqLzZFKqT0TAr03/RX
fHXWqNSIrUzHDX+a9b5mIQwH+6aERMCEo9HJJzzLJaDUWxqSpbJ4TXXr7dJ/oTDW
XzTJCNgiY34h36qF9PwGv9mwiDuCCevCXaDpGShSBpTGdMcPaQgfBBMZ4nWcimNW
0JW7X3aU5+e3+p6EVOI+InENX8LHHlwoo/3LpSTmTMtRzkwyMG9SLEaKPyC/P80u
ywAVtoFF9FxkLP6N7etd3/1X7o7RMq9hgLO6lcb2Aca55/YVlyE7n49xNv+FnA94
aBZAmf9yi7z59spj5J5XUyUUmTwWlGp28aPo5yhte1ENIH8j+WpEvryauUXibi0x
iQGstCqv6KFm0RLD2/NCfZqc8AFlafcg5y9NwTJx0276siyffemdCTaUJp0nvKnD
Swv7tu7+od2wldWCs0lIbb2OSjTQQrzXDngr87w+syMQgtUDWUws9otp9Bz4x637
ybDR2+QuyDpSoVcVoCqToLBydfgJSBCp8qWNXASwz2Xcd9o/JY5cOlCOdlc855V9
36H9u5sA43axL2zkecMA0uisUOgVcmXhkYBb5a1c3HOBJzvVrQFzbQPAGzNE1f9O
MGEzBc30zK0a5D2rxY0ef2rvyjAvEsPMeHTAsv8EcO6r39G3vbCFOwkN47By4hoS
KaTVIwBpramAnnlccdYr7oMJ46Ru3+REPE8i4zbDgVLInaTqJ2ISFqEr+wHatBcr
uhVQi0MhlpAIbErwGhrI4Wyw3mTCi8aj9Yt/qencF8md4FwoiMZ/o/y0CORqN/wW
QoIYADvae9TGYcMaRwUDmaB5IwkQOBoLWwIrPG75lrsz6a683IEhiLDuHjil3+dN
qz91mUgy1Zeg+o9b4Rhv+gDTpIya9nsmdARiazikvR1Pbjc1owT+qKSaE4S9qQtG
PLrUYc5M7LJFg8sE4D3Y9zcNPXPmhcAoTXBG2Dzn0vylEpZ+AUV+bQb3G+f+2LN+
kyp1h6SODz8fnbsHhXeK0ClejksdrJBhEAyNJp+WGykMAG/P0lGiWtpn0I7dRfn4
pDB0x5bTZBWbGTVriP1eSUDA87ial7qeenwu2eY9VjIgfjCLfXpTygxiNUyPr1WL
3k0Y79D79raVjI02ulq6C1a0Z90uXZT+MAAi5eZ1yGboADti9KcX/xJEzN8vqIdo
hBZrRniscQJ0d/O5l6cMB0vwtvsr+WIka7ggVVWPZRyzBXydB3fqtEjgbYgtD0AS
mtXcHPKtLfcAJmiC9zGvn/0bqdTW7sED3u98ZAiHyFAHb5PsJBGiabCYiPyq2bJq
inY7VxCJqLuGVTn4es53nAhdtmqHEWI/TYYw/nPakiBv1hwHt0DjXqsofQZ5RkgN
sOy01vUi/GemSBu62xkwKv+H1O7KqN5QsP/gCltMy9CBciT6YBRd0gmt14p94U0E
UBHfFpuQK/i6/9ZeDYQvUDQf3LR+Z1TsZNFGS4oCXrsmSgMKluBz9JxWuZMOjCGX
1wK8Zw8zuGLfWP/PdVC+TB9IbiGMQ8RGr4cmp108IJhmjV0NH5Y973pzLDI29oAL
slIgjRp3RriheRG6Nrh/eJ98xktDChfDZ+FecD+CmaZkq8WBHHT2WFjy3ILzmf9g
Jr+bPRhc77d+b/Ng0a3y/nUc4necioHuTwtfE9Sd7TPiNuo1hoo4dP2dgwpzY4Il
rJYtBbQ2+dQWAX3l333m7FJsy5MZo1LjeHeQQC86PlnaNdvs9XkVM10J5SNICuiG
W7K5q1GIoYPEmEnroCxFgNUIeIZf+cbGh0/KnwRtPaZSZ4Rl3HvvnsPEvGUsXLuc
7bwI7+Jwxp/NlpMpngickczbopflaKR3XyfaQTgntk/XwYTydYTpMoSSkCy2WwU+
afDgQbP6NbC0HFb0b2GMJF2U9mYoZq7z7S1sJwWJs4jIkosCo8aELr22B7sfbsAQ
k5XivhCZQPjsqB9cTkCUPmHt7mhUrX57VvnAQzu0d21RGI2BA6pt6vsaqQLMTql9
jmktO4j/ftarZt2KUYds6n1upjKRV0ocsCh1R9p9DIDppmn8j1/fj5ibsyG6Sj3A
M59u02g2zvN+ZcExPGL6JiaadRdxxCGLtzEZmAUkhkcv4YvHLOQOW+mzU/HeDVuh
SeARYJ2WNqaMaRndg6/eVZ6QUethU6AHC0DtfSaRRKQJ8JaxUrJxGfPuZN7qeWUN
i0kqTkUybkADNF6N+1/+QEmzKRJR0IiR91C8sWSuSrCc5cvj4KCrEiQJ1u45WPg2
3GkAhe9VlwkL3s74MWMk45kqwHx3UQXqcPLXYbIlTQgEaKaK38R3TtOEehXUbecr
LslrMWAk3Gn2G00nY9qf16rdcO5eDKJhJE9T7U/Bf8Ook0MkuaMVTzvpgbH8htNu
XyT00M0a8QlezOpBJeyGIvKRCqwkQqpDmDjPBeFlU+tJhSfpfPN+N+y6VDjdbum5
iHPni5Jns6byXBOPHJZ4GRp8Rc5wUuH6kirDY99OAd4yKZYlHsZesOoMHlzcozFg
`protect end_protected