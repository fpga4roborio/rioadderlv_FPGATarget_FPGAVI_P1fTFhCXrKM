`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
ddtXksX2+yylW5zu6QL2Lhnb2d1sD00763mmSITNX595NcHTEkwn0zB1Dry37fOW
FufOhVzEJp80NC5qZ/+F0Vk7Ik02dIR0elf3clrjeJRK85K4e3Hoo4xn7YbFUIms
l/8VZSb14+JVGURjfswrIyCUotIzlzVYZ6gzoZwDXIi5gQIBf/gI+KxNXPaKV+PQ
Ufys/12rjO6aI/pPlqSm0hCvftmBcnezN2hk1UeXgOIuKZnogjOsf0iJVX2aOOWE
6pD/psybjbnsNB6kH5uFTA5frkzIzkzl5d9+YDm9OyC+k84E83I/7/j+rk4L2dah
QJOvksSIzN867/4Qt8qYTQ==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="MvBXkzurAa5VTw+1JJ70nePUfoQXBvZOku/SMmg4TwQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
oRtzZL4VJ4iwysPsC8SXYCzXS8Fw2gtZTOskLcDV+1B9Nzn1zTyNtlo6lNICRmmK
ZRVu2BmCc2G+fmzynYlNTnSa7C0Cuel6FYpxCBlOuk3OF2tzAmLAuDyOH3Z1Yjzk
a0aHuoCdIRKv7BrZCdALt03JeUmXKPdOmIlkVGFl8yw=
`protect rights_digest_method = "sha256"
`protect end_toolblock="Jn9CQpRhJt4rnzZPRk+dOpzAubz7omckX1MrFd4p81o="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 105904 )
`protect data_block
gD6l00tciPUa6pDNTk/+tzLxvdHE2s3DQL3/JqqujQBC/Ei+vcAB8wM3doqg5vTg
mdfn9XB1bLOis2CVSfu295W2DNwHfMSTc/8BhCDRnTlLIX0UCJs9Za0+LoM0rMrV
T7EjVWppbP+Em6PkVKCwlmIQ7JKaifJ+Y+kjw9HCGboYo5074hY+K/CBbfsBQY86
74rlQP75eJZOYXSBu74adXZq/kJ99CoqLMczfMeLx1PIuBt38TVqwU+qbkA03QHd
B2luSu0QChW20G/49f7AFfr/3FS55D7OkWH6KZZwowEBau0QFl5VJ4JjWMVI3djF
MQBhTA5FpMiVVw6kbKiWDEbRMqPZFgWvYfw/jeQ64U8ZJpN6GkGEstgzTJYI3F6y
dtk1fk2Ei6yU6eWZ1D5pD605kvKPcAS8zcS58aPI3oBI7Y9fBEfxT3odifrq3Dp/
irHOMFFlIb9PRv/WGzuj3tnN7geCK4RvFbVs1Csurfzv9dR2EQEZxkiXgAd/jLjN
SrlHOydtno5fp2vi4an7g5eue5y5qgFpTOadOPeFFKs2KRrWky5NBCurLodCCjPW
3leBQCOqgAZEGQv7Y0GqCSFcBV78y3SweSGG2bAGBhKMElFFy5VEzVgmmt6Vqmto
s4rGRNQKgi6cv3FVwcaWBkGn54UGU9vEs+TWvEdDWq2Jmswe2hj/fX8sz7Hl03n6
n6Ebtd3ceULLETZ7N0H+tU3dQPICwo1DEwVlK3Mhk+nJmSaJ8MmU2p+q7MShbNgX
Tz0yGvmdfyFY9GR0ngCQ2xEV2nlI4rNdV69iBAm3KJ5YCslPsHeLpWosWMjcrova
C1YYZ9znS5dftyK3HuxaINdLsNVYS29d/Ofq4sf+t/Gugzg+DW7Rb+TTMEqNoTYG
XoA0KzeYTnhluGDBvM0DIIvsjPTsxsEgMM/RYwkvrYKr6HrINWwjlCvpPAZW+zh+
PmWN1OmM44W/mXB7J/nMHzo3EWI9ucGxtKObq9kxD2v+eOB+QrWxPbYxSpwoJV97
EaRiw8PyHDjrAwLimvU9hdGwKrWOrbUuhoGEFwW3wlTvlSRKDSQToM4SblBA5YPb
SzbJ24YquwsbViQcjlWgeXhz8jvSLVmmYWRCmx9kS/grSY94ZrFwxI72QjIcQd/y
VStIplKvfWuI7AdLTQwLJ8TWLZyKm9uijlakKJYtCuiU+ouNISaShkBd9H7UHcVK
6J/+GekH54pn1I2Fcrc+iMNTAF+jFxGWOUxYDzlkRHYPFYlVo0vcfXJXV3jkEztX
YSZoEvl8nM7q+g3Vpx5JVfNAAYIUXU9BEUKwqIfKsiVxoPwvBrSxwjIO5gl8iCbm
pnPyFxtBPLb20VK/Pf/uAULsDL2NZk/zvI0fNJFSIftuCj5ztjtIRuGD7c7kRYaE
uVEL8+M++Ig7sr5A2kTJYRJguWrUPwJ6vHlcT7nJdZgFT+chfJg0E4Itv+avt3uE
ZQyEr5VJmBqFFXwJMj+S2c6PRLmdo9wS5imMQ5isNDFmDIPLiaNHGsZHY4MVyQI0
x74QBAddSVybO92psfXWRraCjM8XU49szcd3+pvIfRiwNI5lOgJEFWVJYp9cio7b
x6rVCQtHuEmtqlv+IPWydOi+n1Ruv+ptsk6tH8wLdW856ItISnaCi5CXfrFIPnxG
2AXCIfMyUCKnlgUyVyYfXlmQBe4T6rIknkKlTvM26o05kiF6gkR/LHW4H2aptNRQ
sGdFqz8gU7gDDYNKAL/WavGJqhCI0NZ9Ob8/wsgzyva690ogVfejcpI/mJK7qQrA
XkuOYrbtEAblhnGRkJCaevAGJDtFw91dNAQ/WTx23WGZ21F3IpzPywsnC0cQuN0W
joEV/mFv2sA7qmQVcr+h6yMwpYAO/rmWoV/KeZ1VQla6w9t3iXqHR52iVSk11jOJ
Jns9TVBuhSR9MmwIxyrX5A/QHnsN7P7PCe3L7zHvzpTR0OPF4mnbACpjuxGtwpTh
ncmc4VJiZTnMEbkbDexs+VhnKkdrb5XltV1UdwXB1IuoJdRSW06ZI3Nbe7QmjV9/
9bkPaSztWnT+jRT2PFnFvlve+SUgiUtCeMqbXZEnSMQMMZ5YWiKStnyhIlfrlJtd
dv0a5NTMJ9C66GOvonyVFMXDiLLDeKcuwhnByLBOVsJIbwiN3I5kymFAcowP4bV2
fuvGT0RI1xUGg7UIM6NjpEKeBPNKEIobnSY/oQm374X41+bueF5+0F1LPOPA5kK0
N31C90YWxikWw+R3VGPR0e3TiglDhJB1guhdSKAvMw+t2C4ZehsGr4adAxT4/gBi
ZyeKBgleIR68leMC/nJqF/+K0yyIvJFOciR4n3uOx0KaAGvrlqIgT4KH6sWsb8E0
+BBH6b2tL2Qcp8RNxO2wyVNBKz6cFZABYvC6yG62Iu111kMtYPb3y5kA0aTVClEB
pKXJR6qAcVDzkfTZkyQkqpcs/nyDPU31mzjubzna8QxXppJwf9z5u+RhBwFuy35Y
VEeTXC2fzB9qM/AU7ZLTRPGWpQlnlEcvKhgRKc/mVd0EbgJ50QNajOmagTEtof1t
k4foIIonnohF0uaWt59QPUlZr9eIWt7UDfaVAJgOGJMrtzpZ0r1q8RpPzQ0iPCj8
lSjvdd2VwUCWq2WmWONDoSyQVeJ4fv7ptY8Qzxwuf7V7iDeWqfRzWa7EnAALI9Hn
yrJCn7rjGLU+krq0STe8P7y8Bvyy4KT+eUdRZPkPRWaBweaD08QT6I9//RcS1laN
GMuNZ8uGyLVjdXWPkmxmjKWTZcluD6WmyM99u+3hb36MlwosIuzwKPcjihtJUEyi
ONbhnszrXxYyLq8BVqgMEzMuY8cJ05YEnZVIuQr0ZNzVniui/h+6rtwIRqayXPAE
lUhWp7AJfrTzf1/YbqqzZYO211aV8P2gP/n0dtgTgHuaIDxUhPWnz8bioNu7sMGm
M0BP4Eox69+hMGmJ09YshfTPyG99eyLnK/N/UyE22DYipWSBRR4/kFLP0aLk/iJ4
jyHSjh/4LS01XcPxaCSDB1nE98x2AgqO+/U0OAt8Ij3L/QJu08FJIU+iakl3Ib7m
wjk8+0d4ibUewue1tQOgVSZENggUW0luxQkuiDzZc7H0n/pin2BJbc10JRNV+0FB
zQEAjf9Ys8wESsENEN4D/vewcHDs7hRQ9sBomvFEU2Y5GNAa6qqUTCMiTszJwLzd
pCZiMvbgPYEX+ssb0UUJyPE9gJ2wCR21dh2xv2pE7Dq/yl1jWKkBDR+7Nya4QOY6
UyRKlTJ1skqNNz9+GKUJMZJg3vzn0haQIFTnrOLBuoFfWFeli2W12afbwlzNNhiB
F9eIcPvkGsK2Ft/jnWCNlVSMss0Y2oDdO8y5TJKQJ75xQjk2iqG0YiTK44JOfHen
sSN+8y0FuZ5UASsUpFLV6aRHz3GiIPBisMgiHskgtYhHgqb11CUIBOwsI0o05Pq4
LUznKjprUfrCTGCDwFuagDQVdIxBivbZKQh7g1kNmWXq796gRW4mp34nL1e/fpw5
ftEwLbXmaa3T7irUbpu73jlzDAIX9G18LdYcZimga41uSF+q6Td0Wg+TZYI37C+M
vAd/1+CE2gAKAkP4eQUqvpZBwgAoNxpKTrewKhzxs4EgB+whdZkIxgTQlaiTRkcq
3U9cVoPtTKMjeu/VKleMtQlLxueU1biYMBv22cCeN5NOt/3zKbYH2tuP8Uzs8K7u
7cSRRClQEktloOe4th3fYBMM/lS6Fz46SfrmmxIjO/ds3KHuSMN6OVwuNzTuC78n
q5OAMdqSpXqF/hDLRqLJRbUeQJAmncPibvb7lUr3yyUMSXqYDjcgWGY3p6AEknxd
kFU7dIn64DuaoFUVMeoNfe/pSSHXi2vgMjJpjR475lRo+qfJdjY0OhQImoYI7emU
kIGxPoYnWDWNc6GGkINlyOWN368IH3LT1mJYfcbZmltSx51CjAWjr1hXiVV+xOLG
nBchnY8cMjwIbNFMDND0Pzj8nLQZSRujrrls9neOewbLhJsVwllUsT0+CpMker6H
ZymS4RiSZKnsGDSYmnGTcsxLNuaAerW65AthUaCI8L04aTcCp7lDQ7kJ/HWWkIPf
2VtI85QlZxC1aoL3CrpqEcQWx5sUKaudAiqNOVzZA/5X6lY8OqVBeCHx7T4ClQkj
ek9mw7U/iqAsebGhPw9iLwtfr1BUIeykUZSZBafBpdV4QJKP/n6VHN73uBRGYA+R
wkShFkx6go0YSzurHS1x9PQ1+lACvSqhpy+8d4lzlwXEsSUjhtOCBb9zWmWr9fe0
X5MmmvATUdp7un+dNEiqc0Y9ozrA3TqCicrsg1Xdpnf1qYY6z7tDVErPMK8w10vI
bYC3ongVawkPgroQTrstAwdx/OGRc3GlCz7JLLoVVdE4s6l6GJecjnbcF1MHOCww
meNwpjQXR/qrC38KfjBsdjNaBffJeFeCHICLTLHPY61AEuKyJ+cTYdpGRjLEaQYO
Msz8FSz6AdgKlmoaET4VpkE3MkigPqZ0jRRpQRX97tHfIbsyuS+kYri9+ONlM30j
k6LFFZWeHSk0RsikotwtHnTyVdyHnE1FE9mA4W3KnxUMWfxUjY3q3cnhfCq0sp3Q
tr3rWuL5NPwdaZ+M49vN9T8Nyba+psLalmFDF8+7yB4DMLdwM1+h1lRzixamKhA9
AIoCrqId9jLP4FVsl753MNcST+B8XFe4HLWP3o2NHJIaZ/9s8QW6YkBV9cSeuR3e
e1y2mAWjIFPldWQv5uZJYXiyqC1OXV5ZRl2diwXLWxOUK3yBbNmoJE5VAQ3wdtj/
dFwT8/DlNftDDEOY6xk0nqQFsDRR5Cu6SX7/Lj0UjEEhDGP7G2kJHSDnbgc6gYMm
VqQM+pMGTNXfiLYhIVYtaSMKVueO0qnh16eG6uHk0Dc/R31eINMudOFS+cUqILxp
O+c8pC160AcX+9oqeUPeRWpFDMX2jXksqLFfaa5f00+uNAJ9F2z/KdNce6rp3+7M
afyifjzBvqZ/0SQfmNnY3p/H0qcwSjn997EhMzl83m3jz9mBM0LoKB00G/ydQCNa
sOUyHSB5IwA68Kb+6ycslpOdW/Ce7n2cVBZNQC1cJmCjb673iK0ca7zbekTACsMA
u64Ib2xrCN4jnIKRtoSwK8QeCRCIpdDFLvfRjhnycjIoCF6zso7JM01tcEB+xCWk
kRP1eV42vU7vrb0SY3ToPcrCQxVRnvPdf5BxxCxzZhtFRASWEtLH0031/+XNrDyc
2sFvjqDllZo8MmS8Z6lONKsH0rUbI1WoUzCCAJERxzCUNuQcJ7XD92NZJ5tU+c5v
FF5we7LReSd29fL4lQ85LWluqMBtPore7iwcXWPfXjJLE0bP7rFi/0qbeZj+bwE9
WEujmqwrDTk+gv2QehyY5kUey0+x6vE/ttyMlpuLMxoUh4L6AznEWGFhkaZMIOBX
8l1vokLXr+GwOmzF021SLIYojc6UButQnWpUFlcp9lIY2J5xbD46Pq5BzcJspCgF
67/LIXIlVOvMOQiK6ofe/DijS3/SE7fU2mwHm4jXw+N58stmWOZwXo5BzTBcA/Jb
xJNyIxK/2erEaZzcc41TT1H/hqqC8+Rm7cTabRPz20rScx3dJ9eUfvzkzhfq84yL
0/JW/9CSXdKNdRM0UCzcxxIDWoTAEKgLepdu5AfxUsuD6xOT/oxYgeDZfwmNak7v
5gkHve8C/7pCL6QFyG8snfLRnItJXk6lQttRyWZkTKCIu+JX7gzpGN+Wj+enhhyV
ZoTJzGgAziy0oMJVKipndSBbJkohrwK039Dn180q36l3YB8Dj7bm3N53OQbAN8Zx
Kr2R0n5vC7qU3PI8Oy7tPkXJrGgt1n/S0VVYq3pkJ9KQ+MsOm3M1PiQC2GMGWmCJ
u9ApxS/Z6gcAFFqip4QLy7rLbmUmk6E1JEruk5joIHnhV+p8qUmQ+VJDoUeDHYB0
QR+wvCCvgU/BJ6pU/ELaRetVJY/fcCOAU182RlG1pi4IH/kVzvWjzOD33uvrHCao
JXArZWwNJYA/PfhCvZW2o89htj13buRGrK9u6WHPILxj6BPqpSM8aIunAJyfIYXB
me3Lw5zuwY706r6TfZRm23Z5FYfg/8TAvP4D1kHFgdAWWX7ktWIbjNdaa3nw1Bl0
fS3R4JgWA2VxDym2/no2eKW8Z1FArkLPZdYxxncjBeBJGmzS6j7e3raO9B+MWJGG
6Sf+ipc9JL4dA4P2R0mzacGhj8ZcNxVSK7lb/TQAeHSIEJFDCkIrZPdJWTWFVS/q
IRrC2/4+6MY3eMjeCwFYGoIcIWQ3GnyIbZb7LK62qeg6Bax0fPxYgORtqeuxB9qj
gHmXMmuD2nPqF+ZQvMVPso2rxrU/LIeIO3eio63T6W3afSdXxvxNH7G/xhp6J0wL
d0FXSDV+aYRns/hpdvffbstv6XfmrIWwO1vCTRmCpBkXLpyPvbKQr1eINUQWId8r
hqEMO/YQcYK1Pv9KKog6BPRIqzme/BV5k4mCRrWU83TncrLYS9gdHc8EhTn8qq8c
mCNM3sxr40SmhOaE9e8nJNvPI9otMj7hxBYQdC5chdKj/4NioQ2PB9VpAnlx+Lot
sP2s/9rao4iyzEfCSVJIm0IRVTDJE6a7oq5ZwYNjcfwIryDIsD3MpEG6RsRCQRyh
oMO9JXPba0tDVzE6hkyixgc5LeSCqcKr/VUGDOvZ/axhBSk6lcbqGipOZXOYHVNq
xK5rW/luH4wzD6K4B4xSzrX5MYtXPAA3NAVen30dtL1gk3V8jlBOu8CXJC7abj6V
TvgKbnW84qbfPea2VF7OVynmk6fiBQ7QRTua038RITJ5LG0H9pR9KoqHz3Hm5oDg
UDvl1iEGQSZvbuPzcniohNE4aOHIYKNjpUEwQskasAt96JjmTGn0I3B4d+SQAdft
JsWkNsHvo6CK3JUkIFYN2GA4vsXjt/eMsA8bhim+qgdZxPnaaw0sNHHaNB3M6dze
Sx3nTth5YsNnANJcacWgE6nc70j9PDMGOgYHzlThReFFWMsSsw4/L3NcRBO6bbTo
0DZRcw8lo92vjpKXWI5MKAosWJaoPLiux/GJwccFJauykMu8GvJU8AkuMMRiC6XW
WQPnQpCZL73q/pcxrwhZFhayDKepM29MIQnAHVXqZvgDK/I4rLqS7vUhcu9a2JZz
zIm/KkfjgJuSv4SETuxShSYZDNEKFccdKIC6qONJ1Vhe5AjQrv5b/IsfMjccRr4a
RXbL0HBezTFW0NAxFz/mPQKChaV+gkH+Ssfbip7qZNE9B6QGbnLX9+24nysOrkWH
Z0K9r9ERCsALuehlHq3/KYHDCNBLaMdV6tQAZE0Pvk9dv5Ae0cZxKxypbZplJ1Vo
HHlt3qMZrv8ZfWXA2gZJyUk/38XELgkCAWp6sBSEgBGAQOnszgpFNnw14v5ZFPdI
4hXcCiRA21XaikGyHg3rNm6bl/zgFvyE69yPuFQYDblUPueHTSO9Fe2t/NzOWKLC
vFnW/9Y5ncRgdmXNAjwDLswJ1rjr3bXS0F8wL3Dp2vTs70ZlBy7ZDwq3SZI9juFz
nMX1AOISIe7TXC1dlyJwkG399nPIFlltdBwj92ZPZCnAwiPK//nQl1nyk8d1NZW+
RFqGZyRCYr58qs5XvQ4mZpLFINWbnkrcO22HEkWp5lKT2e2Ld4QuU3YH8LmIYMg5
6sjjZX2B2lTMde+JFGAdf/68t1jemx/hB9sTo7b3MQ9f8rEFHizfJT4nJsLajd7n
2pwbmJZxBYQfOqO8UmmnpsoC6nUds6J6i4r7V5Nt/YbNSN89FNgaPlSPzJDWBbhy
JUGofriMbau4GPJJzR3qe7Y63sv53PG2CSR+7EfIEoNClb7rdQ6VJ8pBi2Kwef9q
jRaV7/nxrpnNg7SVxOByi5SenQOBFSf8VAjp6EIu8s6sdcU2zMr3QNF7tYH6GVP9
8OeWTHmq4HdOfhXYO9r+HCqVUtOItPyNya6yuVaPJBEDoMwbz/vI5oEzCkr6vtkW
QRGabjh3ttnGfjD8UOdaB7Ojv0V5eoQwCJMvmFhmDTQQxe4PMTZu+Dx9sITsuICR
xDrG8GZvsAigEz88dQYl6uM5aOq7itNEKQgIEEYyOCy5LobyPXXvQLuxueFXYGsj
ia65rZpebTjr7BQWfScKoiCIRIilqaq8XjHZFnq+9JVGGXw7yVSi8FxPgf3Ct7dH
ZdbXQDwGwhPU8y1v3ODgjAmCQJJwFwwQNzStnXAhfVjZXmDKHKW7qggVPO5EJd7r
/T79e92fiSO6YsNrPLbXSs+aNeIW1o20HG4Gzk2NFf4PeM1+hVngGeVvCCnVKjCr
Ja02KLCxss8Z1/ADkeM9oE9bJhpJnNOidD5xpLLQ+dZ+lLwnFW2D25NF8li2ED7J
90WuOGUkQb8HaDMM9GgqQh3/Lhde6xkeg+4yubHyJdRSgVNffpGNesEwp30qvyho
ASEPEuW4Gn94KQyYGBzlNDNgmNTAx1IDEul8NghMvPVkfa1YfNpUuIv6nr1BoDEb
21H4RSkOMLIcOtZCWgsXY+uXadpdl1424Wi3O0WF0ZETUrTDVzlnSVcTtT2WjSNL
8QCb6EY30kMhv2V/PLXJezt/Chq/Bfa8gByc/vx032fokMbdyyrXbUPUOSuMiabD
fXvh4gU14NshRGRzbLAFP6ADW+gQopCjXOYGjVCNWzq1EbbOUELZiJH8nuS1a0Yf
4NKQwcBqSmAQXptGqp+DCnPqLUKwmmG6w4lau5a983KJ0oobh4ndtQGFRSFNQYY5
oYp8ijFH/qTDyD9TOkAKNCfblQF9FCV3G6+zj8RzbYLGBEwzf7uqszUKm8cS6YLN
1iq7TxDY9kM+ykgLWBvAd9p8K9IJr8URZjszvlLJP+v0D7z9h0dJa/+DRT2ZMXPh
6nV5dAvaf7tn7HXHviC51jcd2O0n8izJlXQ1Ir8rgD7aqItDQ9YC2klkppCuPw2Z
FtVC9NnUl//dR649sJM1m0/H5G5k3sDM+hj1dn3gj0anOeS23KTRMfJyI+NftaZv
OxYsHdU3FB3PewJgT+3UJp9/YZJwWE2yKPu7bgQvE3ESmvzC5wsP3KYwiZDJ9Z/+
gDwajaias0QRUBo1mi+WdVZXoL8h0md2GWBFf5l5fGvRqAsr601aj0xeFH2A0GPs
Ygo0sPUFaybXbCqaqh7s+6DVOMR7ABoUSTCq9HQbkaSrNGKo7MwAkV+7udPru00J
5QYAqqO8/aTJvyoJG7JHLsr4qWTlivcBb42OIPSrJrUeu4VUmMrnv0UXEZEywWo0
XL2DOgOFlT0V7tqRc9vteFMMixnweFE6uikdcdpXJKCmbojTEH/HakqFgJmxqAuH
LRRkTfHyBBrpUM+t68+QFkA1qGchjyTf/GGTfvD77HViI//2vyp5KiZr0OcBel/5
L2qMEGRLyXeYzHofwJ21BuDEyx/FJfm9JKZW5f3dhw8dOn/a5RFCXaOAY6qlEmpd
JACiRLWvb5BJbnKFT5ne3+rOIfd3pHH++i67pQW0GnSwwcGDe4RLCVOv2G5QPm61
gySzv2uGnwX3cWOju0F0wpz9E4BfNy7GxWdMczYqVcaC+Epxg5xOU6M6IsH0KTi2
bIe+zOKrAMiSvStbgdJlM90LJy3LHaicdoN3kz14GsQxcGiEF2Frs9UGLT5aJzet
GXxmJASHGGWhmI5+zuFtwhgijryGTNV9qCp95GTFcVea8VkOf5kSNQlrifXpSQLE
IiC8pr/uhA455HL6UzGXNvu0gS6ZG+dSOCya5fA/tb6s+NeJE6Wzo7Tbog1SBiHx
nWlXmdknBQtzWrkjeSRvTlZuyYd5vVucO31fC6EHAJrz7eEqqivwTF/nEDmicJaA
7rN2kjXnquo0MrhVQhvI248NBw2rdOuEx9Zkz7DTHjI036Q8qzgVIMVYX8GCgoYz
sO6dsJLjgI3L6NEw+2nsYPPq9NfoC2WBGXIlUaLj1QhCBsZaBgYLByR8SGhWW/mP
NM+qFrdoqP7aTIiaz5qwyh8TyXTW0KT1u4+fpxFeKmZNsYxeFoKPEA/aAHC6vH0k
Ylfwn1THJXWMqZTTnvS4jl/1SU2LKkcQTh4qeiQYu+LCKp1+HJlzK7lt3GRnvOjp
ROWav6TvkIu2WeDnVhXEjz76qXq8Whp7km1dB+JF+UJSNhESGKLfrXNsTZqfadXr
FQgN10Tyx1Yd50/zIuygo+tQUhnubOJCs6RwJ/aY/71Q9mei9xOIqMesLkKfY2S8
cem524k/WNQdnT8svXDtmJqRv0nWDP5SSp07/Syyr/62rK+ioFXaGcxr9O0QQ3a1
coPvqx3MPUkzUFaoiiW5s+L4ZO/7XcLTcIoQMWkEBTJVmqRJJRAao2p9UQgVA53F
UnA6wvNmEF0/UAkXSaMesOOaJCdSsKoeC0SqBfJReM9RGblbRXMWneyXHryLrFAj
0VoO7OX69C5bc77DOpFtJQg+bbCvNEH9KYI97a8grZPtvKwJ2Zy/MJSDA/Caj/oU
Wbk3mDSTT50eKUPTItw+jo2WQZWhYwNq0C7l/ukAEOjS/fhq08ZaH+RFYgomTS2q
Qz6izw+tr4I5YobWi5EB4kVBnDp11bNUUCgTSUOQ1axXOCvMvKwjVS4c42h+iHEp
PplSXKPvkunMjl+AvJ1ZAGsqDRhqjtAWExcDMrY8KuDHucKR+gqjlENoTAkBeFLl
vPGxXg54NbYK3BJ8SKPjv4VQ1sKcabJm3SN+q77kidKJsC5IIsglk1w9xbMrfUEE
G4DXFOLQGnCdzawz1zcZl0G4izdrCVp5J4SuX1GZ6yfVQblBXS2isx5BTUpfIIZU
VKL4hV9OJVAySYd9H6bkCFGxSs6qBeqgeaDfdp0gqCiIR9XYNF9hednsEvurZTvT
Z/2BV/bxIXZTTRh3zqmNZtfpEsMcQE/V5dYGiriPgUKdnDIQb0412vKIAyiwey8z
ZHrfpY611apof95TbpAbaQ1oenkk2tNfRanE1FhEJFUWZjsfHq/8H2ZvdsRIMQra
vtVjmlHOvtFoZRK1NKC1hWtVk629m8MT3Cq265zasOoanSN9sopCO/T3tMSbZMmw
Fku1tNS/XKrgwZ1XMJRhLjsfAvABCQWyfyppToScMrCQsO+lMQYb/avlItX9Fzvp
hAju1n4PL6ygVfd3lme1Cbizc54IE8D5N2wrwiOrCp9FRnodd9KQ7kScE5trxP5a
pkh2moUtQymce/eRx5oTyYo58YCWIYVYN19mUy4EaWuYLGUVr/nM8B0C7uFaaW1r
LNgdTQNcd12ANd8R+4dnw4rPcB9Xd8qIXfsw0MEX8vfUrorAI6OO6KE2wybwKZ/p
ZbACwBjAyXKjnT81Z7qCCGsQXqZXMnFQ4H+VHC19Vh0dvRmdN8sr7M9Ht87wXq4k
Ko5Y3BP3on1vSuwF8KYhQejq/6Au5w9ezxRLxTuVtjSWwQx4SU8IGSARWycB19rq
dQH8qtnpmV68xFjfsuVU8SeWyXO1b4ISu7BKVwjnuBtkuMfpFZrD1JyythloHSLX
Hl05/DF7SVeOz7P3lUMGs7ItLRIG1qSeypZX4Wll9L1mbnKLVNS38OljlnOXOJD4
kHz2WjsntcMt3CkvsEj8vigmrhj/9mytrIM05G+M0U9qZMN7bHFIGTVcwmK/62Tf
r2V9TOCVd132YPb/acY78qJfE8Re2mpXN1zpLgbPpgtvEQYR3ZWTbOPBdgJjVoE0
Khet+aYaSVjRhl+BIqfIqPTRAX1wNOHf4IJSi9bfoy+hVcNoRVFp/BuYz4A+k23G
9jXmCtz+GSnk6b51JiCLoSieHeuQl2rbzHplOudLA7fQGbgFvd9WBH9MR3X7EQzA
mBm9/u/vL2vG3j9m0NLoUxaxHNibAwWT2CPpIo4jWmo2v+V/iuQ/BziQeNh0tUY/
7dQwNctJtS1T9P+VdS9TfL4D0PDNnz074wBNtkI/rOlqlWvw+K0jbdKUr3A2y8MS
4GS9TYtSRaE1eNESpOhkO19H+bvmxKP9JP/ULChLp18kvIMuvmtJW7N7qChYZH77
UUiTeAmWIcw2wo2m0Q5Hj1SCugh+OQzFNtowDhXQxUC7oyeLiOBGMHMog1XAMHmG
T3u7TRQXhK2H6kVSoCZirmFFFlnIA3wJm9uvHoE3TsoMBWk+/wrewF6b22WQ7x5d
byXXJXJmggyec6Xg5X42rKjYIDViXw0QQ1tO6PkVZ06n3YiSuMzLSRMReMHwxmau
beMFNFoDwG4UMHcitzdfbfVqm5StZkxqByRzlBqt7ZBj6HwnskGKfNydp1I8cVCf
fZA7Lb5Kxlo0qlE+4LzeIFGghPh7KaKS6i77C8TlOuuB5tJ49Oe7RG4bmzrCnpvv
zNTS0/tgCHp3n3dzcaRX9oQg8cda0IU6M/SvY1lv6zO3JTa6s+LQbsA7SNhBec8M
EYqtKC0n/2kRu4ki5NBTycqtgLRYp/aUxAb+6dzz9ZPE4wy+NPxWaA4/84MNXi+T
JsbwsQekwkOBcyCsydfMZwO+BTOSJGc24bDmqAJ2O4KDZWdlm+ALB7J1fnwvO9oo
TRkW8wDntTDxGTswhYwrXQSbCnflDGxr5oQ+oqpfVn+EtoHC/hZiGOXKc9a8MZVR
/0fLb0I801WEdNuTy4OFR2xIkqIou3KU6aMXMdt27M/FP1K0N/zhGBRb4VFY/jDJ
/zyikbqsHRGqS5ZduTyoBu5tmZ/Uikn+Rc777j6FhMqb8ByPIQnJBBZGEd7888XS
6x3Ai3mq3QTt6K8MTePk7OeaZ8AjCv7PBr4qhbgLeEW1MmrZMQtYXNYZE984fQEv
occSxty+va5sC45i1HnVq9BH/DWfbiajxqP9loj+s57vGuIR9xvsVOvNr3hn63Au
sR9DaslONgM0eNw9iFC71s4+EpFDLMXvhjqprtrtPJo1fw8N5SOws4EOtXi4EPHA
OviRKyvKWhnS/4fopaMA7T3vKZ4yuOA/aDhJZkkSontM148QIpulUbR5NLVIZMWC
gwbtrR/l/RZERFjQrTMgg/ItRV+gmCU5LgxJfGEHVtfZPFQ0+PcvyfdylAK6PV4H
wP4l6Zrpiq63dMb/iHi2fqE9iOFkGXLJp6ZlERKDl5YTJ7YMPEV7gl9QlkTX+fiE
ufARVexrmQh6zftu3x2Im4XhGnka/uZsbleOt+feNjk9gNa777d0mWKp4q3LdEIp
Grgqo7VTSpMYnaWvYZDpPzObNmizCFfX3hUMqqd5IKgi+Y8gbcFQegHMA24K5jNn
cfHMzS+VX9y0TO8UW9gKFRqAMEkRJ/3Bk2FE5DYs2Czxrcpzv1+lHNTPEDO6Dx+J
x5ZK25cptXWKjpGK2dO/6+o+nQzVXGC8GglxoCOpwDHci/VYpD+whnsdbBq/qO6x
16nBSFBm1h14QX4j/ouwm4WhAwwdBRDNjtghUCA0KPyomVUkG+rItzkEmKvO52oH
D8AVER6nY12BEWxRrBbz3Mo9yMhWQKGWSN7BMVpGiyyLRpc8X4C480MAzAlrXYc6
pSBk2j/5BkHMOkvjFsLlF0pdjnAU9mNj6yhHETWxYcHW344NglJAKH/hIwdhrDr/
CpDC2qjXGUfg/5D+noqTwYP5/gBnYZxTTtl3aGDf40kB8O6IPYEROqOuQ5SUGGc3
o7FMQrTUsRYvJ1d8oy2ZoB950rCAVqQ6jjOXrsNqIUovg7Y3GHBBVPZdnjMoGwoj
Jeee1eJaiZgiZpfP99CWShb0exOYSzI742xSAYAvuo1R2CbYvYzKj/nUTJHTII9X
kKBJkEComf9GriTpz0F5INQGyhCnYKPlNG981fmCmBxsXEUtFJEMJFM+VABVJF+T
vhDs8uUdSre+h4sPxUyIHO+k/jqN7TwXLQ7TQhS3KF0tss7cniwVZDqgdevhRTuE
R20+B2hauTvIRykAooKVbV2OVgy9gskRI1nkGxnQRnVTyE1n51ULriL+M9m77IqW
CZFb/luMKWUDEhrqpnGKpyF6HN7qszwilzlKkUA40ZSzYrySgy2J9cDGntxkMbAT
x5kr8UhKmlAy7YcqePj/NBk4nvPRbW7qHt2BOdwhhTdUM2VbTkJMFTlWuiS8jTW4
cpZhDveOcy+PhmRvo6ViFppVeTHP83XMHVC1jThojJ0qqsjlqsDDyNNrtX6fY9wB
9lodVozx+YFbXb2fZBlo5t9McsRIHfa6iwq6cvMEXrmTbsx+LkSO2BcGTtSQg4o3
ARzO+3aX6kUZf80DxHR5oNPocIKZfco4Ys1yhFZws8FwjQBZrHgvxRmEdRLQsI8V
rUDkDFUsaHe6uUks52mi0CPub5XGrNrW76QY7jdcM3KV4eu5I+32zIHaWN+bfO6E
+ouSy539wmr2sJfV8Ap4xwERmOcpqdyeYJGRxTTwTTmzXcx955owhfAHnlLE7eJ2
q6Fbbdafb3wFZFON8yQfXbtSipcodKh+AdlyvRsOy1brss09rWfhuSrNCTDv8g+A
zGThmOrjm/o+GZtp06l01Td+yOmJy9v2dLf6GuHdvO6jVX16XPeIQ2YfAIMAlC5P
PEQMu89nnimvGZOpSCnyXmGXFz9ZP9ku9A47gYU3G1TC8+ikcF+rsWnPRgrbl30y
0XudxkuZVWGw5Yh9SjfavX5bXihfjVg/nynqJA3c4bp7jRi3PixD5kOLVX55oJQt
9O4lKJx9s3UCEX3c+VRUHZ5EBKv5KrR4MtjiWVjTMfaTTZZjHtiT7FgNt0KEFb2v
gryNVwslEIjpee0Y8BAxXqiRfWv8bxOFo2wY6NznXwb9WqS3Kt0e5omHdbSInQNo
2uRIA2HYbUT2dKc3iXX5oQrZBZs0uWAqPkLWH06uKtwSysI9rtV1CSsp6GiQleOi
pscr8wXzIMldKn9PMiWi70raZfYrKC/taD9HXVtic1HmJHwLv2LRoMyzHxAiubsW
+n2XKiwVchCZuGgajGV6lFAJt6YUnQ3obyWOMgsfoI5nRzV+q1HdoPSWHZAYIhTz
QjiXOa6J9/NEBeGMaFsP2uVeerm5XDdi6QG0Z049xOJi2CtjTnmiE+L3urWxbtNC
fDJ/CYFv3peWJF+UA+JeXgZGlWz9vZcmJr8CwQBNf5dlMGi/KgT3OPqyXAF5ug8G
M/idMsu2zheGM86qoUheV4K0gUBDnek+J3XqiMCpX7E8LE+cA8/M13S94YjfgcGK
Dv5lC6MPvwHWw8Iei39YK0xt/zePcouovDbKk6YhJgD9gvAgv/6HqeIbNLSSP4aY
YK5kdTVtmmS7Q3b33XQR+Eum+6Jj+ihToyWJphfs5llJPTyKSi6RoU7X4XBnJI5C
g0g5DAIdy6u61TQa54iTbO9RQNiXpyJcGHnuzmlGNl4gEZUmyRJnerRb9a16mVgj
Hp0XJN8uyw5FLQNKZXbqXvAWk7VVuF71uYVhdlk0RULDPxElm6tqbJvgcesMyVmx
Jf3mX6mQD3+pxLH5yRUzNRRCof5LRlx6CoW+4tsbONwLHngRIKASBNCGsrBZ3xW3
9S0xLHlirDDsmxMLe+zM7asSqCtuNqe56r9anYzEdOMDRZgMQ3Ndj3XVMv8MxYWR
A682EirNos4vi0mutCLHM27XR2FrhUGwoO7cDRb7aQJtPzArF3ivrslPqWmeiLzH
noZUpuE4J9ZWAG16w9AliqhLgtyemZWkrTydOUs1DvkvcQpEkzzxDNsFLUh/Qr6Z
qCmnXl3HLlSrpbK0fgo0wzuMEjm3LvMrMro032ayFiO+4z648rmgSfKFVjvGkmeY
+0W+O4w7c47rkF6iVtlWOu6bxk42y4o1PkFR+pZU5zESWmlVD9o7O5JyFJh22W3M
txG0Pd0+HqJPc1yKdc/le2xcV9PCtR6jmB4Ib38ckwz63jpUKhYvanzdxPzUrDBl
ae2U54+3LKjXySOUtPBunNVPJZqJ6adgu6LqNZB0nuIshKja+wkYw+bKWbxtscTQ
HwA7+44QFm1d2hE9p/FADzjvlXHaiJR6w6/n3ra/QcUewujEFEP87LdRukeOYNon
9Jbjx8u1jLEIJV5nPZBXsd1vx3Ocf1MPGZNBsWBQtlDujNM/0EyV3/ArumO9va5Q
6hnoq+BZk4g/bIOkZC4K4Xjzpt6PpbgAPbQVj5lhPhAgYuMzw7NAOGQxe9Gnqu8D
7dA9x1fMihjiOMQBekSC8sALMqyWQIUtE2peOYeJ9u9RIifR6/I6cElsHGQ8GIiz
G1yAW+vT8+En9680EQ1mCWq1pCD4vw2raNEB0yApPe7x07yWpvecfQbXpe+PnTI7
HGzxP7E/dEEMnggJHDXEHqE9iG6A9k9P57R9T3JzWATufkL0HtBiynIBrKr5JpST
rlSVZCE42p1d9g9PC7zxQPmRi3pVbg9zzT9X3IpzVjCKP/w1h/CBbv4Pc4XOWKXr
I6MSf8hQqQuDDH7N4owg4P7+/5z5to0JJVCoWrVOqHEa15mt0VKmLvkrQMEDmaDZ
rNRHs6xeAYCs3wGwZZKGK2cIB5cPc6LnOISsrJ4IcFBuNXww+jEHUs0+d0GCHWKT
LPRn49eKVnOT4ZdfHxH+3WTYTj4AwEHwT+V5SeOfC5C+iB7yaHZu/1aCIpKPv/0Y
/ca1PCqmmBRMYdwdkqUNPXRh11DoVPMPEWWIlQf6jLG4T4G88FG+kZf0CvCWItmH
4HoLBo8KwNuT3tuAVOlW8ANvNTTkNCdOOF6OFcCmp5VBhBMOzv+mD6AG7UH55Seb
dLa8CCJzPAXyhOk7sdwI0bpatRSE4WOYW3bJgaE9X+htIBp6SNf3iovsWMX6Z1c1
Gz/DDZ7XDFOrD1pEwrtpHkDlQRWuKd9oyNd3BU23aau/XXNZIwvM5EGY4vS57E7E
ShShHSSKOXaqkfsYf3bZLOzqq3U1aHYXtyrcseBrEtaFgMMHjHLtk7dKVWP2K0p5
jwSL6/jJhBX6zbRwrhmbx4lCmXsQKzy99whjjfGcKhHdsCTSbusei0EhSHN062Tu
9BDNW2ZNino+h9bIPM5ucNuMECAHK9cNbO70LPDjLmlZe25jKfEAl9NYvHU46/Ql
PSrRq64TF55BTm4x2ANtdSCy/zn0NN4JVfkNX4fZjGKr26oYKY79Ss0xHUGoxpjP
GscGvy5bcLCwaiFGSHBaSs84ND11QxjDtdADCvuzTd2+EqYh/x7MMGrVUoL1YqNQ
BFapseJVv1FH7z+q6NBZ8KwkoIFFqXvq41PkA4QXwwk+wAJsEj6T+X7ds34QYoZd
ft6p7dvDD4m5Xj/ty2U62qwZeHcgRYtg+oUMu2VntbehbKzrwF1pTcM2Dut0TYqb
F5FyS3b07f7wxL4DgaIAe0W4iqoXrOEe+u54A2KMzGKm+oKa1tpDfm5Y+bRjEbXb
KNgwmnScbEbYJwfelLQ0Jz8XyjV09poivz7T1LTmAOhO6fIu76sO8A0cY0cerwHZ
er+M+fmUvW9KaYsMi8MM7EkUhdc3fuKrTiuWLONcNGIhDDctgrbptgOYfdIkPb+O
rZ7mfDbfAbrA46LqIWdGSQgFmuBUQDbBFR/Z7Jwb812TGC/vB8e8G03kpEFOVssg
VEXg81Xp04xdY4IROM171V8rKEKaOuHHxVp/0RBChBUJ9FX5MQzGeJntpZdZmIRv
LEH8eP4P3L3PMnSruNwsqyLpLbnVzMtg79ye1fDuWnh06zPlfpr9iTCrnOdHXyU5
VKFcsGSWX680RvfF53A2ILF9SyfExLEX/in+zZE09z6akpNiu4+5mXlzSHFWvbG7
RPnrhSzrvuLXIsvq1tgp3gsBmBJq/RKVIf63JQ8XperGoxefvHKgBxZC+hmJE1/x
3qDBFNaj56VeXVnAd0Bu684KydL5bnoic/QGh+lyqrW0uoQ2X9HjCs25k5NH/eq3
Az8u5Nuim1qQkieyNfNi486ny/AK7getWdt17n+idAec+afBKfL0nZwvGSGLcU1Y
EQ/4IMERqvfb0bxMOdIny+pBxPJN7X1QTfh9cm2K6fARV0DDE4xWDANaMXC41wHX
o6lE5LwbXGiQ7FVlJL42YnLnj2yvFmIeZTaaMEAkWUs7QUQjvFfh7d0YhXL7Gyqp
jMgEX2cN2rDK3gadKOAnxwKUQGpkpBkxkVjuu7VXCoDT2sdkIyoE2pC/U5DkA+Hr
gAIOzO2FZoE4Jbsemz1w6HXLM3NPUQ4nJuqH3Aqdb6O+lZM9tf/bYgJKovn4npHJ
kq2zSWWIxd/yEYzKajVfeVCQHquLxto2Uk3oyKDp+UhJdo1fQvMBM4/WofFgT/c/
ODcNzKhmjS5EtJJbcvGeAgVUFDTi6dvK7eSE0eYGMy24L5zkKuZIAvb+uA7o9q1h
9K5xTvBjfrLyeE9T6QEdq2SVOH+1xjbC2szJIaMOY0Gv1RDo9pDKd7fdFEPqoVVl
PJbCbGR1lJuuKDdDKVmJv/1qeQLoavxDcNUffSgaAlhvDzPS3gcgak5ZLxVAHaYH
SGkFxEs58GCqd1kae+qXJc5rGx29z4zkf6uxprEeo0FBWp1kt0Mrxe3wHe/YiEQE
XR8o9JMhm8ATdjd7HaRwpWvPr4aMhcI03DgC5/bbDSX+yteTAsFJwszmYLk+z8Vp
QNxQWu3eN/RUXNludfH2RMboX6Je22pc91mnDa2j34znVY/scxOmsCFByy7dGZDI
YLPMb1PmGIXs85bxywoB4cvjpEy6yJHuI9Q596ErEezpSYwpuPDMZ4zstY/FUjQ8
5pDZ5Kqfk5CVLn4/VPxhzyQXGGhS/tcoyfX+hnN7wygk5drnz3+ZZAA6vH7Fobc/
vOXGYOfFWpXG4imlBfO8yHlCKNN/MnYpvVYdWHin0NFWFb7VkXmYzTjOLoDfpH0M
Z4v1gCKbIC7QB4g/3hfeMcH4rWCLofxCPdTB63+yDjlJ1DdUL4v7yFRAaPQ7rG9o
kok9ajPvLONDaPl7bJNB+qrTVXV4KDSOclA0Y6y3vHFHp1kTArfmmHvgpCMiwc8n
ZXHmQeEe4876qA558ZYkUhCjoolv503c54CtKR2RfKU1+aLZthPJWeozkaqXYTBs
rd7SLJg5mUFyz6x+sXRw10O731mBjeBE4/936aIBVH7UoNoayIp0zIceBl554lxm
8AnOZe2iMhSBTsNnMWPJjNZ0wK4yrvHU7SdzJ0uscEQGLYv1MUNDRIMNstiTyxkG
2Ea5Mhu+cihfcTvInMfOevH5cU3CIXrniNd9aBMoBHcxy5lR5vcNT+cuArDMxJin
xINLPlLj852+zSqF+OKdqCcmD2jiAk+YuxpHRRsI9XEt4VXMOaXYa1hfYyWxEkxh
qrvXzMZd6hfWn7r+Gs1RgkqqFSumiYjh2238bmZmv7f/xtrMHRw9hRjYaYeKhSKm
EhNX0rWo1/hd6JWz8PbhVG+6lZpFueGsc8eRbclBWg7QbJjviY3+3b6FTnyVTaAA
d5GwLJEerhnR9vDJuyZ9jN4F0R1IZ8WCEfKUQUc+2eGnNM9Nygbhr+w7R3roybue
Rbfg9dH6GCxDdNDKzVrXCZc0rf4OIR/1/HG+m97nzeDfJJRqZwhvdMgWjMYo2HUQ
HHY87pOXGJb5gOeLKxH3Fc7/Dr+LZ99VZOvxhk6fC69LZoXelfkCHHEWw4SJnSdt
g8wfwXE8os5KciKO0PlLIm/r/dQy433SG+Xem0XpecazutkIgRnvt8awYntvd5tV
wwXbCJ/eKGQhLCvIwYXOgxGM1jXl+hhSNvaHJYBwlj6rCsAKG0Qg7+tO8M/ppXLN
KLuoA7BR91VEHogzYLrP/bf0H33TXJXeMZc72MvCE7RgMwHsmHbmFU3kPF8coXdf
OsQwUeh4Njt9+KRUqyV1A62ZlyU1QnLobXZZdF38pXtT45Z6FCsqbVa9lkxQxYWB
//AymGFh3hTpDC8b//PjC1JEtivI1baABUytrEmaSwxLCOfLN2L6STNlLFBQxajf
cQYz1eR0k6akIkYKNYfHTBmE/0BA3GBnnTBxiGyE+7za9fMp6MEBGP2yj/cYc+z6
sCgl+BoSonlEGGxQf/db1S71dFU6VkLfNCnAXgAgXSt9l3VLX5S01vVjmEF77hQS
i+14oaAwtEvsB4IhSWwoCEMr1AhuDKRjrFVhDWZy5O6CjGkXhlVGRBws3tNn/9Iu
g9HHvFvmAeYR64pwBcaet9HO7X+eli2gkKEQvG3TmHG7/nv94bgf0uZNU5swMMWO
f//zkLU6LLtr4eNsKxVLORkYv33PCA9duwbNqwrRqxfO0Gv9cDWVd1IOTMqLSMfe
6a+zofhQ1k/EFjvTBliVEFVLyES72HfKQT798TexbbpFh2LUwzB/jblnmnjDOxc+
7UQk/pYUpoXKsVpDHud9ZFZWrIqZtmWV2hsf6DK4XISyu4h9tQrgFaXL5Q8tTDzH
7jProXmNp+7DfloRe53PaRkZvmHkPFNktSi9Ew2wfSzIBOdr9flKZcjb2huvldoc
70Q0krp7vUBbVldB9uvJNeKGxENs6nlQhHN0yJ44+3JPIpBKxr97H4/VRL7e7Spf
RE5fCqTNs7o06n1IBYt+jowa9t3AqRcUWrfF2/PAaeJC8bG6EKD0f+hMwMQheXJC
3qaqbreORaFllgOVEcfugUcjB0AOS6sItkJcCOWM3syavB3ijCP+pYExDiZ7T0fg
UpE3mknlN0Ry3jtZOalQxPOBij6zYJG2aHO92e1nHOb3u2MecwSpTw2d6xL46ue3
2yJxtH/MhofRki1LBbHHGwypWrsTfNr2oaOHyjxLlSC0HtPgagYSinEQ6f9za8GU
3nTXOpBHa0+Q/W6NfFXPks7A0EvLkj0b7Noht5WJsM7mNuArhhPYBbh9CThGHiBA
mxY+EbC4puw6bgy0BxWH/fCtjgVFB0RoZwLDPvZGej+whoikHG5URQDMIDomTIJp
EWVmmZTzIFZLksoIMUQltkoLBWkGSwp6kbGnJSQ3j1bGkJrG6jzHRShqw3hGOGa3
zkqEF391PQDpKznP8NSQvtXSh1K3mKQs5x4aXQqIewWSiuCd7oc/RniGA7JZNmZQ
kS5EZsGl716HY80iebJXSow3xStr0BnMetQ63tCOrYlO/xAFxBeTUzd64FLl+fjN
mQFKI3n5J8OyUfG0FKOT4vkkaBs4qz5oOSquMrUjZJS6crEYHIQET8XhkMeaKX3B
3Ye8BTOh2l6PYFKP72sLmftpKHmUdI7fl1u2gF5mPtWtiU4SQQnk8i0ARu3QX6h8
xF5fpeE6DzVl/UyM7jgqQYyh2Qh9pLHcpT6wCZyGmfX3FvF+dbykR1FufKhc4R5k
JpLCyXINnTZwggZYoCH9iODbnHfa7AM1Qf9I1H6WqFjS2XUbboky6gy2C4UalN8n
6OWUhId1sy6B+DIq9J+aIwiGFVh+Rd5cJOPMGj9KMrs3/E20o8Bz9nOwRuj+PYQQ
gmeBSOP/NoVTZQa1AbOl+eQw6ZAs1XI6Nee0Gw0JawhrKcMLv468T1mRpmWV9keM
4GSed7FXKpkfUmOySl5c2koeBfUPzaZl1w7kiPe1COtxw+MBmw3kyvTq2aTpPT52
OsYEbnbLqKFkrfiQXHJM5o8QkBOPtO2qZBk7BIjFl0dhHPfQA4O9LV0ctxCIyTMt
EQH2Xu0RBL9/GBwagKBNbIn8Q/CakLFlZhbUTLEMAOokEKUXBhVIpOGMlxh775TS
//e494ZWPJHRy9OIfDjpY770p3A0WiKzgYjbX9gzLxHp+bHrU9gbXzlK1e62v2M9
q+2U3piRaDIyrOTEwpK583HJqXIP5f3ooTIoEMAUjJDohsMUXRsWnP78nVaELybr
gXzTJzR7tx4TPWyI9w4lWkz+8Zd31DkT7VLSPZbz+ae+qQ2zJz07K4dhBGtAC7EV
cd/nbfemMTbjusEMTFpjdAtXs0A1Rh2xH/vZ6MYxqlHHKmwSTf1LIFCL10vp6Z31
As16bhbJiRUplZE3DRB9GwHhRxFN3nkakWjuokuuFXfp1Jv1HBQVZZTXFBegt2z2
kIzxyhIIC8clwafjnsqIKKEmfvzDxylmWhLL5Rf/pdYG9q+UfSy+uA0LnnyxNh/Q
lQUtKepiosIpRKHRSbbYeer1IjaBoiNyPehb9jc7tEVjOmTLUd2p7XafXl+qDsNc
JknJ0L2z8ikVAc2LBohmZYBX8fTSIPj6zYvXh+4Si2aT59N9Bd8LrlUeb6K0b0xz
qCb4MQFqND5/KboX/KTCjiOFAFGBf7orRKbIJ4JLSK8/OdswWDamzsO7O8oKu2HT
cA8+Xb6O/uA2wmCn393PT74ryCmrcANqqH36IjZ0Poj2qMQAZtwXm8RjTC63w+FS
QeDeAhg0JG6Z1bV83Pbzlh8SY+zNli8BsZKSaRVc8YCrRZayObgUY16yieV18UGR
lGU1pgbPTEF+iGaWgSVZQY13NPtLZV7SS8eZxx3EwYROhHq21sD0w/DTvqkTgl3n
NsB7MD7Aovf3IsiaB678XtUlD8eOGB6GD/cFjtq0jRsamMtsdEfkyL34ArDXrqME
vInwcg7y1gL2WUP3Q4fJ2GYQj+5pPv8Bb6/nACv8jQaJy4ymeYvo7R6yomrMXM4h
VHqAkiAk18zqJwHxnXik2sDX7Gf9oWZodwm6p5WA+ObnPIbX1TeS0NkJUaGMPsrk
XwbAeC2mewGaG15OdCkpe8j0h4jUBcwp6QkvbFjDdDavy0NY2bg6+OI8WSotEcXB
B1tFYxqvA41ROjPVXhgA14K3O6URjJpq6W6jH0jBkhXYBvFUft2yROU1JkMD+4pc
x48YRyjHti4VN/Jjcfp/s4VfXSM5g4BvCnGYeRtrYbYxT0Hh+qm2HgF9MIDT1xVr
JjeSkxqPnxYo9wI92uJHbyZYWVZjwCwAwD0d5vpp9P44Segjuwg170CuaRHRnW4r
Vb0iILvX0kFE+Ruqm2lsxDpAD3QObUPvNt2dUXx7VCaz3C08cGwfOgz4HCBBFMv4
WT2WvL1iDbnkwhqTmwQ42FL8tW+IETMnIKK5TvBJx67GkpASCBQkesCBuEEuf5c7
TIG2yhN5kkapMYyuzVmY1qRPtYTb8nqlvUovnGj5uogsfBgfgNyXqs9So8fO4Va2
JA6MfQU4+8XBR6npHUNBpFZF4KAnUPXw/cm3B7vFPioX9kLzTWA4VkIpsJe8rqOI
vchgb80umUvSSSA2pwPAkr9nshQ/jQqQ0PMmgl53Urmi4oFOLYUc56mI1/mDwxFQ
SX3tc+2IW6gdYVygedYgic+zYfrbZYfS+fl4tL90rRr17wYzUZi1cNnZL5Mwf944
8SfkJs+FzgT1vSzDWHtJ7OdgH9rkA6xN9j0zVnfLG/DwXH7SHRcEyYpjwkRIk7NL
t8b9aKsWWDgE5mxwGjkekaKi2a3B5BLQSX5MD3PolTqb3MGCr6qiwmt5NR57ttlg
hK+AayNQ6YeXCvhSE5bwLcg+RjradYWPrYHWyE2DFoHenv5rdClj7+sdGNae6H6z
VfCcKs4bFxzRBb64qfSjE6ehC89m7IuNStTDecwmlrJtRnI6CBYSX5q2PHGi3Bmj
lokPXEwSFyP59/cWzFM0ZDBpWc+L5JxN1KOi9oswHu7g+4hNPNVLGW00hBv4A6GA
DDns9n/yiBAxbMDc0CgduJjTUo+lxXdCInWebDg66RKGovCXJvWfNlAUQyXB6NpB
GvETB242TpMDfyFh3xkBp1hzRkgtrzsq4IZ1CF2v2vVS+rZhWhVTUa+iLJHS36Tv
bA44dr7q9bj9Q6DcSKHPF8S2fpkruPdo8f8ZPVWVKvlq/5li2zYyIytjt5S+6hjv
FXKbLkVsDSZp3N3gaG5M2zuv1WN+ACrlAPDAVj4CLpD9/bihU8Io8ylSs/1ktj4B
ONrijHtkgO8RDxu5oEW9HaEvv2g4/Ej5PWVUzhd0M7cPF5w5FoXJlC0YmXPpXizj
T0sm+DmbOl+xoyYsKz03sT3HYyh7VLWOwjnfkB87kxLbWWCrGjz/06Is+Kpk2Pbc
S/6ACllMJlYtGW6l6sVv88EBAyCIe2JHSgGJXo08NMCHROJMghce6GWTlJT2emmb
m73lpcJcFvGvatgeiK5SYYYr3AcJIK9stKQsfI1LLMZAs5bMcIZfNZSBe6XGqvgs
Wrv2RjOJTQKn76fLnEan+3AXGYOAKy6BLo79gNwIqZG+kc4IPJKvRI/kzPyZ80Fl
EX0Awe3hwNQ9kI4I3N6xqmZNrs2qx6ZoS93aq4Pz6QGLHB0AfIepWyKVY7H3xvG4
MTRDoYuN26HtXOdOqOALiMfsC6OEBy/G/yMY21m6i2Y41qr9LBAWFodjk35f7gc2
IhF80OspVFjDgvEld63FnfZjYlTZoGpkTy2pEOOZWTkKHIhTYKlfarO91brHNZNN
GCo35BZwy+U8PZL2wxJmf8+ac0v+GIZnE6M4shL4PjJ4S6MPvbi5Rcdnq+j19LFb
71f5gOFt+8x4nmRJ4+o9Li3YjcvxrQpaB1PVsr4bP2UcgS1C6dChEaxLsahaII9k
SsS5UUsPR5YPkXyEmkKoOWaAElTpdpR10XOTLYqp0phrP/aeSiHTda+Xwx3liobw
4CKfrTLf7QZ8rD3OpJgbSzxLFgChvcPCPoPWmg5s4DCs8sIZGQs3tP6srx53ERDK
BePyTWWkLq7CHm+/qEYY/5ssZ07oQ9SH8dX0ABDVb77Tx1xt1oZl5GSDzCu2HjGA
AD8LqMYe/Ufb5uZqEIsdQeXWVZ8TuXeW+b0+fKA9zC6r1bx5ejxQSTAXQo0/Eynh
wFfHBM2pmMVcAT6OzpWqM02TbYHPMFfR0pm/iWtXI3RTMm2qWJhbx7Wtl6FUNCvV
3+IH5TE+IsFDu3VzflT1T1v4CcVRvfVG0MFgGIYuigTItUaa9Cf4a6Z3d8xIGmxo
skleFgQdnnLSzoCkQoj0p6UaXkbNW1dl2iVYhyNEe2UmNxc4hbyPN0V1TmWaE/wa
8gpkaMFZJzqYm02UxLja+40hYBi6hj8y0xvJ1SLdzSxvYpVF0iJry20k0m3/ql0E
iBJqYocdsyoTB4eaXeTuRGQM+vgvXH+yNSdJgOD6MZ4zfQZoYat+/9c3FXqlOpat
WqQiEKDauQvM8/3st4z1n613OLV8Um3i6fM1+UzTCWm9oyYeGyzNUelTnYG3QPl6
h7LVY41m1uheyS3lRIjZ08zIE5HxdjPhS/DLwrGya4cAG8CuSmeTJ+UKk+AM7gJg
xbEphtvKlMew8RR42QdK7KhlBr1Ax8hP7mpLoAGHYPZO1nw0Tykv109bevfAcBPU
DhYzYTy9FV1vDTPmLvNGoc2ZwDW6sFRryx84bfmWN1sQ69ZeWzuoO9t+TNmbdF7Z
t6GNlS51o3UqIdIqgYkq4qSkZtcc0Dq8659e0pBjETKGTPWPXxCTeUTefAB2knx7
bZlKhc7HcT1CbniUfScvI1KzcxYWsvlR5/TNzYSw5i216OQaqcFyQLiEXPQccxLF
wHLMT2Rzo2A1dPf6vKhN7T3EzvPoD3zzo+e13vkYSxMC+pM5KYmJL6pxUkyB9VVa
g2EAsoMU0Ewrxm/Wrz44mOuH1ASSSqAayWPqQUjMZlci8VtbtXqq7e/3F6hyOx4H
u2zLsgMFHp5JDB+9B4HznpIq9Nr+osl068/TOSoGMSxjoJOUwkkAo0FSNMouAB96
Pbb8Wf3WL02gqZqRA7YaVEJ5yJtN3yoR/199Hu2PSV7aX6yVdwsxE+BsDE6wSN5L
+ZiZovYALr7FODztcH7kleoN9d87b/XWRVNqeP7hEH0VwyDt7Ov1Up0PLgluCP2n
OKuITkLhVWj2Ko4Ut34m6t9QU+KyIxnZNkCNeN3xLzRtlCQL4/4GGlEEItw9kdFV
ZF10hwjDjkqrSBb6kj10468Ll10E0nHPD7xDSxorfAY+/mp8Znbe3NUhAt7l0L24
OygUO57Cxr0TMKxWR9WpPHZBfKD+yMFHuF6pePifvrqFUlRpMbOr/dPUBOReIEa1
pXuIKHo71J3FNdMngy0Vm60q+myTtDOxDJCPb2eRy8XMC9KWydi2hesPwrB2a8Nc
JacmThak9dtBknnBFoqpbWhHRfXtx/CcDkD5SGhgJEpCoBN3+gv3SDxX+gqT4MIa
n08zOOJGADhaZ5ZK+ahZBbfooPr/OoL5NdjCbBC+P/jaxkrpfNB7Cqka/kH7u8Pt
9M+hkbGobbT/6UEamS3k8MXSOkhvFJH6fhlJLxmxq+eq0BDjQTAUuAP6uoEZIYyw
RsWUEhv5pxgbWXKLGKwVbH5BxGhhWRgSUE+7l7+Il/5F8KPX/fym2U6V1WYnnq9m
ei9pMjqyLELCW4euY0hfXb4BsmKo8PTlt6h9tjDY/CptHT7mvJF9e3dThF/Q+nEJ
qYsRettd0vhgDzLgI03TyZkb3g38q7/13S3w3kkeMVmWVnrRja6CsaqqcQ6MRjXq
CN7qKIa814GBe0vPku31YryrcWgiy7DFLfDLitFQvOeG/nFDIJ9x/NTorcMn/emk
GEv5FSkLpXiIEj4/wsyb9Qi1Yfcw+UGUwUNDHexGSrGchS1CKbzA1nGOX/rNDzOj
udi+Mnq8HJmwJ5a+SpEpiIYR+dMGfWPksTHDZihqzL0JCi3leEhrs03TSsDJdJb4
ryfax8nWmVVuwQv7Ikgck/0By8CIoQW4rNwelMtX/zADSNDmHXqhCrv/bEtqjusF
ePVlgFmqFNWra2Rbfjuu1SstbxNtJC97BmOpRy7QIzCd6Jf33d9+oZ9SFooPcfM0
/2Rv0cTmVNrV2NdT+NIBeMvnCdv8BMzgsknahVLSeiZoo5Z/CSJ59YwuEniu1Xgq
rrRE0PL2qtJk2CspKBvx9B2pm5NuqTnuyZTLNxg+y/a+e69pG0eN6hHH5KdDSAF/
tipNFx0xZgyq61IblR1P5N9oeKsXQnSz5Iqzm/+CM10Ndvk4Uzk0qtHvApLTW7rH
Ho3sFZ51J2NekZdKvyhgXgZaZtQtHQK+ZjhUMpgVxitfvYt/gY45a9NuG+32DZHb
Wk78QmxaVHNkv2v5QuT2SgZ9bNOhvIRQvSGvd7lfY7ZJqlqxWwvqig0FlhBzJJ/J
FHJsK5W24iAbNjZG16Dz1tiqqnBXJGMZSjmw/cuYmg6HM1uekQRWp6vHGovdLKO5
oz5dZ5PzIgorzll9I68Ll9BQ0AUc2QDosVlkV0BvR14OcWG4Be7M4SRdzH6zXDeq
JRkOZ4jKEKnlxxgbwvVM15hsWcDQILZcBhIhX0f8zZIdFyAQ0lHYIug/xuaYggaY
jBeHzMO9a8zUVQvMcRO1zx2ysz08942DsIu6obTvWf/YONFG3ykUMvqq2sBEYpjo
vPRA3REy1C4x7GL3H0YXLZjHdiSO/aOU4aLRAmxNY0pldcz5jNk4oDEkP0/PDTeQ
ED657zpEk0Ka9FIXPdTTM6JNRxX5YNDG71zLysIN8CatWgz2Uij7k99kMkFLIip6
rBmY7D38SyjmY0tWzOU6BVK134krW6itmMzZAV+NRqqHnWwrHAc73ileA5HAfINv
bgSepaXOTTqqq5+QrjIF53KOvKkdETCxt1mVeGSkvjHqZjgrxxG2C77whCYXC4jd
NwJ/zaj2Mke8JgbZDPCEHvfH7e/I/n0SCsDT6SV7Tn2++aHCtzsz0hA1gTYSQ/gc
SzbbJNoeuw83Kte/AXfn372Rr5hwYEMqALk8A92TLCT/anM7DfOXlLemkEH+FLn6
OfgC+Z6mcGxe3d6Od0r9wAFQEf9OoG1lpTWGLbHDuWveaDK09624OsKTec9+IMw0
C2emBFaq4HMo7r0aLkj7460L99CLpbrLUxRvgvMyb78OfZFL4sdAgMhll//f0nxA
VeGVRQ1ezaXnPr/gsyMx4q1k3Y17vi5aWSS87ZuSalShlUd/aIcVnjT69A3dswPZ
Cj2kemYfgZEWixUIaCRvbGV7ytaO6qubzb9borSvnp8Q46ci6VDbe6RTBzqSRXaw
e0qdM6VZdls3wg90IC35QejHHp47JkHFTxO2cim+uuhJgCY14P2RfZ/XW3G6fhYN
4TqMrcG80ZdDTIPwZNVgRa52cq5bsf4zWlYe3oTyM6LQD25wrBqxiNu0B1ylPn2s
yckX+RwtzGV0gve7VGDxNodXQj8TJILYGkUW6HPrGCvHF1yCi1RSejN2HeA+AVAS
3DaIaS51gA/Xv0I+5ggvq/YBn7bVanM5OEXqctPt3A/8+3Q1yGy2pAmdC3Nnt969
fHPIezEe4hmmFsJ6YIE5P7z8TOjbUja8LyfsYbRZDcMJFYW350nNxqzUTMI1hBkj
MNRziML0RFHM1i4o2QR6XehYJlLVC8yuCccgnOGsmWgiT1Kg6AYbTyXIBkpZMFz/
mt6RGAnljGviMRyMs00H+P8WESnvDbg0p1ySma4ZO0s1J7Ix3091xM5Fj1JgWHfg
Je4tSlPlWzS+Mc0l+5XTkSRN7OiMpLjsddF7EwFKIc2qajwl8jYLAjTpFitAwZlI
JxKeaUbScBLw3cC0ZYWZlmGj9xmjWQIolL443HNr9peSHfkqUMUi9lrcoDBC+xgH
WLn1/HtsLfd3dTSfpPg7SRBiMa7JeDLp1+cQ5+7GZjxegwQ8kRpEHAegpqz7M4bX
YQLGPMrFXlee4Fe+liV4ayouZweTVSJthjf+obHNnJkaO9ERxNDzyR53I3pfXdQa
HQ6Yd5YLi0x18rRK0eVpCkrMxs63cHcByD/s8G8Qe/ay0+qiQbbVEc8RD/QKX5ek
zZmaYi4w+Qo1olrC/z4aiSMGkBZcIVxS9RhMRKeaHreyEWPCntSagJncNB1jdIEw
EzAXAvb5+42Zs2GIC+SBFW1pJ0g4Txdfo4XB6tepiQexur6Cc6TuLvLWYbrA+wXr
jtUt7nrNep7FyVfsWTCzXin9cII/JQKUz8i9G/o2eBwNCWKxzg8Updl7htrsEeNM
/FJXTA1k5Cjpu0J41RqYgAa8Vm8sSgbd+ePlG+Lbp+9QmTM4nVI8+FO9atV18FSR
l6TIzLDefkWcsFA9Wa2D80uDNVaH1pI+0JXUA++anIIVE899CL4RJo0skBlViUEj
3De3vl/YDUOfPcDu5wsi+W+o5EEGKBSvSm2xpKnVZ0oahENldk6V/Y+hHwss9MKS
0x8LAn5RzFBPm6C0ezHnuiBY10vKX15aBo59QvIsFj6gIjHPd5jyeCW3lON7+sCl
1pldHbYzWvCgzpEEp9ZijRd+zKchd8CJTt5eBhOYMq6T0TNg9IzxrDQ8TkwywrFq
Z7aL9CLrPzGtcOzJXEdV3vzEN+pmuPMYJjfBS7o4r5PXa/dy5yzTmm0nFxIZU38A
b39V4brHm8SbIpq+itZ0Gc0YwmBDO7GpA5KROjCM/Ww9yZIeXqN5P2ZIgzDgOoXw
jOBZOT94jE1QDFgmVFA3aujDFkhMbo833bqDTLA3RagUrR8fYsTyNFazyEGLNu3x
JrQc3x0Y1SmUUGlHyg9O+icxQfMynDf27rFcCyLQmeYvUkl/QTigj74pgMjGZsQv
ire3R4w6kHZ9j/GGu7TWa8KVT0B2R+8bbkNAjVLITqmMHR4kCiTOX6es4hS8L1Ws
pOT/5o24QecvlRwYc68Z4gEk0d9j/ApwmZQoC7IusBc+a76qPmm2Vnekhdn3dHJS
8KKy127XCc1OslZwAx7ZuAMhGzGq+iPp+dmzuqmnoty3YLkQl7NJCAC0URXUHfM/
qfAJXpvkmYPPBsd7pTufb2h4e1Swsh8dnOh71yw9lbfDzncWc4xQzni8GyiWNk08
jl5Ah6qoRlIgnVyZuNesU/eY+poi1PwwNcHMvzqJD/rHnF/xfp/04b4dvcO9UZHJ
bDZMnG5DSAIBWY+fBoaJOSmKkuYVHp5WHpk23DP2BVYQX7ytEjTVQK7YYre29Wno
WkuSyy8pfDWhfL61534TjC2n2dOnwo6oIFr9WQqAuLzv6iiBnj9nHWnpPFECfU3I
6SKZV1Z1Qku/61t1el4k28cVvfZIwwXsMMI28CoYeDb7MMresSFrklqOALt9DuyW
95lORayAlhmU12nFB944SZIPxuwRBmeThk6r/uiojjRejCyDs1tt0bId0YLLgu/5
hkM9ZOFyD8931HiPx40BR12L9KWdX6WCfMo2FEpHUtyMzIup0EZJviykcBysfmUU
OtIsTdMMoUOLmrBQ3z8BeqlGmzfaIQNz34sXNzueCvW9dwB2nmqohGOcLmIgXWk7
DvQ+d8p66XmaxJX4SkrpY+9YUbVka54X81QlDA3q72REiU4PbelDNrDGI+n60ea1
cgDkutISjtzR5ddjvArZ7EYR33XoDFAY8Fu65IIR22qEBwwetr8LUWoRgWQHEzvC
yvKTNrzFza0IdkyvnK1dvmRvg5dUGO7iTqUPzWbAFX/86Qa3sGxvQzUKjlqLTPRC
C7vLJzd9/g31lDLnrHl+dGPuQlVcglvV681BXmQd5SW+ZwSalKaduL7AqOmvVrpM
TcUNxWxzPFlxLxE/gtwyB+iLeI5U2QYalRlRX8yBLBQLBY7E7GFQOgH8eUw/lbSa
YUdlB1hnL2FYh9u+T/QZa1ExLjW6tKeh4Zhr6GjrOslXdYUsX6+UeVcfW8WQ5YYf
+A+StHl9A1NVcj8OouvlzTBRNXcT9fwL18THVQyvVCfP894WynlBR+/LpJ0qv7jr
Yc7ZdNYzZuiubcPv0oHrXJX8kGD5zdkfn1gKrimezONM3iAcffEMPOTGxyW74iJH
w5JZmkrt5dI6dMVqSv6hZmxjkTl93oxudJwuXeP4+zUFYe6Ny/YGmuzg+5rhPcDk
KlLFILnB+NFtX5/9wJjhGbVbli3BQN9t+UJ5glvZahAF/WRtKNsPMprs94DWZsz8
rVDsweUAHUa7soTFhWZrj2EZqEcvZ09ceVFpYxHY3qnvS74nZuaMPgWDzsms/TNr
/fJkkT5ROgQVRb3WWAvbOV4txNVwr146E+tHy7RRZHVwaEs1UbGixOLr75Y5smvD
1vuZB/Ci4GzrHtUnhCQp/VXlLlFKBxIk73PqfJA6NfQOR3SiouwRabQKcS1NtEnW
gaFgX5qxKYxnSFmKb9AUgyHVMFvAT+JhzxxxKMojGViNuWg8fdEjEGQSNbnzFbPc
ecOJTDIGbEmxmEz8ffMiH83cmnIwcVQSOppJNQgYnQonzmkkuO7zpQn8WFl8X6jF
iLKSJjXjVPEvpSmxipGiggpJDkZ1wv1ufD9QNJObyB322ETAd07Xc2OQCgNmdWDk
GKWB/jJKD0f88mtSjniyog6kJYaR6hmotlLRIe7CMLHTL3LUyMVyG5TnVVwPWrwZ
yc+7U34FR7KAOOLDUMLdC1DFU1HJnVV5JTKNByPf4jubX4TzUqaUZIdHQxVN96si
dT316FPNdZqO9/hzw3MxdU/1kek286rEcH2CsrLDWgglmr6r84GsBx6Jvy/vI/VN
FQN/pEvrazUdmZkp/gfCY77ipzC2LniT1Qxex8+th0u61EwxvJ+raouK2WZcHwKx
Vom3G/jEuYdt+IhIiorxBQuxCmlNpnsQfThoEYKt1ilkXoGZRw+3sbQ9X+yU0Awo
JueA/Twin/n0wBvqv/6scoUFf+Hx4Eyqf62dk9WQxRMvTRVqeADfz7LcWN8WvQtU
xPs0fujILxTxD8fV8dHYubSOpw4y649KjMKTGNVE47Z6yY9/J72hrnc/SoUjCR4f
EHLk32UPvPRmZ2yYJ3rrTIMdte29UGfNMJWXXdQmNZZXmtZQJE+60RI1ssiEx3mz
/vPugzL8t6nLgqtJ7+YVAWAKbb+zWkBJK7H2UjAUo9XfkMfaEQBKIBIdm+tvpd5o
kSi8hQl1i0U79qQhlvQRBdK62T7MrS6lTDc3magfq5p2e4U1xiKDmjTDoRf+Dsuq
L7EeCBMX6vGd6gDuQA2HFNIMDVO0YxipXUfWZOPegbhhLdss1KweYZENV5LM82T6
mHtKdIJjFZ5S5NiHTnptcJ6Sd1CoH1C/uX8c5aZMZxTSmuj58xrkvOsRHOHLqFAh
RwOUVxS6ogH8xoezltjScJd96/TOEqVeHel0GJfMfj5rumq7GZdSGNGmMKCrDcC0
6DBfzJXmNlXl3248XhdLSUu+o/n6RjAtYQMkHvX9UzOm+TiUwk96W3+Bc9jhIXP6
Z7qZVYpCx5F35sI7TA4E7seLUlG0UVnvMthWOz2PTZvUB8j0tKDcxuGrXmexw5/V
Mw/8dIbaeUpILdVnTHSYU0rigSik8b0XDqsTmqPdM0yAJjE4Ra19XYszy3UwkIxS
XI8PDhKaZ/QFR5Lub55Rt/LVe+dTIiPikf8R1JXbjbi4Eb6CA5p9vl0yUBKuSvIh
/SqKVxdpgk/gZZWvGNedH3D++SQ8UMqimLbuM1ar9pTw/oBQ91HTdqH+3wHqUp08
rS+/ZFiSs+ITTwh48GLKsNWN2J29OwxZBk+/J7PpfrgqdDPYAcvsRZHXEQYPlDo2
8R5Y/l/g4XFaMEXZ9MDKom0MibR1UvYbUVMDhq3lg1Hu6STTt/5JXzg2t3Jn6ya1
USVypij3hyWuDI9fv11Zg0Pz3rwTynvkTycELVfx5x1O+T4+71tujzOGpqKp2qY2
TKj4p6KJWaj8JwMyFWOCylfUMmbkk/2r0vcZoJ9tirGf6TNSnmVeClYCuVpDv1fM
YOt/NFwerdciqgabPfpqMVE4A+Py5xvJOWlvz5OegBvg0F3DSRosw2DGpdKdMv/y
lwOD0OyH8oqtVtkdIvQCD6+KyT62ZOdpUsHpQyEzVI6HbsFUAHDJkaC0IsOYZSeO
FdNLNifkYIJGakpFsh+00xmWEuu/Umy0PrjHbe8dp6Mpq+YHlqSR8SJeWC0MAE97
Ysgt2VrCOfTn/Er+74W3xAaLGEKHdJ25J3/6Q4D0HkBp62E3nhCAWA/6C3gcbvFO
jT/t4w0fF4HFIKVt45xNG/OlsBUgHGujJ1vdCPLdN36F+Hji0X/Wi4roMqYUjpqy
LPoABymxCvhG3yU5jfoqDxmt1+vm4zDds/QDy78M1LkpU1k/LpgCzycvR3gec9qN
B5p6ASPO73TUahCD/aC/F6VNnezizZlBXHZKtYCdAVzl0/BYZMJ3LbqdiDErWjwg
QgTwkXAEICNZx2+Qpn6Dtd/sMuPfeAHC45ybRr/dPY7HmxYBCL0tPqvMFGO33bpc
UJ0cBGPZPVVTxmGGx6bs3uTsVdYognXYzBg76w1YtzLkTFD2ymVob94YPai+WEFh
OlCEOAaePn2+oL+HJA92w7L5kWdVtedw59/777yRH6bUvHXyCRIO08cCHQ43f8mL
CkI4bPuKwxIN+f+tUQ3q1CPWW+1bZIbC+iKp1BvLvsVaiOjlatd6M4vJ/3X+gWpq
8kgT+9yVQF4b/2GD+yLXG+F6Jqu4QL/9mVVTuQbjSoIs11+n0UYvazecKHb3FTG6
vZntLYceWlJ4JG/BLwvGAFKrvkPUZndJJtRycQ9IvG2VBk34DO23lDBFzpvG990R
FrPNG0bItsTNtKw+Do1WDetqIJpXnOjZDydBQ8wRMv+8Rb26VMv0aCRUOBhruLvS
K8foDLOBT4iTPqcF3IFDPIVxuEyQRP73pAryWmHFPF0uMGljTaJEXPkG7gGBVGx1
eG/Nim6VNPqowrvPjBB+EGpff/+V2JcWeW6iLJe3TVOG83a5tiw2ehfrGehbbQk/
a3dSBUpsa8sEHhOigTm/upCrJzEBScqjcRJN0FXOzEbCgmNpH0l+iBnfCVXAccpL
4eaaUYi9EzdBUqvN0nF2jEnMrHGifu0Yu2scmJqvV2AHTDdhp52CcNv8BbBxiGYT
H1+WHyE04FF5oiD1G9N1KM/n6nda5jdN6Ab/kk0PiQAGCitZMYFLKiWZxKfR7Bvi
41RFFAhXnWLFaYP9y25Ojww/4ZwqLN7OeZdGcwJVINgA+vL4W2UaQuIcfql3vCXj
vPo/hCDxrggIkXcOjlYxqH76JdzB/hxKEi/PXgDVIWxFfcprIDqx1T609aK1OHJG
VAuu+zDf1cZenMqkmxsI6TOKaROdO1KZX6aoZSpYKRwGaimppzjzCW2uPFbFFuex
UevO2E+jvDMljkjEro4dj9Yk+ynTF/kuWlcGBA3Dm+QE5LTQrOcaFtHxdQzzX4mk
VSSM5o4mg1euhAk0wSLC19sET0M6RdFupcWEavIleWIaWJ+LIubyyHt2DFy+UzgV
ROzvgdUfzZRj0m9UYvaI7lNnP9SUlFgP6vfCM6n+SNdAJi/YGFSMM5Jo7MuKRzny
kglpiSRsJCP1zRqWHFvIXAq7cWvxL76+Poc6s8gFXO6Qj9nXOaOORlGM/5/COg7G
+5z8YB3NaiUkvoIPxfB7BYhlM1c9/QWEooXDjsGkVMfRTTiJDvhfw1vbRvqzCjOV
UXhdulFmmATj+MBQCSYS5fjZb9290i15o5RKHBjNr2GW2EGK91ie3BTMlvztINED
LGT2TNfjDJ+cuN+n4AOC3TsnogU895JtCY4f+WxOD8xeCs9bQzywoXc4o3uY4kwZ
QhBJJ3d7kvVqNJPJ46mcU9f5NkJn2MZW07uwQ/8u6dVH4NL2jacky8tdZGlzzs5b
LtLrPZC8xtZVVnVGij1eeQphVLMXYP1+/VygUtD8cdymSAlYuku/h2dXGYAUniWk
1BV1xY3dJ5UDqzDHGiXW6RLfHkORzp+Af3dus6lB0G3eIYguMg1Z/x84PJxEaEbh
FPo5xCneKec5aWI8cRzuWjbeElqqhkYZVO6sfeBEdlcvcf539a3kWEADa0q0YLT0
omR9+dbN0uBrUgtap//Lzf7+QXxJusBgNb7AKbH/wD5+s7/UX1n3yrlp4adbdFo8
Cz27sKfSycAxM65sTeCusvQLScJ/x50LCls/qWirXe8WjvnC3xfAl+Vfz3nIPLcM
YoZMp1H7mEANHCBAEZueXWWWLH2IodrhvIoaOgyyHSRK2tTQwT5+eeB+bDjMYCnu
c8jYmgGY3vACoPLtM16G9Q0cSmMcABo52M0Kw9bxouWJZcuHBSGrA8fcIOTUpfus
/wYfWqCX1c+JI2EQ6jGZdaDCdZh1GLp/lhBsmP+M2ejAAj8sioiG4XdLkG8Mum5/
pnPc5eRQ5WkLYNqGRuSWFHksU3LTSIUKN3AUV719mbS3ALNxayOrQzNH8bqaMED2
l8HVpzHhfjgoiL4fb3x/bZNhQFc8CIBgE8ysdZb8H3feserBtSM3CfpdEOVpSVdI
iwyY8JWEuHqHoH6dS6Q6B5WeXkoa1viOkpP/fkfmZzW0dFFm0DPeIGY7ci4ZSHpS
BeLdk1q13vr2gLtIqKCJbxJQDmEaomMSiSo/Lre4lKUbYtkJWDUcOFgMxlabxbJK
eXtVp0PUDVcOhTa5w5bieI63xw822N5sS7dX3nJRfaiC+AvV1JWLPkSfL6DOqTTw
J+wEKCtNt0FLiTvszcCptcyI0Ltyy/zJR442x6ZOFavMQe9wmOMrrJRpG7c16xrY
1pTC0owdpRHwqi+v5Yet9BWDqRvwwQ+CmQ2GCH3DTGZQXauxv85TWRxeTdQjFi/5
vZdlt/iZfB0VbtPgkdQ2veVobyd+T27GO52pZIrVpfRGTRI34FaGgD40XIAKPSbB
gj4/1dbKVy6ZHKXiZcsd/cNBKH8pRfFOCXSSZhukC4Z5VgMImdqrPlTzzebl+1jr
rHXVVDgi7rgqZnaU+nJf0IQOokDEhBgv5c2isPGw3EwLfng2io6rh0gpesjgXVK+
z93w3SK/8eJS49YKWZbAH7bx7ZkhxWUtIwqQ3oTWWHcF/cNXtBp0Q6NJuL2BZecl
q5S+0mKTFsMJRy6vxeEILvsMCsF1VpwtLM3B8sGyWzsee5FMOT5hVLzkPpl5mmcJ
gm9TXqjy5CdR1uyrdilGbPvWTDz6Q+GgFIIslgUY9d/sif86Jj2UI7jZEwLpnDDv
AnARsPp1fFUHUFgBeJT3fBhANIsG4+v0wCaaJfAbCqHBaXfX7ecsb7gScLQ79hkq
oZ8AGYxZG5vTD3CddPt53p54vqbd9v/XvM53RmNhh4xy8aEeS9LTZ3rfhdSkHi40
7yx8Z2UPHVJ4FndgyPt7lL3+5zGvR/NIO8vZa52BrS6C9GUQk8pe8VImvDZi30eZ
7LTpV9m8vADhhb3S4ByN93dI3f7Shpqo9MJG8OkDiuyEZBnWBv90BvocQNS7Jsiy
z5BaTL3zcWcsoF7zv+z9C48C/tnJTbUZFv8DNSh0YYJ3MQIAjnDwp/6A/52rXhL8
3wryFCkx3amvelld6XoMg6IPVV0QFq9TC9s2GEtktHOX0n6zoKqWtplE+0u7Bb0b
UgkUCmhMPVTsDLxIdpcCqeYNrZdoFdijgwxb0f++s5Tisv+GX9tzLhasV0tS1fiS
sQ/wjBtp7k2t67MDVjV2t/JUjTUtLrPDYdQJfGw/V9IA+cptajkbzhj/8FqOQ7Wb
meXhibOajy4u0ePPQ8RCxbq/g4RAW/awsmm+VtFVIP2iIN24fctugQ2pTLLY6ZsT
m9xtsu5jwj8bvxVQyoDN0aFOCQZHchA2+YKBvprdWWO3g6ni93ECH5eB094qIc23
5xinculj9nJLY9pdbqbqMM2O1errPAOaF98BA/ps8d8qW7sJjYHHYDRXdtjLR1si
dZQoXTqAOkcX12dNIN4QEl7g0LR2WCnxAF7bYEgU3Oamk575K7NsHZckj5Kgp5Uh
HabmvKWfHtPbeNu+P4fMDTQe9hBNH65c08m2lxILdsh+W7cLJmUhdY6Lw7JJGnzj
woYrssluPIOd+PUiLNL3Uu0DtaAvXaH1rLdL6TzE+ZbyIA5K4GX4T2EgQJZebBI3
32RCqxEWStlNyFO2E+xFPIUzl9qqVwygZnQjwEk81PSo9aD8IVPX4oNhj9aibTqN
+i0oizEvyr2chWymbGGuUnlBvGrcv8z05F+8PP3XfQFC+rpHB4mxdoE8aBlmsuDt
1jfBzm+tfrM95Vz7gyvV79QdtJV3omKIZoGbTEDZcE1/ZBMaNOSSFX9rYhM0+12m
/C8XggG/6S9HVzjmM3zwcDDXUZ+M2vAZAs408LfRoeRTpQnZd5him8DY+CLBJ23H
VIyyHUI9VDYezG3vR96ar2AMNYNHoxECCrz3rjMSDtVh0dKMXEUhIBU4S5Yui40J
adp4rdLB/2dSbXfGr7YEH5zzCcZ39/YR4az9cexMzJqs86JFJvaw2mgLqq/VRs4w
0+3Y9rLS3/cceo3gJVqvqI0jqyK57saFr5BG/EEkqaO8ttVHrl1grbECLhspfiwl
tnEJHF+wl22L1VJc6WwoGESGMfs+os7Q6XmypjjtNZcdLVgg4C4wd5CzXOLDff8B
44J8AbhVC5mnIlepyTm7z3BTqAmA8YwRmmenrk0UK/rcW2JojhpSNOh3CFAwEIq5
xCnL24eK1zXftlC4iK908qlxPc3EYQXSNcTAK8E0cHeAfQeH2FWSoq8EpQemPtCc
/ssBskJU2waveqR6MrFXIBPY+aQN4V9bZiGr6Jx8zhdTS72mFL62r/5Ns+k7wozN
g9H98puWV3SaVOKP3ATaI383ANLz+TkrEDRKN54fMnuS54MkcVbrjrkj7ZfBQXl/
a2pGZswH/NvvCpW39ySBO6/rfkJd3+8Iw1rI/3txyTIvbNrbuETEx3chLqMrAqxK
1ixLzc7j/W0Uef9EGyrUVoNaI6qrF7Yti5ORSTprPtX2ZbOuV2LNxdpdcOFcpLz+
tO8foqJfDQVc/6u0UF8SOGGJVM1BsMyobAukE6tbxDv/Dw5Me3BX3qL8MR5sd9nN
Gl6GhVbC4x7MLdpJ4AtWpsWbqa2IHOzw++X/IL0fXQP8YxhV9TWm8y4nSzbmyq7q
F+sL86xHZziULefeJ3KdrwqjXFoIDlgRg/9pHWV/TsxkVj/fsEYs0sUE+/+F0InB
dcnFBlEiAN/h1APOjUWLpEOoooDWhSapP6oIpXICbdFi33dk4oZqqV3v4h4uGoSN
zwjFRowWLqaWdTwOh91Z/0ey1pwI+LObq8mQHcepn5g8oYxNGHK+q/ZbbFA5XRip
x8PApNoI/qyastiOj90+kKJCHivetYrtsQTkQ+V70260exledjocDaZGmIt/AOPm
mcojhl95Y1H6h/0U4HCSy8DXdBhGtp2Z1LjQ+DQPXvZ9j3rr2WhdJMzkVYbtJ7lE
dVGAiGtVRKAsfC/IaQHrPsRbpQMMxQzSEWFPOHeKYcmgbsfirBahiQs5QaG3/otc
i7uvgivJhkxs+B/1T5wnmGoQbtDsjHsU2ikpegWHpi18vwlBUsspRbujcw4z1nW7
Rdo0unC1YCTeZcjnRN+p23eP0QWG75KlYC+9MDLBnxXd+kEmI2e5U737/ZQJyJ8F
9CjqiIeSQn830gyhR2btgMGjDVBalI9Zh100ElF7BxlufEfw6/y3XUMDEEncU9Aj
U59b+Ru88X0aKetesUUGxqR4pVPFrFXBS5B1Cdx0WMKy4b8JyV5XjU9VsKvUxMnw
tEKsb8zjEaZAgIFbdZV9C4TviuwgFjUL47fO9woHD5AG+V71hYkuetH1nOiDV4eA
V+RyRjd8wq/E1Zw6YXAb3PFzyZ/FPB+oNzSzqIpgvLs9PTJZDHsHTJ6XZi/2S92k
BjP6mc/tlkqjVBHoAJdozD6Y7ymLP01N4aNMUpuwtGNE6/zqPiEnoesC01YxAl1W
G68AxAi48g5khfpYt2HBYDoV63q56wyveXetMfgb1LChrB4ycvgKMildxub2QUgl
yelDDMweCZeG6uF/GnlFLbL9mW2msgf4bxiETUl6/n7bW2QwArd26fFcFyybRhyX
42DmKaob3wo+41zx69usLPVkcvT2YwMqt8mJ32daJowgt67FHADDcB/p+064VuzA
98PldW3jlCBqgfiRUOr/xvOMYma0xzUG1LYWmoHsaBBkIWxYD8JpQqkH0Nx1Jj6D
vvpel4kpGWHbly0loj4Ud4sOjwFTHAgidpoajmuORgLDxiBEe4w7QtOqVxaKzS1R
uV7QuY8dmLEv9PzKUkg4hAMkSjuNfhlhQTzyY9GbOr/1KYt4sSYHwYX2WqYUlMGz
3X9aBODdD2mkT4hzCCU5T8FOo5iGEcYbo2ylkXM3rFWTD16IXaUycaDU3lgJB6UH
RTiv8HHQrCTtIjHw7JqP9CDsL+Wi4464ua8ogfUfK/asBsRazs1JpzKKbIj6O2Z5
/UwluT+lOC2F/3G9DBK2Ub2WePLMeZnPAv1pAgCwXgcBqfdCKZ0EGqe9ad9ApZI6
tYwTqf1FBMz1qfL5gikWJ5f1zvEt2RD3TxyaM5belqD1osTwX08LlKEBFKtccoVA
dlSbfwSfQBZ5PtqNiRkzSe1SuTjTukacR+wV8snih3oW2Al4kC2/cU1PPVsCTj1b
RBe9gv61TW0BpQYMNY8sgDqzf9XFiCaLTc9+R9n+3T2uL5NyVxVQQGt0xfBrCZyx
wM4yu/QVj+6XH3esxZCmcFBFYu8X7R0UgcPgOTGPkAxq6nQqtjK1X4/prStwl5K5
u2BzcZBHJCDn+DYBW4xiA2bK57Dq9G3clIVVQhGHj+HF/fWs+BdnEQg2/YBbXK6F
Y2cocJk5PBbAxr86sNrMYFA3sD0zzVvONSfxTOBSBYovfJSvEWaYTxODruUwHSr+
TGaa0fNyNoBgIo0T2Fo5A18fw+4O12roTcstLiFjgQCoXatbRvATucONMKzIcXIY
NgB4ALjwixWT7CocYqWpbSHnPsFMBaV0s3KTFHw4vedo/KRsSigF7z1CoUQl4GKe
bWAxNY0CwNDejVBDHOjZ8SlY3QrzuWaFwpOD7VNMNMZth63nJcOUgkouzZEIFrKq
u3qFiqPbZ+U8RMobsWS6ovleMHeWqFGFyovg/CSiTJfoI3wKK+Z6FTZse9m0z/Br
1IwQQhjpaDhIK+8b7OLz3ZoAXCk+pIj0aUDc5Y3dIWd/XdiidCsB12bNCrk+jZgX
ccLjWLjgR9h+UhgWGlT64unP+wo7TE3Pm09GKX8Fn7vOPlE4bupzQn6Xyg6DBRYC
hSwLufo+fYv0xcfXtqjo3PBEisJNS3rPnOTeB8eCwDW2PNTvr3zZVaJR77mLPAeN
UYE6Qpi+TYwc4rAvYqSnhRIbOnHaiyyXq5q6ScJdumIK/t+0llOGMAFaIFaNa3sJ
BiD02xBJGZr0h1MGfj9BXArbFu8Aw6Sic5tpbSROzTp0jXJnp6sC0UQlgwYqQuy0
Irg6FUfkBvc5MN57LNViVDEGz52DMGwxYW/TiCTgrsLKRWqqWnmcy+L0EHENI+78
/PBJwZVH9/6SEi+O0umD9xfDJoGACsomHqrImvvKyH27Hl1eNr4Fa2StyqadWwyf
63VJ5Pa+8dUy3HW33SYTRUWhyrMEGwtimQUybTk3hASvWbgtABy+FNlLh9EE4u7G
fGL2/sVKGwfhtqbeYu7fe/0zH1CSVcJ5CPGHr2MCiQnJY/gcdyTjqs6l4vryqDjd
siVQeUl9iH92s0kTS32Vc4jSQ2afhvHqLnyFWWAjxb8GpbWhcfBC1G+2hVSp8MaV
PY+orhS/Bxm1AaUZgo5SiUjvdIapX7F1ABMFpQL5dBSNg020XdM1vMi2Ce7cBHjd
VpT7H/L0s3U/Kkk+vBG+WgZL3SXOurJ23J+yIOJs45eTDplx/rMjZQFrccPWfdKt
N3vTdkC0ECqcb+eKzaxNdXm195VKASPoZ0jcjhlejUcwBEqafFjX2KrP3jARaP+C
RRdc9k3nJA4lcRz2Q9fQbjPrlFdHRwu1ueYgmDLWJDHJSNXTCiraN3CXvyjZPm8c
Sdw83IDGye0XXmjEGvj3nXO54hLTyXINPW+EuumpTxUm1v7TAL8HbJCTr/oP6fbs
HKG3V1XBtvAcNWZXQZ9mIls+9dgVFeuWinYmPWn6wd8KKDm5UgeDLu1f7KkUnRtq
0hIT93TAr5ERWYW1rQEm8qWeLm00jnl+XBhslg6Jfqc6CTwAzy4r4o2p8WOSHjaa
VaiOf89eI0IOMbC3ta0wS6ar4EUFQow0JclGNNi7guhPTyV4lCEXzEBwM9N2bjk9
SjRXCIy8/Z20BQk28VGkzpIJuxw4xjYX5ohC5yYoTBbXY/lC+KVuVd74wmZkXepn
d/wO54LamWnuJskFZhxrlEPtrnKIgsKaKN1qojWhsd4lXEDO0j4bQRP0EoDoaChG
ZjmLkXY+NCv7ZSFqcTZEX9bkud4vPxhkkL6Icp4WztlNy1/kSZexy0Sn8PC9S/XR
U1QFiGMSVueyt1UndYMNaLb5uinFbLmBi9oDVvQ/6tw2NUH9BOw0fNzLeuCdhXNX
2gAOwn7kagnzFD1ph+Z61jVJ8E+03aiR3MZRzIXTn5x4z3+OSPPY9rGSCPmgdkOH
nPoRjQ/OEZGKnMCgB98DuIcwKHA7mbDbyTn44YaRTwj9mysYH4vDfHMDDqoeIraC
OlpE0a3DmBY76KWbKEND8DAxOIYcjg4OltE/c4m7jQRA4/jnWpP0DBh/NafdUxyF
SK2IUpg3GWZtvWV+vzO5QKpgnksVdce78b9Jwjwb5O5IrGL5+IrlbXb94Ahr5sxG
FFeShTisj84IIEoSONT2cb/tA4SoHsWY63MG+0E0iP+EV7cA1P0AZP+Dhz1FsTal
urWG40xU4V3fm8yL/9JcujwkB5jJ5qcwuCIO0A/eaeJaHsNl9Snn6nOWzgFmbMN8
33EtvyoYEeEPb/cSICKXHL2nZnT78c6B5MO+7PEPPgSSGmNqSDArVOAO8t4NEjG1
BmQ50Gpcc6vXgtBc2k3rIjdTWRVNhvtRf5W2rrFSFT2zeqbo31PL8RSu7E5eAtx3
qGg/d/Se1y5/4rvlN2tG8G+5CTJCgCF3jbpT7VVb5Go5xsiifZfFfxtoJ+Pyl2QZ
sDe94BWXEXWJF+JYt96UuSSh+3zkV07iRmDV2L7KUW3Gr1xJojtqqFKEeZB6C1+Z
pPjvYG9Uc75mj9dhVJ2iBTXpRtVuclwBsFgdYMQV7VGKnRP2AZ2pEUV7IGEfx8gn
O0tjUjVVdfnk3/wFtnHerHOFjb2yFDdgYKJ0Lvud+ykXTk2Us4Kbiqt8ZXLNiGPh
Vuhtyn9lr4k0ZH4BGlxW74+AICs2xJE+KdB/a+lqgSkGV0iPqrKUGpDLnmlIumZ0
wa9Ugfs5lypoAcgydhyUm9R7jhgVcKteu3gUfdIyhXdoNPKexAlFV296DnYr1NYW
XaBQOo5WrtgqgcdFluhTk5LDD/hoXUmXxmjzXn/2dOBjfDjTDfHYvIsl63QQVxu+
bQ75hAO2p2B8ystcyFDlHsXSDqWrLNBgBlFPsApzi2J3vCxt08/6uKxJQPudG1D/
8pj/iAQT56kGLsO8+TcxFSfKXQA00lE/pitj+46l6Yt1S5W4rlEQtUgt63AnshF8
KKWTtBUEkAiZkV/59hJ7mKVyXUB4AKz9chdHgIwTT3DG2I7cq9jdCF1oPFiTUC1B
27v/iRonZo19ZRVmR38Eg1OEN49MoIRr9lmYDw59WpJ8ph6yIYxuB3o1lg57ZnJL
svMFL4btrXSP9IsIYmvok0hHdtlCHWXlcuF3uEQq/dVNoN9bZd6N44fLZEy1ZjSX
lJbJLKLXLbWk2ezCOsdoh6M2XPJcmlf+SD8hIywI+HQByuJtDu4+cKtnNlsY/58C
NWzwfKFkFM1CuKV9bAYrQlhYhx0UbhwtB82EDnDZBD5llyIc+jEh9VH2CPCIlfvM
L/BR7Z4hbo5U774GHkPYx98s/vFPT2yQZ9CF9R+LrZm2AP6Cgi39Gy9Tb+EjYUQ/
aTvotrcEZAlUfYf4+q3Md6U7T7KUE6rh5Q0yAA0nXSutgl3bMRAXps0TJLKIbLpI
86JASoXOrG7ssAmyg4g8jHCDlKx6lDt4A1QNvJt2oL7ww2jN+mZbmUQ43AGDc9bC
3KormgrzsV8FZMo8XkXmAxxZNjlCOihOcoenrMS910sLnbopCgNZpE0yL+pOKvGZ
zqxZnK7s86EWn/uHTwx3xMplQNtKtHhxFXZgT8j/viZK7od07VCyX/uCUHxRGkbA
CMAXUSNpaVBQ/8zRjWTRwKKFETRurGcwQncwTEsrYttbmu2qUWDIrGRe4ebaru7h
VHKwA2tejzrdeR4d7cgt47TUNeh/uS5j0J7akr87MElo+AR5zeWcSTkWRXEJenSN
SYIfP126M4OxQmtanpOZURFsXLXLLi6S3LotbY3ZQZUrNLp6bx9k6yu+pG7L7v3W
Bf179DuB8HeF1tpLs9uwARg8h71smAGrqmn5iuVf+yvckuruBvNxDKP6ZOV/O1T7
6fRLXW3xGMO7ccmjtK91QmnIG+ClR0Lu/SlX+9pSDW90wRIKb6AYHUSOlE4yHSIX
HUiAIsBdH1PRDfqJGpT30x1lDxPV4hsWJ6XwlWL4AZ1iJWnv6bXv5EP8Ll1q0ZP/
Ix1/6i/oNDJrsyNxWffHcU/n4ciRte0hUDz/u0NVnAnk96wOUza77e0ffeSg7sYX
8a8ZYO7YvykjkKj0Ya/iFMK4TGkIam0KypozSSZPiYGeaAhdGEtJS1AHDDZad4RL
9ghaNJmRNIMNhhDAcciY7oFB609jk6bi1A5syibDGbHrPQ7i0OIdCKddQ1kDKZUM
EHGNvm3GBqR0xrjE8SNAg7Sf3OmGkZYWlRkldn7Q9I6mHybcJjMB3jic39Vn01Ez
DHPbHFzxHDwFn8vOGIiUAya9mlnjiYwt1bxzlIUOBqvoo7NXZ1+BrTeIOu3BNIhy
EBOfMq+UebtJlLlLmmGDumCTNuMXjOuafsJGmCyaFx/Vmu4SOIILGWSOh1YIbBKy
7qYL/e479+eAPZA6htpftR/lnxnRd8bLwLgqYfpYH7YWsXY4BFvYJ0NMuk/hI4r+
c6oBoZRmS6/b9tRfXD5LFpuWFh0I9yTgs+BhYV/BvD7pblolj3oNH5twdRm5v2bh
dhFQweAVOkvG9sK5bLqsbpWPJA5r/ClpQsgrhNJN0S1pugW0UNOmaPJH1pxydtU9
apP6rYg4KuaNVcnuQdg9RKNasotk2Q8YrjCl3c+KXy2YoAALIDFjhL96NX/lJsMS
/S8vkpFU3epUs8cXZ53oGjGb0Or8xue/KJTY1oRhl+AU/FZ1OZErFI9KraogPZcD
7X281C3GGMBqrgIeJWBO9IJgtNefC6hLkjKLrN4dH4j9yajvPZaQA1mn+RhAqPrl
Mfw7GOUgx6F6PvnJc68hqOyPYh7m2vfa13hb1bBv2QUlAfFh/SISYEIOMmdW6G4h
RWwruPnrjrQPUmt8e1olrUTmoibYOvoBi2LaQwDP2UO2U38JVnX9tO4umEaTe+tt
Ea9AWn04NK+okNiyc4ZkQI+fTewv93f04+eHBbl+z/FZPf8uTOrUkQhXpUmdy+1K
5cRFdFmtyfCazst9gaO5WF4l9QA0kJmGiWtbXOtdrKNj1a13NHElw1+6GAw/rXkM
XqlmSRJavkjkAcq4pA0M+QNmYDdxrTSAvA3m6NqiugplCdSWzQMgNsF7U2uF6Kti
dsL9rNFleqZkbTVBJmxqv5mB9JFdujg5g+mrT0Gm5jq/yKz3zoCZB8klk8qNoMA3
pfnTICh522arNNHShinDX+u7el0sXouYb0I/XolJDMWJ/OCB/pmQfl7x6QgHxOnq
KOuA60GVMfqnKwzQ51Esv1P8QD42uCbfEqzx1d3TryL/xNZLhsjysrxyrNLLkztz
F1QWJBVgoltZxV1OBNV7ZC1QmFcnE1jCHWpxu82D+dEZR5lwjhwGhedYLBweqy77
pnMsSUz1/WW7qrURfGH/wZPSazP9OUDkYubz3ZEZPEb1yw90kIaggNgzEEGH66nh
I5nZG1Y6gpXBLA7gqVtSKNad8U9icDQ/XNHIvOWN+vygEScMW2VGaosR+SWdpB01
PJGlfA0Zj3HhWLx+fG0IsqUzCP7kSwE9MrzGrtkKZPWlXhXb0VUGzN6GkPYL2daL
qpKKNscE7+D35e9adeCZcdKbSxFK6jBB4KUXMgbeJ3kGS+2WyrJK+lENcZI0PkMA
YxqcfZOI44a/OWNVWmPa4SIEWDHVSr5mtOpw1Gg1dngdoTnZ4fo6578Jy+E7DrnP
FtYZ1wCA/qFDZB0PLVPQI0tHFlIRzskyB23qoq/Zs+WRStIY5sTEmREN+AgCg3M9
xgPyaR1cKllnGbwGsGstWG1GWpnrIcr3LYhP8MAdjzu6pF8pnrFNQFEroeuSXEp8
heN+KYnEfDFiRn0J2mDGGQmMFtUJROWE3muRVCBGP4oZeptLuc/ejiY9eXlEmeyI
7cPqC44S6CReqYc5c1kf7u4g1c/nJwiZPh1mDbknl4x45ah3YZgug1a5lFcJYGmQ
gmOtyilTifV2osnZ69cPNvMMBEvPx7XMsiIe8vGUgz/pF4ltU+gSufX/4VocalOM
eoKfePTZmq0O13T7BP+hFun127V25s5uHJcIQ4wXMXCg44R7puc2tO0Synf1+QwU
3QMsGUgNFC8bY7PMcOyRK3vXxirRhpMNSovtKgS0FtPQllzfjx3m2phjXYQa75iE
fy7me9XiUqdyqYgPGvcGGLwMiuBJilTjJlRI7K4LV39aGWWYj48Ww8V5V19qQLFJ
1lAZXRKXPfc6W3itKaS0ry9OYIabvPoub5iBlL9TRmwWUek6z9kBsTJVFpOKw6V2
66RcmdwDVaQ2SFV0zvqQXWxW8qOBTCgj+0B/cgTeNUSiquHEuCxq7qGI1yW3Ou5s
H38tny9U9HgKUbsAuDgX7LSCaaC0oE1cHn7lLCOPJ0oigECwqv28wcqpBC1mkSir
eF6FnDby9L5rBBIlcms0y+ACGDoSlRvBAutLy6ufKiGdAPNqoMgXLG+ULlXgqv8s
PyXCRD+zqfPMW1aiSng+bCwLTuQm7CyA/7NtpLajGGlYKsX8TfRQQiZuRyUAEhSG
rr3U9pclJOSsmuMYYwV6Yywki/b0p6Rq/aLfhbkXkjWozSZCEvIDJ8CBBlm6s5Uk
h5iNaRN1E/ZbqPqFwqG+zSqSK0p18XMtzxSjnc8WHqe+sEimMW2Yhuj51JnVbvl3
UJMA923QkciFZKL82wC6MjpTNxx6RfWH7YIQH1h3O7UU44nBx2ICToD4U2F8XZPD
Gqy26UJV8ypWpZzyRY9zdmgb5/2giWUCzdBrW17xy2QXpc0fOe8NwqDFJw+W/+dN
w6y3KYHx/veDld7IuOFSr+TtBCLzKP+IuykIWKw+FBdS0dmoycwB7A7D81CJhdog
oS2lxf34zS5zYY3KfUNn57kiI5qI+mvhYROwGtqwmq0yVuLCsmOeoUcWyIv4OMQ5
Gdov/yWtq/awCgz1llJqjxBuUQ6DdqwhOxA6gNZ6ux2lwIN5d24p9/UCMiY8qBdU
4IqTzFjELmnEBtKhOHHVTSQhrIqt39RoDuFN+uGvvDe4u9eTyM7QqRsr80vdVEUT
KiktZzcXY45zZh/yBazD1TtH8MC78scRb+RgCcx/IdIw+cgyvkl4yIlJkmbG7HrI
wld0N5RluoXwZnh+84FL7/iHIea2Xg17XylobFgv2pQabAo1qtmWxksH/lz5214S
adPJ44KHCrpynn9+v/bgGKQv/OdPebgYpQM5WU1mcfRMZN/jLk1CG2BopAUvkn28
BGKS2F2y4+GAwZ0TDjWHyj445kVQFZBhsKcsk4nxRLkL5O+Kn8DpO6d2flILnJ/m
X63bhHnylsze7y4VF47t71Cv6TeEr1r9CPgHgEhQgSdyH09akJLaTkqlFHrP3PJV
OPvW1UqpB0FBiCnD2OrtBMy0HpGVp0LjihyjejbWpKx5w40ksdFMCzW8IIq9VIXV
xw5lRMfF4/5muYcJ99qOUxvHbrOG9hUqyvvJJ0QRhah0BYNRy9ZudFmKZem8wexj
DAzK+CzH8X2d/lrsNbSrmD8Ty8z1Vv8XX5T6A+l6douKM8NXNp/CDmUHZzNOtDLb
iOrKztQ+zA42YmKf/DVm8J0us4zQ0X6MLNYiLrDANmFECx61+enJWXW4dwu5ARMd
it036wO5J8itx7PGaS8s9p2PJACFuKXlGCcZ8N4JLovM7Y0eOak1mMkH6nVE+gZF
GRskfkV/zTQgFC+mMx37uF8aP6uY5lzyf10SFH6WyuQj5RRwghA7XqFzlNOUWbb0
7CDT1Sr0q0KlwYfppBC2Tl8fbbFOdpurQqmrIJMRN5yL6LsCQR3iSnrQ05/1+FJ/
SP+MLN9TK1+aOmdNzb42ktETB8/zo6RyASCyqmv3eQ0wlMORKf18SxZdRWtS98kR
05CLUgTu1OOt5Eqi+Hn1t/u4iHIKQubclpPG8Tg/v7GilKa+Qo2XL45wK4QZzNTc
j6pI1hPtmDNDE4civlTF/x4+mWyR2+Qt5z1ca0u4MsnX/M6kRva69ZFHyiVl20Np
Qj2gvVI9KxR/0DDpD138n2q+4KI50AT5WsI764NAJyysneyqAXAoj4DLq2PBzRl1
Cm3KTFR7Y5Y6p04SIwOHCFBd/lABiZJmtWseQp61Jy6J+3uN2Dwu9QAmam+i1oga
sCWB+BD1ud2+vvEn4SOQfTyMd7bjWpvcEoyUusUkB/qwBhr5N0L7RAz4/9Uzq/Hi
F3R4nj8JIbXv5mt8SDGMGzOkut6aiK+O5QvWp+3dMHWUwL+u8Q2wNksiCxDtkMnQ
CRVYASRbLM85MyS8TJPy5hNQVy3cg4P8qBQLJHl/RjPHjdbbU+8T1J1cbAMpcLur
hZy5Z+oHxqfHbQnfLp3fB3lCVtnIWBQSFmzfzpUjlgy1J4myvEGSJi/YQwarpPxq
pzh8tJMNWXof5DksLRsLjrEItW8cCkF9VTDfRQzKowqCQPffZG8D4JngqUBN+2f3
5WhhxLRPByMohUsVGOicJ6ZxT0HAeUYOZJbbqSqzeZWbB0ZCvqEfa1fnziR219sa
ovnby3QlfTQwTDbDLdNkajYiB6chelmtxNkL/08yfNH4ZNPQOX4LvA3k0i5gXhyn
YllKA10LfkESq5JhP/bfCCR9+YikwIhjZeJWpO4ajAJFLADZTV8/TpKaXZqT8gAR
jnlP0Wplv5oSZyyka9ZI+AEj3kLVrzM/w7guUoPWi218t9irDUZGfzN1il6F8MgX
CJnyBuQpmqB+VcVMCIZ2/aQVo6BWwFF4YkfJzNJwF5C5sFdRneu/jykkPQpF+db/
+loY7N9fzYdH7DRy7F6X5xCajrgRvP5XpuxJYJ+FcgF9VWy27ByfapoUx6zxgn0n
MhmLBIgKNTZUeh/X2OFsETwHry2cMcagiZoXrYYT6o/QkvJzwfA4PswFZYR7C3na
GsONV/s4Pjq0dO6XQnHJvMksC7lY4ys7iQADe8apUOBLlHNIuoZ1fP7Jin/Q05R1
x4D87pdjlOKQJZ1bw/gCPj0hJPnvnnd8hILO4lnozA01uXooy7S6PlgFbAQRe1HM
xB2UKsNW7BY0sdG/lvJvmslju1UGzA9bqMjVez2rRZtG0cxM58Dux33ssYzGgxDN
diokUvT4P9u7VAAbDUHXAIY7Pmo6xF9rjwDzdvIGN7U1pBY3JkrIW6ByIUji5yP+
kxIEx6JO5wF9oanLGUJSyxi+br1m05QgQKT97SgHUJwWdYDdaV3OUQU4aLk+zUFj
NorXaF1RwPfP0gQd1VwzO8k2/k7E6iYtAD1hPKyeMcfx810z0snPBBa5lNkkAZeu
/I/YuHJRESOUvCdL5RnTduyE5BpY2xoIHjp6h6H2tNfHFNUD9ETvgyhs++idila5
EmsTyInaO7/61WQut6ir3cSDympsLg4F/EpNLSmxVBLRaDV3oksL6q+XcC3IJBob
GyY7qzq67ftZ25vzAC7MNkDgnVouATsNsWlvn+DRTXfR6s4aVTecJ9W8RJxgRg4t
L6mSh4HbhU6LOXYdMZsrqSm0vQ1lanAhv5de2k7G7CqRRJQcIf2tDkFXGLhxdcG6
sqo0fnojKRaewUxNzsw/XIa9VJ54W8frKtUQ0J0ikrSiraOlOMVIMCVswKQwjZMq
CFUNPs3PryErNleUfRzLlzcx8MxeU66Jpzp/PJRmDZAJ1qzEDzPm37lgOoARNjyw
GrC+s6HDCaQKUv+qdHYuqO2rCKTLWpXayfD1M9INuEI9aWEXKjgfC/XpSAD2M6+q
S/QcJlYz8v/u8VcrE5tEIIKuZjsM5PLGbFirMznKSAijY/n8YPcZt5pDqqsScR1O
br7dHv6qhhJeM/IurLYdORhoACUyNDLPa/qcAxfZhA2lO3hoFrN/tMemPhjPtjqz
ddfVlqcLKP1pdbo+PE/m44oIo2LYvKQz71Z3pAe1Tk6lhZqzOr4+lloBFSf4POmQ
LckJ1fhqTtd91OMu6y5+9itv6TL7ny2MjtaABpaOZPMlPWdY6uOiN27pSZPs/6NP
RkbxA2BzEywDkAfAuW6gV9pjDYSkkwqz3SdfgBs4DZONBLuMDo/p0oP03l1Z8QoE
7uX5mds6aBli3lAjEuGF7Cqz/5Ob0RMp1yh2/KWwuJebVVVv+y812iHBx88jUBA2
Hw+RI9srCbOSvqXeNbAf3wO08gptDY1LVuVpDjdm2UtXF3bVFGk7J2dadST70tFB
vfYQglY2GZuS6SicgOm2suIvfIxquxQX+c+iwEpIueMYFl/5/RCeC4AKPesT9VBR
Iors7mk+vVLN979cXwVflf5+eqTUwdr4sDuzbEhOCr06UyRTohA8KK5M3sWV9MW5
DlYGVgNU3l01DT0GUFhQ0/9mo3Z1SxAAonaDg1bjtdP22+E8nXybTCGtFm0nc/iM
9lff22oDLCJIr7MtU64ddHo4Cb7E1tgG5Ls4qLvLiKy8/QLrms1PMQsP/10AWO+C
aYSJO3Z7un2uPsYk+lVDNV5XlyPrxZse4GwhrQ6zTT1UrXxtDwCZ0sMFCbA0zobM
6dMGrTAOHVu4tdrmRJ441Y8q7Gl9QL80wwq0AhAE/VWj4dBtjyqwYRDZ4fGQgRiN
O5g6Zt6+9BCVfUWPH25s0U9ZOaNLbbjd1dwp8NjjIEDLkU6iwpb6dEQm519Ro/Us
ObdN0dwMVVy0/FjO0zK0rYlZh+QzZOw3coWoLaYKIwOf8qYN0Ncau0rBqM7ER7Jf
LipMC0jP6tEmefMFmLy7Wv1dBIGmvcRnZmzTNP4feXTvNRnNjr5V3mAqg8NVLewL
tk21JEmgcW8cSmGv/ZQhiCID3G/0BRnUUL0LZ0BK7grA65/eUpUatvM1DWThTGEB
b25zrVvqpi517+iYyFrdSBs2rnBonru49HJeVlwl6tJ99sN5K/O+I0HMmWm3+Zil
6vfqhMjfuQIkQk6AcERvHxrrpjb6Oshv4Oe3PUm8/tjEFFZMIDrCVDlEpwc7m3GH
azXM7aaPDXbfezwV3h/3wIWn70aWRc1E3azGTkzUYkrMAaFEFv2LnQ0iq+DN7rAR
MRrJS8NPQQZ5wXQAG5gvbPxQEGOih0G1NAS+6FcFXsCazL2qOTF6A/Y3LEhHyASP
aHo9Gy1pU1/t/1w/0+0xvHXvgaDPE2iY8nRfoIgPol/QpOma8ACm3bimIJ4T8pHr
bpRFPcTmiEZGkuRGnQmnUrn5Z3t8PEpwsLpCgd9TP3IT3+JmMVu3Yu8Rdg8YX3vB
nS2RwbfaSugFg+cEGu5ALFg8z8bp01CCFpzRrUyuDD+JTfzqPzNUnqnWYXRAUdnS
uKGPUQZ9+4LbD60NU1cukPqNYYbg/mtXESa4Lv+gxG5vHwYSzxhnVFdpaBelyGeG
wAu1NgSLGDZW/kC2zZblfHqXIslNnbDJxenR4rPKuLHF82iA1zH6xpja4EIW2e1I
9apzIv+0iC6H59Udr+MqO6JAtCDDiAxHOwxNkW30DIo4sBaP8csb+VhydGQ7yvZH
5szNC+/85NsVldo95eJuebSvOGsWzjgASk3dxxqTPsgX9qE2BsSgkv8/xcBqSeeA
BKa5AiKyKDbhE2JLG2ADUO6an7vdnih+px38S8LkI2ji145Q69FRZdZYyn6GIHgS
Pg5SsTdYpz4hxNGL0gKUxovLBx8BtixA5IiL2Jd0tqViwVBZVJMEiU2Xu7lpTFVZ
/Xk7zcjpC/5XPg1psVDprNo/j0gUDVn4VO9cqEUMqX+crN1XPR2/Pjf7HvcNom4X
aDjSvjp2IR2kk9b/itbtZCFTJE+C6g5a+4z5caM7R7N2GQsxdn0ZuEO6xJFs8dLs
rmzZX5brt89Q5IzqgO6Gl5i+fOOpeyIuYnFJDgeknWbTcigaJrWvWI6jDwtMx0bM
XwRaAelKOB3imV5sbK0bXUll3eO2FAh6qgfen2x3MesRqRyCjFptSTfGOmlTD1Cc
TlfWJU0tzm84RkrOLtnuP7Mfk3P0KkcGZpOwFiP9NEYwB6s+vbJXIuqb7yZlLcte
5BXLSL9RPpC/6sEsi/oXps/WNDY6As9zuaD3vXRS7ObU0U6s3f1lDylNdKvMopVx
LZt5rmoazuNRHR1/kJTQjWEL+Ul0CRgqdOlfyNlexvOqUHykAcQwWxrhyqxALlkR
2H6OyWJ0Y1iV5o4BPR7HUNzzuWqbsMCbRv/yGubyBp8PeTNOCnBnhlgIkag2al4O
0S5d54gUHYrKjiZauz3vrC+OHDQTRmoKfFZd9qp9+aJQosVy8UknobWutFyDK6Bm
rE8y5Of4ThOgCCMR5LNR2BWO8tjnXZqA6+DIB6LxUT8C6JBJSp44I7tx8Q1DycZT
+/av+m0cMhQq7jYGOX95DL72KTfIQmaRO5BmoYMOMvHirPfGsdNQ54xcjaaXkZzP
N5TayTlHE7BwF+23Qd7EoUmdxMBG+ebRpHmL5GNZf7PA7hHPpUM0/1nsAj03UrOD
+58yKveXMebbhHIQyqTbz/tdFZ2ecyrI1pATVsfhqReSNIpJcFPfSVc1CgnlDCit
SdR/AvKwZnwSafs/w0obh9yZ2wdaWj66MEjUm0VcpDfUOhmvoi86WvLcXR5hUb0R
zvGdv6TGttRstnAsUpH0JXJvhUyyA9s1RJTuNaanSWp1c7cuq1Q4Z/EkMAUYUgr+
j9Yqz7/iTxAnicQpqVhInZepV5Pu0KukvsfrnMHchE6nFsxH01/rLP6xlo9vDcV+
222midIaeFfwNaV6cV+Sf1EpKPtn8J/oJKTLjcbooA5D+nVW10qoY/egr+YBsPCY
qdmD2IwRshM/PLCq+oX4DjgUTy0HTXqiakOFcxxp8wC8hLmXnwEMXU1UbRKzLOv0
JlfOxjkUBF49OYNjy5pbpGxDo04U4pejCAigcZGXI320Ut1CPpHhj0xXHNEA12In
A3LKdw5vKJAFPsnClC027CQr3Zn5lI33C7rCTSGi3NfxIRHKm8pMpXCf5L+LXoIu
6qjOHibYAyKwNAvcbZWmFw49yHajtulQUJEQGlyfTW5CzrN/vrBC9o85Wrule+lc
okhm+5m2zYbMLlSP6Nr1SDczBe1QWTwx4qTQSz/V1cmjCFATrphLbp7SuYGHd27a
oUUk40PMLxqRhHzw8DL/kkz7/k0zQ2aaBoKi+8Xt01QeZ4SdNECrRauxJqJxVwcY
AEgLyrBGTFYZ13QevuIi1DdJv8m/snxCktxI6yufG2eXN/7uLU5BXtYC2I1FWDpw
9c2P5xTvkKprmGh7YdTrEO0IOfsGpUON2nnS0CPc3an1KsN9KDzq+O0Q+fnrwwYA
GFVN/QtKzfA/U4cyNBIAl73Scp70Sbl+szmFxOHEPolzLfZhMKFCPRWkkyMHqfMN
1J1lTErQGFYUJDCUTLJ7cFcb9OYys5JBWP+8A7YyOKLshEbOBn9tdpvWvtiYGrh5
Ak85/1Mmg8eai1jPoE9sN6CWigG/x/7398azAGR9G3HHkWuMFUhfq02PdmQfxR/O
q80uwhDvbNtfL1fDlGZKfWVwFLuouHJR+J0GhEQkYoeaF+pAb2PCuPsJvxKVEDFk
xWToK/y4UJCoYJYtovBkCm0+DkSlz2FobmgXzme3xsieXA5Pg5hL5H1dNTL63pGL
4zhYHHVWGT3raV00d/QLcoWkyk8iV/cpopZGV0SedYqmCinslcvmh1EWBWtUMpTa
NjpFccZ3TutXVDL/jMq3+7ZoYs/oZ18bxPaT6kiUh1nDvSzMISS0N9VwDwzCFrcV
J6eaIEPEKf1S4NfcGUYwWCKqP+PLjj38Vkt7TEib393cT5rvyvnUxnvQFRSL5K+r
hdyVDlteiPpYGlmXsIbyZ6ySzZVqjQUDmDIUIu+KjE7U4BEnBVD0x5axfB0/Y83n
KicYqkMSPGr7svVuAoNqvpoPdb6PnDLJ+MlOJC075xdNKcrcSWxqPK5Nrsvq6Q5V
3iMKzJFBu0EErXiySbQlZcnZin2QEPjgouRoZFUqqK7I3d64ALm52jLS5bmtK6ED
iZap3zjt654o+6Il8K9AQKqCfJXoZUXoZ2AutpyZ7fz917UGzKmcbWfH67Z/Bm+p
wrd9/HWvnjvH22xNVfcz5jL7pRAK2gXVrMh+/9tofubOzU8kyQ+ZKb5GJpv7vq9J
/hKgdrTCCV2uqdmdVuJMaXLHX21ZqQZcPhAn1Zrv8Qn+hQTGOUV+DbThHaDPrVxR
JEMZmVbIZT6hklgaFcxnWtM6U0QgrlUdXT2Ojwpr6B01XR3f6FgMW1csNarH4DvE
yCo4z9r56QQW4NGAWHnMVolaX41XtbHhe57Xh8p87BLNTS5UxWfBl8awFB46Za06
hzwD46ib8VF3cexXlrxv//nrobJxix0lBcARnRka6BYCJPZasBl7XmLFVRRf8/kG
wiQqNw0FqJcvwmqhitJqgIpNLXBdYXuWoE2zfp0RQ8UOcEo0dh8wgpPPLEmkslmY
RXfD3la/lMb7S5YyhLsn0fZsFD4XEJV7qM3aQftlmw26TYrpFPspRwd9mjgPoZPD
Ds7reQReTMooZdbNpGlIR8IX+2eDSC2sfdwTEmiDpeJi25lWawtbcelAojY4oszG
t7i2pK5yGr7YJP6rDpV8JnuiTsjQr/XGbxT0O1CdIF8yKnxDnudv/sbdS9/P6AU9
HoUkfthTMpjjoOAKoYHGqlYyM1b535F9IO7dDgy49nYETtjDp4dew3eMfFvM1QN4
4Au1sIyHiWbzN0jkivs/Pn1sotmscO5Qpk13CfHvojQFKfb0zeOHEXCjZ5IkEz4M
46H+1hD76AGq/0udjf/NvNU6BKepjxAaBMcJr9w+/fX6E1/zamoQ+Li92e/1oul2
BlGMZloeuoDdxuqdSemJ62WEPb7C8jJswfPcUmGSTu5A7AYiJ9NGmVxISg9u8rNT
heiPEJhHFdZjH5B/z16GkszCaMkN/uGb57BlrRKXlkaZDHphlAyzrHQZbsX/rzo5
zEoyjdXjKpOFUug7FTy6s35unNGnyaZeWXPY+qeclpQw/wXDcMDerg1K75CtQBwM
z73hki5f54N0tGqCZFEBqjHHnCFAhLOPBSnw7jo7Uwe/txWyL4/VQ1kBdPp/leaN
7ZSouxh1J31cAUQWm+nEejbJdh2RBr/wi2L0LFQPTnWrN+1ZMAJU9KyDPdily/lY
H9BAmeNB0AUtL/vQ+govsSKaA6t5zCA/IuhQ7nfo5HHv7jSijPNvkC3X9EpR8r5q
66Aiw1WK/wz1iE6VMwbjViqh60YalLfzxPYUOIWiM7UKpKX089PlZGmmBafGBwWT
OOQ95CTM8/YBWr6quhs+vQ4+n3ZFc7H24kGD8jy1M4DC3/xgrpB5ZEvtSAMaxkib
W3ZoGMhFWDLWwuL2ZHgyOwALnljfb9JSDyEtHi4jjXdDv2YqvEbbDM5oNe/3mvIG
NseC6lAcE2EmichjkBSdG0qoMvLsRKVBo6wTJXndYbGnBYkGwrgbjqjWgSRHGE2Q
5A+Hl++t/3MoCoJv3n1c1aAnu9mru8Rn/sQ+tgP3BdGZhdaZybh5tKIRJIi8NpZW
uaBzj803H+j2B6kstuL1YFIJjyXhni3vvC7Fh+DURLoR1EWw4nO6mTUILNEWdTXS
T93Ca9uXWkLOR3lIXOEAeFtETz2B98qwsuyfe5R3x84o+xsgEKwRcenXIDY1+iZY
/jDoP9HSFYdgOyzFC13cJJ/LaKOjrIWxF/RfamwhhC36w246dZO0rjZ5QiW+0DWo
To43yfyAXdKf60RHFL0y71HHadwc2eqNtjH193Ua6m00tWghjty6ZqC7jV/rX689
/DndgWq5hKOKI2HVsWElHVRPWCmZDdWG/oAzdM5vSwKlWl66/ipOy//iFXXLsl+O
qAwqc7mwkuLTkjOtSkZIUPNfr04xurwpwG/sIlW/qrAhrNvyL6/8xk3zmAnyNPth
uuzM+ITzFqvUMIi8QkITdCzx5fAy3Y19HXakkn7F+jJKLBf/g4VDa3b2g0XW+4hY
dgJ4iRWk6P9VC7oGfWP4/brWtB3iJASvD6YzG3wkTBTKdsW1HzrTUxJ9ihhtohka
L3gP6d1E2aXMjsmMifCigH8fcoajqkTysZzrOfObGHJ7VUzE1BksBsDXy0uApTXm
KD3EiVbCd8O1u3pS/xRhz994EdgLh8gt8F1I5VJjE0ibNYOTU2mzsOOUCihzkT8g
elJC87KYjCBOzuahqz8yUP/zhRF85oGkD6H6kGZVrB4eSFsi9h3Yy4pkJikdDPh+
OrOlLMVg+Mqcpm+L0+/k0ad9A6xjCooTmeBEJvvCb1nHvVBuBh4unqnEhkJAsfLL
TOdhMbD/EPXoBh5WfDSlmrN1gI94JJjG+P0/rofbNl5Zp3p9fi+dcAhDje6BdUmY
BSLdwXRZxPPKg933uBWqf89miutkBxaOONEkK2hiuxvcXJYG776sNB66DIIjPi9v
ln7KiLngfobKFI+/elAr4vJKevTygjc8VhXFAZ78konNi7dmuGVUIjLUosnm/ZqF
B79KRJ7EGUgOxxOEFH8WP67KS7KxlvG/U8RKJgZ6MGg43ppDm4Xi1TCf08tamgJ6
liPW+ki2bmzYigNgiVSRYhUZDCUFPRCyUP26mViI3Xbwch5XPfePug/6NtYJTW5L
Bwd+wXu+5K/qzYa9Rhr7etAhra4ZBy5o4JAvZU1RYT1ZY3W/AF2gI7H21V7Zvn1F
z8EugNTN8Su1mwsTybXFAFkn6rtwz+ChbeX9+BnSwjPu0HpIcLbMSQHV5EhRzTzA
2dJ6iRjmTq2+l6xtdEr9UJIjaLD0VFynVU5nfryhODWfHxv8t7cU94Gc6Kb6a6Cd
YgGzD2SvIN6eL53bu9ChkqPYnvoOv3P2LihUYPvUvdGwL4pDLQYnt8EYtHeKt3Ot
E1VRfyplWlXVZSQA+1H8zIHDinkYLVFmF8zlt6U/k4dfphJIqKMmiLXipnQiKzAU
5U/kbpow5EgmCdBicSWyedGuua3WO50jbHBBoya1Dz0DJibOIbUdHFbECQoEdNni
aA9Q55D77ZkFsjLzV7y9oYYdAFNdbOwi7G8dK928k4tyjRBRUOhE7WFUM6lIL2rM
RwfeBhVAlg1gpkYkJkFNTMFzc53a0CeiGdYI68Fd4HzYVRlOch2U3Dlv7tTXtomM
6TThbTUoeLUluLBVOjn65Mu69YIe1K4DBG1FXJuFo2ibj0xb6f8lapkL9MVAP8pJ
Yg1Dqx3OOBw9ZYKTMTY4QnHQG9ddVF898DzdhIFMGdCic+WfthBtk2JiLzqIH6RL
/O9sltspPyvasWf7HOmsIOwCMGNdV0f/7OwEgtv15SfaMT1cRXcTKC2JM6JxvVYk
xEL0BbvBlP5eRgq7c+otWzccdNFuxnbliHnnU8lGfQi5jFO9BMATfUq8lWIgBdaZ
ZrGuEvAy02CeCrTBFO/wadPElc3qss+R/2+4msXrxlKsWjhH8Lh4+T754ZM8fPHO
A3RcpQwGY2Le2N7XRz1WR5CsN3PdbiWcyqKUZRAPIAoJSSlj2FweJofA8jBwUXjj
GpV30Cg3LfAzxYDcrVmYDUEU32LRiCucV+QpJQeDoph4ouvuGX3tU+APa493qvzY
go4a/Jkl12ee1zOT31Vf2kSQ5u+4ezIQZJ+8WQDEvEb7C6JvHiz0lgKaDUeH0d1N
nsWykKFtTSdZQ1iIdQTj/LayBZmPONV93Op4DaU8HQcAdLnCrLDpNuipVa+Q2KMK
2tB7gLsITCxq8Geqda69D8eeF4uo0AnewRoBw9nLjA0dVbQODtev1SjMkj055+na
scnYzReDwf12Dobc1WqBrMPCx9LzmvB3AOyu2PrNi/xOslPAat2aPH+5yLcJR0zF
P0W2q7kpTZgRZzNhp1LCT6uSrlSyGxo0ibPu2bgNM+9QjfKsY44bA1pamv/U2IpV
sEEod5JxdCcu0gNrKeSiLbn8m/GcGgLi6U/ujBtGfiwzmay1AjWeng+/trneQz0H
8qfDNZlIkSpO2/OqEvUx3Z/mzzu9yLG9sk6gl66DRzazyfC2ijnZEMLjKkZFJnch
C4Lba1oZhYfgyNYmPze7E8AXe9Q7GLXChO1Zg/fqMbRsj4LA3JdMZ7EFJNNWFk1r
rseqO/LSeFQygai/BWP6TBdg1P9N6fGIbxmjc4mHPcaanj/cRXT2ubDtFODEvISs
S5PXaUvXLtNrVAHQ/9vWgtaMWQNdIx64Zx4kHBGtQ+sSHRyAU2wJTTcuKYWH7IiL
z/66zv4IU5HI/EJRFphp542JLh7L+sSbBEx6ZflQ3ONfKFmNa1sPJyLjZ5uDscSZ
C1Ie69offmhCJciz5NXRGVAzbv7LFnZqelfk0ijxzrrT/Lyax19qPvpjPjHkoCBW
xJFz9li444FQAHScaWYQympUt8Gh+ytMVJnt9U14nmXfGxu781G4PRvCD+1aY8O/
L/hYrAHD3FrVlZmymWHY/sAqW3HN/wqzUwwnY/JY6eBo5S2p1WckNiXVxdNxKM3h
jH9AtlSKMl6rLqVEqs+aD/P9ISAhQ0PveXPsYediQSDPrMcV93hchLNXxsUlhANj
ghd1AKDxt8fcriOnMkcLK3fxPikJ9wpzYN2GO7u7qiHNpclmqQEiWzocQuOhzVAB
LApRzIjmQS6M0LuZRakpJ0WYI4GsIVQUXgPOhkOR5qEp76KkbEFkhM9NAWqC4Eug
csc4lYtG43t+f/R5x0kYi7X+KH2dyMTk/Mpi037WaY0bSyINISt6ngfEg6+HBp0M
Cp+HGv/fkEQa/gaykmqiTaSAoh1E6S+7hbAq6V+CxBFj0jTiKXberx/hK5PPjogf
yyplMUO0o0qvIKrsj5ORWPZ9Zm/vKTzQVODG75aJJ3w+YbviQoqdoqjTon6NFdVS
FoUESsxrFjx5QJWyGDvFzHREon4PBzrw4P+NTQ04MgmHlvOxOI35+lTk9tmX3vll
7tzUk+szCxxYmagVCrB0ITTBzdlkWxEGzUbVSwqo73uZE/unMd02cua81zBBgJU0
N8/hHHL1txHvzMM4cHoim7oomgBBeY/1KMuNYEzmkaAzg65//foWxaxIhvhdZtTK
Ur4K+0swowCn9Hygb+MxgiHK5+EKn+NJDJYktlymWQwNkVOY6jgRJSVxs1glan6W
qI+XIlxVLbXsDUNmIEPLpaYBpNwqWwfTqtZIytUeNRxcJWGHUW4wd9ULMSAOo4rL
TlzzGaTZwiaPmX9rzZAscb7FrndzsBLUn5Gl9YS4UYT0rm9CNC9hpOoNwC4KDIAC
DdLiHjInai+fOYxztK2LguyvTnUy/iKk4ub29P3CMKZOUMP56cfedHchW98fCa4Q
agW8l21SOPBQOHM0N2nRA3DFuKq+KtrzICsHTO51exe/VirIYIXqG1eXcnReZ+EU
AqK3UZYnMfdhU1lD08fSf0V3GsAfqH0/vv+kVk6Z4Q7/PU5oXmZqLKbhZoOTuCws
QTu+jwcS+81xyjJNzMhMinbvKaUrF0zfBj6gmwHkzVqDiCRwud5D8Fu9EMQN+tpF
VKsuB+jXlZwO0aPWTvY/lWhinJNE+MWHWgce+ptomQ56N26BpfK2HKIm7ixCWGza
MOcTv1Z2wUl76ha2cxW11USsN3TUACXyPnRRy5zxbNgVgUmWDvAJKx5tt9S4gIoL
jAkyc6J8k0K4233pmACRKVvDhE3nfhpDrpNJRBI31Jp2Idd5o9kpG4gl9SzSrU7H
hyzEnx/I3vF3vSg3xUZXcy8Z0mBVjFFmfRLJvwl+Z91XPOo3MRuXp7TAAKr9UzQJ
rsU97kK4eE/EViTUwxrPn62+/iIhxERvNi/rCtXi1NtvORH4Pye/gJ8JzcxyZrRy
wVvFoyc0RigLysORWpydY95IUwFHdqWKPtkh9Ek94T7QICvtGA33+j4lcAOv+qtx
mHbmN47JsCzi2rb7m1ht0eJAGTzzmoqlyPWqRva+/zClLQnSoLsWXORKu9WFXXWM
p/qECIhBPNONOcJ6rov2nJtFq5dF0YGrGyOG/QiU92sDRFqouOQLw83M5GzrkLDo
J1FaLEWA/Padf//3UwponDwi6fsXrkch+K+Kh9CvGACwtyVWODujX0A8hJC0b/P4
OV4ag7ECw2Mwb85O9Q++mgh3uMym71YZsdVDPeZdzPzkQ6jomgqgNs27JwOp8xCs
x/5CSMjweIFYqIApIP3aM+TD+Xw7Tuc/+eoi47ELLIBINhlbAT6S1qV8pB9TVenC
fTKExojSnaUkYdmiU8xXWFyuzt5Cri6VpsoC2TthyS31RR3QeWDO13nXOQ5RFvLj
uTZVEN2ClJGZ9aOY4BxvFv6qmpHvtSmTaUQDi9tsSbWc250zWmxyWMEJi3VlDjaH
I7fQQwfn9RvlLHspz4Xk5/Bgf8FrkN0wlk7kjAsjQDzJ6nQvVRjwp6EaOYf5YIRB
SprzzegyVZQJniKURdIHpTuvPHlEAWK8Fdj0Af5MIs4CB7YmETnxWrviX2yVe7eX
H3EDNk460V9O0bgr1SROz34e35FfiJpTee+B7kfFJLThR4TJv6htn9tTrDqC7pmf
3Ujq42Xc2zB2uXvWm+9wfFgqHKApTduH5A0HJgdCcD3EDme4gA+fyAZpccgQjmXW
xsQP5m3gb1M8rtj6Xbg6YUvTZ1EcekI5aH/521gCYi+4l0yED4G2m9A521nM+WQJ
Kw2WKLyqrYDwl42H4+uGGlp40BRhhNER/wHNuAja5mW4R7foiyEMngLt7DeQLcQC
vPIpSpqyeWLS3BYCJY0A6ixeGYEB/Gn/uD/6mcabnjdkRn0Q5nEV08cHz5zPGcf2
/lhbkl4HYiIJtc/WdZQyyc6nVTyOswRfTGKrn+1OoxkH+TWk/AYFToD4qLwmXmkj
r0Ex9aWVWpiejCzbxX5Srxyl9f8HS5sgeFNn/6K/bvluu899jyk+atHF8pYZBsTl
l4eCDYHszeOGCzyIv+TzUnaYMdbHpwbTWKC3qTbi9o7dyF4YKVPtprq4rVhgKFSe
Uu7b4PZeBy8NsW2HktiK+j5VZdRwEYi0+U5oAwMFUx9nJQLsrK+KZYmvNoneZaKu
V6F5xqXgsaJu/QLIa+mlP+C4cx6y0DEN+C7nvA/fCqaHNjTfqSn0jcpyF8TnFVoY
SSwVn45Cvas5CIbzaDI3Jw81CGdSM7iIwoEmH1Z0f01lWsmOOnfakg9XepwjiFQm
4Q1TPDWTw+SyW6Z8Qgd/24KAQp04QXNFP9Z1wBxzp6orIIiilt6GK/g3r2YweTuL
2gP2blPCUFdurOGtTvgux1MSZ5bTYf58QKw+Edc6971oF/2ExUvmiGctFeATe33o
j90/JrdFDfHoP8z1nzAynLMPCCVqpFPVhxFFmBV5dZtMEj2EEXP9r/UYOKfiC5XM
66wOShksHzCch8TY20ZG7KPvpgM4NTeSgslldrDyhkhQByW45kTJM7cCy8Gln9kw
RDPz6lLUBz6jJa7ELsLX6fJW0uAhleyZYkST/LpfLDsBInmZRrXfVoGan0b1zTN2
IWfYH87YB7tv1euFnO2SLhUcw+FdBJNz+X+LPMhnRxK4Fyt4vKYB6r8v5CXBKm6u
nY9d/fRjP0ltw9TiSkIywHKhWbAX5kWfdS7gAC+IjWHex6fcOmXmjmyZB1f0pSXi
BG4M81Eq9WdPttRtXtHTPGz6RFp4zOT+yNEwy6g+i+MXrVDP741SYP0SKCk+e8+E
ihQblvr8cr3od0rLkqH1ozpVl+DY00EtmRsdJAvvH+AnX3w/hiDeOxnk+KLpJLD8
Piq49e5+Q89telqUI1n40gPIbl65RrOZQkSbfH5GyDwn9Yi503WqQMv9blXnar+g
9+lB/lE+gxY/bxfY1Jhqa07wNX5Ny6JxlLq4mLmlaowbaqUw5F3BZmUu11uoVbJs
IRXwe3tG7JMOXyeSrLqkrJcdCda+VSGCm50qtHkZC/4XrGNJOUbpTk3ksevMNNxy
rGDDL6tJSw8ExnZKvCcMKkR4EBoXKd1S683tHFhHgduvCwV0w8yEQrT+aHVfvNa5
g3lByfe48E2uKkuGU7pUppzacYg5DztJjtjQEYOF64sCZf/2UaoJSde0SpcFTK3k
wxkokoKpiLSHTAd0/bJ/Ydv6KkiETFjXhEg2izmiHcBmbVHnlOYJOq2agWKtuI4c
PtuvRaN4IU9vNaey+eOYsVWVUH3bGKDwEM/iVCgj8iop1ZilISOX4CqL5CW95q38
kLq4jfd/78W9AUDYsnY9c2LH/vI2VJvYUDGVclz7PW9P53Lj/mj89np0a93vQqaF
3U5vatcMwdpGZ9HAxf7O7DBCud78i9tuWsCAaGwB3mlX9IQP/JAx9ayatFS6iIS+
Bcii+mG5o6M9C1urIJjWtyqA0XdA510rRgK5h3HpYoG9WKnwDV6ePFsKflKR9ue5
xprPW4oAriDjVfp9pZ9Iwqo1yu2lPEtZmneuQKjgscz8dxTev/kP1N04kwaeXmMy
+FPxJ3IXE2k4Grpl4RqKauwzHezTVM2vSIz3CDbyFa0UBauPulVYg8UKBgf8TpOK
M+kJzV8DldUVRUfYeUnWarbUk7yg+WUzCgks0pCzcu2YNicYsYnt+jUPmyrjAukO
w+hygPVCOpfosrTIOfh5PM/86SG6lPfyJGGsVrWn8OAF6RYDWrFu1lwqGXUPA/oF
GFoqclCHO68sWZhWO8DYvkzmOR9Y5AEv+5HPEDTLa6keDwQD1VygnwT2BF11Aghu
H6GPa61xWUFVBZluFTSw3oBURrDm38FkKOZWQB+cwX2lAJYcEWfjOYYvugkecefP
v6pwXDABhjfX17XE8/JCZrDSduHAS7Ad601W/drdB8RrPuPudpetKabbJXg1zWLz
/7hQ7GWyZf8CHRR428qgOre9eu5FGuwpSe2bAicAz2S+UnpVU0pEoriekhoFR+rB
IZMcodLsmfktsnkbjcenORmyO9WRbJU02DYOpePCGfZrZKUWZzFFH6R3ibM/2OKZ
6p25TZag8kbuHkRc8nC7jemLvCI5Wz3BHHPB9Ray+6zaDCUOK3Bn30WDYw2bjFXP
Rsr+0cslI4hNvIzSzGs6b1pVKdGJpUuWLBZXXAIuercinqKzUnqkA4mAcW8qmT/2
Ln8Gzwgzu/x8E/GOtlPOV6Pq9Fw6JsGF8sa6JBH6K6K/ftFYrzVX7yA3GzzaWbp0
3NSj4MR0nNRfUjaAABbQSiAdbAku4eyYEceN83/0GvyFWZvdNq9ea8MABVn3O2im
AHC73wB59b5rPCSLlLrnfz+N6CsIEJina+PqkbBhdBTh17fbO0ZMqtdUPDbt//3p
xYhTi2aP3XR8QjRm4MUKmBKrqvTaZUX15h0hC+Rv7Bqx0uT/FNyYcp+iGlE0UFuc
XlA+hOig2HMcYtMLKaInwCPGKhqvvHDd8RR2wfl6bd9OiRHSKXw4Kp+NjsjdZwEC
sRiPoqN8szTUxl/bIz2D8H2evdoEX/20AHb44sBVp6dV7sDeM0/0+X5EfINMe750
AbfVPpEkJu+Al6O3Vx3MJIa3vN1Q5UP0XB6GtY3d9+WXO72CqtI/XfMD7ptsA4HQ
CxwnbmvwfduehvbFYgiPHY/x8ukM76bYN+RIJAdAzTkx1avpnL98DcvFdtcv9lXg
57kw8lWQNdT0XG92DcXhcQPg0xcuG4eiqRNnVBC2UTmApaRy5yJWjTqN62iQbno5
m8v8Q4JDBjJ9Aakvwuwti2lK6hIvusucfEX+ZnMmPsp2vqvyJipvKd+RDmuSYvil
MIESZV0u6jwscUF4BUYE8IFwX1UDgDPO1ngDaFqEiTb59Ju5LV/hvpi8fFnV0lxA
gVFkr1b4QNuCx2teb5enOtGL53D4mGw8SsDvd9HXqp6K9bmfUICiarNfVUtYCC/U
ARWZ+v6p2sO7sC1OFBVq3VmIc0SF80gyeJ+mhltL5mzKEiML51TpK19tkQzzBEUa
uIX3ZDOJv70gJf1wdTTFV28yt0nM7kK75/OfygcTQgkBzUXGMZAudk/vO/r75yaN
BMYhtoMnn5udzBZ2NwiD75/3k2tn16u8vNBQI/97ueZA+ZKKbfYnX+vRFWhoDiKs
WzeylcOQBWwGuuiRVRbsM62W4DV1rN28N1iMwLzgK+jhiRC8b2RuBF7ZPmg2bG+t
39/EyETr6xjEeC4xZUKgmOSe79FJnt85XYuLKTgebeMgnewD/JCKEPZw3XN9RuU8
iA2Bp7aXEgJJzog0s7YiAD9OxbBb9/blxfhOGA+lJCl/TNU3yI72ngeprftMuQjN
uBTzyD7fYlrA5oeYE2/eB8Rl7PJe7SfDU8yj8FXR8C67S3jx1VgoHP4xuEkC5tQh
smEHQIF20hHOW6Y2D7KotHsWNogtcZoi8i9BK+GjBhXKsrfcMPlN9Q5FXBkAdG3U
2V6qTJnL7YPwuy/jM+72/iBVTfuUTHGW3OVzQTGKreVBfBw5wUGN3nocCyYs7c3d
Fglfy8v+z88TTCx0RbzabHN5MxekexvBuzv+Pa/zEPyOsVI9Xqjj7IQ1kCej7Pt0
uyNauzzkp3gs9ao35ep0TsEqhYqjnLeXKGI9fB6LB1rM0KZra/M5Hh3JtigZpX8Z
SsdZm3L/LcPNAm7Q6sj+MFcGVZ3adyyEirVnTutQyoSA8ZlR5Pch3J00+2PKw36s
i5Mcc7tSFM8xrLn9RxaL/upW//7Y6i3KIQYGlWgHomYMFwbubVnu8k/vvA1t7qDe
UIALbK/4rfll58hcYRxoeH0/YurPL54GaVXK9NpJSdeH1mrDWY/g+0Em6kPefGUH
DLNb4spHE1BgPUo2F+OtYJvhnKb+GqtbLZ35y5RoI7LQGaNfd5IpH6M+YUSrOVh7
ohHU6IBGjgqnZxa+FOALu+TfscyKNVqhs/Jn33j5zZtxg+B2g+mfjLs89m/JhnRZ
Kg+D8JJaWgRbWkJPm3qmpPVgB/A3nRdLy7k8xXD4oGGWynYGnFXu//GHeX9Z5GhB
LOJjKFMoBqGijaj26gxwMvc0FgNbcThKnQjgwrWrvVsAp9yCu4X4JcgXh2JYkWjM
URpComcDAxjgwZNAcs4hJrZl9TFGEZffa+mbNqLzyYPOQkXNr3t3LCTj1scEsBsB
ytEa19xDkhcyRIti0BnxW6i68EdLFHQsBa3A2Nlp2TrcVY6fPGiAs/P4m/7sWmgD
R4tPdRF2xpF0r5ReB73sr04AkTwnk4siHdfnF2JaBvPnCPiC5lwChMpz+sUnp14v
/SfyRczH8OoAP9n2qxXCmoeEAd2WR8HGCVoUnMG7audk4aJ+O4QsxBx7RIUrBXIm
q5mlrGvNYKmbkkR2BXUeQVpO4rAgGEDvtVkZeWM2gIWh2jh9Imbsz39FkXa1lKV4
EH+qJmHG4lKRb7rZm+DS7HQLdBu4ffxYcnPeE6UoDPnGaLBoC9O9SYOKuF3R02U+
HeFCt54KflzZsfIpL4urIGvq+ZRbwXBi6vDksx15R1HjSJlfeK1Q+9KZb5A+O95W
qnMgsq2B06F+jpGqoErcspU8nUb+KsTsY9xjz20ajc+70+veqwQrXGlt3mgcmK4X
na51xkT1njONL1SZ/2zf37Q024zvOCZeXq6WJyIHsD+ZkUFgg+kWYcX2K2CIXDlR
E6I1o5bbDxM94Z2Ibt8wjg5xA9Jyft11qxxVZPKVOhD5Im/3KPyvsBYbtc16xkte
HYFxM06ZxoqoA+zCXIlOuBrKfXGtC2jieoKpv86ec8LGn2cEdb7kzsGMeemeoNQE
I3dWYXYalZh2l24gvWvNlSG56BZH6Kqk08UnaySWvldP3nDrAevTuB98mzckoFd7
DA6ojeCwIyDyvcajPkYoVkGkGjymvm4ZP/wuYg1ocPCylu6FttGfzOEzoXCRyl7b
cBgtSMnZd5k+Kl7w03+ALW2RpRMDBofYVaCcw3nUlcbOF2HT8FajJD0Rkp3rijLD
cbbj3lCnMSPUgzNCM1BKx6VjhgKKtMYN8G0oxtkFrr2s0+LX5EJjQYIRHOYibPU8
gfNAWNzk+wwa9Xl4NZlinZX0igiutLFJ0pV8orA6J3F2Gbd4QVpU/pftDrswCtc0
wf55bfPvj2qQbQRlM2PENFnJcdbfiJskz53ALPeVugHLVNHIV/iwQEmvJIeds2jB
3FYhqjzamh2gNUu/nS6aRNfXaZmDDXW1Mx2XxEyE6mgQLCYwgeQOG82uC34e7roY
KmhHd5Tmm9v424B0zmb4IWSTWVDqMS6zDaDvrvYGl321smvOpSalYncIEayhKfK7
9Xr7/At8nYHnkvU/ikG8joJDkwWJq46K4s9TWWSnYDtOIntE843l2vg71oOMmnUJ
NBSxILFQn4LuywKGRfk03AwSOHhnN2zkXkjyxmuLqeYwj2t7JR2Yw8VaaD+BejSW
+fEmOjxyXl6Qq7T1OOV4nenKqQ+0DjMTPXEOzD1nZUcVPAmTZIghCvDUXVCwUhEY
orFF1GS3rsc2iifJlqfAmYEe8HyX14XK/hfz0HFDQLG3RXdjiHtiQGzSMFC3G5nO
tUM0X6y6fCmYvF7r5DERFd0NdS2FkUxFDU31I/eBIblZYwdeVEHEz88iyUDcoh+j
lMuE8nqjz6orjay4tWyZbCFhYgqeCDQW2jBUUOyZTP0mPIjRU5nP31lzkL9Y2GT2
FQ8LjfnVgzZzxSG172SouJ+HkV/2EM0sQgklxdW8L2RHdeJaOUpXaCGc1il+lB71
z9bv/iikJtep4mf0GNdIdvqyJv4uav8YrfQc87o5Jy/yU1LtnbixlwxXgX+dh0+b
Ey6uPu9CWn2MpEXqXjzqv0xh7cXG+LXO82nhBBvRh1WcNU2rzWStFaM++s9V3aTE
yg4y77b5DNJYBZhCQI5uqPIrPr7M+epNh357XokOv529+pYdYOxs4ZteePgHSH0j
VruI/ruMcTZUmPtyZ+Y6bEJogEoilC4Ti7g1XIc8oJotFlwnRm9LXpaNbvXLsKkR
DeOu4p+92ydVyPWaRXQSPdTtZYDX3qU6FysnUuDVhgCk8IiIfAT7UgSZJEe/3sS+
dnHI1scmLbqy7ZY2rQU3QD+gTVs6wXe4cYbzrpimsYBEANJYpPjyIZdmiCWQEJ91
CNsCkvg53jT/JfLt7grHdjqOZLXFLi5Hhq31YRllsJ5k3aaYAzG6ss1zuQfIM1mC
CkzSx+27DELPKwM/AFAy0pRTe5ixW5/3OklAsG+h4u0izBNf46qTI/O33ZfSWdoO
uJpOaiqnAeMorhZ9VVJXMUzJM3RsS4fxDzkY/NCKb0LzfvfA28LTvkV6odj4trCK
dx6HyDdKw7YpnPW/rGqOA7Kvm0ab6O8De+heICgNRNrG7eMfnMyg39Mvmp+sfui9
OPsObMAiEeKJHU/PxCzSjs3PKS4HQ4gt566yD4CGOP/FNmaJtmCECTGXyrJXMdcz
LvtyLB2OdXUuYaWN3kAp5svjz6hcJGfcmcM+1QibTvsb6tuhuTOK8S5LY4y1Hf3v
cOUEDr5rLF96XECXiju8SEGskzzMlevO77muhcC/PlWNVUIKC+tGfbt1tZFoe9Fn
S2scYVMyOIKBG8bDhsv5g8on7YLf8kKbd6hH4C75q0YJtTUkvPXzzpWJGMDpNLJ5
e6YyrOmiMJvb1fbHLZPqoJ1+QHezjEXpRRngkytpLC5DaVpItG2rrkpyCTl4nDM7
0RzhNLkYD3C30MmqQOBGvDYe6HwSMFG1YUfWZMluQ8FbyOqftP2gGVkSxBkDftoL
w+pPWTdy6ASwEfNy+1+kPUZx7j6V0QchybqnbwQSZgAGeLqljL17Y3QkOMtCynad
EB+pRUCq62WLOUzuG/O6icCu/uTmjKM4E4j2tPm/AjW1jx25JEX0vab2lGdIowFh
Cqd7LZj5oZe9DGrq3mJrVmcfxNQuWk70XkS60bz0Jtpq78O2I/X0ncljARJiMfs2
5KsQNhiqaID+T1R4zvxhR9G0TMfuS9jOt12MgRqyNFUsKQh0S+kjzqnt5azpKQz7
j8liB+lhpkvX4qX16jUP/Zghi1lvzDyNjsQAie2c4HMLoR4XmeKH8QB7mGCKez0z
2XoDJEBk68DolNpITsvxHZRXAf9BQ7FwoqTd+lnJjmusIBXi2JwMG9AGbdM0HsSO
Iqyo+poIXMlNtAUOhZfjdbEGqE80CWcOcvcUmaugLLeXqVX5CJC7M772DBY/3A0S
8W76IHywXYMf2Kkrfyi7IztxsvEHukSMhVSnuOlAZDbMecy8Gamif5r+CPFaOOXN
AjbAMJ/YBxkBk1dqYTczQ8viSa7U3Bo9Lrct/m+aMdcucK0ukK8AkESATHvDxooE
GKoB79NDPuLVaUi1hB6J2umw2MJSAU99vWiJaunL55DjrMk73JrTBRv0lsfGIm/j
szElClsfs8DcsII4quCZlMgbuAMiuC/8CAtLXUPN8SrlJRGLQjlePWy+odnQZoEC
4Y288HH8LWRVRyrtaRtdlKhF4C+nqUlRec8WTa7lMONO8iHE+JlcgxYkBl2KtVWZ
1kVjbzRiYjc6eExFYNxMLZDiEUqYQLv4FK1nSnV3jMiTZUH5+vRhqYrd8hlxGHdp
7hz4g5pvtPBbL6y1xxKeRQgzfaLs49tGEA1pJ26QfcnqaABZwJgKWuG4zBGq821m
NXwzXrBFqbl1SoyvV6RnQe4xptktYdYeAob4ohfZZVBARNgwBfO6MWpWRJJ1xPGe
IK1hZNEpLaYrK2yQByToZscNNmYmz6meB1ShEOfoKXLKFM+g3NM6UsqefQMLdpt7
D9fqxp0NN3xVqcDIzFw4ZpydJlsGiwZdVAUKaVbKCvl7MV7CC9gtz7M97j106E/Q
/TWfZ5uRKM0uuIinAsGg84PSmbfXlHYlh7AEA2hp9sbTxycH5Mo167w+u0N8qB+e
/RAA4OzbuYQR0l8ve1xqJRfA1lJDVBuMtlkw1l/lU4s+46YtNm+BTChTJABBpnOe
qvGNbO8B96dyiVRUUoPzNwckNXc11i+KX3tvHkpWeaGTjXvUXlWzAclGUpZz3C0t
FlmcXRKNk3xv4e9Qb0sNM+RjTZ0G7rFr9TPOw98iM2XnHjYSY+tBV+amx+8gONYm
Yk+GcsCImMSuL9+G+5QokliuPw4CBA44ajhrOX++VKa/2TEaUoxeagCkdeUcMChq
m5AIzk02wUI2GME4AqqFODgLq2GisPXI1+V8HeDpklTJrmcBJHNHQgs/Nr0kCe2I
NgXJXbxXdNAZGzQtLtT0e7XXsrCCzhVziqmSz3gUu0gru0MyxUuqApC3Yy5oJGTo
uOa01IZ/lfeBtGCH1yjysdzJWm12nKsmFRjFjfjJvOeVFuRRvoP8qc7GQi5yrLhk
U30XcDg9RkXRBLu4uWBlA0Tu5DkqOgQYMUex3dJl708wkKV2ruJEMcFzumCDse1S
02r++gISMobRC4s5XwQ//zxEoQC/E7ILmI1X8VrWXbgs+noQ9sFJsKtycrOP0os5
Q/nPL/eoVWF2UggME9kZYAHBd1MFSD2OmbOnx6/kouohfeO5UOnoiu2jQGrcVszD
F3665k797wn8PnPNIhIZY+M7Qb2grg3r36BnB0FrJ5sAAQBZ30WYYZvV9yFTDrIQ
S9CSviGms6fOBq9EdqkE3XM0Rvx6DnuptrocuB0pf2uC3m6uWyPU7s2Am44qZKjU
Zja+XMp5qPvPYgnfyYIa8FGylw3QMJHz7je0vl9Y6WSEXXvVm6CXYcvKmfcoNJJs
WfsKuQP07FZOWyGn9m5FUolp18AyZLQYhVlLF2Ij0tz81xEvKxjJ7ONo8GGn0XVh
PHq7Z2pbkyvy3x4Kp0yPHZ3Ho15g6LlD4wKIunhFHdODJITgVwapVSLqphDpG7dJ
wcVx4CYG7H0WyxTlriPprSPY/dxse7IZtrfR8aobNJDg0r4MiIbmCT31UxLQPiUD
apbrBLPgLbxPr4bCaZ0iy0E7lnIGDMAk0F8hX/NscZvN59uCXwQbMehSO4G3pB8s
k125JzyKtoMsdzAABshFVtHa3Fxgt+CfGkwW3HD1xs8bUYvzVa15TfDn+YPuYCkD
5572ratMDYQBfkmHoBbPGJYglruRsuPrfdjSU7XHNrkBrcc628iotlkA1LucKbcm
B7pCiQltGl9+xq1FkXbLUQrfsn+qZzdpqKy1QOSq2REE/VxhraCj5bmpQsDQf/bT
y1NB5uuyGkBwQ4ildor59nv4qO5eh93r95qPJsGC0eWyad4NKlBbYIw7YxfLVbRf
lJZ6C6q4Op+I0PY8cE0XwQUdw+1xje6JCvQ0IbniftbNyJo9/sRyA0EMzsCx5UPk
A1b/E9f2gNrnUMJ3JXXWEQYCCavoaroY8V9HJiknMnzW8Wm9dW7xEAuOYUsrRWYV
Xv4YS7zr7KaRhxQmzUuTixPlIJsE5YZ2r95+F6llCqs9sOv6af1l5Hrc/laCm/5X
UNsm4Ry4HFN8VNNl0FgSt7V+fpgDtwGBcHAGNoRdRdgZQAlPMtXpUYoJMW69Rd7a
byQEb5LVSylGTnXszpopRguXKuF1QvFjE1g+DRtB20j5NCwNJrCj08amhxdcFW7k
n0hREh25mwFfz4lk+2kcGpoOvUN5sNeDgBkhx46SS8HEtBVV7+Iu2Lf6U+YyKk5b
ODY7rLzk6hKkRkTwnSG4vCGHV4xpfp6PcUKbSaPfxfWl+wMi5b17LEK1LI1ebCgK
vDU8txMamQqJ3aWnFC3VQptlvVLD6oDhHiUlFo0MrkcBOGghk7q3jWNyrqH3klY+
ecRIcAaPrXh70s47i5SEeoId00+5PPTah+aa32Y0Y2rsdhoiZZA47jrxtc6q/OGo
PMtdJnf++BEoa83V39smkDpB1AzZMLSNtbRZgvBr+HQvOcy1jSywYd/ufD9sGgE+
Q2EZ3zyxPGULbGSpNwNZ6r/rqfGdLyIwHlaMhtZxOBt2v7+ux5eGV+LLHPU7tiCO
8YWF/k18XoDeSYd49C96gP8ZOMq/xzqS4jr5JyrArsLbmCd7fVb0I9gCXlkZKI0o
1vtjWR7fVZKfJcrByvs9vodo1q2s65zIoEpXolXRqD+jaxxeSai9BTtLg7Uhs2vA
riz8ptctrTG3avSmzQEMcq6tSViM4HoHuhRSy9pgxg+BPqUK44mY6vftlWQmjZjM
PjaN4Cf2EFlTPTUJMb5AKwsadHYcqF09vYXPS8Q9lobzDfb+vckcj53oJ7tcrAsK
oeDhpptWxq6E6aiaXfux8SabUWVifGGj2MptFyKS1xFxo4B8uVhboqMHR8ik2/5A
RxzJ+kIvwEbyYpbO8PNv+w/iUeCmFcL1ygS6V07xEuyPX8DmPz/r+e9bwzoENF49
C42a4wxj+MmHEE+NkFywfj6SLMadrgFMpZ4cfVIL2HqrY+Xek7QLXGjE/OPU78kd
0AsbZApG/xX0N2ffXUXgHx26I17dYn2Q4mKNktlBckDTcGGxN3y4j9YtxTPquf+7
rP1f7fX2oq7aMbW5NUubRBGkX+N6lh8OksvBS0fD8pmezabP1XwS9atH27Nll7jD
UFn098vQ+yCKgpVCCa0ktKRNmJUGcQWLXjrOYPemDO4pQJJiF12hfaJkcqscdR39
fSCpxZv2NO48IKd4BonMt23KhapTl1QY1z2H3ewjlVVUFu+Wap7KkT3RdiItof/j
oTYCOmDHWSP/1VnAmlZYLS6UbGOT8jC4Hk7qtkSboCpwqNm8SDtdBbthBtcZidZ8
r7Gnt1pm9iCGN518wUkr8E1+LmzR1ax8CqDQ+Kf/lT3a/JUBxgiFoLwWCCldS2fO
S4fKrscn0rfy/A/XtuCpog6hF+pNIUdeWboEDt4ciGNSVk1noJquy7/iDfs2PyXF
jIAxWHSsX21JtW6xW0buqJOyjHM7E1gc3VFrxobhFGtTH1rHCVBz9PYtP8PNZ5tO
5eofNBkp5pA9KR4wRu+4ySQQCX/tXTfhJIvA0MZMJm4x5kn4B75i1GHceukQYhDS
wKwlaidUXaCcW0yIAcBfbtPyKvJUSgZ8tzdH9ZA6X5/EO5neZ5bXpqpxtsvDM2Xe
79GjGnBkssyacVrggFGW9HsFSVkFTXwKLcqLHeTMhAuL3A16N5diYLDJpr2pIi8T
NWRxuuvJwfJsqFGBZAJDemOxm/WSI9AR3oV3aesTyKQNAyP5ULYykFabBSbaOeua
2E8rQi0z8EdkVB4681dWz8TDkzQxGTTeC/pQcfnOYKizeN//cYnzqM0Jf9DPfhak
7p8v02bN3Q7YrLXmJXc2EUkQLU9U6OrBHJayDbX7bLNc+OlLb2k/1TvD4yUhE0LG
ZjE12OpuUsmD2sgwP8AqGk/1bQ15Xf3QtloDaBWGu4vU/XjMbSERPXynQlgzsZO/
s8717Mpzd9S8TTXIdrTMjZm45tZQREh5JsXyzBI5G7Tf0pdP0QpxU+2ciKqdxzfq
RmRzOWer6vZblrz9WBAUsk0KnV3D3WR6fXmSre2ajIbYUOPDPqCPEJ/OgXjvlQUH
hGsc1v8VJ0fvccFW8vW7LVrGF4NbxTdg6IXrTi3uCsOQ/incZSU9CdM2+USm6kmp
lDXt0wH0k8MpkvAsWIF5a+1nMFql5TRLENn+1q4BJkQKJJVtW3i4/7/hv/hO2hD6
wdrE806Wy0uZTuIjLACH9BoIXkHdeENKO+0jS2ezSWyMOyqBA/f4HUxocnwtRr/6
3t1fhMb+BLJWCrWjfQQd0cELTuWh3frcmCNixC3D2KMMEoOnWJmB+ObgTYBah1Ob
xCtFC8rw6sO3P014eUmEVdvLso3j6ZUySDhW8kHzd6UY62kTEMCYUZQLVMWfJAdH
ibgnMDCjQrjNmAUIAYEZa8I/8+YsUGDjoRNlwDQmcIOveuToifeOJqO5YZ848AO2
zaNTkVWfotEWRBGi6BxdWxaMS99mJTK5bN6q6HEEKbViSJjJ71/SQZ7efffF3r49
MNILnMEphwid9e+OD9tzoe4oakIE9vrCIxJLCybr4mYTankT1HToFv8sxg3KtNrl
nLXCw8AL/vPZ6oW4XPnHOnS0sY3MC0e7wkqhAHfc3oyAJOi/Yno1HxrHkcVHBubk
DoTl7Hg+THS9ILFaPnt6S4F9tOMYvnok9NGUXQHoxMy8M+sMxf6HoYVnFU0bNw2I
wHrDVXL2MadcLoJ3xBlX7mHPBdEHBJNTxyznfK5tRm8fsNSnGxl0RAhS2CELpiiu
N5NRtEd80X6JkdK2Rc5Elb1TnKI24M7/8Jxia6c4hsgSsO5OozYjMd95e7FN4U4P
OcjV72nKsq1eoJm2RKygQD+7L/65MChp+Z5O19uEVPR3BTrswXfhqySXBNRrfqft
5C5MZZbK79IkHjSoLnEioSUyJtQSZLQL8sM3DyyEqv7M4+gOH4xcVTFXoBaWZSNl
Rj1N1UXBDYr/EF3Chsk+3oWOIrrX1/X+u9gKkx2fO7u6Vy+Z0bhOXbU2yJOovzvp
Mqw6D1qNfMy+ZKPF1VOJbC3ufxquAn++fcD2icMuMNrXUVakV8fV0o4xS1nOpmO1
BgW9E8/b5foNS0absg5eX/Z/B71JiHq3sO8knGka5rLThXoQ6zEJh55oT62HFq24
+K1HYjBE8WhSAYW2yztVvbhFkem4F91z6g/wQENYXdh6ZBsV53CVB7lwA1YF6sL+
+TkwRfOHY5uTxr8d/DqVmB0uQqZnyfevui6NY8G7Cqws4IYFfMSNVdAJfHeJJ3O5
vzX18w2OWdnCNrfz1P77NaJUOKOwFwSzOCoV3KsMnL3EwRLU/7OIZN/KNvxKHoh7
al4H+ahMXr8Envrq1EROMzgLebaXYGpKfI9YhebDkGY7l5y5aBIbFkLDoYgMRfUV
YWvi/05Pi71l4ZL31iOCR5RYEgBc0tctHUNbGjKgSsmadM3oNWSqxlFT3MCjNnsk
NeC/eUzahi8TBLvkPxJm9tvAT3i+yfjjZmbLNaPKW92vOkdDX4ScaLkdrQBoXbUy
NXv0MqL7zI0R5D+bW5Ldzf1EysmMkDu4uYKHyJ3oJZu32MueONHnfxDBKkUXjCHI
Ed8HM0sZUaJhVHqf+5ZhizAFq7QeGu8+VhW1hkICWtDbkYWKegB0/sWCT+tz5FwI
5qlqSpD6l+GnE2uZxESSJBJGFZzN2v7kHYWq9VAy0SqI3aRWgalZno8+uw8+H5hd
sFLZQ8pXar+VnZii1rAaekcqa3IFEmj6y+W+0GaB4hweXy08tUDT56nC95TInw9Q
ooOT2KLpQSwl5xMxDyUWfuYfTNL5FgfXek36ZFdydDBGwnYWyZB/NNy5OVPXjB+W
mo2/UrbF/jPMVRrjsIRXHEhfxmZ/FMrfzd9DSdLJCQcaM1JypdPNrruT8v4VEYHa
e56Y+VAMs6vSusy4tOn2IXlZe+/M67zu2pFuqQC8pakyMj6X3I9H047w/ieaG3Rk
+JK3qMCfIH2Zort91gqjSLpm/wyjATJ0tyjYdwVGM7kbapYIqdlOMrctDH11L9CZ
4wgF3aQUMNs75+FRjO6iZE3pdunSL0MkH1LfVq+8Nr0fBvOKIZ1EWK5S9giharM4
vPkKkca2m/IzJTVd5d1Fxmk9K5fyDY96Cp0qVnqst+d5bacROKAgxqjw3AlqT8nl
PE533MOXYTr12SQfTXua34TXzR4vH7KBJ8JSSvW5aWathnj5IeDAQW4Gbn+u6soX
8F+fOH3BClITAO42bYko2zWvdM/fTc6cjV9YMJO5rqRzvSvDNA+ywPjwozwldq1v
PXlaF/W/1uoMaN+6sLaPat1BPbQ4fq7ybT4SHE96iYLJH+80o+bdknrgeNDWZwN9
9kFJfg76gUrRQHjC18T5bOFGmdFYKCKNXNWp8Jlohw2VO6Tv8zxn/ahgpvlQuOU9
33m6TD10b8bozVVbrzVSKvSuD59gXxkWpvKLJsd6cfokoXiQdngpT4wkp3ZsM/aQ
s/0YrAbGQvsfMSUykEDtjHa6NH9tJTrbkVTYy99aUeoHmR690yZCHA+WsGz8dTjm
dtTDcwuEsE63GqoBEXhPilvSnPNP9RCs60hgiEEmZ+DrR5hxSZtcK72o5n/OOkLq
fkmwjT/f2oyC2KRdJ5j7LRXhZVDOmn3Zur/25J8fFdPF9fOLAc9EKMdxo6kzKxjp
lcoADvj2xsOK2Kw8dEQAVPl1Bdx9pHrDo8+7ALDB4T06JS7f937v3ilzWc/o+SwZ
3/oS4VItfae5jv+xrIkZsE4O72aFdIVNyNM6VXlhWXN0CTMgeRR2itdjkyir6t7F
D40dUREqyWm4ITSuakwe6ulqdwbMPoWUhZ48yMW9o5y4Oh1A/MvrwMZ3YABW5BRa
2Th70UAHNd60AKdSb5H3WuxJ9QvV2fy54OrSJj2NYWoEFV+AcEaWCDBjVTdP1DhM
Sc66OhSc3Cib2UKCL8maqFs9duAjdstCTr3r+F2HtK7v4eMmmRPAzvPZY2z8/s6M
yKAK0OG/gg3lbUvbN1vVLUoel0wQAxbJLSpb9XjR2w+RPTusAvodN01x+A98nwF4
IgVg1A1LBkJZR+CkkdJj3FzHURC75G8ACQntpyMTGoEo6fdlP2JBVzkvZeku3k3i
ZTgQ5MJxDrx4+fBlGigqTAh1k+6GSJATyaMMz16lS7H5QRj3Y4awJct/Re0HYCd0
WbGKXsHz4RnM4QACJp+xO/hBef3Q9J87MSXLCS7vbRSkH54M2qzWJef+4vKVJtpy
h2fVTfZiDmLeFQQ1gHnj8J6Wt34GoMzR9Wav8j+WilThz+pYw3ZGUcfxzeYkssA/
o4qh31pEWJJ37bTDeu9bdj/hMwl5KiQKse+q9VfQ8uOloX6m6fPY55nbGeK8WXOc
AEqpmgwPWG+5e9/sUMWyhYffNwTEy9ln8n3nqULwNbGZAO2SHjGl3Y8xTutnKZfn
v2A1GZmJ7/Hjim+0ezWpGBU5aa4Oj7xVPL/oG+DFA9tZUGzDz+569JAp4kovKDwe
el2v/+YtzJqyFgOeaMFvLrR5rcRkxVeoLyrsSeZODYFQnueo0q0Sq01CpOcO+qc0
F6VFOw6SP1nwIsNgrkdb1LVegy4E3EUV1C9M0kii7nR8JjWxnHUcp+wjnto0aBK9
0Z1GEZ+zCNkI6IAPFwNh9n+L78I96M8pzDgXTd0N8YPAOzcpKxFXOWsHZBJkCahW
98piDqCcs4BN8lDnKb5Kmq16HhOAB9zh17ZelnUJnSQUThKLLo/iQN7pnBVhlROk
81xe3hhij9hwg96H8R0eZ2BGzkLk/oK0NJshhsDE6K6oudGDrVl9ZXLFVCWJMUnK
OGVfu1+dqPMJiKJa50BLCLzX3tUmW26kdW1eVxHtnVAfal5xYUORIweB7eHZp92n
fli8tLKi9XhfdIs2/ChAmnAQpfKd6pQ8BuhklS9H2ehwPO+SyIyJv+pwjxwdnQIR
e6JW1+9pN6kn996FdDbD1di+BEZxUtx8NEZrWoQF5X9ICrg2Mxa7HtzzYEOQObxm
QwSUk9fspDAsDfQfucD6x4FTKadWPoNlWPnGbpuL/xfVIaHBu8tiOv2OD45sqkyK
DPTOMB7arywrfSOG6C1wFJzdYMrjLwesKZtvaeYa//9UjhMUZGExYiOaWGYMbg4M
3aPCBYGVGcLS59EkWATiowhNkf6M/Pn1stBuT6Sx0E6QZoUXS+owmUdlgy9PNSN0
xTpvS62kxui4R7TS6JTzFPfk6Yn9JGoBpKGFFJ6THXX6axY64spnVwLCxM+L7sRR
HbY+Br/EhsT7Cmb7BAp8jqxSq4mf8GJ4cEdnw4U5P8OgQQCtBmW0raNXnhbnkw7k
/48UCl7RD3h3l/FpKozHRlledbfIT4iTPIXgEij+XaOcUA+0ypx9SD7goeNStins
EFH2U+0xZZZhtdnUJEM00KT3oC17ijfNLKJYLDroLwV0mqrYZnsY3zmojogZhGZ3
lTENwdPdErm+spFJIRnDe0R0kVDd4LdQz/+sG4tZXvroD8u2LrUowImCMYuPubd/
qElvwMKD0/PPHE0IH+j4FhBRXVSvAcdXIfALqAogxcWfFswD1f6SXFmw10OwMw+k
rreqb9K7Qk1fl7RVgZGK2jIOcbcjFKz4UCynuSXRQnyI5152Pq4aWUtQLlNmGP8b
t5di3tbWTTY5dwEKcWVOmVilp64PbIedvoR9Pfw0KwLD/Hexv9s1FRDBVlDdC59z
r9NiNFTvUGuzYCTwJXG5H+JgJEZ+Wm3scc3cZDYCLnFyO1sf1CX8+8zDikffLSU+
tqpY5kySzBrVP8QiTU3/trEM7PWjcpKMz7V9XjZjyJnqZMAsw31RveC8NX9brCN9
14EDgM03lzbDv9pl9d/Q4zijr+okK/j5PrLkj3JhqQqmCBRUowtyXVM4hOpR4TWH
S+aohK+d0T8UFaZegSUgRQnDUsmijmdakPvE1YAgVOAU1DopUvkzYES+zos8NBIa
3PbGz60akM/La78CZHLMxfbpIAu+IPMaFhoqphcoDCihdYokTwE4+L/bBaPToAFA
8XPgcwGy59m0S3u+/X3FevBvsmtitCcayvR1SivSb4at6bE0HPCL52Mgu07s8H9p
2QqhuMXMLdrhCQhR1AE2EVzzLhD2rHLf2l8FSREQpL9OCuybpUZjR7Pnsow8lZBz
Zy/jnKyfJcljn1hzVB/WKz27k2BNdNAuWBEzuKMZ+Vtvyj5iWbowrH/ceQ9WRN8w
W13CbU+gsvNvk1hofgVZqLfj5ltygQMzNHzi6G7qvEtrKJIo02qUqUD0LZcfwqkQ
opyR4pPRjmVrCrHrQhVlz8PYZClFDQSXvFl3mBxklZD2OQqlkxjNeDAnHFiMpT0W
TJRkCXS0BXj/vB/yNcamx6AfxzIIF1jcpG9Xc/7P8cYArIWZBFei6FlzaTeTNW/h
mw+p1d+8HQfOh83lwRLquEFEq0ZH5F/4QA1N77DPoz8U7mL4EL6PJhRloI/lb9n9
OfpMlI5V2ZWgVtnIRrYlUoz4eQtC23vTn42gQ3Sslj0h4klu2BC8E7Oi3Qk0eEJ6
dkrwRuDmWKMP/NyD8XGYW2oTd0vvh+V9B4Lu8H69UoplQQRxXSHotSe950Cw5suZ
9yXtin/Q6H7+np7kP6vcdUHteJnVQR16Kn4dlmBw8uO/2IMejmpGSW6P1hpYqi+4
r9jxOlwYL7CipAyeVH/pLD8WbiRT8fkL4/gEpa2Yprhjz3StMthyIQO/eL4s4ugQ
6jHReW4yIh0kTu50Pn/ROCJD56ZXkJ+OY6B2NF23/m9gcRQy/Ol01MRGmch+ubrG
0Q/82Aq7u3jvB7WTEBGoZ5Ql8HKEicKsRcstuWZkmQj0xHCZSvpx4cYcZApa0eK0
734MftxOgNt1Q45FaGtahHgzMHKWWpx0t1S8EorkTPmlT1O5D5x4UHE4ZJrYgqg3
0Lkhjuv/Hk40IiiR1R0d5wQ2RPlcQs6IlfGpBbbgwNP24m9WbLn/MdGs8PklDfc4
szgBa84ug/hHGjZTuDAvXwQA8JnGhXUtwiX1/GAVgAsXDaAKQGbR3kAY6vzKuwVa
kk71IIoqnpypcNOq39yT+ujfrQ5CVHNoFsQbHMaZYNWzSP9lIylD1r36fyxmk2dr
HpF/tXfzohyVSYOwre1dnJfWFqfWcVibCFYNCJ1+mySjnD/rOsxaB8PTrVu8bWAf
8Vix0p2MsfP/pA29xRWIXL/r1l/KIHxM5WRqr6r6bn9gxJcRM7fOYZPCCQviNJ6D
CheDg387nLZc92BP5DvkUlfzXc2zFnMFdfv3IAztf8WrZDRjVYEhcJ8b6yfZFqKh
tKWvhNXkicVDcde65ranCpZH68pubu+S2Rj4mIOSirpQfBNwZ6uYtq5mPHxyCp+u
59yymOTUeiwSd4+TgxwfIGUdlmtwaZ0d0j3raoFcQTS3nofarzuDeRcXaj+AlNFZ
tOfUAWkclRhLD7x5dao7fFkARrd9jjlRmP/EFSXQygUXu8K4dqGv4/78ZJCEZMh4
Dc2kxJ/h3G5ezxpUXWN0XCdA3AW38UWT06t4CVVqFvdyxGC2uFLa4+Zd/aCtiuB5
rRITQtOnNhvqFrh6ZFnp6beKR2ZV/xIOlFwqEhMV5XlMhX4xoUCclSd3VYV857sj
lUAVdyQ6XowmSq9I0igjJezA3J3uPFao7GwXUzwkpQRphl8cdT89Gn/nO9K+P/YA
DPlY2AkwC1G+Beh8ik/TBkXMHVR7TkY4nuyeKiQ5zWd6Qyx4S8konJUOv5M98fDF
BE+byk9vDWCG8BSIkpwXEqyfpAaerOZuLdE0sV2Sep519ASdmFDncOi3rMI65yRt
hulW1pMrChr7CfZ2XvnSLbkJjrHaPsQ3j5gC+yihQErrrqsjrPUEBG5wrOfVkdy+
N/GiHVxUh0qqjpplbcs4OYfFGqwFuMiC/ea9b8SKz37UXpwPE+f0ylmDI1jCPL/5
E64t/2e2N5kNwL2EkbJocKRTmvM0n+zvpmxKuqxHw4ohpBahP5e/wx7xpcDIPfAq
BZpW49aVo/fmeIj9qTesckhi/x/0wQ3jGJXw7Cb1JeHvYqPF2Zcm33WoVfaViMmF
V5XfOPZAlPtvejeZYAho40km6fEy0JB5mjoMyH5dcirFBwOJFTRsD3NOopoWkOBT
EM6x0UQo+zvMANHdNIkPgq+T7FXT5bi+pIrx0+Joaqic77bnLSQRJFz8yzB5AxrD
6UoOzsd+ryyyTc/sapFd77DqyGUQCdDQ39A3+fZVjbSoZpA+4uVFJ9JwBdflnjCB
dpY3QAgeQ2KHApLHrmjT0vnObxrDZVpKV8gT+ABZkuOLHoAn22D01dCp2ilMBlCA
wkyim6BUYSoH6F6KqiVnISyPZ16QEqr2GxZ7ChPvHIJ8dds8kDJDpCAVrt+Z6wq8
sQq02MmvM5/J7XPqXMfsdTMw7jtl4vyB7QpDcVW9wbsxkkxqgTZ6t4djfRyK+d3i
BXTOAKxEHrKeOKKs9iwbVSwNG2rAZHCK7nncdzJmixYOHjrcI3EYkv5CWx03mkrO
q1x3EGiEHZ36vBUrG3FJcm3P67w0y3Fq00CUFuLyxfwbXpHY0WVb0/PqnvjeD4g2
PCWm2YhCOrqyYkjgCBrOine/fD//XHphTaymUW0Q+XdRrROZqdGBck3/m0EGT/NL
0LmYuLR+OTGPuQKRxroBJvN67DLWvkBhOSHW+ALtByCfCOCLgX7b2ibp1GfMe1Ln
KABLFOjba7zdf8/U8VvbYsrF6CnPx4pi2Yg0qT28r7frNsgQnkkKgdd0Gt3oMDe2
fbR+8lreZeJ8c9U1IH0XYaU5SEPwsKbdf0yRuDqLnKkix0SQdQJDmH5lpdrsyPCf
KFVAx1jFvNiv0pMyQu6lcLEVUFbMEIbtpm4q524a6uiMXnueoxLMAami9+BggYp7
/b/eOjVEPr2Lbz6Rz8ixr6dxg4MV7Dcbo/rPMZ7P6dH9CwBcrhzfE4evWO7t911N
XriiTgaKonDCkQ1uaMC0OeqYr4TxBua6uoyFK47Y1fDkf9B6opksQVPQYafMuJYo
0pS4SIkSU2XSCoAbhiH2Saz3JXsxz1XgLOicuGrgO44qrq1hIqvNTi72htMCy2mw
pXCAw3nxhW6X1eI4FXsdhCrE4TGOK2FoV39TB7OC37lellBJRye13Wzou13nmegX
eI13oXUgDvCU11qNDMPSey1Z3+9T/p2hGNmwLW1sHFnfRvfcVf4vuwilbYyturFH
Bo8r98rVv85ICbXE9ratcZj1ynyiCL/xvm8LrWx0s0i8IXGyrM2S/eHP/TS59liU
T6Z2vVpQNUzA41z3s8uCHm1pb7crL1Q2WgnzjM1hvrdvbm4hkRQzbnLCx54/8QuK
MQwmm6NXy+8Lt8gWfO1oUR94R9V8AKYLAgGqOLHRh5z6DjMRzHd4FvDPteRiCVZ9
hKn0J2f4Wq9yAbZRpgpEP69quRfhsmnOkuTBiXn/30M0KZXroxYWuEHbwWRy1GVn
DdEO5s88/agiCRALLTxygz/GCra1eNOO4EficdqiyXq0DNluoYRp5FTN+jrwdoVk
FHWFO181rsTSuoFJUWzC1SGafrfW9hZTdMQh09d1NSVxHAwkIDgPC3tfXd4phvMl
SHVJbQyWOB1oZQ54rozMhzUiMBnMKxkchqE+bq8h2j/u+xNaPfcQXxqQPAHkamyW
NA0Xbs1v9OOWc2q9ms6EtVslzFtRrWhhXgTAmRBJADKkIwl21vyYAlAjtsk9lYOZ
eDak/xT3k1XPfsZgJOiO1T3lwfFtmgccsDOV+nrZCw+wGFgT995VFPZgMOuY5tLp
XFTXmWOaNb8Ym5XEXErJH6JJ60ZYbXItIwC8l6Va1zwHTvLffhkNeAtKxfHv9403
agS7e8l3UGBDXqoNfzmjkoI9WU+CW55Wc/n+E7dq3LerH0KWrpSJvfPl7S+hNo/p
HDTZTIHQr+kUEshEBuAEK+F5FD3V4jIrMNKqFfB7U/ZutIMwl5bKXDxlJy+1ME0k
KRJuEUQAXVXdfS3gaZ5gdRmWLBMCvtwSbjm+AsZ2yfQTTqlbu5FePo+yo5Z5nytb
xGkpoytBsh84/0ZqaewEfPVRfFELjtHu9YeD+KOo4k6nAg6LxUhw9rkWZUptPFvZ
W3xBAz3RZh7y+kQB54yBMHEpq5+JL9V+5jlY8YjTZVars6OrYWsze2lWen2GnQHF
l83KMFhY5p59HtmLBQqnRpsiJhItn3kfTBJtMCHe7lNfEfPw+Gunaf74c+I04ya9
ton7+CQbFWPxyLSST5ExGTx7GPo74nSXtU/MYX8CV3xHdAHJ4XHkhRxLHZ2kH9i+
9Z0686QeMQN+49uKvK084WqX5TxW8PQZ/ZSxO6bzRfRgfFTHoDs8RpIVMmONRFbk
wEPmXDd92oGozNreL75gixh2XmvkXOx4ovqoepXLXh6Ad39H+HWN3aGqGkAToS9l
WG/eylK0/CAiiUuoWi5mbpH6VHroVnrYyzbE1omQXSQuMuw4EqtUdeFUnPfu62Pn
HP+QGNAEfOmNQ7WYsrtburNuBvvpEHYoiSWnZxSwsrA2zQYy1DOvUFIrYP4Cjqrf
589U/+KUMxscW9aq9UuquneoGUBZ95jndr77C3OE1lznge3KJPs14qyeWimePd2m
Zp14Dfu3jZaYU0zyZcVfon+ivfvXYlIf+U0LBz1IbDArCFQ5znF7+AMWkwnskcM4
VQxQcJyr5Aq4Tei3grwJMn92+HltDdEXY27AfuRHPpkwlIV6qMNLEasJFDYNXcfi
koIecvNT3/mecjpVOYUUTyE3F3fzBmvZFJ+xNQUNpnB3XvLVUxkrgcEYxR7SzwAS
wSCmZ8PFoDhFiXUIy+NhKTNE9gajWjBeatoHEqBq0kzDtpQBJi2CF45svWW4RrGf
4tY+6SybFC+b6z9Gor3gR4X0NVlWD+NNbcOdJc1iqfc1HFLFvdFqgYDfMMdfWf2m
MQqdWyo9Ik9dwyyLvQBt4I3/I702goZZjoW5xIEAUj6O6EI3OglXrpLzGgjlCkH2
TGFZocnkcbVCshvLQZMAqwYFHoyXlo6wCdXwcFZyYndPBc1wP8IJkIHEjjGknMpl
e8VKqiHz2gBL7T8SJZ1MLOpkAzJeLTethl6QfZsARcakWD64lHf1c+NKKVGVL8pF
or82rDwkUajswXcLykS5FhrH4GbLOY6CJBmzPcouln+3nXVa2hI/c2l/x2bzLDRf
iY0yEBvyekDRmAxFsulgYV88HYuFrCMrYnNTYmA23BAyO/agzKAc8hrL7Iri4jE4
ZPkxeFX92ZUca3YpeBuLkCjY5Y2kcEHWiaL+QYSkVk55qxay52YTqdHfIKVrbq+i
NvH6lvjZCi14TOMmMz5k4evg+pQrkaQ8jANSRBnnqqFzHW8MR9cqf7TuYHEXC04l
9pijSjczYtQiKsx3o6bH5Rdf9HGhcdH7s/avDiY/wzxqRSs75pt8D0X4kHuzZFIF
iFW4zyw9NtoVsrwICIPpqln/zyjy6E2XeLM87GNnNpNdYyQT8XOOi95n7r8qTZEj
sYq1JswdtbeMYMgCVnlWB6fEPs0Yo3zR/TKjN8mt4MdkjLDWHpt3ElHpJC70vSMm
OJTUtrYyGmyghhUxf8g268J5HpAz5DjPK9F7wWCeTimRRKEQb6HV76cZDEA1vJ2F
cguCbnLN0SPZiFIAwwqogHQJCrqLtkGdYC478C/ksM/HNjubCbgy5haYly7pNvex
io/KZ9mYhTCfcqifb646qgEHyJtvl4HTwkW0iUfuiZnONw59NBIhZvgnReavUQD1
5ird60iLcsksPLJm/gIZ9QJ/BzGJorjbSJKamtLdHAOitaYUbjvbbtYNLRSIzsQc
qsQgXLEVUC0zVL9NKOlwBOCQetetZiU9Ta+G49GPBiMZJ5lap56qfwVws2Ej8woa
oinLBeZ5dsmbQid3oMJ3wApafm411D1OLN44UTrq3MziGbjEiusbvjEeSnbRwhYv
f2yA/2eaiRdX2TH2uWH/xCjKj1tBroZX0S9TyUKZ9KZfNfjWYb0xOZgC6iZjLQKd
9BQ+SqbLqEBMA0oNqjSWKjC1/ZYwDmDmJrXfLffkdrknvgfUUFzSyf/prn/SzF01
76H5egeornKlZVjGSC8+Lcxs40NTKn1Y2zxHpTxrfR3uk8hV+K5jDr/QrvHD4cSO
XVF7tX2jdqS7GAtEkDV/T1T0BERjPq/LpaZle7Xtoa0M4sH2ZjN7uHA+YUkcvLJD
yl6OxV2m4PIKTPaDnVHfT5CMFh/l8+z5kzrEE3vzDY8w4CJd2qt+lNxIOQQmrl81
ASTQPqXLoKefYiI8ItApjFYTMEp5BJmyY7Q+Q9v9tbuRFUr+27I/c5vFheBu7vxM
OR3KDMzGIuqmNii/FukwfJg3wmRON+rzp9COG+rb3UEPqBMuLykGptUoSE/ZmLjI
zLAnqweCjSHNQS3ateuc+dsgNG1ArTfgq/eha5LJ2LVwl9fEKIW9WyqQMgj28VNp
K74Snfb/GlQXdEKCix2qivkY+V+6u2HSaQfB85/uA0nF4z5/Vs73UhNM8Z8xGxF1
1VQgiooGE4jsNNnipB5UNBHARSPdnSjX6iRavTSFTVvXka+8D2ElWpUhwnlJrMh+
uOOMs/HzRoiNCUSmk4RaqSPvHZkBSVAH+X+7GwFBYAEXdrk+6osE/vv1XWq7uCSx
VXnb2UBRs66TTr0o/0BiTWUH6d0sGA2yf6NolQ1gXdItLSZfHL+RsX+x/A2UwBXR
UKjaJEIEXFSty64WT7grF/Mq7UuC9fQ6JPhECUJofI8iFG+1+shWIv7Oya1RSLkc
vUKxR5KgqvfFstK3nnpJY5IgirBWzVkg7cC1eAl30ho5cPZ4X3FZlnuCZcmaExCt
5KgoTfxCiKo94LGVfKQRQUBAm2m7EfmXHz2u+gPyGWG0p3njAS6/e0njpt6DLweB
zo7dJnRqL6GpwtU/+KBptGnHTAbN21exIUt4xoo4ISd9/gCtsvpDLA0Tr/8YGPbz
AypEXhnpBHBFmL/ofv9yxuJfuA+YADuq+sL4nFa1qssOsyQvTdm8H+Kj9CzJrFZs
w+Gbx3cf7aAC93hkijRZgZS8zH4a76ySIUJGievrmoOnpR1fem+ray7Sj0i7Nwb4
Dcl5j//k/lUG8epl3gtRARv9+DmpnC/JeZdaX88vnYDQNW4oz/g34BF58troL8SD
AC2Mb2G5DsdFIIDyyw4Tlcs2n6dTmTd99ynL+dbuXwE3sGaGsjJvKaik19Z2VRJ2
ZXHxlnqgEG517+zcX2gUrq9frz4/oa4HpmU2h3u5IwSfQieeRgg2K89EpC++mxjV
W4PlUrzcGBHX6qDH1jbNsMRI+QF03LxRfPvZEg4LT80xpD8tj9n9IA6LTP8Fbpq5
/fHoSDm8zlM2zR1OG3BU2GHSO2mQ8NeLoG9o07w6R6eydS8YYNpCnSYQM+jhkpAz
nuJmY6LC65Mf9XZh697pv+wwhaGGvfyZrEkVl6VpIjPqGAblFEPj78kL5xktwLIv
6VqoacyS/MtyKEprBDljOC4nka8tjdquUMtuV14gGYXA3bPIWzT9Oa/zLIpKvF6E
VWV7GkT4p2bzq3zgyd45RQfKy/Wc12XZhpxIpMy/7mTm262UOw/6VXQlgsWN7rWf
rmfP/XO11sW+nhfF2Mtix7x9PzUcYVgYhPGC9pfUHcmBWJOwbfkZSpaiLcFqximw
HMqCgQwCQDX3XAHZ1M+qPfu6BMPjq3DKlBp6Yr2uAbUr9Hwe0XWg3vSuY96O8XFn
2umX6hxp5bRNK6nt8mMN7kUKwWrNuQnuyq4QujG+z527wOm6kX/wi+XYJc0CXUVj
q2yOzJ303tmAvZiYmkE4MCQUtfIWWHP1ez6RA7739M6Vxx3mGa6RyELOQfeha+7T
4tCChVCCiwdlgTNGV0sBTG+okjqmU7jxXpa1AUbTcaakhjVbvAkxs2u5TI7Gxy2D
TiZ/QQDB/6jEV+Fwl+rHNphl00lIBi6I3FcoXE+Zj3RKP3RyuS4MDs5VdlzCTxrp
WAJqV7/ZM6Ub9Gi9yraCdvqAmSt4KXWAdhj/SLXwqP7H9EWGBDchgidrYuqevcqu
RXerq1TJacE8S0OrIOI1FXlM6/+g9BJcd8uWsDeJQBqsTJiPKqmYHRwb28tqzYgo
Fo5cLC+txZJYXaU9b3/tBFKEiwRRFfXDPlc99j+tbEZBGw/FzEJPwo09BCItZ/xk
cNc+3fBcfOBcuE71QL4Dz792lb0dtmlT4SOslmtnsH0/BXbLQ6GFTikeTWP+ANsR
2AAB2LktOOfaM4elSHzUE4wnblOSUXLoSRAvlIwqaLZsTquZWX+buz0qGhQ3d2nY
DIRiLD6l3h7YYi6sh2vP85JqplBEVe2ZQzQd4uL6F2L0bYPDOL2E5x9M1QIQaRxA
ZlAxUiNer4gaevBbBv5236Wdqcu7xAAiAP5tU/F9zlgxgx5JFa1A9ybWjtr9sjsp
6g9MvpL6dRBR/DVVaksi1RzgYMhC8aGJAe7Z5h30qqBur1jN60KSK1xrw1bDv9+R
o8dv9UtrNntKegMGOxSYYoZOXcueySr1WdOjgW12OS3Go/Dw4GdZJpHiokQ8bztP
x+0EBajskV8cE0TPHi5cxLk2LuZLSQWff4xsG9ozHWo1mVINOGNz7IYZBKbzkjDG
SrzEMoUShGl9ZRgT9Dn2hGuKHv6bATOByjaa4RZ4tpD0VaQvz3mNQYnBCGO74QzM
SCNlgPE/UeIuFFipcGQpBpvTZKrsTABTqn6klDn6lDB328YsbU0slk1t13MR5WZd
7fWA0fSNTTiOrRT/Mj2f0SFXoo4FepPJk8W8ikc4e4VjJEGywRq8on8IqHIpNaJj
rjMUXrZp9H5Z8XafHP2GjCZQPc9RtEvs0zcnmAA6OAF0fFYEzRppUNXcUXM94QPy
f/Irz30ZjFHxf2alfNHxI3Pw4PCRydPlpRwEWAaMhXHE+Jjbzom/ubwydGHu73Kq
FqwVtP5JhBf2TyzrzMHjzyY2aouSfmsVJhbI4F4fUwf1TdC2G7yfBco4uBvozT3T
Y5vSjbEl1cU2A6snEgjPmZcrOHl5jBsqOKYW1u2QyxMkNXhQ6J3unWbVyV8xp+/W
On4mTJUXhpyCTT9MRn2ki+ty0uTxAKUg9m+GN1ThcyXsvY3NX2yut8lSXS4odV6g
PYx7e1Ywd1gPMy2j0gPfuNAwY+GY3cZylB7MWEX6nmDg48Ed7gLs3BiQFQt+xyGp
F98+pmGRwdA/LkBwPeBkDWQ9LjbcGbjMmjU+j8PH8Y/RsflGTDorPKhvP/IJZVfv
lc4DhejBiVxOI7tM2hIIeO3uYpvUCUAo4qQgBMnuYIj0xShJrw6HdF/cgnTOVU48
HX1qD/0XfN8vuqLI97BXAC+kXpU8q5Gk8xiGvAWJeAbk1NnK/2P3gVDlQXPLbGOi
jbltlQHrEX5P3uwb8bY7w9hbNgx7UiuVIWM6L2ntbQJFlak4vS89QrR++fQuTOar
uiM6clR5WZK05cdlQAs5+MGFkzsm33RInRBoMgW3wxplZizkVv3HxyvgDYfeYQea
qJXNkb0w/1o5bx5rjSNafK8QTgZjaoAyrviVd5z30KBTydfYyteETwNdpyPWGRcB
y9TkJN+yHOrv5T2TlSgElbMxJLrlx1ySNHP4EVcQu+mOiY/DTwnTQXAk7LEPv/+T
Ny6uvzhEUXpdqsZF2DBqyVW4RUdiiNz3x21OSP2neHjMcS6w1AkJ2ebJrTH+Leiw
QPF0cjU57do67oWMf5qULBPKlWNW7UA8CP2RcKHvTcnZ07nAMea2YyZwH9Esd3q+
0eLYomm3PIoNofDrPS/ifCNVRBqq4rLO4K/F5AC+O4H5ybiBHG8cBtOHRQyhDBYA
LFltNNFxA1AL505AfSxnVx1zvNUl+Lp3CyptuJmb1R86K+6t/6ag77ROOzL6OB0y
eTEwBRdvKOPoDvkmVl7OPEckSlR/BCqmMXaJDCsnrdIBYyKIGU/x3fvA/gNvBy1r
Qu5bE3B6+iR+Ge1f6tGC7bQ3TCMlctaSZYVeVJiA4wS6Jng0ALuihatHSFm5RLe5
SfcstFuPqWvXsy5ub5cC1ZZ3Hh+R1GXQ5aw7UdraroNC1MuT69X/88Ra28MaRAIK
nyjFy/2ENkseGjy3zZoHfZDiKKlXm0iCkSuhzVxBQ/5wMsTD/tDkxrUFvZFz2uWR
feFerkAUCM08TxVMt+34oV4UzgjPKTkgut/uThW2ZvpAe3N7RS4r3wbIkZ6YlUbG
oUfk6c7SEMZNlopnLt2dMi+akgh3xGfk9wPQD6ilJwFG0ys37zCMQG1b6G00Rmlx
5Lbs7VinoFUZGaEyTWea3Ae+HcMN7KNx/P+vCi2k4oeUQ8ZcX7gzgwcg3oH4sQ+Q
mFn5tFdIC8fBi2q3UiQDh7P2i7eH+ga2MzgQVCllh2+ua6AWVE7UhfvdEDPpN7rq
YlrRNUAdUPdpbODUIwvTw+RzISV2Bg2pYaz/TEKUrS9LEyBX/pEyBLij1xjaz2f/
A2X9gitQO8d+3SCmaG8sbNqat2TWwgzUHEtZjmFss1SIU9XTad0nOk0P/5X/g7dM
nU6F42Jdz3n9bat2y8lSJuziOuXqPB8xuiXT1ZC3Pk4v87crrxum9gMTgTqm6sto
MeRwek4l1+Ohn5oB8HK/MEqK6wdZF6JfVJobckzNh9ECNXHQ/BHrQGlq7g1INt95
A99cxF7V3uQIb494B+mKJYs0i7S7S14K1pqvE+z8Ktvkj7PIWGWwFPs2E4BxuTRa
71FMW7YCHVgOpVcMOARv9xEnZSV38zCQE20c/3rra2ajhubLfbse/ysJKdCaoun4
1PmzPtgZT+SVcY2mtwWQz4fmIl4Ikd8i1eggpzbm9kj7z/ONmrv+DktBNF6S4iZ+
afishU9lxdyAE3Z0lnGG1UFB9OT6sfIIC1JYuIpQb42DuhLC79VSCo/vJADhZERS
wphAZsxy1+Mfjf2DJ5YaPzjX7xZK87OqsNHZleO9Ci/qmTVIpm1M8Imd0oMaz9b4
8jb7X7U7QAa9wLPzC5xXpm0X4qvFkwsPJqSkpQi0+iOY4bMHMIE2vy0frA2Kx5O8
54EfuSx6QFb4247aUCNi7DeDQtH8hfI5UnuSp3pf4VXbnjCm9yLR1FN8nkqDuElj
vweXR4jp48x3VsYoP4rQhNwIqNM0AFdS57dJ8Z0Z3y5+YZ8DML3TM6FeDEBdQacT
2GU/KSLY4G/KJYKZ4VhszrApZdKJBap6cQUI7I5pDlmPx4nZQNxb4Kh+3iKtJpBN
IylCmCz28/Xp0j09xMOqT5KgYiVIrAdbN8Q3iaU6CGDM0nnS4GhgkPFTnzSwpIRh
RumT/i4VN3346nBr4QYb6OMJ26KE5hr6Hvm4EjcsAJj3nt1MEktZ/mmMRLZtQhGV
A2quS/IvT5QZOhUgYqRbCMV4KoyD00XsJXBIw9bqePajg7bXY+h8vWqOrZu2USw7
RUlWuWoXqI4/gnr8/hqY595Zi+7SFz9Xbr+iQzXupmoFiYEUghJ+jZBUTOYZCVmi
vccx/w36KqBgePWsfnSvkOlIGz7c++XqWrwBG050T96JFlAre3zYRAeR1eN2E9Sm
o52QTDqfWpxLiTHlvS7ubPpDqVUs4wMLw9sbO4q0ioTtvABMbEpqI50Ud0Ir4hAO
elw/ACFae/JAVYzq6eB/zB47JxDe/fVqR53VqzUmhE4szbfUjYv3KBkXZfpXHkG+
Nh6Tp60fY7xIyNUUSAk7Kne/wIGd5PPxoT0oEsO+dEextln9EzEOJFnTtY3DKLAJ
NdtwqJu0IPtDvsebR+0ghoxXeiK5gq2TVVjnKdXOW5B+P1nl9DoaPOxGOfOdSWLY
yykw63rLEmlYyHa9H4kV4BmGDYx4c1x1BmKjLPyXg7t435nYnvkFJHjTB1snih+5
lCtJYMUfe1r0Ood2vMK/frtIsnFJTMARgHz065MXkIvGdjC3OdOadi7uveUJWk6u
k1wn+IFQ7OtHEVNcfieolKC5J8BvvzyAdoaWDWKx6C8/3bEJ8xLBjPO/59kglbMj
HJLRVyPanvjfeLdnxUkGDYEV4QGIIOSYJd97F6Yy2oxLCi+csYbZl6pz9uyiS5Bu
N5HZ7HHnTkbOUyK/dIo/uZBxSjn9HFg2T0NVjbFTQoPYMXvb6RBvh8nPl7sFxLDM
tAFGIuQzMf+/BEPdccUMaiUc+g32V1ZhwiXfc5eUli/SsQRIpSZM8Oo/Eo2i4Ids
Y8sfvHNUoi+69U7D6s45Xld83mzRt/VbvqDhsH1ipK923JqEyyPnWOGDsQd/EvAa
i0HVyRmKxbilNUSUnPUBDEHuHYZNYJIvg9AfDWoMvu5o3bL2m0sr1AUmjNr3Iksg
ZJnTZ///p/pxSFwKdoxn3VNLfU+112E0Iy0ChRP3d9BYJWCa5sbkU75n2NsetVvU
0xbPqvR8gZiKWWKoAu6LWrygFZtxa63CTiH6+mOtMfhMHRPcLQIeTC2M4luHgJay
ZquJMdoSmYK71Cz7IV5gNFXaUhXW0b9PQSxwi97thUZXNoCAIv1PAqSEXZ7s4uCZ
rqcJmUNE0r+Cf/5pzehIqFCQWDaU8ngYOu2R+u8LTVb443ajCh6QD8QBJnXFtiyz
Pc8KUACjTHE7LZQku2WKbztK74/RKn5X/hPnD/F2GvRaQd2QpegGmQdRHrSriqra
QL47i6+JA8+zMsuadVcS2XX6Qedj2s8IsTc3h79oqxu4UuCqLPQLJ0pzyUKlFHbq
qVOhEr9T4rho7u0JhQ6yO6smIeWwHdOSTR1+Sko4nEXONqto0hlb3gaC2mcQ1+CL
1eaQ5GNeqsiyG7xAAiY1NaOyICFPS0gBut204iJi37VR8qNWGHpwL91agK1zBp2L
Kf1g4j9HNRQ7mBm9nnRwko4JLjEGWUaVD5N7w9mB395fEzReMqJwQRfgefduskqi
YGhmsw8t3rWIqQI17WDY29XtSPE4mrlXM2/Yv/tgu0mEK/9RFoYrorkW2uhYa2fP
O0A7YhlvEIU07Wa+s4l1Z3Mscs1wrlEcGe6kAndDV+DQErCdiIo9SJNuQFtWU8g9
dmEPio4KnRoC9HFK1b+dxj3SJVCK+rrAQnpmJhProwelE2AkL2Td0IvLHjqUJ7Yh
1GNuSmbTQtB8hvYYOsvFJM4mO9XPn7Es57gzWV9bGJ9mlew20jY7Chu0G+1YZqHS
VJb3ZmsorLnWyyMA28p4X85QORuPI0BSM1PsIhV1WXdypqHlcZVbd5Z0FvgYC7MW
7UGpVhNvoZZL5BDZRUEpwznXcobhmlL8yrilnhdcfLPnf6r2us1zszT5wYOE/+D6
N+9kv9r7scWMBGjJuPOc84p0AF/8FMp6G78ej42BhDWWA5QC0Cx9jN5OPLjwyuMZ
OJZQzqJr5SWw9RoGnw7cYdWQ9QRHjmeLIb1WXI0s/CV3ElMqYy9dIvthS45HvjLJ
4hsM4KUwVxbZWv2H+Rv/pU3QIdPUWGi2wVes3ViC8iKWeTDZ9ETpbbESNIYgPiGT
VSK7Ck1OA7li7IK6GOA7iVaSR2OA3evHCggoOI01Wt7luVRfhohAIn4YiWZzB7A+
6MVEvWn8nQeH2lAm2WNnzks6NXJV4WZ/9deGlS+hYFCfnaeJraRCalPqBpB9oRZB
fUT4sWjKw87sKA9wEqConSYVsHOQeOm0Ga9t+emL3ep4qHZwfMgEkKf0LWRVkWEK
SFyHdELI7n9SMfHPZSuFEPjz+M4ouzdPURJDsWWTlT+UCd5YHa7reVYI/riTA6LA
+7Whm4rvVrYLrWg6TAyEbvltRkYXnMP3jCuAU8ua/q/IJr+UXEkuszqRwXmIBjTS
GPPpr/kbsbWsCjQS2Lo/5mnK9mGjfeWz98i5dw4vhE36qBmMj2QjotOF14+Uh9jR
/cpXJ6XkQTJBK9B/Z0Ee7K68glz9aS2IINlQhQ3lyd8W8ArazxPK+8il9LRTDeQ+
CMjOYkYlvvVutNmH3no0Hl228/dObzTOHtexMtKzzWXO71KmZGCWhqyQBHxGvC0T
wEJSgqn8YGeF+H4awGYDTCEGFuRojnpW/R6YwgXd5IVaWZjJxP3NSqinOoQr/tLf
UTOM8wizuXrs70o/5r35C+YgZlyY2lMYH65XQZn48cTWC6UmSs4bpjYzTVrG2WG0
J/gLNrPcbSqQLBVgxvFhAhol6LXLcPuUqDrmzy13TdccaKChk0yFRkQ4gpWNwseI
NchRAnY0Nh9u+BG4LIdjxWkYz/sLffqpGPUQlpO4yoLza3GHX/ECk/d1rFy6UIS+
/7wK7ynS7DrGPJMmhu6DPkCiCWWHdyqlwLxyt+Of3LpIoRbXATKC6ILD1OgWt14Q
FuxdAZsZs8LoTkNHciBewykouvWhRSPN8QHQMLVGltBWFQO0Gg3z6mXxX6KF8yTp
MttTRGLQzkpn8nC+iw3Di4yQ15aH4ZwrsVIhkz9Vgp3gsPam+3QJJCtGtGT50d7L
xlxtyaNO+kSv95fOCdW/nN6OnOJy8ME4CQwQX8pwBV8dvqiaeAeh3Xiv3dxvBwAE
/kDRuuefjZPj4NJuqS3+FHJE+zZTmqeodRXMEhTJhS5Fb2mdXGPGdvKoyM6CcGc8
OKeyq/R7XsrY1uTSUAQouMKCdZStPffDEGJx3+SE6O768OuaQ0TQj59wT8fgws9k
C05KHKZk4Zz5CetBJWAAASNyZHQY19WLKDRGmfPx9/qEShqEtJ9H1SjPHujSVz85
kFkc0+4DC5AMbbLnT6IGPYzZfjWGqVJhtQZp3tWSmBxGF0twAPiqsD/LjpDdGMYL
8ts8E2xfGGMcMW112pX4V4QUeagkB+66h8NVfHBxZ/oNByWrkHX1NQjKCU2TVzKH
3rzSgDb4sSTy85XGAvplbKNOwCRTPdtTvlXKdRBuiU/1cwl6860vPN9+cGgih9mE
iCFD3Aji+1mLZT/ZmGFe7B2eimW7ff+TIR/hyA8MV9w83WoPEgEM5l+qwt1SUgct
FqOyAuxRdy8zYX2AL4UXzypkMnma/Mhp7dyZdjuMIXNSZePhNPt5L2ikBj2+L4Lm
Q6MYwZgO8WboPJw+9+Clc3ZUfj+y3pBfzuC3VQY3NMq0THTfPoL+82HA5CMQugWC
4pFBKY2QlxNCYtBDn8Z6HeZSatkweylxrJfbQfHZLRLp7gOZm9/D1fMH+J00eds3
H7n/fyj1npxKpHeozc/ICyg9MJbpLrba1W94XCw5sjntKb/mf3QBgWIfIH78VZlN
Y/M/SvD3oHBVpIDJWSQGZa/BbP9MRZgkIYxO7xPFQZQe7bnx7Q4H2SEh9UbG+EbM
y77ONg3XOUuT1L9epygdDZ639flnn9tTX5XAKGLAuVoBARaq4M87awXPyOXwqSoE
rzeD+moIDQgvrBXyNJuELuejv3RV84dtEMkT7BORL3COCDzlk+GG+ipv+Rfs3DMB
TpY3aHa/cvFILq0/GBtMpXAV6CggdiFwd7oH4iOzKzooePyuSy2BmX1vtugd0U4C
7ITpoSmrmZdrzEyxyM9FAbRyMmE5XixtioJgc4aSQgM7U03EdGmG5PD7R/A0rmt5
CN3X97XTBrESfe5F9wby3/ijOQ2I0mW1Kj997usBqTjxqbUoUKeFrDpuqRR3QJE0
sW15J5gTbk1MWa3L/6TW77VhpJPtygU12BAqlJXYD6nlJ7fiHtF2Wm6OPhAkfUcD
n1kIap/+FPO1Iv0Ky3pZdK4L65QRxZYVSlViTH3TlxJSXhCruZGwVOXGZkhmdfpJ
4vPVPhrorLM028k1nW3H5GZmjoZa2BrUEjxkEdh+nw/ffzfVrHMbmGhCTMyvHgkv
t0kecy6qnqMr6Uc63+Aox01ipj8haXNJgWosHg8XBY8d8AQyJBEVv47J33kmckyJ
inIpvFho5ZZWpC6nfhADmrGyw1wF8Mte1F+124BxCfY7CzMtNNYSpJlEA44XVlap
3gNh8NRZ+sh1L8oAE9kVI13UlyOwCtm2uZVlM6I46ISKTOA0HpmLh4Lp55Goxq2b
4oiWPDAho4X3EtiY6jp+TM37vqPkjfFQhT5dnCpuguiglDSIzFXIIyv90b82NiNG
RgdYsXfhmTQYbjP/Td5xPeHqnHZCKrYpFUt9VURXYx+zQblRW+vm/8BEI3FMKpFv
ZQPckCLzXnb71AGSzIXiPScSJwExlyTUgLZ06AdJiTIZYTBcPPxn2WH5SMH4tVRk
DXQdMjHUC0krPwbJAOsPAd4C44q1s8ddbBoWf646KuvrKsjAf36nvZhGh8WtJLId
2FtamfzrzBrpXsCzyp0D0doHFA2zHGip5rQHAFesUF8kVWpxukqTntvH98Wt84vk
3fvLhrfESdTJ5Y9OdsFBJJiqBmp+9jjqzNz6BDo9Rkyi1TOUNbfIEwOUXUowUMb4
VFuRCirjdJxgYb+N97PKYjXpSOTDsGs1bRYM0Gsrr18wx+1LF/YqkhEABSBto2F2
rpT6Y7vcKRIkjnkzuKWkdnRGzneOXX9jnnYWmdzvxgIotJO05dP7G/Xx9rlRI3yk
yIkIORZYWVmqRpn9GCpFjFOjYz2mbB4Ua+QjYzDEUQ88+3KnOq+mIHJfABfD28hR
215cxMtNcLjTMhq8Ii/e+ia7WbhK9BJbzYTasIPYMabaYcmD/+K4yaClBxp9EP6A
pUduRs/RDiO3rn53B2UkuAXHWcFz2YaCfO17S3lAdHaqvJnAkWNh+hBX+6INQOGe
nMInZzcZMRl913vPm0WHao8jwW3uJtALD/sM1Iw9ay4kSvWzRIaqpdQdO/VHepWw
NuCYFu2xNXKB9CqbBw7fJxGl6brTs1GfqX0HrVfCxx09OfJcgN861+KGpfURCYaF
VLzWdKiqoqPf1x3sb09rmcoLSE0JaVrL+8+t2eOtn7l87FXIMw97BPY0v3X0paJT
XXVbsRyD+xBtWSE5agPqjkXQAB6uDTgnSuqU2P63UMsHOpWaD1Z7OjEL4P479pBM
5XtxfQ+SZnFZtacuAwNYLrbftk25cHdBpwL6CbzfC+Jhc/t/U2GKjcfEeIPHLaQj
R83jxvQNawqhXIHHvjti/p9cdL8Fs34OwyWSl6hDK/i44Sj4Tz0/5kW3VpbmfE55
RPDZtbO6kUri5lLRK95BRncpHGxT9U+xAt8GniuYR1fQp6PeB0MA/7J2UP7Q3jaa
W1sZ4KKyOn2/l0bZVxSZR2AbqjM28IRBFvmaVejSIne91Q3Awl054oQAUSvxRqeA
za6cNhaA9B/88YeepbmDhQx147DWo6kOvpBg6m5wb9AVX9oq14M0Bp3QA/3qNOR5
UedZoO7qIg/jgoL+/15INgWCfOAmezn+2am6GCElfXwFIxzzziJjsxVvOWicQnws
Gvs301iyB25JgRO9Ls4bf7um8RkS5ZH3tNXqnx5Q14F6F12yx/1525FvScC9tXxG
qPMiF9vE5s2HxN3gZdjs4XGAEQTBjyKeZwr81x6NMH+3xE9CtTpPkfq8T+vbRE4R
TlKQ/Co6ch7JVoCiAhZpHBZ/18+Yq9S7GIrPdYCSbxA2G3eCpSJglLxB7m3j0a61
5qpGnU7NtqnP2nfsqunlvT/YlosiBIQoEp8JQ/65f75vE+IfmMjQSgndgcHfpW54
JThlpeT4rSjgfN4ujywyugopJhw7oZh5FgKlT+ALQEQzABVCIjQrDMYN6+CZErKf
N5F7Kwzsu0ghrV8Jcjd3ykzQvIgN/eiHvtOl8HK9lXmnsQJN1P25pHAmORPRGK5f
cD6zAuA6nE55tL6zO4FRDMk0mVldo3gOuoGdaQXIBhkgSqU+sBmyaH8pqSrRMdiX
2riiiUkWcgm4vLpxd/hyap9Vu6CPuGHHe4P5aU2i7K6qW/CZ9TinlY6Is+MelQ5p
62xDr7p7zPQfekOkVutlqPVjqxQ3LBOTkA0evv6xLEBn4A08Ja/3Vcf1Vu1wYN1/
a78vyyohddL7uN9nwRSczt6t2wZlCJoBEhlJEgWk6kwyWXqsKsG4vg3HGYKXcbTk
b64iWZn2cYiDa/mAV2qP029zOJPKPeBuEX1yjEp+qcbmynO0JAc/QpZGFnd2iHfX
R9LljY/wGe7ENmj058w0DhtyaoUEIF7o1cRA3L56iP0Tu57JSUT6/aCE75pPAY9p
FGyR5A0p0W79yQvmd63M67n7Z4NFq1hvR11Hc25ZR1lL5nFefCEhR2Q5n6TxpCBW
87KMIoDl+GRCC0piciqRxeZDehfUozNHIWrWAb7MVvARRV8mvql6wDyogUpESSF3
cPmWI17KBYs7ca7wQgKcQXBTnrDt2vtRuc7AsAVB30O1dXPZQrm5s4bHO55+ThCk
bm+WnGbT+9vyWBY9c1lRjX+SBcm4Yrb8XJIhbRPGBHYHPojlkjJ8Xd0VyybKo/YK
Bt37GbH8dVYigwM09RF7Cj3+ZOBu1VTMX0eIaI8JSxv9lO6/DhwdEoiISLYdUYrX
htpqW8IVTkYGXf25YpsTviVB8lg8xieLlvczCw265EwHiEHfR1tuRUSLxSIoIwMe
HNaosAqNYmVtgyvm0MGp4x0EvyCH9wQznI9e216133TG80ebZwn5ESAw43U8yJ7v
hcMrmNrJSA3RyfhKTrJJhVv9OUPRnlyP+fyws/kY//5d+AJ1unU/Ybx3QMYd7CuE
j7ZxaYATlhCjIJA8BmDnBjL2B7nbLjJxXKFsETTc8rzs8KXAHw55Im3swx0Vn+5o
B92zjvFItoj+iuU/oreW9ZNyOBSiby9DPz2+ghlnmRg1cHqKN2gvJcKW3Khkod+1
1QaFpiMXzmKID5naHw+PWDm0iv+dH0ePwC7jF5KPOFxCPRdI5TcstzVlemBMKoeN
n/lBUMYqsKCbuPB1F0GBdFSOamLRA9TTEbkDs3sFHO2yygz+6qespxGGYPodxNTT
qDLN+dUD9N4KDf6O3m/g9isYigC2+iGhBCekpezigrliinhuAoCO9h0NGSz28ho6
uGQDMKexAq5ooNXiMHsY4HspLUmWP23232K9cgRLbgHFT4CImuO/3JqjVZ1wntOp
NL5/0tXCt9fscIF58KXT1lUYtoTGG817gLmYcLPUbwFiQr+edUfs0+NuYJRxeiYe
V8b08NS28yL+I2apTrLloU2BtRYmoHNVT8eB31ZBdp/STtzsm3zIjq8wqhUgcdgA
kv4lQ/gQA/vPDWTkgm+BhsIi9JjWYaFDXrj4nq1kzMpgGsJS6UYxI7/OUPf3K5rH
0z6Ej6ZU1qkbVEsHH/RMkMeyJ78e9FSQxg+5FwSO4LGA+KJAs40yJe6Dj5yFxuF2
QXf3uyf/R9xOlP0PENIpPvAoplLzimPL55VqMRVcEAwOcES41Trob6ZoWtI24Wtu
feMTcfDJ1w1O6gndQbKriwObN2ItjoaI8rCxZEh7VefAUxolHdgqy404EFOp2aOm
w5GfK4QYLfNsqlpqozGFEHupLH7TRm09avpIFE5DuwFgqgoydoyjSnNpjb+yJYFX
mqDCEB64uWkVlKmXW4xyUVC2zwWSeiJj8p8tGFO+MVSuTBX9S2muzBh9r/bLGpKy
zBGTD8J1W7lTNA/FtJhffYN2cFB27NC3v4ZkNwwaSh2DkXlfID6YNZs6vYuweLEK
b2VNfSi198zwclLFgjI6lTVj2pgBkFrBZ/oyavAQal7Dxp8ciX+Q7/qf/7n7v3QE
AZFf5mlHVL2+LSfqNnPUzI4nF9czTBwTB2/Zs8b+tA9FoBH7Qg7/3OwOkw3bg6v2
4G2ogCSrUUaiw/AwCAu8kSU8erhhR27BKqJXpsHcRqnTlrIQl4Z0U0UEukUnTscp
Su7IQ07EwQwwgulnVYqA5CnU3YMa1sErmhF0p5Sbz++IslYeNLpbXMdDYzUv3him
h0n88tLwbSGRiTveogeV+ghvCyzACh2m5eT6m4MufYQXADBYts++ETnOam2d6CDz
xpFnFrNW8bk7aPkYEO1tGOjla5ZyRiBNDNn6IZ4izscogWpU68HE6Pr3VnASw2LR
rz9sLplS/5/31Q7CseZnL593cZUGnPpJwi6tkw5knFQNvNoAI0zmNrS5tbP/ApKx
be5mr4pYHZTPT2OnS2C1IIkytA88+LK5KI3T6emrU2C4BFOUl9CguPBGw69gNH0n
wbwnhKbetbeWBH4phSdP5Xj70IPWk2qWwRbwwVR2+ZhREL0G9ao7Sdfpz7UoMmpE
8c/dwEOqN+gL8OTNzw9/NZTiaiAbzNYqM6NHbIZc318dplzwK1+Jsl53IIJs6EoO
ek5raDjt2dFqiZtaZnFAm2VoPlCHEZrbWZhRbaVx3DGW+AAaTpJgak6J7Iq0l6jR
DGHGRqpF4ojDcQwsRNWohAiZ/Au9u8cVzS3aWOmWjDa5HBKFM8TIVqFcRRABPe99
D5+TNWpbiAoDtKP1DoouoDuWyPFA98T+9X0e89l0aT2htiz86i3xbioMMj6LaaEb
vnrPU7o9MJGWlCfXDgCLccRL8uIka0vpd50BnmRuXOXenBpFo3yJrduCg11LSN1w
vGehq2MP5WUz9L+ygNFJ+RigztzXBntY6Ok6Yq4HSoF31XMKM5kOZqJzWMRJ9mdO
ZtOUhYA+REmhTixw1/2201yPorTrw3foPDEHUwvXF7hqvrAcQEoHmFq0F6fp/0k2
NGX/rTHzpA9UajjVQz6un/W2U38EQCIXiF0Y3SbJ8RASzJ1mk029uavjVQtpwRFX
RRjjvs0GxY7MKdzol9Yw6Totl6Z9dltSzVUyzKu7d6keIs2LxJ0Gc5A8GdN4LoHI
cHuhhLga4oiFDKz/LzryLfeqpA14fPMLcpuR/Lz+6m/mweZuTSGcpOvYa63aXrRH
RqhR+S8fFEw5A/UEwqhHQS270JFgtcr+0it6AqM9XQA57GYInAHdepNgY8c+lbyP
CKQ7A26qREHhKchWD290s1uZNGgc18nXeEcCLxj0IYah3E336+BR7VL6Ay8DwO4m
znXLX9yc7zGQejVUhaXNav2r+h7mgyuEVz5DAK9kkTlFfrLdlXO89Bw/tQxWPR23
5qAWwfktpbAuwdvY8lTeBjawIgtEJdmPvFDRO+5EX56IYcddwReWWP9cR3FbIInR
sYENWhZCNWRvIn8wKVgRQKgHCfaKdgcA4iswgX5DQkpPlx7W8bIaMfkW95+ZKuUq
zEYeoLE9RBw/Y0F1TsS4rEWUtL2+5ukUgOsYYIwBg6xUVVC+YHMK1bjU9S7MiWp1
JpLDvFA2pc9tzE2Dd91hXqRe+m0Hi59ZsTi060xN3EBXBau94fbof4FP4fao9h8j
knSrSJFeeNVEvQ+b9wNDgQdJAqU7wsLwPGx2T3kb1hT2n7mv+mm7qTY4g8BuUv9+
8S/OjrWTlKpD7092/equP0q/aReTtU1sUx8IwYdU0WDJ433JJ0MYvOAa3rWcqz2u
TWfpL8Ylg+1ib38cEa9NwPtVA7ahidouiIrGxgGoJtBARoqi5K9A4H6LsFfdbxro
iNsIAqNIkUZU73KAXDgcg5VXbHpKUsrvoeNe6q+YCOolNhtYTyJHQ69KwqvBiuJk
HZNtZoapR7BWGS4qhXvkZ0vzdvbuU8jekKlBJ1SFC5GwY8tfWvTs2Qa9YDzHAO6h
EVj8OJDxKGVQXemWsUJwzRt6hAtXeVE3av2AzJWuMrDycdWlPixjPWovxkuAnHdh
rTUFA3ZThYuw5WI8goGNPdsHOQqGQpS9LIV+lX+222lBM5PHOuUZGD7lh0Xh7zVN
qu1fmEjwmo3c/cDcWBH0RVPzt+nBLWLrRuIb8HR3xprx0qwklW2V+3zA0c/Q757C
lZckVp2VfPl6MXMUTYwQ+VJ6dH198MaI/Xl7V9EMb64/7tMcmoxwsmxERCjPNkKw
mWp3xaUf984d+9L6PYmzXyh/r66hOZtIyxwCmfdxiQCYlje4nnD7KCMP2qAqzxSH
vgJa2rYHeVAwgJTGuwfjCwWuWhbm7hru9aHJ1rDyLmK7+l8ay/9gmAmsMg7H1lTW
uKP8zVtn0xmMEiuXY5WQnEBU/wDO0XnrVWqloSJ4ka13mUnfalS+PAfc8Vgux34P
fdNXP71+qVdkmWvrsl+ruu9OMK9bHLlvYMTL2w/Tcal3WMb4epkc1J3YKXcvP64z
RDbZS52OfWi2qjFcx3dyd7JUIIWkljA2ZZzqYJ8eP649CfzJ06QYDeejMn9QOjAB
yTWao2hLTOFoaxNuGuEHCd9l2WWXu2dJIFTAoPvbFbCvRrtiL3/RukWwsLw8rXoS
Xf/F6+ycWyO1keG9Ca145QQ7HrI6EmxNq4rF6/7xL70qdlG0aln0IzYo5gt4tlb9
GL9GNCEFffgDRypE20E7sGFT6Tw9MJm8i7oEUyWaWgmMqhzVytvPA5+lnQsDwqiV
3ycdqVaMKeo4LqtOU32OGZiVP2f4rH6vHHs5CNneVy2zm5Ek5iDmb9yT4NgVZ4/A
JefxSpXSXTc0Lt00eV/7iktnkz2NmFfepN+M3xuIy1WwHEQiDviR6YJdryDskUZ+
iKSiBSrS7d5D2TU0HlNVCNXj0n81KZxrARMO2zb6hG3eh3LmseOhZ9LU6TAGTVqN
dZibfm3fq9ve0pZIuV9+jRiToby2e1P1JGZn+Gcmjh30wCFaa63XqOMvEF2egIBJ
foEdnrl9POiBDaisYkNUUgRczes7KHBVBwLWBo4nphHFZElLOinF4sOSJCi8UZ90
NeWFxESPqadYJ1pOqAMQHNTxOGXzljmkdf9B5znRfWydoAfAs2IYN0fJr7P988fl
JaXHoqHu1SJZ9Y62pnm2jg0vBKX5CbgPr9+WjKkiq82yP3uP2xjcwl2sm13B8Qwy
qDmQirZERlzbpamDhhRdytOry4JqpSjQyeTJp0Nl27Z543LEzWbxPzteiKEwrmd9
t95QUeOsspSkvQM7aM26yPR6RhpH9dRQ7yDwWCwwDAYBhYptCN2vP22xamyNcjrE
qgYDq7s4/bY6NwfCjyx6hhIxkjVqJhpBeziyh2/jWdmFLLQoDdqOP/UH23TF5vQQ
KlLbEu8O0Vj6MowRUHAHsoN1sym4utOYinhabdksaoEsmvtvAuJ9Ao2cSk0250nw
bA6A0Hp4KM1l2ZI3Ez61ZI5FJjENvAEHJ8f0vP3UNSmcHxPPKTl/IsmfKK5Fy2qy
fpG95/3UnejIU/RfTwRAtBV8wVFbsRc7XIAPmika9Uvn64UQK+vdjmD62TiYA9eB
wXKp7bqmWAZn+B1WMBtiajEw/8nsk8uTddwi8DrjFA7NtQ9/7jetrl3/bnBV/sb5
ciZksHRO1ZLTYKXK87MZalAlOxoyHaEGfg5PEaJzy7udfnKJLo+3odf7+k623ASq
xNMKVx2pJIdRXjLD8G3oKtnII0n7LnjLtDtfIfFJaqHje04iubW9CKwSzuqTXIgp
z1pu/7HG9o03k50vSlCEMmVXVEVfEpK1wLJd2kFuu/rH7Zt9eQART5+deYEN8VNi
A1S5T7qBFhW07WUyFfOoCbUt6JH2RdnEIccq4OiowLGbOumlVlplnQoMXsMtdlvv
CB5/b77ZS+aF7sOrgfCBwImXMEHpTKrF35mhVEDZ492POuyGDKG9f2jHErKOp5wu
88Sg43PO0eb33BtlayN4gH4IWTh5OGlbclr3CO84CShHpT2ohnn8ZvdiPWBlwH8E
kv1ovHT6IjPT9a5QEf0i6zxls7WBKiZa9FuUldxZVotAGm30Avy0ApvQytzp3DXx
8aY+udJGK0P23WhQns7CGMEyS56/abJcSLsBy9e4HH0p2huOOzQz5JkRpaQYC7Y5
KldGaO6gWGcY/4xlj/OfP61s4NFyqfz7HIbVuYpvvAU3uj1odyRrE+Yx8z/Ka/kp
x+2sZZ4Ufx01gSwplEztELtr7UMY3vcWPHniZ0LxvPnyqBFw8yzUMt3toa95hRfW
TZpimGmS9J2gpdXuViLGLSLWCYMkS7NM4GisXZZS3A3D3j8+itW0mjhxBtStpVHI
ENhtLWOljJSCfX3rMvFb9GM+PWQk1Ii2d7BSNMAUVULk5VoOTHfiITmggxqo4oVy
6QehsHlX1o8zbqYSGWExwLm6XBS/Khh2rr5V5N+lXgFT3XFwz7zdNr5/X5/6RzIx
O0TFUCkFbxaaP4GOBF/wmN9w/Fhd+Jtdm65XRZFIZhOcxvlTzv4lbSp6lwUwzYlT
fPqkRATR1ECN9fW19jdPsU5dpghy1zQ8sNUc8hcM/0DavNaF5B70DAqZcuHp07ap
YrjMnOhME6J6NU/l95ZmO4czcBrzJFAHZWNf1jjEd0iyEe7Pg7wyjcVhzBevyXTa
OiDTEfSnwaQ3gEgeRl/4Rh0LxZS0kPGN/IR4XaksBTH2MgkLveWHpGEN3tiIH5rU
r5fPHJ4zybetIc0QaBV+z8EIeBkWqBShnhKO+OWmwIHtYsUJ1d4o9odD1YP8pyuH
9MrKfvKOe8IIpoRbZF5dL708Y+6egHB2GI2iyhPspg7lYEBZ1JlocbGDcafPkV+r
NT2syW6faysozsremJ97sgLF22VmGT9j8+xMUj/HEYyr5Y3i6IDcpfbhxxtqfrCz
3xP3E52kLbVUiiBUzqVvS/OPG9ZrqPaAsoVx5DN1+T9+urvnI2dfxp3dGDSDUyGj
KYNgDOn+7w01AWhpBvRDMsKk8MU+E2NNvok4Uz0Ujqhb851SUV05tm7lgzxc2WUU
4i7zgBlr39O15bewxtPuxApwVcz/N/5VHoinhJdzveFUfP9J6bHpbAJWig54liLP
V+sye7BLReofBmtpf8UUAvP9EUDH8egBJO3ciSoh0Nh0RWZNKV8tqQPqNfv1nYxn
TMW4rEU6fV2FMKp2DWEVTfwN51PaHQmLnoZm+LNCwc8iePclGww1sPSZBIfS4v8F
gmeNeHqFVcYGrlO4ef22fwVAx+1arwXWJLhouhE/4Opr8ylxtmGoZ+HkvM4WzXKq
rT0e/LUaqrTO/MN0Yg8DjESrPpqmaX8xyci1yp1e6uYO0U77gnnZRX+MXs7kagqQ
LNPv/UiYwH7xXgJjx1rts9BK3Je3pWi2pOGCxJ0j1L5WQZ8TTgcrBFbjuIf2befi
4vDXDtEH/H12C7t9oKN6x/Ya13IQNeal00dm9BYhr0Qbw0Rb37F+5a5lapC633sM
JbLvRi//zYESKqFWdRfqlFoqNjnZB8Isg2QNJlrbE8KV4woNwAqDZdZwIEC48sZo
4EsTxxBVGAp6X0R9aDV9GR4KZCWFLnrmNLZnu61mhuF83/LUdrk1dohRYUOPBieT
eqMJIG6t/Uge+QCl3VYDC5ObnN12azDI21XBI6WYl/K2wqIeWALAyK4i2JMHSqKH
OsWEXtDg6RLpcVoB19vKta741p4+/6qMZzdiv8Uc/A9aKjskUP4tncxE2PlcoqqE
ecsP2rFhG8Ji0oTMLoq9y+TTIk1M20rygh2Qi4WCvVDXNdGToY1FI7pM4ZB/EvNL
oYsOhRrM0ykipaqLucMn+DC5hUHQVP0RTWsVauTLQ3BHbHy7gvGglQdwZ4KF+2Rp
N2YDbzceDej4W2DkpqEuXND0mkVIL3k9ubpmSgr13vbD6yL4CdnODq5WlYr8YXSQ
coBlgcWNMmlratP69vp26oe7DLNXneVYwn9VyXpxNYgCTWplPWZ5tBDR9qUBSdMo
dpKqtZTBsfe43AqahegNkMhsnTkkiEMW8UNloiqIowPd2LQC+7DvrVO9Qee/nZG9
nervHvJUe94I0hOs+G8iL+Xohp60pvQAVcrM/GDAH91XlrA/zzI9fBUdeGANdwkp
XM4sTE38kfTOKv61mlfht1dEhWAQib8COsO5VRGwslJpSU3QJpvUee3MXh41gA45
+nzt2pO+R3PFSl5l824n6oTf19nOsazbd0Dr8Z29CDbjNM1VIqJTA0WCvEeriuFd
SYgdXXhK9EvZSwcMlTGu7CUxbd3ozWxdnsf4UZ4YvDTicZWVbunfGBL3VtMKAOv1
Fj4maX1MACxhLh/35owkRdchBZ3dX94nFBgPsRtOkXWldwrj9VA9OrGvxIDNb2N8
YtR4lK+VnGlVcJV5zJsw8gTgvFz/LpdtkIZUek0Nhxt6wcqay4UUi3hMBdaJ7NFd
sqjmf1vY12br5ZDU2WTa/wArD+ZIt9kusTl1wbO2pYxhREAM+eM6kvpWyXrQrc/g
7jgJyawP48QD8TydcHHhlTg7y5qCDyQJ2YdimvA6IFmj46ufbo4Y1Zso/OrIcv3H
SrZrdTQANuTDzTR2UY0cjilg9X9RgI7fLE1K2cz/0idVZy7BYXjjLuKE9zEMl4Z3
rGDsPGH3zpDweM43zdlo35MyQZBemtVC0h7E04JPfSMoWo1jgSSCPeRAAZBfwRiM
HpC5695DlkhcOuMMxYjEr96ZwhdCPMj7hSvHB8gkmcv7UoSPO7nkH6bwLc581eBA
ELlVyhMtVikhA8wLhZRAwMO6zz0Mz6RgeoerPk4vLRx47nExe4/okr8a00CtoiAS
RvQyGNEaZuD8eHdsCm/1z0wXA2cwtN3KH/nhZk2wtUsHok+5O4D5JFPIpnt44JpD
kdLkiovsvdCjyOSfAyC1UBs+f9EhQWa/X/ygyL+ozXEvBc9YorNv+vOwiw0qMvtN
cln6pXH0yr1SHjN8rYK0Rcb15g2bDwzZKmtcGATspnfh9xtingS9De/JYByp13Yr
YnQcGhqZyb3h7YbcxDQ9NLRHnUAZtXjjjF+tTNoLd9sFm9l2dSGtT90yKXFNoBo4
X6R0N29L0hu+Gfpic9ZA37/H3n/owl4VfXcZ90Mt0noSgr/P1rDnswGxNlXxR2/I
252m+0+wFqnEGK4sMsRMvazxvc8NAwhQaHETs9gHtXPkdJoGpRmzU3a1QfT4NpcV
O29xxRwTEZw1zYj7Z1g4O2sBQ64kZ0Eiipbp5R2mvzxH0lEXZr6ESGsRuwUTHglM
snYClf+z7YiGK4uunxNvIZZrQPTERCWNA3UaJQV5BJxBbV21MTBwXTHYVAPhSWam
Lm6bOtICA/Jb49DBOPXAWR7nMSEQXx+gijQjQofbey82emYMHi15MQshb3p2Z+9/
S3UXMIyigJAoruZAD7AhK7FxDgxUvVjpiYblngOnURBOfz9BvT3vi55dN3wssArK
Nq1bMCGIaAhTzBGGoI1v2YVEsKUpm8Ux+RdhBFoE1HBXZMBDc/Gs8zhmIyuT1thF
4mWSAPuB0Mi93mD1ZlWnE75Wy+uXEorHf9B74ayT17DiskcrjPKcPpUx0NibBWa2
ORYKMP6YOPpDfVIAe8h89R9vJ7E7NraGdyNwh8XrmeWVC73FO30no/V1yr1zTsuT
8LgrmJK4SaU3aAKY7ocHehkbDuMnXwf1olXi1c7/QYMbylWhgxId2rFJ11JwsOH0
n1p7Na79Pl63nC46xnyTFLa7y2EFG0DqGCYLtftoM6R8cnwNxZFr/ZY/nj6rAL5F
U5DAGg0GB09qEPhiv7vIQThsEVUFhAcYR1mTVDoxcPtwxSQDhWG6ErtjviSPhTOq
bXKRsL2hMmuZ0JgpNeZvLGV8Fz1pryCQPn7v+biAfRJoUzEbUHCeexbpUYg73APF
ZAcSErgjwoXXso6Tn0YHnMoySqMYUWYlQX6lOPTxVFvBgsX7evuimjgkHES7nShp
hFaZO6HZvpN153RzSipgDywndqf1SsxvkeWhnSSdpzWzIb26csqTVEfNO8umyq0t
HuZ+G3SPIaNAXwGO5ygJtRFh6UyrRUx4FNkhRo/prIWGnHRLYBVAxhYai1bMa0X4
laoxuNGhULUXWHcOnKdNRLsr8+oIg3IFV6wVrC3qY4900JknnXO92NEBMWCfrY6B
CemLkpIdLZP2bA5spkoEOUKRv1AD5QsE53GLFCc/+bPIpTgfG1U1+lo1zxbielEv
uOzqtoRHAY9VEroF52qIjzMtUzZiF2Jhqoa23RX+xbGVKgKWYDfXkk4c/fQQmD1u
YfaRjlpbcL5DnlUFkvo3WvM+HCov/vA/QL1thsomOFlVKaAfYmy+nOjJkf5ZiFkf
zfpBo+t2S04dfzvMoI0H3QqFQFKDjlaP3o1JCx7ZN+MLyZ0DzyFH2uTszVuLraFC
lq9irvEnTVcDkiNvQFyt+WZBviI01vWAuky6aowDcRQVPzgoRFLpa0rPMVUIfBiQ
ghoO0DmQcHBiNg9pWn1lnzD5wMqLHADuIE/hEm3PTNu7xfDLSKLiji2/ezmO6Y9+
TFbCQ7F6qiQsFqWS8vFPWm8fXPE/JwHaR9FAmUH6J/eP0RZQHLnSDI6gIQtWvY7O
S9PsZerh6rFoF8XzhOuEDLHS/KfEkR7Q3rA+FzYiTA9Z82DSs4pzPP6BQcf455KZ
RfFyARJ9YyqyuplzG86Uauq1JVaYlcXPkzf1S7ASs+UZrqvfDckwuVDVtAeyG2Rp
xgrZJSGWv4cLHExHoQ4GFiYLJN5dQW8c+AEMHAf8dbZGp90q/6W+OCM1q3ofblsT
K9niSmarXbbBBuOrcLSAlvw9Azk7aNl3EikwqYawhVCfO/CZz25lavhpGRfBSkJD
oHYysBZRLrcte+i3m9LFRE55EOmXxTJjMRo6et7AfEVFmzF2NPWuGcBakkPIDPpW
qYMRiyNcJxCBsPfT5+M0GeLw4BFMvabk3056O06zbIgRu8KGbHAh/aWn4cmWhE7Q
J6q65ZUl7Er4/BvWId3faFC5BHw4aztDL7jQIgwUCCs2Y8xuA7M2JcYcE1gsky6r
jnvNP7avDookwvdGWPoPwpHKcWl1mqCV2vr3rtseIJorBxbKTCion740pIQYHaTj
/Mf7kzEy964Yv/cIcBMI3PRZgKhXA8nm8ruweerHBht5jhGC1P8Tw8m13bG/gr4g
qeYB+dwQn4z8P3Sk7J8z4sJob2uaZnjdBgADEBjB2fazZO87LudurHWx7EZvmeoz
T576nrCrfofEVL6X59ACT2K3B2dnwK1kkMEcLXrhVwsPcn1mh8zUgtaSzMXsfX2H
9FbqKZWfhD2PE4+9ZUmYcbR7F8l57U3qhYGtXHjoSxur7efJvyVjNewChpSMqLwa
vfA7s16Gs79gBw6J3hzZNywy5x/r/Nyh3svTfCt39rXcNIxrs7NtRqgYEWdA6ojq
oRXDPaMejcrOtZf5I0YcLhcUygGXDK5mtPPXs/LOLXnyHiaTHbKRK8oH4TO8bJJ2
cQyPfJcyCEuqkKvK2IL3euiKrYvVKMmIjfes6i7plUXXBfV04HeryI66zIWIWGOq
ycEa/jwcfxT7JVYocsYlbf3xCikP5GiVYiGrHwQERtJWpj/imaI0s6S7Zb/5kCjZ
YjT9jXkUF5DtTN+Ex3Z2W2Aog5FZNYzHN1g8r7N9wf4ulgFap4LgKMVZ5zT4rTCg
kpPZuBR8uOIToiMbcF9kgYOyjaE0Cp4t36sELiEXOEQgnWHxtfJmPQWgniRfO67Y
JYPc0zJxgpi5yA+u63/EQDXqzVZAYV55RFMDBz0Azf4skOHQrWSe018Z9MltsLa4
nf9KS/MYkIgv0s7Iz1B4S/vGw9qxcb6X2Ex1Bu++gLhdwJKxaBEQM8kUJxdnFfRT
jE7pGCtEAi3FRnNrATzTP+D+jT8lUVbjzgVq0lsX2tksVU9vHTJ8LOunoVbiAPc1
J9uMKbvRj4kIHoWbg0WMaifmLAitoGItHtTQOuwSb8JAwnM9pLirnNZ+dTKJF535
1Levw5A8v3vVi+wTac8J6oZBLHEbSFK2QGrcsKYV4QGqlD04qgoIfj1fDg1+x4NG
jpj5J2K167k+DyRraH+K+DGevJ4TZ72elBSeg5zeoHxRFP0thchz0rJ24JIM4EA+
DWgq4dLgpJRQC1A/aGpk3f3FfYc1aiA/ceqiHffOaHNXhMjJMS5PaAPeGE3MHEDe
SirODzsNPq39VXAyP85361M1i3YfNtNBDOWrIxkbZCCOQ44LGY7K8vlZD2VjZGOT
lX4cOzAPioSI18Cu98soVguDno08U/ybcxLjgmOdrM5olsayvzCfmIQfQwx1E4IX
xfjWX8OIEEtFcOTmv+yAsv8hEWBFvyV5tuJbl9kgdCCm1gxT52MZm+MrT+EzvXDy
n2Ru20vEuR+84rlhbegolms8LPZsPPpZ+JzggcfMzDJZ3Bo+GOKHftdi/B/B2Aj8
NGqryT3AzNUg9M1tWfmx3Gz1uebphN7IAg9FR+IME13TC9y8W8w0PUmI7y9oZ5aX
uTE/TneF1iG71kFtFKxJz+qC+jizib2O1ndQNZg/Vywh+4DqpVmL/xYdMMCWAJk7
URViIQXzMpNQDybHlVXTGcM5ZB51506yAA7ss0s12TjsU116aWJny9g1R5Tra6n0
dsrclesGo8csdkDJmptEiRK1d1j+m/tBi1olzuUsc5IHdMnJzzzbtFVhS6/qYrfF
pnELMw0fzysu28cjFfn6Zzr7fpUMNkaLuT9uF31iFShE7A/xoNQC3QIuKdOWuGfK
eyjz1ehAjsaDCDn+ndOAgWS6cVUA2HxC9BHOyDoNacXlRcEOivYlJHTQq0L+V8aK
hnxsGjZHjlFriLgAViulUlBPwARjw5KSgr5Z+Yd2UnH9ODCDVgCwAGINswsa3uao
207r/egoKl134VHRZQ/TYQ4OGzd0ouLpXAq81j8iMHqpggMngdyiZueHbnz/qq9n
aikcJVOIIxo0NU7FLnmwTfkSqiSlGXFj70P9ufgwv2JK4XVIheCpUWaDLYz96K23
qpeMO3vaZg/hD6AFMP9zXkpESgq+EOFCda2HaOM5NfceBcIH7a9w3VmIMderpG3H
1jiuGWyFZ/13XMiKf+6Fb4bVHmN4QPUjiB3UGT/pNeUtmhvYXT7AoSkPlm9yxTU4
Y/RbfXuxMYnoud6a35lyyX8uupeoS8Ck8LS9MHi5hZp7MtLOKT9D2ieD1OK0v+tw
2xEFO/7kvFFMGl+Df4sQi6c+GcNGQdxzJW+C2jiNW5ARGkgSwgvBMNetSDi9c8Re
hH5s9ioMO5OPS4Wk6IkU+UxUshT9CmZjmjC0QdAjq9hvyY0E8/5O8no9g496LYlv
vrIyQXcUkKHeu5YOADsfzt0AF1DGseFGcxRfUzY3kb9H5Qzx0k2J1WSLgZMDOScR
W3tvJ4r/L7cWKl95WVZbPQzhZ2gbTW4r1rV4oh7Kj8Vyhv/05X41q52TFah0jJ2Z
p6KIDa+ksqKBIS+PnDVg+yilKWOPd4BrH/OpP3p1OM3CkFPmJeUP33otA5GRLj9X
/7tIIw+tIIMhQv6uF/SxgfHIuviNdndrVEO95yB0cxPhziTEcdVfo0pvQT+v85MJ
CVL0fKrXdM8VOedlsb7gRexqWi7GsvCNGIM3D2NtvHyRRqcKj66DEIBjHsFZuWgC
ZgAKEgTpFvy5b+C0C4bSxotVlHe7x3JXgzjPC6/Cpz/qAfKsR923rFHPoKyH4lsW
g5f86s5EKqBhF3F7j0We0EdFSSwW6ok+KfdZTR/26kgSHAK0BGoVSW3bRZ5o3wre
vrmT7BJ0t8fjxD33arGeSRh112rknXsQtkgBOQKNj9lBXyuipzknYFqQAyIRhGBZ
GW25wm2jBVNcV3DQS6Qyd1JuyKSRMPmOnN+PjS4ZHmKbwwegEWN9j9N9SJhGTU6I
wYBl7bfDIm5QDbSjpF38rOrNlnZ6kwif/3+fz1Vg/zHzbfpvoSwW0DGcHkXs4SV3
NvRGEkBaQEDdBvUxoGR27CiwRuBC/AxaeiE9PTvGcbH+X0j0AcPY1SbR0Lvkfb5A
4p9dbtigfCBcGmqzx+nI+aLInH5EfoEBARWcs+UCaiFLZzu1y2SWOlG4LdAZvVJq
vqVoNzbHr1pZnJDXOZTC0dMykIk7EHnboBRqpLlWHv7iIv/5r2Sr2HPaeJ1DZo4P
8SawKtXSzNa2oqC8onw+44AIE/inG/bdr/xx6mZoPM1iPjI38ilPghqlPSVpI8MX
LLq1C6K9EZ2iu1p+7GNTNvekt7/4tGm5ywwg6RWDz1ttUBi+SdUiBdvntNM+uOll
mSf1wJnBQAZPZTwQ0ZCbaaIUPau3MsoNjnHJkzltrLX6FTK8MHkExbP60bJWNSJT
7LZCRolVS7LcD5GOZ+4xYdNe/KE726M/M/U9sq8O/qtqeWqwCo+Ez1y7pgihIkok
/lrnI8RhGUYui8noPqRCvWKuS3Yr/X03TYsX3LU6taMcbexALadhEYshlYHx8R/a
PbwTKt2ei5sm3qk0UOqoqEZp8kE5CX00fvY+Ad/yO39OHxdzNdQBSJQIaXyz/hpC
qjdBYkJvI6MjQJZHSUrSdQiRAwnoa5JHjzAz9kGGdlN6j74fn0pxNoFNF5uZPwuk
TLad898MH0KAwBlXBaSkY/X8aLoKLgGy0QasK5K4NdBX6+xFvqXwci2FUwmuyyNT
CLm2WZrs/uZKXi+ikyR6Sz5L9+mz93HER8tygR7yXkQ0jQKZGbQslVxPeY4z6Fy3
x3O9cmIGlcqp/E4JmaF24T2XhsTBB9tRK+/N43NQ+tEoJNytRlFa5iBYsYj6moNA
JLU9fcEYvLtieZFFSG+ADQkz5Es1B5dz862BHKJn6CsUL8oA7ehC0SkyMoBXIz5b
ztGjlVupztYNUd0ZNXrmly3n7srObGLrKrYFwYHAnWW9tEBuXt5qFRvHC9YlD627
zDfiIP3BpIc4qVFF70/iP6EeJzWylBbKIHi6idZrWkqt9fyb/AFVKQ4RnevBzxux
Gh0YOALR56lv55Q7ZpR8LywhXX6bdYfaNz62kSYHK1uw0O8xIfM732TcIPPkOW9r
++htHBIJOrR8zgXNpafjvgS57oZfMX/W7CkdOGktVxOWQjygHKeaUO8MpTFDlcvs
YHENFCAdImvZ6fK3f5WFfItRHcIiDjNECLHHV8w0ZeZmgnvMBGaSQcOW9MFBPFJ6
P4ZxQNZw65W1WBtIml13C1TJn9kfGFUImfrzz9NbFiXVPGYgZITYhC87hssIFSpw
TGQJzQPO/KrAWp0Mm2HTRqVS7I6VvBKyDqDVNOJxBVAYYZHZZ1Na7sCtNh4HtQwM
NbInnT1WAQLqJYQdpbwsrhC+TPRnk3wbG8GoGSE/3KDpluAPupdTYULHM+dtR/7b
0XpMKiXdHT+HeYhvRbroHK4x+5wdF1yswRyg2pFreJrINL/4p6+j6H00NZSOeXOR
KK7rTWKaYQcoeMbfznNAt3LZS6OwajKZ72ohsWw45ZBTRFZvPqO/T1CLch1Bq6l/
g7V40Ai43corlsQCXlsFqLGmHN2XF+NSv3KEUJtKHzEaTZvnSy35UsuMtcKGMgzZ
t4FeH/+YP8pmVo5ZmaGrDPzg6aGZUHF0y6TypIqIPasrBTckZiMPjWJddHhjbvGY
MlJboISXbJZBV/CSZONs4HhswVTqV4xaWdbxz2ob6bqqXcGxFYNHz6lroBBtxz6b
540TIK1EAyjQhac5pNm1lgOs4ngIoFDdf0lgX1Qw/1NLLyjfvn228Y+zU9kmhroV
F7VftxjUzNOH4cr1CUimnvqNTNIylM+zoEXgKMSUrSxBKD4lWtH0zOt01wyoaX47
4GOatGsSnryFp/2/78EwWGkGm5BuXd1OPIhZCTk4eR2HGbsDFw5EfYFuuR1I/QiJ
Ktcza66sKDwguw0aWVWyAuqV0MV5S/PkzNUWyGXbmeF913mtOPrp3XC0qX/iOPcR
/sfuNbs79Lsa/znMB8HkJNRLrhBzvvUcGDUzfNkgVC2UL42ABNwF3bMX/sFUP7sb
yk74AmLfyC9n/Bsf9f+TVib2G3cb2+LfFJv/vmIRSEcqRgv+hksLBUnhPslBcRe3
TR9XVipBCjlMuyTRmUpecFkx7zBruJGcCDdSKncvT7Fw6gJjYvhQRSVzqEZwGJWv
rL6Vb1Tf+G1VGNTEBwaFXZMJN4xRze1PbMmgm8a45xnwjUuTVbujfP6OFxX7P6fG
cC6oTxgrlzmNj7nS5mCYFrG9LH0sSwJcahs1g50H8nUYrFM0QckxEjtxhvx8NUEC
E4tJc0BrPMYxlEQ4V9p0I/Vul+KNn4FFsh+NSnr79d7czssKIxhKsQi9kxdiyFFI
NKQQ5C0guFWpKj4j7OpmBoAjY7oc+Lb4sgRDCz+mJVZVc6WeLA5YtFFZMCBFhnwf
+z925+09BJh5TgDAJeVeJI/BrWnWtgavUzwwip59IVjgzhF3TlMePJ0s8HXULie6
VNCLu9nZy3iPilIXD/cyxFUoS5uvZu5M997KjKamcWmIXwITXQ9gqXRykwIit/Jq
72VkrzWejftGNhnnCjzm9/UMr6XA4gHXsc/mLcELCBfHnnARv9GkFK1qjSbwzhd0
XP4cKDXZTlh+ao0SzfY20GmBaFbI88TLfdaWrx54WM/+vidg/LW+SRW8MpJ7+OhN
OG3a9TVsW1/4pTGNpl/hotxFweXyg4oY2uRzLND48kAQ6fE5zm877tc21NTpg/TL
SZgt1XBNpfe77HLe1aZVnqZKP9Vb+rdaDR8/8xvLP0y1446RbDoz82SBbAfoEAPz
A9YCUWk6cJTT7H9NZ4oiCTCtohpfsdjKyCh4CZ9eg5Ddal2OdDVrEP/Kh5w+g/2w
b8UfhgT/MfO+KCQBrwcmJPkImpvZSEE1BazXR2jkrrPxps9F6j0qo0n0m/9Zkt2X
lZHvH/qmXPqBNN7u3RWpKvBJr3UKOkafWfM2XC19iRGRNk7YQq5tH6CqUcCpHh01
ub6cv8nQ+3QIRtklp0+nM11ptB6xzbhVzrPqGfbd2CjxeWdCuMcaFUr72M+Brzfa
dq5T2lgbw9TJXsaE5wBBHbPeR/y80kW8PdtdvKdm0WIeJU7efc72lrQ5kE89FNQt
2+ba0X0qBpSrR1OXnYmUe6+XgTmJP36h8omTi02XsVThRHPTHaplbNxNqTxKcv27
UXu3Cr3H5LTRGdmuLMRaWTaSpOfFH+f5excP8YOHPBcrxb9EYxKRVXJ9Klx4WPmZ
vpG2nzAeyrn3Yts38ola/GyJ7Za4ickuUkbmjgj9cV+tJx6lZsIM9p9Qy6HLJWOz
Q7kN6nUI1wLk0DoATyWL/z8w+EXft/XR7+6Qdy9vBVxAYvw1smkRVPigSKWTK/o1
xl524T5RfFQVNvMS4vN6NeTpcdLRHJDg7UNeYHCjC3iUJqbTY0J0n4NgKRhqrQWL
EOWJlMKYT7HyQcf2z1cDJ9yI7RP/sPgfk53sr9yYRSy/YsmO78MDh1A7ZLlVN7Hl
RannrQpyPccb1m+/AXJCwakPAGBs5fMp1j/sAnvrZOrL/vU8B+s3d0ErYeZ+BNO7
SLhYD/FVWXYfuPi7bl9vI6aJJgy2xbhINg+fkLK2UphXbAwTrjtFG5SkePg3Rao+
KMXR3ZPTbxgfPXCXf12kXQnqCktiiiKQrXd9m7ed/6gycHaPJt6Ct9Hsx27uRr0W
oIoNWRgriPIhUb1PIdnTtf81locUJhcxRp69Q38pTlqXNk6Gu/tlFNxbB4g8mgMz
wppc7RWpdPf2EoB7oS+GuaPXZkCJCaZvH/MxIQLcwX2kyeNkn4uhohKUjqRllgF7
4PdrS8KybmrmBThFOipiKzTrlpaGSBhu77SsL7sTT0XKVuSBdrj/N+jHy3luAgH/
lzyAsOyNChJiYSWdRNoAntkrasV2qourDEYMW0IFJ5QG6XJPBD6HC2lrmMFtEPvE
hqa5M+FInNeyA5VPjQfWUzlB1weXCSGqykPZE+qNTdVqveA8hCMuLuo65y0um+7i
UjbN9hIB1SzGXcrRRePAyhKgEbj9xxqRQ0MyTbL4QILQi5okjTIH8OxjQOhvntRr
B0/yJbOClgvGVF6vsnQ39yjPEhKdCKiHbmHKEZR7NUUTRNB3o4kW8F67hbaSxay4
f2MOxEf/j3Mxso6y0CfctmJr3ElLYls7IP6u6MSWa3ROozUnsDoBEdhqfm9p4S/w
lXZRS8rkjdwnQq0KJ85pBpj5Zi0B0FxjcPrSPcrK+E/z/8maWRmJuVdfxq72AnpR
CkhKsd/sXf3MfnIHzcU6oPdB0RhL6cCK+QUAcLBX9qxWtGVglE5iwn4YqhlgdPaW
LvyBUZFVqeEAM+b5ZdS9+c2dSSDQFRyt2G7KNfjx94/6aL5hN9G9vyRgy470qaZl
rAoWzQsvY7PyKPM/TbfffIIa1stKi8Vkg+OXUsC+dS7AjjP0eHu5zpMVw0KQmaGz
fxWJnjX4xNrUPjbtz8D8cgvRbgf6Wd/mbYNT+BKHrZxR43UNdKRqSCG7h0nRIqzc
BpGwrzuV3UuXv3Suhr47+qh5DswkCITmL5fWD1WrmwXgkvxuGDHls43Q8nL/yuDq
wyJc40lw+7mfk18lFEJmw6DUzrjaNHZWowCaQ2H1uWAokShvjJXHV7IQTj1lZHQK
zdGOIlRsC5TQVurv1QePbdSa3YWzRqkTzr+VPJEnp3+v84ADMGXEe+Ms6xyqUTq9
xzkdw6p+p1nvpajGwilpG/67UtjQhpyqLSBVQF2ehbXrfzCg0uWGfia8tx1Yeh80
Mk701AZSsCRiTtvS7F3D2xBDdweqNeD6ZqT5uP1b0hBvGG2ZkAw9n3r2xPB/R5Vt
FJEA5WjCwW6CxdkgRmR3vlL2nNKsFOgC4J1o2e1kcXcmTKYwJyc553MiKDfNU9YD
WarUpumMraaMmpWCdzhHOgRIrOOpB09jzgsT9/evI3XG4M9r8DqtliR3FJAMMLzR
M0w623TgFBaPJWtLEW3oVj+okF6D18hXTTSHTSDmc7Hc8nrpDoAk4Unk6CmTYpjt
z2HvpnpBwNymNcgnpmJh+OeD1HZ26cNTa8NIKp0UPM1kQdbLf6TRljGIj9MamlAl
pf3VdbDJDn/L11RaJm/xwhnhEDcpHAb7IPBMfphCeDMPsz9DFsQ4EkVc0LsJ+gLh
yesZks0XZUzwMuEOVbo/5vPoIAcl4CoqhzCgjRdXNBYAbliU19/K3aA0QslsaPko
JdG6Z22mSjs5DZA1phJ/vhI+tKihaZS/yCxtgmqgo2iGlO+vh5Sg57Yx5S5E7C8m
Np0ChsB80be2l4ZTbMTepVptCruZfCMTtmTlbYswE0nui9jxWYm5HdpKus78YuQK
Px+UNTwMRnOz2ET2VsDvdCGnHJJiq1YnQdreH/gnugpkplcnaK2l1rGFXv9/snoa
yn6JKRehCnnw5BsKpir4LkhusycsESN/S0xABQKIvJ6U/t7ZANR3vNMl7nlGg2kJ
G1VP8euSLbq1FV5hHABDTc+an04b46CMW73QN0hl14X3zKqnKFO5cj2s5lrUXaYz
vGSBtYFe9NarWTSdBa41O1m52WvQIu/HQPElxe6b1g3ycUcjEDi99uvWeCPWWOp3
dJPEyiPlxId+V4rXg8eFYSwoyito2jJ0p82gcqXl1wj4CMK+5BtwqG9VG7Z1T1+P
PiKzGP0fL6X2ocRFb5vzn+CvcTONKWnDH3uf22y5PR/CCiPwYqUQOXTWGOU+ra1g
pWjO/a2aixruv9vOvc5grlc8bKIrpk4AmDjOppy70zOVtV/+XswwsQO/3Ze1t9aQ
OAu35AEnruAH3apkKwrDToCAIPfMHsqfrcQFNx3TpiSrO2tRtxpOvCEr8Mb58DNX
+cwQHRLFQ4EAC8/x7g6gvi5KRtzakYr3sggKBqd8iLt8Ve1JUk7+pPYL/aZQlVnJ
pKHJ2sFUjBtFvvWq+/XuHiRLRjEmYlSNdekHGX3Cx+e9Hrs87dXGYy5WLfdc4tpZ
98tBEiOP4HNWN7ecMv/4yhDPU3ruKYm+WwLOwfAbIxkrPaQtxUPXUu/a2AI31RgF
PZ05jKBHasi7v3wCtxgp3LK0ruPDgAdKWd5KafBIykQgxMGCBTw+O+tkXZMrNffy
jFLbyNp1h8fAn0ja+hciZ1nRJMH6iY/bJz6/3puPsgHNk0eZz7o3WTTaJXIV74sa
ADBQU3Uh9P5U92XV6HG6iRzDlSCkqY3MTHlPyYiHzhNGytRfVfJDsIFB4Nahg7vF
VAEPDMGTaz2PssNUEV9nDu1mThW5StS6skjxee37ozkZ8gbm5RnToJlNoAfh+G6E
hb9uVXcneZFum3f686eywBQc9JmB8nkSsw2ChkeaWRgl7iZ7O8+QZsUDh0FMuGaY
vfFWIBXdJKPPLm5yr+XhDq6ty0/I8iIvU6f86wRrGxXP0M2k8B1o+k08ZWY5IYDp
BVLPw5FYEI47jrSXwYQvRIhX+MgqETAqUCpJpyZh4cdWjWU01HA3B62olv8GEewa
ui4FWPlUr9uyunVetvrB8k/u1jrnBmI7BRXp2WG22FJ1AR84s9Dod6zGkJrU3/sZ
SgvXOIRoRiBtAWzqccidHmbJLojc5pTHWU1dwY7TR8rEofUZtZJAb3H518fYMSZu
48SN/Ds7yG3TrFmcngyE7Dqz2lcRTL6loWdVT8TeWgd0yeiwFCTDJv7OnjSidNpa
TC4g/oP/RXcuX2s38hOO8+uNyAb50wOnqW/e3uoQ6F7O92JXMlWUpruuYXH26y5C
t6JXdIONRmsfGHtYexUCU0bZ31XNB6cXPUrk3RnwOsdKneplwBXYkqSTdJqI4P7B
WRh0UQzwVkGzZ+MBoZGmOI/Q25nn2UJ4vbH+O70YrzTdIFDZY6vN8rcyNx6F/zlc
bjvCZuCt463uuXiU/drACvMt/Rdg97DyoiCbutC6E3jmNqz7X5GJkJ1r5l2PkxSp
mUt+PQIgMk3fXq5xhTSoDVelyiePhe7XGw8CZsbBWvdzofzPq0y+LE1bmle8f6S0
HPclTB0xoglAvCuRFa/WlJQ4VlDp2am4LYqfobuSMNfY0WLeLDzb6EYCJlvC75EP
rOpgXexvd9vdQuzQuVl4m26Y3RtPKSebsrPjHaaF+ITwOpT0nhaEAuzLK8/A9eZQ
YFFswhAneccYJP2YJHdLBguQwzs6dDhqqnaM23YLLpw9gMDDCwPsxJ7SG3+dHix/
Gr/Ij9w/1/rrmgc/IsvYYvP9GJkxdNc01EYhQloOztIB+5kJZbrYvGsjUsD4VlbF
b7gz16UlYicHqyfjUNGKrPxnR2uDUiZHNW2eNsbNIDe3MVRTYyB4i35PjJX6apco
S3goa/LtU52iNAVEBYRP8cT8KRHCEY4kHquQFS7uY/FzE+ON/tFeDnBlDaleqh8D
A/WT3mCZGpPXMZ55KtBf0VL3otaCR2xT2iYcrMWeKfJ7qyMk1xespcBADbUBZtjq
0hoX/uCCyGb428PaLoLDHdQkkuXeTJfLeR/PEX62D+XJwQ91T1yFBreH7jYgtYPI
tct2zq4QSnuSgWfRcgutxRZawVxlYtbYzomY3ie1dXgsYJxmGZuZzmxLyb8HPFuk
eEWWhcxRSdkfvOdkeQ71/fHTzYx78LX0/b9h/GjNLOp6eOapC7CjXeXIhnAUQTGw
AeHiGZLjHCMGjgQvJl29Qwg7/dSTcgtwPGiVl+yRHdNW5k2sUy9PxWnT5F4EUCTM
KHOQODDHMC0t6B7xSeSQeDqH1HnONNUborxOyLhhak+xjO/LAJPqGFuKfJLDKPwj
aRkoTuN/6RzeD7XnlZSOvH6lvaDdVjqyMSfL1CwhdpvIaKy4l6QWUUF+j07vYaOS
5A5JJos4esaOb7Mr5aiS0YmbDgC94yrpLmNy8nCfuRDllT15jNsmlAFrOXt2JsqQ
No9K4yvpADY3wrmvPAe/NezRmuSPYMpt5U1d1KLxgJ4DGmlalKy/p0QX0HMM19w9
Zg3UyGsNaA+MvtfkpPG5HlewiF9VuGqLTL94pdhDHysff0woJ4iQF/7uiQMx+MRt
3dNtyqT57dvh4BlALQjIXa6W+9f9ZMSIL4GP7sIvA2L/bdrB9V4pM98QcxnOE4SQ
9SVvssJtJ70mX4laf7r8s4BVpOO+2nw2HtTEMTnCtKsVjn1N6HLSfzWlZ6nmC+ZN
HtTHGjD2dIzmjv2YC35/7bnzElx04yoPRDeqv61GPQWeBo6EjHXP9VEaGZAWMeaq
UUxWvI8K+6S8aP1Ah+lj6mmHeVwc008Hrdci9smtxOaDK5skyZ6qWmMf1MKSEs0+
wPIMsyVK3Fm2yEC+ibJ5DvpNoWNDzdv//Hr6zUzvqma5d9xT+Qxq76Je27sd9594
JWjSilTEZfd2/X0noYWbSZd49U4Dl0XY8mrc/guUeY8NQMxjzM2nMlUebix3VkPu
cEc2k0+p53B0QKGy9Mnf+9LrJ2LfCNcAwnLkYv1u7JXb2YoanAUgWsQrngvCrrlf
nsv4gK7gnX5un/JuiMcvZwMBWICY1HB7c+BnKc6HHcnoiiJkEW/g+1D4kGUOFY5F
qUOF+BnyYLgkMgFwuUgIXvmcc2MKsydvr7iZ8YMHh0XJXYkGhuqh9oYZpWzdbJtH
/SJiVB4uAS7WmjC1QyBn7t4aFz2KiNkBhafbeSMGmm3rw6vpsiK3fqRzkz34mkC5
Xc1W7FvbfAO/sFp47PEpZS2U3FqEVm7FU6kXrT7INmCYUeuVwLQ6jprfkvBVWelb
VOU4cRsKCpNx6A1CGhckZiQSiAi7ikC7ZYxN4rJUUdpR1wTWEztJIHRsbIzBwI8W
3tFxuBHn9wUi4O0uUIeKxYCgUo41PA9tn0+DfKjzMT2vWhq3WZ69eAOPpMedx0So
f4J5DFwtM45V8QQCjJLUYzvBaFUgjV93MX6kStjO5Rz0RQXF17Rr+S+FgLm57Csk
PAXOHMek/+6XCXoqoqqWyqu6QkudcMDLjZFdvFRT5RGK1mK8soXLkc7ueJmtlK47
fw3T2XT5HUQfrFuKLiF42PJzSKl/85jK4uX8HfgQE7RuWNtr6Q5KWGnPyfCFqtla
/Rkb2epjaz+MEicdYivAuSwsIVaovKbKZo+RZSar+AtxQqjqzzG4zytNe+SVYmOX
NYLgQxBmlFs1eRdFzzTbCWe9nMJSD47vI+gqaAufyGMV0JsqYn+8M8rlirfTxi9A
A7m5/61T+GJkS9OFNDsy9SyBJ3Y/eENd8og7UeygcEOHOs1fPG0pekRNHw7JCx99
FfzhVMZExo64h/dykNC+A8M1sXN3tmmwWBozQIuCPeDT772icaXPyOdvVrG0BNwH
AXbPPJCxljRX91tIQUHIApxfMBr4/JnmtYKnQsj3pWg7I/1eJRuyIy4Wx/8LSnhA
OOGc4gJQ46TBTK30Q1nyh0FoJbGFYlG0U4z4u/FzCx0U6CM4KjmHWxDeVAURgeNC
wHZVTjXfFEfQ5b1eh3yxlQ06CzuIZ4X1FqfbbUjQ3vdgYnW1GWQUb2RXNgdtXVSN
yE2o3xUm4/BSbHbl1eez/GR/gof8cL+voChZwREgGgp1kEqfxTC601CeTus+jA7+
rnP/v7hPEcaJn5xtlp3xKFlRWOkq7meMUQnMgFUmstpmPBCpEeKqir6vLPgOa813
MUeTTjDQPiRPkPmp7qzysfhPVrrrWY+MYyszukJ+VSUf0bmzOctbB7dlT9WcDtih
lDBGoujjr2c8+Qk5I1tYgvlFCZpw/2ew8XiKz6i+1n71PgViaRUZfv6tPFMReDIi
dLWtKkRs/PNBwM7XNo8q7PTS4ibseOkXdNQpRzZawi2L/7ylD+VVcJ8xNR4/zbhx
hDrtxYB0EiNVuGxO38Xtc1xOpBN0po3bwQSKDWX6caoWCWs53gimdNrvN3bx4uW1
WrXJZqEMxdLVcJmmvYpRtK/UWFWHnQvlepYJ6FnGQYZ8ObrV/CeX9DbZuGbwy2qM
XB6Mtp4ryeHM4kF7rN4TDiNdx37KDiaKCJlO04hABLyt2PBrJYwq42H6itVhP+Wr
OXS1D28AZ10Pvov6sKnEjFdNZeRFjY9v0YYl+Eh7PS4NhSdrnnII6QEWgMNJw7cW
HVvA8AzB7alPtBN4z2iWImAiSflv7v+f5OQvLNMcF77xXIk/bmsUZmK6kQT3/8sc
NzUfqVIkh3hHHPFU1deUyNgsXR/s1Gw1NxzcedPp7OVb48d6xyCToATqi3Y6eZTx
DO0HSfcX5H3Nz6Lp2iLxPR/GmpfAZ5ouxxMDFS2MdO5vmqQM2H8WGq6nUDvrTiCE
0GoTAWFab2tpos0vCEE5CZEOoLv3yIQO3v7f32nY3zKvGeaElULzq98gdpkTBiy7
4FHBQqWqGI+J0mE9ja1PfqHbwMZFmF/QrUiUsz8Wyn0+NRJeLC7rnCY/pjCivQ0+
KYjWMzO2ItZkPRnJ91tYPmSkQirSaYa0rhVi1n4NxNb5kg1puolFCRwhcM8eZ/kJ
YmEjBqBlljbXOhi5nV7MTQYcCG3nfeErnj9TCv9jgtXe+XZF5m/itIbSqNhDH7Gp
lZH2QVpbq6BKF2bB5qw5tP6rC/HOWjDoXnXaZzB0+3wxhdPdLop8lwuZRaTja3Dk
gpaYxm8GdoZ0Vy+OYtjOrAHv3RNX6m8bofO1cHMELo54vt01fivE4jHVPqwbpbOa
W/Kp37hM0rIOeHF+RO7PXsxRWlRjUrKMTgB1Mm5ghWBSpcN5qorBFaPXcpethVNx
91x2c2xH2EIlx0TpUgB6be4/5Up0Yk7vH9OB1+wJ3e3vacAYeP+l5KgDxvHtsddQ
1zXMZUtKLo4i8eXqY4+3l4gcmbK7KK9RprR0b947li17oyfttBI12QbvAkO4+CJM
1s+pvH7HJO4DFr3y0POXPHW8a4KARwXhUSi8IQaudo/7kp1dekSx+s1xHEieQ0sr
ByJ18CaGN7424wuOsj88VemEqEYU9Sn2xnbgj5WDN2ui7RWHdib+mGb73hoaD058
DErk8NCYB1mg01WEZRjzXFM/amdyJvGxIfpjfCJVsNx+IlnFF9ugDuPZfUHLF1SE
wOC3i2LORqamfjEqzRiogs/TR9LR8uFcD2W73HZepzMP8t5DovhuxgW4U9dQRBg1
saGmNUphRyxSJ3ZjNdwfTwl+qFxjG564b5B6DkID2SCdldUT+21mM+c7Eo3mAA4U
32SmREzOgAUbod0TFy70JJZ9DDOzvrBKY2g12qWe7y39YZ+boY0gd/X1Zu9npKJ7
9UzZpNHOJUXGmgp6f/eLL/pkcEbhGTGvrHvYrQgMI0jYwDkdNS29S7VzUgU0tn0g
tZgs8JQKZ3o2VwTBh6kJLgzoOalpWKXKDliuMoX+4IVFxpfB3pv5ZQEHlEQeSMfj
RSCjsz8B1JsL5WPOrmZ8TbyNdCq5GNnf+8BEXcKFg0efecWUF+W+5tJfx7tu1WmZ
8LBMRQ/Q77Nav9Y55y2/Y6j5IOAXRJGQqtkFWH9cPWptspEcPSvvIAsq2HvMo5te
yVWIH6sLOsFmy+GmdJo87CTsuPRnvrXhWDFS6Sss/NWApbuWdW2Y379Fn9LKcSyP
aMfoMqWu1zlz3BtEKQQr/P2RFYBcB635lgBhh5MIiC3L0qCF3j9gxoftm2+Uk13e
kRPywFtYOctltPm7vyYq2IK4S8z1AfPZ26Md1KXLzIj4XjmVBjVq+Gae9JoQLGhk
j6t7V74FQRjDWITxLLKVMMbFdO8ukDG/aBh/EBWH6iJtz86lkcx9eJ1C7NvcOzWc
7ytkxxAw5obQB1rmCsEAEQla3hhDErqa9JIb5D0SBLa/3kz9Oihl4ylT9vLBAnX1
wZbaw5tDV1cow7jhzLJKH408UEf35RjOv4tYZqA7JW3pTm4TmnRriEAy4EEutPoG
kIS8SA8c6GPUFJDYDfkS/AbXq1Rp+/rHkHfwEDXcDZXXqbgYBWnu+smfzqCCileP
kJeterLrnhb0NTRKa1lE6FM/bHv07z0u1yczJGw8+HX9e3PWfi2Hr+RzjBalxrmy
EKni7rPU+VbBj3VnB712689qKcGV6s79qbFCBh2uiAXeUI9tsghTQZgCZtMWqmbC
g5KFx8Y8ypK+k/xpMoc7Ms0Gjuw1Zimdl1LELM1KPdfMuuy9g5STd1jV8zdcmW/m
l+J1apRyO2Jc4fUzsmgC86H+d3Dku8Mz//AkBELTg/b5PN3+1Xen9GbuNBu9mlO8
4nv0iOog3lXkICbSKeiunifrNc8KOIEF97KrB5QAizQ/twmWiMQB/j0CY1asqVh6
sFfDFblWlQhj8Wzgz7fpSV2XFqeg8KHTzZizuootEcZNy13V1tflBxuorzHkQs9x
G1bsnuXwr/yC3iBYun5wayUu8/ZJirDs7/z8hMkgnjNCirhL+t1wzNkVjaFa/w6w
YyBpjbctEvvosTLwhs/+YCXueM5Ig7XQA8bp2VHeq2w0dx1igt86rZ1phJOdLxwL
mtqWZkT2D184BOKRvi1aUh4jtx+/uq0MF0h+Pz2JoS817zWCAR0jJ//ozNHYUTyg
AgtzUUe8O/i4ZnhQNf1l38espTM7ngKTj8iKUcw7CrD+LEM8m81RGYBjSCUSnh+J
wJWz20ymI4h+8g8AhYtTzA/1kxgFALjYpRhDAaI/vQhLWYN7WPkU0GgDOmtclojB
WUl+Pk335G4kjspNF/FVLG0/UFofTceAvsezj90aUBc8OyHb1l6azrViBIqZlyia
uriSItgkdER1piRYu/7j2odXiMkB9wHWwJTQRD9YcGm8GbXZ7rsmTloLRwUl080b
xmvIYxBxY6kmgLwk5p06RaMaTm6OZ9aYva+V6hiK1Ddi8I1SE/Tn2xVuoUaLqkGU
sMGPsjjBoRnpaNvmVrreyr2X4XjKilUaKNMNSZ5IauW6Vk3o8gDwuEP0UPMfNgqs
v3ylS6QKhld3tnCghjpBPnlmw259oXt2G5noJh7GreegA5ivmAko0eRKoo5zuRDZ
jGcjGJja3perfjliCnho6riD0m1k0jUK6P7xBj0Qg1La70V1wPPrCFzlnAa4VWZh
qBoMHMwxQJaMZb46/ZY8feDk3vRM+7vUE/yBgcITrByGENxZf1RANVnXVZ3GX5Q2
zeixd825prUKGo4TsrpVsqgyJ+BDTjo2G3QaW0Tb6bDdyIggcGzpJXe/V2kBuuGL
4Hew4BVEXQQr5FoMgRQJFoX3rQZW9et4Uw7ukhkQpHLWEN/Qc/1XRtRYqUpjXlMi
al/adyKLF2yc+qbVupRUH/tQVdrqOGd4EmbfxtwB7S4bue6qnMfIEzQ3TTNfKXCM
pL9atpL35kM0xDkR/GKTR6bD7MPjmCvFVCr0If+47Qp+pGP9rbGQkqmgRHVoqdai
vE4MNgD+/24duhCqOjMlxr/nzUiTI7YLmaf0egsluuQAUtZRH7CkY4yumtjzQ0tz
gXpd1MJ8a2nbY75COriFKzTJkyQyVm+eezrZW1+dhp9bdRPXeVclCKK5q18KWVSu
2JQ+JV3rPz6NkXA/3sSRjII3p2lNhr8d8l1dxE7snc+AZYk34fDQWV/vymTemu7L
7fFwiFvFXUmbBcI8nwhyeSQWTd7wpqsn08ZoXElRcPVpmBTnG6WghvDvO3x2Vz9C
3kyE3CoLA9NUTdS2mJ7oDjdqW89sdN7WP+DEkawFtQ3uTtsZk8sp8Mm5dSQl/Axy
1rExhWNxY0LxqzEkBL9+q4BacgB2RdOROJUMaPU7g1LuweaT2PECvMp9gnYHV2af
sAiyM7Dafzb/3An8/EEhI5JK+x8mQ+JCq+fKkzQ8+GBu0BxZaNFD/Z+c1NYAdNWX
4cCNKnOHs80TvG6pZvUt+Eu/ZMmq0BoS5B7Kf/EPsGBEecRqYbdX01ihndyhOWRt
9AIExUxqkqb98Gs0RG+vjGJYRehpRcKIUlVzFr5xrnWaNhDr/o659pCu3PAESE50
hszXMM4wv19KIOVZ1Rpa5oNmQvMYbcjT/T91sM9uUfBBVdI6Oqnq3muikaJwkkSW
JNkdGb/FYtAU8djUm71ywoI0f4BKyKDP7HwQ9KL6Pt4WzwpaWPKVjIQ+5FMGb6RL
Mty4+AW1aqVpt+oDXhFoUPCGFQhOJhHH3d6vjoXZIs+kW65lqxY4h9yEnfNefXjp
zCknuFJTU/7b0mYmZW2B/kUuJ2lEiXVDzKNUL1MiBiKX/EdtH73dK1WhogiwgQ6I
hAAyji2R3gOismG1P5/UHGu411fz49s3WJ+jHIah7EXTeVerMW06BtpMKif8CQQX
TerkG9S2Ng4cJk7JpG68d5hSTtRjogzCLi9A+XhLAeQK5olv5hdicsN0sSpw9cF4
niMLbir2MYVksbRDQDS+BEf9REB6Dym7E9fqZHGl0ixeCtyP1Lh/V79z4FYPOq87
FgQhC0hU5QFHOHVv9AE9Mq0pE/K92ftOnR7S43W0HThKz41+zd3vH49YU4fBLV1o
16uF8DnmzIyNhffG4pIslQrxtS4h5ROa9FPnVTnhBG6bhZswsr7+muOyFweHLWv/
mALTX2zG6JsJLB7JGqs+X+fy1fTQsRzm9cuXqDfrAAfxucM/d2X64zxP1CicvHo5
JPK3nH2ByYtDrONx32BdF6E69ZxZD5h/ja5Fts/S/OJ622MylwsIjzQ2xogMs8S/
pOzia15dsT88FvPZh7aysYi6oJ4+U7N5yftoDB1Hj1F7IC4XAzmZb+7qcU14D3Wb
5K3bAA9rb1WQ5VaWdacV3a401a/rQefFSVCxAWNUugxti/haa9Cii4LsMSpXyI0N
WSB6bs4H2DnlcyCkFa2gnXMJ8OqsB2Fr6XuCr0fL+qLdcv8qH2Z01ZekR9t7lw1Z
QcZf4Q0U+8QD4ZVlI3HckJZPPmNuTpvy53sdMAjjlM2wrQWrsVZOmxK71rrJTnp5
cgaReZ5G9TJZiBwdy2A2kR2LKzVvt25EUKZaVuXQrUjmFJGoDLL70nSaf7a6nfVe
UwpMPPMf4ZHNK+SO9FYa1I3uXYSkstQaFQd1KXeaMn16g6MXnHa9vjwnDIO5nbDW
lLG5pVT1fBvKDUQB6g1wACFverz8Nz9wBDKGKzOA2eymn8FeNbgutwJeevSfZRK7
/+JCE1wV7Mq2YzhgLSRmzNa8Ulh0roNKoSG1cCmiPmjw5l+XoXLba0Wq8fqJFdlN
5d3xv1AxGOZhA4t10GOOf0Jje196z303SdX90yG48GA2ON8E27D6Je9GTJVDsS7v
ar3cCfaLgRxp2wvKg/LUnJduCJlCKh/O+h3PjB73E9b2Ho9httCdbRRkH6snubOn
XKqaWNWfVhA5+YDPJOGbHDeb9qmYs3rbWZvTBZ9bKCJ0aJVTbvuG8OR/XPHMNdkt
0pu8LcLfLF6SzuQv2mI0svppecq1DLeEl9Lkwm883XM4gLIkW8JshSwz1vmcNZwl
5OD3Op+yflXPhCwHjhiwp//Ts0lRA9l78QXOEAZiOmCDjpPI36K0q5H5YpAc8l+T
DjF/hD6hmYuu60R5QhQYiGAixjDgV0qZbuaPJuO7vuArNLZCch7BMcLHczT/wtt1
CPg1XiuCyLPkTjzMKHfl61hdzf/y9wfooXOmwTnpYhEgPHaYmqUL5Yag824iqePJ
MZAIh8wDFS8W/B9chRuiQsohVijr1ATML5CZAFzJOUABZPAx0h7MSUOx22QzktjM
eJUnlTQz2HGeGtJYYNyVkHBLQBM5td4N7VomVkZEHs75TLQvxy+nh4j/QWUQy/ZQ
7OBmfndgP6RreF6prIXqvIuE2ipWYOQdMyeWWy11SeqTHzRBCYtXYGrJSlBvx8cs
f4FBw5KLhnAsubOw+uRW+HtBY6LfUYZCJdQ2Kv/pIuFqSXXx7dy2hDp8fF308wPA
uSDb9Xt0M+u2LYHv03WjWD+DFf5y7bJG0g6GqfRqd54WKUzS+3AkZWco8b8TLaiA
Q8mXZFG1VWQRcqgEHl8Hz2uPI8bmzCq4PFclfeERfuY6NJygsAXoeO8Xo0ZNwb/J
vI7MZeoRW1Y1yJ1iGRQv0YOu6QMC5/rqBRttLc/9A6jbwflmnkuacqmGlH05mWNq
ZOXM2xfU55yoDyJh4fZVpxl9BxpRzQvzqOOL4VLpxphzrNMmrE2rdpuaMvVCbBdc
attnYTab3QyWuy7gYho+cUwalCJrv6GMKtiHeSlzkF9NeiTPv+4zdAXp5esL6Dci
KMF8gcONEXsXreeRJfFZ9KiWMhhjsDJXytXegRNKs5eEc5pcfs2iSrvIWqu9v7Sh
e6OXCzxWZvfx6hp6NldoHbJnmEaYkd3vUzpHGAEsSSNtitx2EylNjjTDBPRC8V7J
dd4SQHRQPHrhpTlTLcUrij87ImhLMRMdfABowqUsiqPWhol1Nuxx5sHPd0TO4itc
ErE84SELCaTS+gSf+L6XFUkU7pBs4+uX/agaTyYMEfbK2b44oWergNAMrCLFyt/N
mKNzzBoa5IYJ/E7I8p6kN+gF7iRU+Hu9U4Ti288v0vH0Xcqc95mR3lVjceTnL91a
1w665LVRQR4I5TPb2v0KCGOllQxcy24Pvrp3UB1jaeIsoY02rQjIerqo2+OWic+0
jo7hN/dkj8Qzf312qBaIuGfMWrd2SZAoBu350PCe3ZMacXcF/JI8tQpspBnRYLNg
ec53Xln3/ZDmxwWRgbtIJGuYVJ8gby515uY7m9lJFvyQEuWQhxL0UQXKEJMbmG+N
m9vy8I67bJkfH+8bOFTVwFgXJfk9FIvykoOoTywGwGs/nKhc/oytiiEEITXARQP3
7I0KUo0fbGAZ9iRbxDCz9PaSJJyW/75uNOnOTZkDColDNun8bE9uc4eEiYK71Z+N
8t3ju5CXz04xUl7liJScjkMXKWt/w6elE69ZIgMAU3WS9bc9ld+Yj1R4sbHnyUKW
NSkEW66By2m/9icc/SfXt+bhEFyzHM3fr/T614KCxpi3Lb30R1t3mxBatW3UaBus
qE6nY/wwQp1Pn4l3esBxPYdcaeJAtI4p3RPpybm0ptaMNjFIZIA+MgPstX3kmSWB
uo8ZuKrsJvRAhfVoIzP8mtUB9y1AFB/w4YCsdaE+A+GY+F2E3N761k8w18eY3MWs
EBg7kXr6ry4Za5bQ1hxAvMN4gnUazNc+Lv+Y1hfukZOFnIMhVc+cBNCvdXYfy5iR
4vmNlZf4h2jp9LaY4y73a4WG8bBnUtwpGI01vouh4xCRtIoTZbL2LE8gG6JPNdnp
CIwoexRWTCE3Ne5qGHt+82D+a3OmiEHDA4wDT844y2RRWodXQWefwCVoYAHYytuW
wZCACNh3dmMk2YG2t6kLZXiJ0+PXj4WKE4wH9JSwDlXTkAmaVksFjBsv6n24WTWT
eDHv1606Gk2D042wtROW+/6xxw+nQyZH+QI/RPYqTdJQ22DaT6l9P/oWK6Mx47ZI
kn/XBcAu3a46+m8rYL/z/OLOuiePopV0dQ4Poim1QoYkelb5VjV8Wv++vlIkHHH4
Nm236jWOyEIe98VDjMynzOttyzK3tD6EolNt+KsfKkD2Wh6pu3u3AZMk/iq2LrGp
R5g6MFBHkhaZWQWOi5O6FU9+n9O3txv9KomP514aE7v2zc/muL10/oM8bgkmMsqU
91zxGlQL5KpRn1GQMWmYsBrQ6+0j53npuO0Chqtgp0wfpspZwjPNmd9COBVGMzaE
H6iBfnlyb1bOa07/8onUBFzj6th467BB9XpoMbVJMZHLzt//lroBaektWkTun/m4
rxmTZbS/aP4y40JEOso3uKcZHKwgKUnjjQgwbeMAwitkutExHI1o06wZazFIZzhu
EjNXSSjq1QIuVbUTBZ5ypOXpRKFyiA5cwkqubhXefD1u36YpwIxlhgPcjA1nyRNs
iZK56yVUOIiqwCfTjTFLfnd0W3M/7862cHUIYJ2ox0Z2NtfWwPooPTPPbCwldfx6
LCsSPXh2d2mYWzxSBvVVr16QBnfiyT7afsvxQsXQ6i8dfwKfQbhWpU+VNoooEKV8
ngpN3xoesnZzDo3WkUecgtsBi2bY4gTvu8IXztonb76KzrNXSFNp4mcpy96I+qhG
RIw5hcMHBP1WKtM8/0YGJ3m7HjCcIZm8XjUih1uK6bvMmbih7xBwWliQmJkMC5FD
MmR44EhjpTERFV+2Z3EiZ8Xxo2c2VaQotm5okVfY1609gGWOYFKQgfyTSxB9upk6
nLp7rq0XM0v1LTDpJa4VZk060JLjxrZKm+RpUOz3JOt19BCgegKJ/2ptwKrmmQ6y
pG9wyx8z6GdLiRbm2dFAWNAeRZ4N1C3RVo39mZrxi1Xu1yR1gHbqXcQXqazq07/i
eMPGCi2Mr0oeFSdbaL+HIbOqgm60scy9qh4Supvx5TGlmT1XZz7VlIDFS7BoNa76
Eu9VIHAT/hgdL3gKoLjYzf9FIANC30QXCqe35UAkZDs89V0vsAjTScHu1Ytd8djA
KVmioptyaHNwrpcGJogIQEfcNMo2sG3Q0XhFXEuR6U1moqlhJDMkP09egQYnw4kY
bwO1zk4OLD7NcIuI+mWSTjBloCKHHw6wY33xVrVN5trfJryGp2E1H85wEZGo1m/I
0VxOwnF81JeFhPZcapnwT/7lHbhel/bPZ/brcA5TYmC5KcVvghTpxE9bQj3slwQH
CQ0fkeNZv0O5ZKLU3ycZr/CvvjPrll59nx8uVGSmWPldgB1fah43vVhaE2VeMnmk
wgwCj/Hhr1F4QD2Iu4PEi7FCTAs1WQhewfI8q1JrwaxqUWBoKXCFhCBBzRGK3Egg
ssPexhYmfZ7X4dPaNO1/hrxUjitMLQiE4vHN0ClpOheVmtRsmc+4TzF5vPTK6z/e
fzGuVv8oD3Ma1jp8YS87Ona+0x6GXnf38mJVvinm0CV9kf6C9UP2gkZo9PC7q+5R
+4Flr3aXnX2pj3z2OwMiJkmFYIdUpd6LZfeMzazfs7JrB1jCyS+6DaP6xeyh1wO3
szbR7rPaVXJg9yIK/7DSLPXjHaRhpx6bmJUb+N9v5wdOttq0SCmb2tNT+xV9torI
hkuxYqft0kZunTPfBsqE5Ka6dGvYxaIateBsPTIRUF6RWX1S9R/mi2Cv2eRLV8Jy
L71U0ak8kbZ+C/IROUSYApE7VKY+irsvw4Jn/tOtPE9nANxHbVM+Bb67C1QQqV+W
Jx8dtqZuHccJbzCY1f2zuWJmhnVHiZxlI3Gk8lNquPixPN4RHpnEHgE+tt/WDmPU
q9Zxume09crU1O7iFIr1PGyaCWlz0dW3EJq01Wqwe+w5LfU4lk/6U3YKM58yI69v
CRQkNrJhNpLT1mIF+45tbUy1j+suJEITCf6thXS6fn9VEQg73pXrOunSSu9OBrjL
3SbXRpEUfctqzVRA1WJij3ZlU0ei9XwvzsNDRQyiYTu3szvU0wLYqGW1i+S/G+TI
FEQx0l99QyOQUsv8JUrC6cI+jv3QVWVUl96P6at7SrQNnk+Az2RRXi6aq/DXaUuc
W7OcIPGldCkhiU0ThbMiEArHFRIAXSkmZnRbJfWCUnqWkw9ZH8I4BGQndCOHQgVw
HTDrhOCFfBAAOAaxwLC3eKstdMkRA+HIg0/rRad/kQpShevVSfRxN7fB4Y+d8V8I
fpQLmJh35opJ+HTHj1Z2AdGWbv4M18e6qxUgcqaidNIaX+E6nhz4AkvHAC4Na0Kr
vaFKw00dXuw3bBjuPcXH4Uf+6QmzoYPy10YWS6+g7SDDPrSWyCkYrWhDxky7ITWu
JKh4wq22I/m2TQPLDVjLM4+T3NRLKT4gFwGdzkHUscfGDHYBlRdtFHiUz0mtfGC/
62z+J1pAp8A4SLaGDNCV507pP8xB24hwD9/zxTx+unrrgw+/45xQ7WiYh5/4fI36
Tn67Z2XbIvqjnDsx2AYmhwe6xl6QVErOnmeB/UHtii6cYo5UMp8kBZtcRZl9qmXE
QDfhhslQRRbzhrQnOvwK0UiELhQptYaRJLDT3Dx9sv8+ma0iNxdjo4RvPFuPXTDB
gZu8dlFMuWiXxz7h0GuaWDKD2urgIPQrrGKwgOiadWse8STyQiNxRxComNt45WGp
2BFDx63Q9sgU9suChCt+d8WdIGEJXcLmisi4KkBta6bsdfpt0cG/OXig7wJW4Mdy
6zc1ZksjXdZpsZu90yQjJ8Dx+Y0x7RBdeji6Bf7LUkTM2ayYlSjtksqy2keBgd9Z
Ltggm/4V7gWqrC3vowoeS6AMzJ665FDwPBDTZXfTgW7UUQPZ0n1k3AKAgRyTqM8Q
lZyeCkM+zFlAMGhyBf7YFXb8i9dD7NTzeH0iGCLWNpV3WLvjc7eMIlOweARdoMC3
NZs8v+yo7e63Qf/ZgBfQ9FEXBw+qrCExG+v2XIVXXGlgu0zK265FmZIQ45T3azeC
ZG01pvUm5XbgjawV2Vc1NiTTi9a560dtYR7KfebuGeLXDlTOy6YmWwyGpTwgYHM7
oNNhoYyVFBtuDE6Ow0HKCpzaYJHE2ovv80bQQRWJBLt2NfHePDTi334txGstoo1t
vqjJRG+0iiwkWHS7OuZP05sCCvpsBCbV0G6TMwcuXxdkbQ9JY4p/0BDbqUYByvGQ
SI/t7o5ScekbkNM8fOEiLO73chjLR+SLTeDIPrgC1XQ2Od0Rq0Il80+jA6poYu8q
rlYkKkqff8hNI2OQm7CvGTp8bKL1r/ct4qEjNozWVw+TNr+aXYeim532HxibQdEZ
lKWSzX68fY+aODQA2rMNXh2WxhGY+uafUoeyEID8PPKNvKdaeZXiMNqeV3VvoEoA
H1HTf/VZpEZTIWkgEbEz1lm8i33F26fxTfn5SPLD6EToX9pOenBzLDEHKR6uQn/O
69eFGy9j6M2Kce5HpL/HCyRmWk/QlGean76YW3rn9ylL+0ITd4Zgrr1SFzjCp+2C
XHTyIs5P1cOSAMzNeMAxszrmuqO5gLxYUOyEvCSANEqJpHnTUIPF9IJzJ+XnQ+bR
PwQEIGWSU/wYcOe6Z9TeX6QZKQfvUMmwh3PkLtoAAGg+fZOwA3L5yfTXxKTBSDjb
noHyeKrXUSHR6HZ/yPcuQvTD8UlYGb50Oer0mdJ1giQUldKend5rVrjPDK1UkJsn
ZVZXt3ffiFTvi/r6jXUulwgu/osz8S2r1/J/fMDDSeLxyB/A/0REWMEXgymcNBvY
S6MFtIDKySLn/b9QQzL8K1nTIRaFkQldR1iQlb0jO6G0kg4xF+we4gdyohazYabU
FHCHhFNsfWMDawUaf7K6YS+nAJw5rerqRURNWHLpZZEyvhffJkAKLQ4vCJ11UMDQ
Jo4XFotbJILthYGdpecFrWdxPBHz6EgFtmKolfYInEYxGlWwukwjmuo/N9Io0hJq
AwOZEfKCzFWTr63cMgcKbJZrwswbM3v8LffYqkABEyELgO7+eS/59fdwj/mt2xwd
Eru1Nzitv/WdwbFXgomcn7vA4SbTlbRnpokQNBQgr0fo63KAtmE90mE2cG5sZHNr
OxEoC0gDLseEOdZH3T0Zln0yYawEQ1cBhinPCHrsukhhxTTT6w5dgE87Vuz4LDxZ
Dl09400A6eRKXIXbhw3TFBKAe+gGIMcjpE6lqrfECUwblUFfIQJyZvNqOve/adNO
U3BCSuFErtvkFOW2fA+cnXELJzNnG2cvq2q3W1kq+N5dM+hDa0eEwsG6Lc2DOT3B
rETcIP95Prz0KhAOKfOmT06v7D/2w68ZdZIcM5gsBiAzzT2UgZ1nuO93n/H9YvcD
iiEl3FDPb6Bkazrh3NVPL8L8JjRJpzGaKAISFqnG12JACXGPP9TMWK2dbdmJ+mlH
+rWreT9ja75u22V4FoIq4CnyJKBDkTU8jWIMEP5WcxGr3+u8PIpOl5+umPMYENV3
ILidXpTnrsyYccMEqLMH8+tk4PBK4I8JnRqFlWaFBDRf5f9RUbf+x4xgLBoXfjjp
XMaaUbXeKAqQDU5bXBfN2rpKIsvfo/12ZxW+v17cqCdvyjK6v+PDAEoOGL0b66e+
5m114dGKGALkfyoQZ8hygHABTghXghDQrx/4y8adLNFnmYB8kOXchjrn9wojoZ9D
35B9zecGM8Dud+6dZBAiwdqFLEv4VNFi7gCoT8U1qJKm1Cea4rqGXH/hHlc3TP7u
Dpv1SbMEPKHj3lmGeWf3XRsk139p7YoXzTSptC8+Jwpow/TeOSWAptBkp1cKIeCV
YfMcl+oHiXuyB5F6zDLeFk+yPxUNyclf69AJZS+m52B7mUXkh9b8mD7cOHJS6gL4
1xOOLAzJQ4t6sXrRLBWHiXMixoeOTiaTRsA7oyhMdsAmyW9NTy60ZRYqJBmaOpR5
rZtKMv3tFKypHborqwta9Z+jmaHrhbqZwz4gHRRgxTu5VheJOVTlsSPsLuoHg+1l
zhV8HH1g2DwtP3RPUUQmafYZZ8Ko5Tpkv4ztGA0SbcW4SMwyBwvk/x1oQNUJUCHz
cIXpli8Rjkyyr0w/TEuLJDMnwnqvTjaZvS3PI/6ZoZWWvxQP1KeroKvAKDkpKR1I
PUxbG0N25CZG5FnbNEPSIUmLbk5lSPOoDLbFVEnvGiNPWGbAhaEPyD+BG2sljTAs
OxHtYt7F2b1JAGQcy7psdYelAs1iC4StU+bRB5K7OD4hBWYlLHytzz8XXjt2YA23
tp8N3vzhEgTcBXzBBgh5LnuCI8A2h4sjIX+WEX0iQsC+kYK16uvpr5bvmIwzY/xq
lZuiTDD8392PUriiQZ9A0qokcLsYDAmxuFXdx4F4e5U9NtzBbhS9TIPz989yM9XB
GP/wgVYaYmCTgsqwnoCNOQupusP8Q4bDskXJ14O3tao+47No41KOt1ydVmou4P8u
3Q6dpgp0+q6UhpTF8zM2/24r35TmRtkauu+0+myKY17PiqGrAOZf1ZjDdK4+UylZ
6tQbPKWRnVYUmZVQubDkSUkzoMnAgYxRZvquIPVhZBMYYR7dplg4RlEuo2F20dLN
WywfenZqSKtcjL+VDhfdh6SQINZKEQ7F2RNDv3Q22T/SXdlBS25V9oXNopKicdEr
QRi7deWvbuiOijju1ILAyQemjKdtjorwBwmGGEAFV3HxnqzOTcC6ckREkS1TPlWL
DCqrwtPXI/NkzGEKAJlAcfOKW49hF/tT2zbnZFalbblKuY5ry0rKhWY/acj5NtoL
V36+TohpjIY9QLUTwW5SaNydMIvKbi4S/8Ztwsm2j2Ea9ut8KBKhBYeOGxfFC7OD
fBavwnf1ju6aAuPVwq0S/FHmrDJ7qsjQbf4ALAKh+mBG/m/qmG5LEh9rmxobAqxB
88v2qw2Kbf8h5xKxXQDAAaIbEIykn0TpPLayfEtBg1DPhZzMy6kZQn7rOYWwtOQv
EVDbypvDYcubCjZck9Vg3/UK5giWRgpiAz5ANjI6cqzb8vSAg+1t+akfM+rBhrAB
IJgDzd3E0HMBpt0o1H/PMMNo83uLoLJVrggMMdfYJqLIHWRel/UmxPyyeUcJ1OlC
FY3dLHAW/iNQ5yfrIurhzLxf3PXn9K6621VlUxtK34pqyaDFdOXD3sqHCdySSgQ0
3q32ss/Q7XcYFR9SMy7TKYVpq9ewh+KBH1exVIh+nv7RrzKwFVSx9/q14peqn3QE
2wDdfuiNcCzymTWRxbv13g1edcZdaOXENKWW8i41WtFAhgHXMBev9ZSbEqCZh9Um
CTDaUtX7ZDXztKTF9QAHOO1L2fjoPMpeH+cnGh0yM/j5KFtfEIS0J9clrUKG4Qmc
pXHGIZoZpNHiT4sLOd2/f+8Kh0If+EjdDKPb2adzdR0ea+iWawv7IznN7uL6KeWj
vVSGUYNWeq0xMVS69K5f2OE/Jm5D0RfqctJI6Kfuuymdd0FYRAVYTEQZB5iIh9Vb
MWFy4+dpS9Z1M8kUpiCC9Oy3agOR4n8+ZbuJ6V22VPHYPZPrPgdXGGgEZJ5ERriI
DkL/ba1M33rxoNgtqF4c0FktiFrbYjgrZQ/IQH2X08YZ9bicMmuLm+oRy9ww3Gmf
Fj3WdlG+IkzvrlVnJh5pifhj/mkahhFPYOCi9vZOvc6jIQEqz7+KhQ8PQ3Q8KGbs
wZ0kye8Z5tGlc38rAULyVs2hK7km5BYrtzkDzvEJqtGRFhGYQTolTVawTyJGOWaI
kHz9Mi0Ohv+RLTNgJAIup4bAxtiCUrhv08QnsBon01C5rR8aX5SRDZS/Xjv+gFKx
NGkUC19P6Gw8PTqsoj8kNY2YK7I4qWgkKxIhEcFy5HWJQyiQRJ75ApVFBsTRE+u5
2nr3JfusAr88NGrsuMi3Qsj59mys337mSofk/DFRY1tiPfcl939yRjO2Z6YAC4xc
Ja8qFg8SB22IfoWAAoUAdMcTCoXn8la31Ylv1WNuddqKeQQ3vSm6yHYF6dp73vM0
JHhcI9AcPOGKON2g9kh4U++Bp8AlmFIxJriBsywGmkZvRwSs33RiIT9kUBwRnxKl
KzKhRFZU6r9WKRPEQoMGBlXcQFkK4PPyPtxcXCS9Fx+WPP+0gnhHmM9ke+5cwWBt
7ovIRawPbCLClS5bcvNGn0jEv49y8+2eoQD1JOLeNQ61cHv/W48B4DJj2JufMbhi
Y9MgSyrmZtJjz/JDnoFuEUenunZHTaz1dJwi+5JjqKGwDCI2puDv9i3MeY7I54nV
o+L7hCxlmzcma0pfurwLvLi14IEG82Genw3No06EZcsEO+HG2rOs9kzt+3716sZA
kwg0M1AzJkX7K4SJ6a3Knay9lmvf1V30wzvjo6wOW7DUQ7AfmwZUuEN9gJ1brLib
u5iv7uNM93imRXmGDoJ59GpX6v3wayeN1gNreUTbxC9P8chQn5OoKiBbtKBYHEfs
JDJGqvRjQ+HzY9+XxNgGa//ygGTDSZeLhj2zzYY8duy14wW30RlKemRDvruD+El+
4tWWNSZBSn6ktEd6YO4bYcvOqxKW6H0H8FBsdf1cMZ2vcSiwPsShQY+nByrvAyw1
Y6AQDUTuvTA8wFkxCxN++7evzuN2x2KXxakvBK8t/EZrnDxmjU3c3aWeX6DwfOzW
FIsJNa7Oj2fzt0zgZ0lPFBm8jXJe/Gwt9A7ykbvG1Vi6qGNPpLj/fQL6oNo1/l34
4d8TCpUpqJvX+oPBSkJNhLovbKSwKa+h5ls1r2f+RqmEi2ELfl6KzLmsUpflamvF
Wm3YWxHoVEQhwzoz4kQOnUTHKQtbWm78h3dp7DwhGUNrgFraI9/5WBOJFJQ7nPrd
3uGgurDc9c1taG4PLzl55AalQ7qlmPdcKgEDdWqA2AI0ncfnHP9ODraJpcG2rx1K
msSNbnUIW54DsJB67EgRwnbdzwfTxexWW5+azUoNr2WmYqCnUiFLtGVKz+/GvaQ7
TpTSksEvpDerg59waVRr5W1WfGVIcH3Pj/7sz15ZW+JkAxp4v338UtAyBd7F0KQl
DSfIYJ6+MS9q+o17ZPN8/LjDNZYsAkTmKRRF6Fgjy6QYYBBjmv2mWa2aiyOKpnJ8
VqSOnqBBe7/T104YaP07JDH9wfWoWv3OQj023LYYF3kEsE+ZYUyMiTP42ReW+iZ3
xwmNCwaJRF4h6SG/kAFaZDe09x1BijpzoX/sK1lCB5r9aH9worH1Oz1CM/AjFisP
gNzn+ngOkdb4pdXgxApwt8It/W4+VSbFE5NfCHctwfKOtB7F38iUY8aJ5ESybwrs
h54MbzLFWs8bPMX1baq+8WRGi+5WZ1w/s40X2vqp70RxFzeYvF8mpc+PEaoi9d/i
dQYs5VyL9p9pv0GHHYtpuv8snytxTaiElMNOw/UxRVJ8Wl+OQnDqj9F/1O9/+bRX
/vVTjoEEjZblLBMki6bjOpTP1evwpUHMhSN0k/tCAL7o0QGmW92m1+PcW8WEFenK
K//O3OoNtrWt4kY91pzDEDABukCpMCPfTyCz7Y6kapHlcXl2O5a7DnXSVu+pKWpL
F65ZwTc4QEphRObDf3mvdzdJziMObMEYb+cdcfKsCSbpEnxOT2hWe/9hH+jkykZl
frG61f2mL3MRwrv3QIveEHHL6sbTR5QEU8R4/jOUv7WPGNywA/92Qv/R6ZEiNfHh
5nbXWZ6hh9lgoPiZjcknlbdXvdYWniWoSkZrW/iZIBTjr2j0Fh+VgoPJlJeIObHz
9Zq2lCX7A3JyB6L8WD2Q20q2kEqoA9L0cfz1P7lcjwg3P+24CxpuciCY0I79wRty
9gAkJj1+GoXSKsrP7ZMlTL0X3Q6oaLobloRUzmNN3NczW3+5DyrcQyd9DK9J75B7
JOsgWyEJvszF/ItNPVmaoBs99yYuUUOUGwfWigfPHcW1iAv7UA/s2C/jhkVcPJcp
M5yFWIKBGSLzyI5GjZFoggHKQX34R9KzDGoC6s6ZN/2BpDkIMULJpQZlzjRc1+q+
1FXqjav8ZHsLjsRuebAGjHFLoI3mzHK1THdN2ceIU35K52uZTzl3UnFiLUA8VFMy
3w40axEHrti946+N9YeK8DobzGYNhysNe+U+XnY3N5I9xydXy9xUAIZAlAAlyqSU
AEfOYTJbX8vGLXOhwpa+fIyg0vLTVn+nGeKqN0Ot11hn0/2kZz/4vh7gSVjVwURg
vXQZCfZ4lEYRRgQikxww54x2B9Iv6nvZuzTDPxCoWNjb+cHI3i1lZwtgEx/dFxIZ
k4ut3th7U6XRHXWtfgl7/ZvYDub7hkkP8vtY23l87jjMyOmP38X5kmOyZLte4Ipt
sb3cYQgirn8llkvpAUPATKZxx+Q1bdrZwU5L+ZuGxvkgSr8y1ezUzHg5HsLvoJuh
D4QKLfoBfCZX0vNcjtgjjUtVeEgRidAgqZJWQrxU4QbHBbpUUu2HqmcUoDWvg5YX
CjsO/WBXwJGffqoiR3+3pqibU0aPn1h7kW+xX+eFQuPxRhvqz8gNZZyqZO/HHljy
0Hko0GRzRs48TZf7a9yP89m4fJP/sZo1uVtHGOfRGtfSH16Wo/+zaq8wG5UomXY5
n88vCiVFqNLTS2tOWjTNzswokk+i1WrhFtWebOwRuFVU2h56RqT6oQmd2XfY1t6N
ND41DEWQaO0JaHHv2CY5SVoH5bPk8qPlw1E5jacLPzxnD/ZD97/44TWWA0fvN4xY
ion+rBSFsvdyCFBoGuCtJ7+76MEEv1E8JGU3Qlf0hF7VfqaNp8AHm9pRiUtHzxa7
XMbK/sbysGLnLqN9DZ/W3xcYDYP5zTCTdjTHIT0r2EWRKHmKnTQ6Kf52yFjTcyf8
/pWe0QeNZT4ayhLA6RYYCTrRPIqbRkRll0CXMnYX4wurpJLzI3oOmCTLjKJkdG3m
Ny8lbZUAKK4dEH7Ds2ISqdhd/J2uG79NywLxETlgo0nmH3pZ0kPRTU7Q32U3xALX
9hJ75yxgQTiqBJKKZAZVRyZuUImq8I1REYGmh+hHeOObA4h0PbD5ZArwv+/On+rQ
hi4k/IKUO4e5CCNkPriBP5+2ABYlceqgmS4tL3zhKbgUIPBdUwiL0HVCHg8Hnsrp
NjmwoaWj6rvyeZQdlgOOPKTDB9soEZT4rsHLpixfbl7L7rtme2doEJcfL20Ra1To
ioqr2QFXQM1f4eiYuGFZJsKj4rGMLViyXZZvJWVayYQAYCrPHdXtmHXQltiMS7F3
NDnbbJ9UWRTMK0Sn7Rp8o7rFqzubyZQWKsER/3wHEhN2bKtewWLWjtbiJcvIaT5i
V+2G8S17wtMrx73RTqO1HBZs9XwqdiwLwBiwOQ4Hz1pGRsTFuA1GsP4c7p96oxn9
e84ER2edRWKOLL8cw/3n/D0r/AVtLyFzvniMQP5ubdVSOCsThTls0Auc52Cb/Yab
s9LPc4ps324cqybXby/lHvQ/zpv2VLU/PujwXIwB4l3U4w9udGXK47AQVuk+V6Nk
Iz8/8taKwjcpsQ9XzArF12eYrQWZYTiPy+weTJ25ynTz4yfT+c64dZsXtip8LaMa
Z/3G+ngzVKMIaYRszHq77f1B+AqjKRZ6AoTaQ1DuG/9EWagykhA0QKqw/ln0fyZP
4we7InZrVjL4Yk5v0JVHLnzFSlvJDkKr2nJCVutpuDAx1xzvkbzImso78nnZKSFi
d0I+CMT9Z899lKo/omz6Zn1gRYYrhcyuuC60sEVspEDg7FTL0nFAoF0Dx7eANAvb
Gf6fDPRxPT87YZgWIYZh+CtYdXSt1yTVUb6oqlR4065Tl2hBLkR6oYzUtp2zxkFo
QSWS8D59KOf3+qDpvQI7mMISbxqjmCbUKVy5HlZiL9WszZCUYqhQayn1Hyb0N5vg
dtNSIZDLeLqRDcTXxQkBraDPvm6mwfsmx/F/ggNFiJr2/lkBG905ESui5r0i0Tm4
AxS8Oo4MCpu09SwJHg6X7QkHcbtsN5KsrlzA2squ/Ads/PpTbqqjwqa3xJxk60Bg
dn/O2qugmh5IHywb4OJBXUSoIq2Tm2aqp3GUkP7vzvR6iGNbfPRukMsxetp0fQqt
5q9pTez2zs6/vRo9LphrPYsccA/3Kp619W5mQ+IMRZX9E23sH5GnzfwuRSZ6N8v+
MuXDWe5RBkienUnBk4O2QjjB+lm7BZdA5pEuYsaKopV5W4ZcxxGlWrP0ghemtvXb
TUkoZzeW70BMAeJM5o6QHM3tAgl2cZRyUUGBVEao/Zif7ZTO8XimCXGLLZOA9Tjd
EBBL+vFfrUDsF0GgqjqcZIANzqDdxBytUvG5GAh/HDhNm6kkwb+oQsO/XHfNrl11
El0EbGMhvZH5tnf4ncNumcH7E4cn6lvcOPq1lWWSMDXmMAvl4RkBs0EYXshbdCCd
V+p8JFxE+QXAVySS4l8Ph8yQ9m+AZLFazHoEjVBW4gWs8yOWTaiA+N32B/muQu2J
JL0ovQKW86KvH2fOxWUC0r8XQHMJwwkMDouMlD52aL0ZPhy1Iha6i9Fm4FOh0kJG
crP0AC6z1mfiUojbFUv9Ewbws43PgnCc5Gqy9i37SHisYF0yeWKObYlVCZL3QMrw
UxzSrtgHMBvuPoMQDDYR3ygUX2zcJmDoxjHr64VWbpSQr6ySXNgCDfW/xO4m6EbC
dLNEaj+nsio30K3SWj9W0LPJ9yqWB+h2lWwiHiLSGiSwd20Q+ey4W4tZf1n6sxv1
k9mAYAbr5ddHvurikZqwgd7RKSi7ri/usg6JenjaViuAiO3bKPdxIRW3m3mU0F2e
HgOLUNtXlDU9LvO3lj5HT8NewVOvvBOA2/CFrD3cTBO7sznh/abHCBG8qMMcOIM8
7VssiOS0+yMz27zS5Q5KpiaqHQnopSVDgcfL7TdiUwKKsKbtVGZBzfCSIISWD9KE
b7D2WyOiG3ipQOlLM3ScrJU/JUUvAMgGnhtilDsZxR7Th1gi/Z60Hze5bN/FsjMW
BO2wSWikbwYnIqRO2zqvvtjGZizcfp1LcTxdGh+xP+FW3k0XU4OjuY8KcW7UaJ1W
N8byQOeO1ecKlobL3/VuQ2NwtDsWRooM0mlGkXW77Y/MHZdS9PuJa1NyogI9WFss
kpI0dgArePHrMp5v4ssk0lGCQkoWv++JF8/aaUz8HsaJ9h2dcNsSljQnwNqjfNh1
T3p822ueeF+bcZ6Ok1mJi0nK1EFtr/gD2oFn7qppwAfa+hBfIDGpnMh34cuUVfql
F7oE6+fba2UeYLV7t0CCPb2YusM0tA8jRdzuEaohYMMVs1p2/yCLDDESACpn8YlH
CfFLqlr1EnntcQ9/ppVzQphYoUrmeRQyKw6VsADpiqwWzK5/O5pgkWayU5R7UKnX
W4HY9k2G5rYY8qRmzri6QfhSH+OPhmqZ0DQTKnolHAfygI8qofNgN1w/pJd+U/OI
iWiaRvcpYD+JqBREzW58lgW0YZlrXwWuLb39lD8n2RQD9g9uF0KVmWZ/JDNj+ktK
6WUKp2lFPtjo+3m6O/FibBsLWeBE4ufiELKYFQ68myrf3iJu2nN9vj61Is1c6tZ4
5KCfEmS7yVLF5I27zwFf8IfGGdywueRPfjBH6+cG36QPkjN4e9/q64G7h/n2wm1x
xKjUs5U3ONBu3axJtss44ogn5ACkc1hWk26FDe9lbxmCZmVpmhonbNACxehmpDC3
7BnAQiiL+uHcL6Uxsk3Q6xOupcR8hBg2xZFM0mL+eGwrvHax4eRlhyYoNMK2R7dH
7DpP8E9spuncZC0+XN8VVXuBdGRZwvhxIfiYorI4rlaG8Lvi/gYsH+q1UMHgt770
43fJMD8CpS24JyDQrf6bu6Mo+MCdhFQY4tPnnxidtlI0D6vnLlkmu91pKvK0mSrG
UeL7Azujp+cf0Wjfug6oHb25QQCWif3HbZ1FKNWEzVYmZHCe/juM+CiErG4mcKn5
Rqg7z5R7gZcNMy5S2EY6ZYVFP0s8TTsLp5ZNOrdK9TH2/E7Y7940FVSOoSjnD0Rj
SYiNegah4gz+V3U4NyY3nZT4ocbqaMFLPaOGF2fq12zKMZ07NOLBXpto536QrwsK
FUeMCCUJBEPQHUQ3F6iZNEUOrYtA2Br9DyAv6j7Rz/5jNubjKCkioSsSPuy3c1wJ
5SYPXKU9oASNM7OqczBbNLoUTYUSuQWeFtokNWjnI2vPpX7212MePBeFVHtqIHv1
DctckidxgmAWC/4yAPLSdNuzohlC3yKqL+2HClYoy4AVwCjQxgaAQ63dpMAJnSKM
oj70e/wRS1o1QQjzbzqTakMy7q+SyiFcjBT7W7qY2YHMztSfYcNHeR1tXaAESNXW
MIvhEzioI/KruBb97+amM7cBrfNN3EpgQsBGG29NV2mueq6THQbrL3G7FS9+iE8N
wDb3JTcVH3MwudJbjDtsiVJ5OXGolSe/hwYNukejcfpSeLqmT7aU6CkFAQ+w0cEI
noru5PS66dCeRvKw7XFs1Q8cY+ytkJLcCnhZ++5/XwjkA8dkmtDzFWhHKqF7qrai
asSf2WE3uDtLga14gtGe1QrW9qqo64F/KreqlBqFoxZIiJ77cFUYuGxkVJfUmSlR
jcfraF4Yp1Ik7MTuD9cNhmM9IJ8GTuOTpt1DnjT2ey3OotAgWibM4LOyBL6/OZfU
Zl5NU7sXzzXsBuGIZuLQyjsKcHeKp5b+3T6GcxVNgGGvBgH1S5S1x+jjFkj/elV2
nOYrtuF4bpXVr2QbtuWp5F+HHnHLPqIKmuMF/HQl15BSX1dLfeTqMFv5+WR3UQw7
ttNZr5a5nl+pw5Mw4djLLjVc5cx2dBmyI/yt/Zy3eCsMs/zTfD3RrMeboyNdRabX
3lFhl10vJCK08HXiu3s92oUrWQWU46wtuwXkM9tbri0M9ymb0N7yaRUoBaTJgdS4
k6AhhxKP+KOapZIE6DaNdI9ntZETprl1i8ygNh05SG9uA2OXfxXGu+CZiYgBL+uo
8uCSbGUhfhE8yav1L5C77DB6X0wQvfTnwrDYS42OwvWzA9vJcLAkq1tu7BU3AK86
xc7Ck/gsrvzO2cjrA3wKihSOLkYe8+rw4SR8Do/MBlH/jeh+W6V1XmoTWOCcNbaB
xaOzVUWxQKzvzID+nwk+PkfWcaCS/p1EPKoiUJ2cOwEUZkN1jJhsnn6DPE3byUXF
TyEz7XTFwOm58dRwYIXTr7pDoUX3IGDQCzUJexijuxhZzv1t4Qtm9Ymg52DH3Ahv
U8S1nIIP4djBt67c99nFQFECvUTtdFu2rMfNWuzq4vQMVdywH8k8asidmzIgky8v
CEUxkqvipg5uAxaNAevOC/+Rk8lQYnmBx71v1c5jiVnkwuX0ulmANvwigPc0PepD
rrbrc+eKWbWZYl+ffc7214d+iWP5lV5VvzV9PYXpQXKcsZFUZL2n406zpZI5enP0
kcW3FXXXQwXbbQvOnqCLDnGvVa2LfjWsEkGW1FReUDCBs2gQQR+CBXxP2BC9NNdK
YLT7FnjK5x0o0HVPJ31c+9YXuV9gAsXwe/FKqyY/VTZ2S9TGQyXInmITwRPqzUmW
R35aIRsJbORTa3wbOEBGb0ba4JxbDVAHGvbDrd8T7qs26LHbUGDXyKva+XODqq9X
SJj51v7/Eetwd1THNqmpkNikeJ5yfBZXodUhHeJx5riVzuqQNIz0lhwNvCAwwe2I
0+NgZYKcLBB0PNidjQ0XQzGp/0l9COS1YTtvnL3FIkhQxYSEbD4j1GBDFRBQZyos
fc9R6e1V4TB7rhHb81vnmZXA5oQ7yeatc6zsQVA35NjEiL24kz0zeJIdoojGNXmp
myaLsehm9IMZLTwo5jim+yTkvF5QVZJBdisCKgNzW64IEMAE6auYVsHY9opGpOOs
ESeVicAMWx35sDqzf+0w/CvuCmEpXQOV1DUGO8f1adgeTsIx9IY7zVyY0H2mCmAP
n/pBWPbErfbCKySJYxzrJK/IxW0GMerDu/QDJYta/lE1xkg6Y6KjV216X+DvjCXN
t2+MMwyQHDAF9LqON9iT+shcU24LvtYzNTFVb3BXYuxff6XnxiLEMtqcSpJ59dNe
CMMpnnsCEyeHi+Qe4bGeUFZ/oOrhdA/GfeM8qOwHf2go/ykwVMXnMHFT4P41wvHe
UK33BFEDjGyigYaU22XN1z6ax45kIQ7KqCxyYUmgqKjUa+xGYFeCgxtFtWPpLkAg
0BDv8e3N2TKXzxVtz+RjLtHcF8vODVtQTwU7qqrEqxTn76aKh7YaeDjQVixFvsKz
KGoj1iKQmd9mkBfPSCvX+TdUWt7rX6sr0LezfzMa6Buck9YduKxXxnHVxInSB2IQ
lK/BGInJ+n8HqERcXQ2iyRwbQXrk7/4Cpy0VHZzIZqCZoEx+jAhJnm9bcDZewQIA
cZN01iDoXtlw12bqmwA3rHIepsBjzx9GE/ItduRMaUZaj3SN6vHthM3PBFgNEppt
dMKt+5BWII6gmJ1fZ2PI1XC4PuVx4AhGVcf3GuxmQ52cUiHrvi7XKd2YvMUlNk4m
sIKJOxkk2CgwqdYWf+UuXRWjAn+7LpsPAfVZc+HBThUP6LcnbM2OnhckbrJKYr/J
yYVkn9UnLx0se7Ezq2qEuvW0Z2hvZ4FeroI5avAZpeMeTixwh+vMEVNgQNBzTF/I
A/eCYnK5YarpRmdRvfJc8A==
`protect end_protected