`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
ddtXksX2+yylW5zu6QL2Lhnb2d1sD00763mmSITNX595NcHTEkwn0zB1Dry37fOW
FufOhVzEJp80NC5qZ/+F0Vk7Ik02dIR0elf3clrjeJRK85K4e3Hoo4xn7YbFUIms
l/8VZSb14+JVGURjfswrIyCUotIzlzVYZ6gzoZwDXIi5gQIBf/gI+KxNXPaKV+PQ
Ufys/12rjO6aI/pPlqSm0hCvftmBcnezN2hk1UeXgOIuKZnogjOsf0iJVX2aOOWE
6pD/psybjbnsNB6kH5uFTA5frkzIzkzl5d9+YDm9OyC+k84E83I/7/j+rk4L2dah
QJOvksSIzN867/4Qt8qYTQ==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="MvBXkzurAa5VTw+1JJ70nePUfoQXBvZOku/SMmg4TwQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
oRtzZL4VJ4iwysPsC8SXYCzXS8Fw2gtZTOskLcDV+1B9Nzn1zTyNtlo6lNICRmmK
ZRVu2BmCc2G+fmzynYlNTnSa7C0Cuel6FYpxCBlOuk3OF2tzAmLAuDyOH3Z1Yjzk
a0aHuoCdIRKv7BrZCdALt03JeUmXKPdOmIlkVGFl8yw=
`protect rights_digest_method = "sha256"
`protect end_toolblock="Jn9CQpRhJt4rnzZPRk+dOpzAubz7omckX1MrFd4p81o="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 24720 )
`protect data_block
gD6l00tciPUa6pDNTk/+t0OO0nC/UTtBwLB41d4inuAUA3i/ALrNyoJVcBnAmEQW
ptbcNp5fxEUJjnOxnedyZEuEBxWRieZFQnkRdF269oMDC76fAAWMgSVbdZCkMybD
/6NiYKNNW01fGt7O0DxKciEzTxUSlBIqSejgiW98FatvRavmUPyaM87Q7f6TdjvO
mMNUWvaPeqdq+iHxyXnrnjlk6FfxTVpkA9fxWOpEGq2RWd93t8J7Hjk/HIiIIuM3
F/rafZUKYWjf9MpukrFr74CV545PKS8YcAqeGl8Ej58eKgVbJhP4xXlY8wkaiZHn
5kMWllB+ZFyQbV1ijfik1XI3q7AiQg5pHaXPHSvWxtITNc2fKJv+xSb5t+VpWxhI
6BRRUIypbZPvxD67hJ9U/qCiSV1DixK4cMfVwLtNmZCtP3ZNnq/ERXR7QAIWl5SC
wYlGAhrshWYNcBI/H4rbz+lsfi40XvSh11IeBxOLiKEhiIY2u8fIX6q4CpnWjgUQ
l5sOp5RXKt0DLk59u7Tq43MUlMEo2zmn7H92A6AkWKKwiqzgvY6xN+/AQSMYbThu
/VqKDsPCtSqK21542gmG53LcCE/fsB3ADOchMD03FZrkNDx9snB1stbzWRxzQ+pn
tdCjbFRNeRINgrv722Ds9d5wjJVOJQLVc/XxquWKslUXUenEsNwvVN/YHhgfP4bY
+Qcjf9oA7Qjsj6gGiY1UUZDWgS40cT1/xzz5nU/DErJi1MXe01ONyF5RP0/pu2im
mGqsTAZw/bbpw4yrmy/RBL9Jpw5k83e/VXmD//XAWAhNPjcZby3qIT4WUNeAzNeB
Ns+GPSVfPpuIPLyt2RQppcTVtDftaVCBrydsczdf4R56pw7Azh7pn1rePJ5+a28V
YN0x+jLmVDUWq63fmztWjtOd2et5AZqCilxpeeOvnstK1bD17NO6FGIqaW+7Gb9t
L7Dciejqe+vuerJ/N0FJEBzPwU41sYS9dxSWD1KNvpkJ6i875Ni1j8D1O4ek+mL5
P6YH6oDVpIPKwGB1NO8R7ZsA65bYA8jobEhfdviBwWXwLRouW9QJDAIDqxZX7v10
Ia/yESnM0RXc9rIKrkZrVdbwSr2m5Iqh0m/HFcl95L9uo0n11PFn0wB+PCC+3N8Q
nfpd4Vl7hOAHCuGc1odEBL3/+bnyUCbhcJJRggarTh/t/tt0P0PtA/9H8/P8mcPW
CppKksFZkdOmKi8blGXLoR8Li0W0vSjdi4RmAA5MdilumRQHoAGVM2oupoTTCZ5l
4ZNJIr8ygZhmfioQfITBoVkj2rzKZMHP7xcUkNMUyMPTnX2nTgrfcWBet9ju8IWH
bSBGQDAkk0X2GOIHhWYM9+He+2FasiL0avOqSfDgBBuoszfiWxrSQYA1j6MXU1jH
AN6BcDGfCVeAy1eFTbkxsdkSvSN8vxrdsfJ4o8IvQykI+oHUlgSG73yqV+67BvKD
4Kch+CnLqVGQh8YX+il00clXtchf2lyKezkP079MtecxW/EYHh+yPaPcNxkVwTcH
T9uNSC3UzvEoRSkMA6alIOFZt92jVF8gecipb7AnhUnhhEvr5owt+ECwD1Gcr6xy
IqCF/dGL7bCq7k5x6j53nURfwKtOpdDi8CdUsHIku2kmCZLyh/DtoXbekFoaP9f5
9n43uTULKR42OzDGA7Ru6g5jld+f6g7kAIcxUKkL0VIlRO0R1BavYSXTBM1awRpU
Pw3+f0iV4s+NVo6JIBkEuXqFo0nkZpUxVG8biPMbO2bZro3WlKO0pTefv3FjZyH6
GyGtwE6EA+Bmpu0Are6mhb4ji0Dl4L6+OfwgLUEQwXlJDF4nedha6+BAH0mOrvx1
oBTRx225oCg4h3Oyatr+7RhtD6qQBPXxZEpNfxibgRdVLjwxifJteWHizhMJRfLl
DN4UZ32ZeumRDAFPZAxHaMZdi98T3smz2t+FaMhhq6sqT4/kXsStnbd+0SYS0PMY
pITquf4YFo2byG9PkoFJNo0Beag5e2cOFtpgAwpXzgM04fWBxa6ikyN7394TcZ31
/8zwPvwY5VjNCF7Rphdysy4K5dk+QoKXZsbb2a0Y7hqE29vX4ga03mB9PXWyw/eA
TGqtZN4fCG4/p/fIQ8m3WxFWwm/Nyb6RR7g05GPy2ioMQD62lSWX1qoBvMRnAjyc
B+psrHcGkABFJ4GcmNUHqvZi+W/hVs0ijevDqOdXjkHf5l/2TutpOCN4ba+YtQgd
pQpj9MmRpmNjtNDx58sxLvxkzF9eqkpPOj924dMsRvMnWNNV9hOmKLWbOFs1Enzw
lT8+Pxyh1Nv64eaanmJntVWLVUFqIShJlF/ccJTO/A7YovaYCqtAb3DoO9svukws
n9m7CX+ozQTc0B6fcHIY8W4w+r/t/JOl6iUuAMhRsnLbkUo9137bTUmyNQMUpXn2
cl0aNpJlqfr8kmc0IWMb8FUkhorpL3rgYdhk71Z/jUFcR9fBu0hyIbshLL0VjCN1
8PsryVU33cl2/dvco1PSHIocX+0DEs9G5/oIy2p75QcRsnxk6hY1RmDX/aYXWWij
rBDhTnozNk/DFNI4W6rW7NH5W2anV2nVlQOgLhubwQZu8/kQQE/5hzVQfEPYoV8C
V/sVY9ThQEtv7VwH10ZNCq8yK6GW0/IzPrX6BNTShlHPJ6ZOMdMR7ZVmPSJ8D7W1
bM9jDkGFjqNjcrDjqUZO46iN78Tkak8nwBGm5Y+axkF2xJ9rSvxlg7qFISTayz4l
a5CualBmY4BCL4M21af7aBN9Vi4sHR446wzYqhkQ4HVeHoOPts57pnC/Mu3geHiV
ggYO9XQn3jpKHlCqBNdAhCfnwuCMq+4r+tfQBr2x2uU9A/XTOAdC6ogBadhPlnPk
ttlbwt09wWTD1ZYHcoWqkzLO88++SmVfV5n/MilGR31OYlkT5E4hyAiPqkBBkyQo
SVhzPN7GQrAm/4WSm7STihxIZ+TI1bL70UOq4mVXX6+uQTmpsHY3T36ZEVXQcxOz
CM5mzo9NaWlo9RQOIfzkZwYcfh3FmfMCPVvEc6Rhm5aDa3ICb9U1i+zytfnBHs8t
0kYTr8JCWmQvn/vQDBbbSxD8aeDrjKonbCWwqqAGgd98E01yvy5aueMVGz9dD41w
QLWPpPTvZ1E8WpVRGcDn3zMddQ+6HzgHOQViXX0/iYLdurtVAu+lBRRU7jIKdnFV
krI5w2m3vcLJwYClckkEVe6tm3D2brXWLoOhMNqTQzFFsN00yeF5vxCuVp0qOUXR
e7hJQpYD9Of8OAEnlsOO6ZBGezkxP0fhP3F7W2Qt1v+nTD/EoqUYk/YgGNzdII4S
n1X4aBr0+gW9EkTyGGOwqsKhqkzyo5XlPcZftauQcbBQk2P64YeYf/wMjgmR9oBH
cq/0M3QOJEQ/hKOgPEMtouH9sJBhn09hNT+yQE/5mqlrPC6cfyXCwx7qiJLHm4t6
BuIiWN/3Slvd8yZMSym8/ejiM1r9JgM+Y79QZqwDg4+GXdYhHeej5TNXRoRGqG/F
BuSoPYVbDldYVcm3sAjHfBfy+HZ5qgZnVT3TflBxP4m4y7DrM7nUgQH2xQ6w4gl7
xrLcEbX2QKDAZonHlQGgr6XdSCAbfmzVea4tHMqe4D9fxojrm2Pgs6pjANaJzxNx
aFDGgxlFhKjVIsJhQBo3AEcJ2fVEEC4Dbo3DQ0aMPCtO9KuKYPU3cS6wYUljN0fj
P0sF5JhupHq+Zo9B2v2GMQIMb2rNyWVOTIPZmDE1g8E0lvNiSakcuyDFyQDsNXeM
NBhuqzNnU2dTUnn+AmS82YDPL96KHaF8YsYMJLfqgcAEbTlYk81JlqSeqm2m+xY1
uJ/W+yVS4rc8fc8B8Q8tXWrUWSMF0/Vuc04IR4UH2FBiBIi4ULeawz946oOD8uTC
JLBGWx/w5nk91PvFGCXjQx1Hy42/qzFI0Gj7J4ltmPLUpSYL0ut+PD9XRp53vfB3
aQqqtuZPwbrCuWCLYDpzdR6ZAPohIEcHlERpTrnq+l1n3P1rlwUidDQExeBSaSXZ
fuzPHIvg4WRbn7G/c2HzW4BMkg1NOk1pKdjmjBqn5dbUh+VxXfVw9rrUsd45YWG8
lyzI7TLw926F71I5XS7cNTCB10t+i/PHJD6d+5Yz5VcWhkgRzZe2iFBvtXPlzKxa
zYqy2DjrjKmry5/Aa65mobUicwz91rm2WLVjg0cHYZ2KkkRFC1ladgH6vszFLPF7
UG5qFu5kwcOT1R4wyngsoX3emLyyc8p4zYGpb6AP2EGmQPh7O6F4DkwA7CNyCOq2
+zn6IHqh4uLizm9hlD8w9Mff6XTeg/EWPDCOuLfWlIz/2dmZLiI2DaNMTLMGEkjG
PENkOJrEfGGAdq0QMeLFKw7CVPDtikIpQRVBA4TOg6nASkeDbgDo8IR8u9lbvFCU
IaN3xO3xazoZ53YL8xcvgL3oe7AQOORMJGzZr/9Rg/wTEUo9MKYMKTgPXWL8NRKu
8g1LXs3MbR3YZiBf+LV3U1Th8zMQIpOdMA7Sn+xE3s0TTjsFnN6+lk0Jkbh3wiqU
2yOACoKiw+jcD4wqqMFcFUozJTNmlOdGwGjfA2oAHXMCzjqG8uwLs6DRIb1NjODR
eOv6xtEo+rkCjD1TINP+VxbL+UZEyYVt6H+ADtxygstdXVV0cwYRwgLqA615b5Ws
K0STzEvi4T/RhrEiKw2gUmHE5JfX/npGbfZqIQ2lqkekyeDIRLD9+Ptw3uW4SXk7
r9TrdwHSbVnnQJBvcPFXzzCFDzOl9kYNqBK2Cq8WOKPJ6WmylVI96gPIIdob7M2l
YOO7WeJdAtAGDuDthrmftDmXdKvinSbFP7S93mVKdNL0OwQWi2H7ssh78GHNUT+0
Vjo80t9XiG47U2TBami6+WvojXtQ/upJ4VbkB+Yr+HqJUSqq1M5iV2Idu+3G95D/
j5RvFMDdzyxrA1A1WSY8Ymjr3zAskKv9q02V4i4jd3DU5QDVHPcGuVS+PDmJaiJN
UKQQCOQAD0ZuQjYPFpmtjjdgXA+vqjHoRZHRus2s/S38yCotaLpkZfECJgYyrGSc
09o4NfwHi4wBPibDmhHJWG/kkpUEMdIgwhjHraKOP6R95gejH1km1HrbSKyEQgb3
VS8j2RnPDR29GE7f4Ul02MnRr9xoKBC+sFnYSYQh3pdKtRc7l/uNmnQIi8sApVf0
guMOqtf9U7MuVomjNm0OtMM38q+vPD17iNpP+3xdW+zwciqphJUnQrTJAnaz+lSy
vAYBj069UiJ1wKL+OgQ6QYSbT35B+TWLYg6pSXrWCOzOhKIZZ1MpSDTmlJGzwuIo
MI2cqIkiCQrU7pmCs4kusL1YXIN40TmrGKoY6DhOJPYxqd12wRHxvvfky9H1XRY6
TE9olZlL1qw60zguaNuUL/g5LMiESG9AYjZ6PJGDRjurHA7+SzW9qO3VwOoUIcbz
3mQUbLTzClzEOopJJplkdgzs7sDTgtt0OS5RK4xomf6nV5E5YlzKhJffkyYZP7Ld
XUXYZnJJrWRhGCm9qnAKgwlv6r71V5jYFhou8KRiS9+LZeY84a8wcND+lu9Vgtb9
3qbe7tmDpW1yUv9E0vI9UMFsUwpJVV7ak7DkKJOneGzs3Je/1NQ2A69/Kd48qj4K
jRKhSSCT2E79IKnKpLUr72dFhDqRrIxgotcGd7M3fsufNY9lgT+xm+OfGQCUUpO1
iIowF+XeFdrPqBsYIP5oMBl/HRNcTnKNfP2vNSoC1R3DEL+BQNdNnUV84J4q7XKD
9kptaMNRjhLMAyE0vn04/EQHlAezXyQrhNUI7FYXjrgp8ceTVL0bFooiuQ0Lydop
pxiP4ezwMQD3e1GKmu2ko8s8AmvGqf8oNh1kGifTJUHeCvNdldP7WtSvI3C1JnhJ
DHXuKidcR2CVNAHflRb9gcVbVztYbGYHpATIuwKfUJ0lH7YTaffOSl0remS7DF84
u01gyn0zs5KoELt4XkZOAhsZOueIgwDyFC8omPlnDagYw7pT9fzNzeh78TKHBUic
JhaWZh1n0MhV9/IA2JvUMdbTUVkvkndHQDLZk6ttZwDdrQPIMpbkl5fWSoNgkM7g
YfnLEZoHhvYrE1sTVKPPEYC4fy8w/g1yRpi8mbCyMmMINTQDfRTjbZdhbI8Blek6
ubHc/d81aiWs1/K1rEgMu/+/id8TU/i63UZutV/gaP1W73l4yCkANLBrWH9yP6uM
b8SzhXO0ie3chFM87xUy2YOUBq4Uy4Wq5Qry5xOr+2m1zm1Ur18UZzJOib8hWenf
YjL8iaRcPNLDeR0TWIe8h0Y/EMBh0b11t993r8J9FQuIxeXB2KzMi0hpreIJ3MX3
jUausE+JwloXbWp8D1NpNqfSVoQ2GTuCiUAdGIxMwIA/MoJYKxWufme7EaFwlS6C
uJtH2/J0E4Z9InqXN5yPsUIW1LsPgO4HN5BjQzsc5G4C9RqBJQTnnJBE0e7/b82Q
KFsymzrfUwWkhdpTJZHZgwKhP4heuhDv40QYziLgEIkV9f66efZaMbdQa+MstqZt
yLvgXe3D9SIeIZyiimRw+1aiV83gqtza52VJTw5pmBAqt6PvzdpjWpWWvH5CQUS/
eOejKRCW4yuLN52Ivstmd7UN4jnkFvgwNQ0m3Pf20GKdtHlGNzGNa9B1JALB3S3e
2e1G8aexnCUwzSVdE595Ub2zoDlneYT/KepBdVwAHBPWgol9pMnHwZpzVtcgL8jL
pz7HX0OEitr84a4ogG1RoTk1ev5IsgxWFLQ2giHK1t6CgfnS+cwzs8R0QfplLxEh
yMRK6rI0ApIk2HDeDv4hQqd5j59k5SQ8gMZwUBk3grrD+FaMrXanF6CKUsSH5wBc
/F71uiwdFaTmQKhJjHPpzoFayCxdJnbAxScLBMWN6QHGdMeef3OAXGsgwFkuh02Z
2c8iJKZIwum0UV0v8u1rsMLqxybF9XdhMjNz+jWQajrACtihltoPsYBVIl+xaKER
gLGjHb+zDb1C2YPMkyRt3VVzRPbLHHiVF+j3nP7sPOcSC7INFs+rlTboip0BzhWn
b8w8BWbEdaY3m5MCUihwan+/dvN5ce/a7u/BzNsPvhADVT7EnvBOd89LNEB6C2rY
AghRkc0R7Mtu6KkEHknED0dpWYiEKYErHzLpad0l8W9pAb+tL50jQB93GsTL9Mcm
YAEGvkzBfLJpGD/s7MXS5AKIQQ6L36WG6vU1lOStOiJxr/XKKOTF3Q69UGiRuP/m
toDwAflJ393pg8tcNpDAf2S/SVovaJWUIFd9f4PpLPaa8FftGZngQcgYHxOKawSu
kqw71EGy6x/qAH/ziAadLYg2//ydG3O7S8TlkWpAlsl1BufuSKpcE/Vq9cAPm/af
udsopAJhLa4rTnBQfka5ib2V5TMN8hREZywmT4Vkx+PE3rdQCAAcswRCHed3vazi
8MYe6a1Kjbyw/K9dChELG5UDPVvskiZCh7/3poPTn/R66vOEzCNg9rdU1scZOuiQ
xsZRfbl+lezTt+2v3HHMvhzFV9/uozpgcP5llPWbtGcVZK1BrWwAUtsKXrgDEJNr
hIT0krkWiLtUyeYMtujN9b6H8zS0vSHo5jAObwkzMseRMBaPuA7aKaUVgULywPBI
SmX/8K/i9UBPVh/sUttNCkRp9ieU2MD7YIQ+oeUjaWUSUz/gpOhlwZq5McYfRehm
/lospXmvD43GSiqqlFWsKKKWstLiOYZPua7zQyprN+cHpJY4fi5RgkDctiyFIEbi
LD/vUFPHRY6e6VH7K6aQBPrBuVc3DcWydwQqNDEGzDRLpgx8MhQ/vpwXVUoDc+dO
nUcQCI5TQlmYAoBtELDvxUd1T0dkPZb3RfxkoMTYeI0T29EINBa1M5PZ/b6sNGuU
XxGIb82cxZID1owrZAWbKZ5j4dmrGTBlDHegzlet0gBXr4lflEmqlWO5zixnoUY/
PWM2rc29/ARAHgq8hcroPMWOg953vCZvlgwARfb7KykX7jjL0//5IZwi1fWNkXzI
ywVtJnLOZtFXMoZWB6bScpCtZVceMWRdPgDvZWaqN1IKK7zE/cuweSwDCp8hQ06o
wi1c+RJq+SPJZaNRUf2Pv1a1EYwo5qj/THyEttjl8fe1yhyLIiGNeoSVHBJO7HcI
wjdsdULN7pLFpVHLCm8Wjm5Ib6oQHEMUDexGlzXpl1UwuRuekU2YLXhr6Q/35ztG
iuUz95PtScBFmbo2rKa67/dApMgKxvJi9jb/lYWL+kP8MYSJy14bwn/RiPNwzsT/
+WwLT8pn2dyjRM2ecq2fhpLr3wzrip8iOafa49swxmasMMiMCDRRQaQAKbGKYlVv
uZ9dsQRuhfBRACPdmxKR5WR5nLD+uKE35j1bjT1Gn1P928hHJC95PwWqvULDXJT0
lmRqkBWfyBaRkgONAKywYtSIaIpMooSfep2FQgP5RqlFBgfrL1vMre0ZkkaPGuWC
xNKVnxVm6GKiJt7Yl2yfF3Azn3oQxIeQOvVAyoIZHdwQAgDGJmN2EktVt+7iHIUk
86lL+Dyti+ka6JqVyT8+Tl7p/EFrsjxP+roSSmlAjsFY85WxlYkbGGiJ0p0PeVdX
m4F+pq2AT8juQEtZxn9DkOLIb7eeuDktP5eSdfV02umtX6ZfhwyzCDoEUgPLmjyc
GKsk0qe0cVMJQNqFZpdlpXy3iApyPcr3Wb7ysXs7t7I8m6Q+brMb2kRF/qGXgaU5
jPgBoOYr5r3o2MZq9Y9+vW//yKVESpxddnDe2fL27xQRbh/Y7ctqY4n6UYlfjn1h
a2FJApNihaH9pp9R4REWtm887wz1M5RvrrUUWEPxKZEOEEzqG6uzOB6KsPqP5ODf
ca5YmjxUKnPqoJl3OxhH3Z6o0NkUjjw9SUWss7N5cAXWb/1QW7oy3pohb7imDQCb
loxLN4zfrawysoHD3xVIYNanmJrm0ceXBtFzX9FHqxDc09eE4gYk4i2l5qiMUSjd
WVFKnyO2cMJ7OMP7zSY81rFnQ+h7c046TYSjgdjZozO2Yvp0qedkkHJh4O3JbYJ8
Kfl2PF1qAC93Y/aPtjZsICgmegkYJsRMS0ltK/NBzeshpEMxJVD/jSk9LLO08FFw
BjlCcsNp9jaMo4VBhH1d38IGLpzyRJSf+KSrIaL6jKCVP/nmnuEQadZMdinNak4q
CDmOsyCkMQUcMFcw3n2PtLaqgSTdmIXLdI6AELsLckLAWJ7uMBdD1e0voL8zOHlb
thC6B7qjwVQJ4nPpOlQ7hFL9B0hipbGgaudB4+nFr/mvYdIEml9rTdZ/w/BX5Dsp
WOvR2fbq9m86BmN4BUxydtM+NQJRQfoF8fmd77crOZz45U6hr3r+8Dp7N9i0KO7E
X7jVgQVJ7v3M2PTvj8HtJtZZJQCyI1iIITXPLarUucfe9jPzhBUdiM00hCLuKdim
6XmjRooP1qgkjBdbXhxIjCQGVxGIOzsQ2nFzCRrkLdnitz1PRGvR7TAoug5Kqk7T
GRGRdX9GZjNTN8VwvQUy+gSIm9CbKESwjW+iJdZQMQCyCWyAD3VUpYgrkTelR70O
T1wxauwoqDKnZ14f2gOVXs2w/KhrrfIVTT3vBp9HMi39EyQjfcZMhXuCX1vJqjfT
xXrcS7I0Si0fXYoH6hXNPympV49+FEDGJOofL9WMMFVIOlwoiGZgse1cfNKEYSJF
koP3qaDbbqSk3ufJcgkWGYUHfdinAxAWTMUFXnYSV4/qykKyabScktxFjdLxk1PU
FQTaQvwnfWnd6WbLf5FhDa0Z9XHZt1+RvSOt/7zaRVYgwcLRd3eff3WZvjaBUar6
gwwN2KV9YhXZSpx8rK1aN01cqGi6i4JT4IpHw7kZpu7hrtKmVem6dFF8ZDLU1FMa
bu5fsVy45mFmSqjkwkGO+LQDNUz2HoLO4zf7BpzhkmM53apOm4WqJo9jq8kbVk9W
+cz1w8Q6m4mWdXCuMu0bngLsxo5c/Ryo0BKO3HqVQE/V2loUiYOxCBk4ZANUBel7
xdAp3NOZ/RPq4nr4jghIzzCN+7Tgbigoi5hx7JD6OVvmqzQDndGQgMPrJZD107tt
hskJmsHQfSw08HDdmEkM5IHegYzhxciaCbSzMjB5kxQLV9OYmPBgA9BpSQAoSU1Q
wjf1RO6d+pjvwefMihh511XieCX55hbTiyVdHkQ+mC/Cy2e0bm+YYcq8oRlaCSYb
66uZa0YZOQZH94TxRMTLIkMx2ucNqUWFx5SdCFHYzvtODxduEyCZMQea4bmg5nFd
LUPw5ekkYWwJjdiwNzuXwnt4vqvPACPlhx++uOOuM05uAmEPEWUvKdYUGv9XSPe7
rz0C6be8Z38YvKDgBJWUzjqhpp0xMzlOKTZj47xKTcMMcTozVibpf5xSlEfnC7TX
fSzAlXq5woTpzGrIETZ9xkVtywuZiKkH5sD2CLZCShh3xmB/SZCyxmrWX/rZ9NxO
GSgaQRwMWXXpspu3PTDWyxCcp2UJ80fDp9E+6E0JCSX4qT+LveX+tYlPGMUFe1PF
ClZa8oLaQ6E2ybHlxCpgi2F7iBOFe9tCpidxlaHgA7fu3JBHV0jtrhYxco3nAPUT
vSHPHUSP64wmpxuDq3LQ9l5dHN9hgqBzcl4c2h9kHiVfpV6BWVDV0irj/be+JWKW
0bpla1sRV3XSJq+j4Y1u3WftL0Kduex+eu8Miux5uwOm1FnOsfmkFhrLaaLefzxs
/lPxXLDtd7IJS3zw7VuzdBzxcc5fD+Mg39xWdsPG+IIMJo71+t/s+wo6MMi/rhWj
IxeF0rvSDH/MvauOimneRxb2USzRVOT6mLNOigG4US29Si2ZH7rCsI+u2I6YkLJv
cE1erWgsy9mso+oflLNnZBpRx6duaGcJIetskmOmG33Fg20xOiWeuaDkhkMcMQXu
8i2RyCnkenHE6E8MPRAK+MZienNlwQWH/8WjTnBE+EXzI8cubs1BHV568hO0WMxH
o6J2UZlaOQBAxb7iPshAd85keFX0PDOGC5V/cYmTs4IpAR7ERoOD16rDD+SN2Kvi
f+Vpt7zIkFn6qkgfH93PwRGFYKsf4li2Atr1dbFJXvWuxwigKrnVsosKqJtKawFZ
ZATBIibnkQZ8W9y6Fcm80tQAMhxMeiI4+jqfjKtVwjcVb/w8MVyD18lPzvgUsWug
B4Qas8T764tPJhm/cR8Nm9VWmC6D2gx44Kr8TUTX2nM5kOJ9gThdwIcUjeEjNfCy
XE1UUcXYCkH59vkFql3zt6ipuiu+7f2TDiGIkR5krL8ZBlpdtLv8fX31c5U/eTdl
nniKVQ6IZczHQe4ysqoiicAWlAR4hlWNj8kBZKFMu1bXly6uE6wLvkdSO5zqm3Ll
xiR3egLVcoiKuZO9LvUKUqwTfrPraJDXYeYAgyUJSrCC+oKC/Qj3+kLHy8nxf67c
oeSNfLuaObMD1PV58aWq8bbcxpYN01tkD3J5hn04ZYTKqtvVvoOsj8tHeWRTp8H0
Ndqqztq7x1+t9R+MnKk4xTSLHRRO+41ud6opaLqr5Z5W03geneqDufBNF8pe8aBr
DvzNznJYkhvpq0Ar0e2JA2ZAB0dXLrLBa2zi4e0ZWdiyHXxjw6EB5hp8Po73dkXK
j5TQbquUNUcwI0xlGMQSvF5SevTk/F6bHF5t31MNYr0m1UBAmfLzUyhcWIZ0kf5p
ZxtbN4AIFSW++hphFT8uxRzWKEKImzukxrnoLOLMT0u8rTd9zm0wtDyOe10CpTqO
8MGt2x1UXV4OwF/hJ8LvXMsQrbhPCvoLH+LEiF0CkiJaWlvQcqS23FoHm5rEW8w3
qKp1rKQO/L1cDz67RiTZVO/PM/D4C9mC7l21itDVz5XhfPgIv096gooCsDouCCsT
1rHLuG/LFxTSAb9lfSZo6ZZmurwYkNk3xPW0ayWKQJCK2rfzNGze7Z/xD+NHVnfy
awJy4p6pivYX317UiKO46+15Dv4Zin87jJ993QL9PaDbaEhSdbkUm5ynxgvOex93
EHCybxoJydOlyee76/suORWNzlTu2k3LMQiuyuswJo1IPvJDVahrjNgz9T0Hh3uw
jY+ont7MKvQzU5TCPPm2esr+RcLmpgyAB1zbgiSYA+PamFFTI02e/3I1vuhfUx7e
H2eTLSN2lTxCkAP2CnOEyi/oyNZVBFoMgLciQo53Je6Wwnse9nDbWQQmQb3GzN57
FAuBL7sGSPgtyg6opg+qUDjLOYnrrebTlnGMF2OtWlib5PKsGK0TwoehNAjCAhmb
SnyBq/z0476iFYzrGE0UTP9JYqKm0+HDilY0nmS+nCo1GmW3kqf+xIULwKtt6yGi
6W9DjFkucVWiqIs44DfyGbupNmUV4XMVdd9h8Fplw5Avzr6rs63IhZ489imHtfwQ
1L+ItNnzn964X8hKFpAOMX0s14ZI1PSu+7HuzsYwMOjfyAprybH/aRcJDJilz4xN
bLlnt7TgR7EQpYn1WsqR8cHi0NA9wYhsOJGKlj1Jo+mU+cBEprbkB05+EJkPAsjI
g1uOsearYWJgxElkQYSxHJtx+wcYt9YQBjU6lerTdg2iQRUC4WlhzlfBj5f5X/GK
4+K8pDO2X2Z6ot8JRCYGuS5XrqkTEWQj4GWBcUsZzBxxWKccVg/IvOz2Pk6VtQa7
Yr1KigZM0e0zqNa1ZYog5wqL5uXMwKLdk+dMAfrlMgwoFiBGCMJEeBh44bnnJH4v
w/nFceO5+qSLPedx2FLihpK9HwOpDo59IWI2/ZFd9d3HiMPrZ9+Rnje1WWvwjAVi
6FXwVYIulZdbjFlM0xmxWV/2/RapREcxuSAVY2fDhUKLrig0c3nIQlG59XFY1W4e
wuzFppFUS0gqTMne/20nTMqGGSq0/ZSc48nM9Xe6mHxkR4n5SI86kOuqxeXYg1oR
CRW3ljyfBysEQHd46OKW3fK7TWheQlcdWXJrkGnq5pffcv8gW6MSLQs1tX6xXU5d
QD0usEUiZvCsN06Xad2PrkgKA95FKn+M0aHU4YbTmJsPCgfUrS9uxb0LXYJchEY9
fBYU0X9/ohilhajfL/BVmwRFTmz+ZSUIOq3IdFapSmE4/N0NDNcIBel/UlVUIzUA
aL8aCqVrkzySGfT8J8E+dxE1tcQbjs3ysiDnuPlyZUGvVqb7lWBiiJ2GVnQJPhrp
+zS9Jz0SJzMsc0YPyGxhCZ2Iodvr30kxs+NymFioJS+iAAqwEKAAPLJviFV63XNN
JWYf2biTl7gXjXcWr3mG5r4fqidOErz24IjKRcD9miGyLfOlWhNytDTMT9VjN0A9
vH9blahS6cfBP+XPkANUTt1BeHSRnWxb0uVDFMkaw9XuTA3mZeKpTcw+x/sIMs4D
n6bVAH6LLAFnIz6LKcCPrHJcGqGaJfbyeh3L6FW8ppSOEFZwPbYPYnY493t9u6Gn
MrPXTW49yx4cEPKwOEhDghypJKXP5WBYi/XHl3ijWYp1AY5+JIxddRy/znvcRfSA
1JtVoxmOAisnrpvoIt2/KORIr2KuIQzJ43u0funZtjxVfEOcKFBDm30Iq9ZkSjfX
XVI98G6CpRIWYUE12L2Kdfo/ST6K0lFTdYS/+4WwERERI5BFHKmjsoBRvshZHMmC
flPFSq2xhylkWB5H4AS+RLUwHzILZX/wpcGws6qAkYOVgF1wopACrYnPBP32XZJh
7Js/ZyHSv+3Z++6B0g4/hyCGBECzZlB2NfIwQtv3Xq/hs90qyESSLz3TiH/yh0Br
vF/MyW52eK+VjY2BJjmg4VMutmsNAeaYXXKEl9WOQGbWJO36A1yhO3kP1Gi7zxDh
1Zm7NtJlqDcHiMJft4+u7GsgAiX1LVpDpwUNu1iPg7eJVZroLJMwX96cd0GviGQy
/OCadk2rHG8J+aA18CtjgZQhfUMBZkjk+KDVYMiPZ5vp1YajNPZSgh9iqeaOI2KI
8fUo1iF7k+baiItSq7bT+MMn4QK+zI0RxpF4nXyVYVNj1tgGg4E78kHwHv1Xqib2
A8EGl/dArxDfPek1megmM8jOXYQfI21xSoUKX3DeG7h0pOwT1Sv2UEcoXil9dUuj
hHTCOF/CgKgDqA9wObaIq97GKJjuEM+BM+moTiL8Y9I88uD32vyn+74Hzv/NPca5
fxss3x7UaiMoc4N1vgA92+Cb5NQgVzbL6rkcQdb1gts5M/txQTp78CEbwZXa3zDk
N8gGychMJaFdZsga+6xxbx1i9Kq/Sb7FwVdC1vpyTcaKd5m3iHZgU0LieVeMvTcf
vH3GM/8oayuLFmPkgTNeJ66WC8DvkKzX6VN/6v9RsmudsoI0rl9xEZfh7qBYBBhV
vXRX6SwueGrja4C0vnf0pFfVFZ5IiGbtgb1UQOB6i0/O9LSsmcWDYUNzPEZz8Cf/
ig5gG24qaoFjViQ/OqrvXD9ed903yXhKQmlyFVFcRUuLOeseYBdBw+wrSsnm8LkL
mRxq3Q4okroztYjI2abtOF0aOyfZGA3NWOJ9lEk1NzNd6dHaamNDrc+STcqDvNxD
PcJYXtb35E9rqPgj+yIDgkKO+QT3bO9L+eqfkHLCG2v2J+meWVTNzrRomFxL/Jz+
OEPf8nXHwNd9vXzg7yXrt9noUj1qUc04yXrV3FfEFovl/U0/RmfigOaRIuwXyPCM
cTiHqSRyVY3fei95mabMXvMM9oMUPrtpXzLq6dwpGJOfXh7jIuzYE5bLVUt7KjsW
jZY1p5qrGlvNT0ZXwdo+YdkU5C1KcnTXbCmS6WOm7q/Rt3aQ+UWQ8td9A4k9CtEL
0SVKV26oNSF6qkCPES00C8hLF84WZMmVSiXfepWlMQ9oiJRGJfo02ulTyHdGFqwI
0P6aY7uYfkSL71hWdwoPEVwLizGR5++NharVGsOKN3iAfck8dfEsBurXnK+dY8zh
y5dWU0mIKP6jUAyWgKHcn+wVdXEnViFIIDsbyI4gEyoYNNrGBTM39hM1fKNNcw7c
l3wVwL4KPVdOVMkA1UVZdZMdhuJSre1Wru2h9elJRi8zKDLo9o1OCHCNFscuSdCh
OsP6Ve0f2N6AP74Jki6qqvW6FhBVYG/Q+KxvX73jWiHzskXj8zR9se//3WPmOnm2
xhP5/yLCKiDak0L/C1nYmCg/x8g8pguymSXJQJe8w+gKy/syjNkC4oQLJ8aNn6aY
eNOI4/8oz+KknQ8BCYbqX+zk124crC6qSGIg4OzKiegg1bSK9hkMtSZGVGSoH7Gb
LoKA3l567fVoNEN2TxK35KhApDdTMPy5qKxV84pFgLkEkqVpIq+rPTZtTCeI+9Xi
53eW4654gnRQH85lNmclLdO7GZzGDhftZM3ko8jk/CjxJTHeiXqErqhkQLYzJrOb
qYPC3AYnfaLpGjE8DpTF0hUJ6XKuLW40mTnpmSrdFFfg9Wyp3yGkWMdvxV3d+Vca
d1XSHWXOPY6pzADrsKsVoCTFVdIWHZxEB/lJ1Zu7MHKYuu+wITZzIHHLLLlyMPKl
J65/kPlBF0HatuV1rDK2nJRJp2vibnniw2VYqikqdKKp1K4E7hqCb+OMwXemQ6/t
sO8AUj7C/3iF3IINSbJIYx9i4Gx9oNwKHZcHLgr+vF3eVGUs9VEXyMYqXa+GsVqB
PxYlBvrJ9ZNytTGjX3cn5P6+2t1kva1Z38W87YdROqpznp5VxNs0OL9XmwiFFx5Z
6WVFFS9GQJa4/UB3fHEjaFhQcP1NF5PkAhtgY5K3wjZMOa1yRHjcG4Q/JVU7nqsf
UEOXq2GZk77GX3uIUSdRtUDxvMvUv5N+s1FJOWxbAaoexvSyEBMe3YTOoCVfONEZ
4GNxayf75A8oBJZe0VlT/In7ZWq02Wsc+qYi5jp+OsIuco97Pjk6ldRyf12swSR2
3+8TLog8GgbAtJc6Le+jDpfi+E+zYFoWUqkPORIjGqeeUNKIJicfjag67eRQ6wJF
+bUguodsNAjMUjOWtcZLBtDQoJ/kQL23/dHjC8naanWz90AcHFw7GpKfYRZ815FP
uJAb7KO0+zwEXTN6vT6zz4h1avBG1UpcGe/UQ83HHL5pdpXosWl9gdDLKsEjMNIg
rXxfQFM0ENmz1VQjQhoEDQuF9DnTgeZ59ppeiuCIap0ppy8/WEkaM7I3Q6cvdmnZ
uqRY7Mg7NCTclifaNQ1wXnmEvAvmkvcsjlRJ+w9qZS+0vCuFUQINROuPwsQz5M9r
HAdK9crerbr4xmqgId8H5XPSDlivD9bxNyertIwkp1BY5gaREHqyTWfIXFoQ7KVX
Ff5jnm4kBdGSFNkhCf2MB8CDsEF5z4uHX0LPdloGiH61oxgnDqyonhxTUxERdun0
S6CunJeLY5ESMKbr8cbeCmmWsKxWk9qjFI5O0P6QTAIEf52Ehf0DQah1uhA4Lkxr
H3MCzcWXgOohkn02iEYvSQmU7OSCLXhuXZHPMm8UK8CXwD660cKfQEPFI/erBGrG
4yud/ymu19P2263kkBGBYTTVjti1warpFWPcWYJQSAYOKAQuiyp9Prj6RWiyUWH9
HUFZ/HBNqmiKG3vP01hHG/AjPCgUgfNicYW3A+IdtC8qd7chCmUQYWztMVk0ohp2
xI3USDe303QnrnRZRUS2I5tbd/gSKQhkwYarWE6hb6QSPR+P9EbT2pFfT5PA9prn
SJEeuFuYAuZbs/IvfXwOhLZg5lS5cEPKuYKRw7LS6z6Hv6eYwztmdpfQZUpR63/Q
a94fPP8QK8eivlIeLG3QtrZEGakrFyJztp1aPjEMUfuDMUp8oG3DP5cEWi2MeQzf
+3io1RHeA4oUEEnk61xbzC1EJBM4223Zu8PP2vTtHkkovZVCHjvSnZMdrAghKIs4
LGE9bhBziqLNxjqJpFc+iGrygTUqMR/on8gxi65Aje1JQRzIT8YDh5LOGtg8zM1T
JrCtgQj07KSxRg19t2QCkGlbI5eNVSkctpbP9lsEPvBrushYkqUxpg1UOJ9eh5Yg
awdCurTFFQCq9QJ6jVjvXThsy1w4SuBJmtdS7Y2Ns2CllUAPovp4xXpBiJ3p3xsv
i0N7lxaOQVqk3NqwJv8dR7IDr0tIhgLkNJszyqsMWTF0p6F3OttBi7VLthlNOk2O
/gF3USvDfGyjpvlbQGkoY3iJrSSk11FPb3/Xcnfzy3mLD/bVyIlDPTvi+mfvYvN4
49btrvVqYr9kSZOyQT9RvZPmsIrZBxL95iTF1nStIuaWTbcApbRPgLTeF7y8P2V3
hxKIaOsxTbtuTeOkfJ119wHfU4mJiGi8eNcK8BuSHGDW+3PygBroRT8+bfvmQqma
lswq0Gnq+o3jPbvgSsqigY195mboGJ5xyACgsROEsUjvGHiqCFsXEiTvsuR+qh1b
D4MOQXPI3FhiL7RctgzHo+Y+oywC1tHN3C4JLbprHeNhV5/W+leBCWXk2gAAIFmc
S6Dd2t0H6ubHgXCz2DmVVvtlErk8BA7T7u3xA6H4S8jf0TjrCg/81Nw8Fow8YINQ
bB4Q7vvxbAFM/+KFc973OHPWd3RaMolw4EfGUj/l2l2C8XddFVdkMW6tBVxHSYNh
2lyLx8VHZxm+t/G1zvFg9jeqx0/vOT4ILs3Pw8pxG5tfp++kYyug11iIoxBObYJD
6Fjzkcay9xA3V4kf5UsWRkUIImzpQ3kh31ACXJmUTJQ8EAFndUpZbM6MtCdIFW3b
k5/Kt3Ohwy48aHU4fyAhuOLG40xU0FcvVv2bH2WT0Tf5Cd5i8Dr6y/fUJATjWvw2
5oa4cCKOsyHvjFsxGdMiyXxWS/e7GAQaokciTHbgWw2vYkRcL99g6w2EZsN5d75V
Ct3WR/ZzCadJAkxpxgCSjxI6AkJw/mYsTVxkoq43dAZhVJYdTvglUvs2THO12Xj0
BTwSVCbME6jIlnENO3uCA29YBBuUtC76+VNeThRUH6Gr8m+ynlac0N2J8ddIlbIB
ANtU5KaXm6YvpCcqc3lKk/HDsA8nCYPa5p+198lmfF+Ef7F78FNhS7Xe5etdRCZW
fPt1rxTpiGqvVXo2U2XdyBBzWhh5QqhBCK1mIp49fBl2NceUtkhXKH6C+fMF4VHE
dKh8gSeGs7xVfM4x9xB319aVDfaDB/adMyrPcefaPpYELjtenQhbrjJJatLuy4Rx
nd78mZIHSA/Y6ihGDYrMpk2YcgN34coLW4ehWo5EhTKWA6FzfeeFJ2KCOV7jUqCI
f8sCN4orRTSaKdDqC5Qqh5wkC6kuDpgKb7XUPnE/Dc3l04R/j0IuqoRjBDYV1EFv
rmehoB/VV/eaBbu694pPHm5ZqbDugDWdxAstjYphS9yBzC2TtZ9XxPwOi9cgZ5gb
YPcq3ISORHTN4oO+Yh+tVjEvAm5J4hdEqcpx63WHf6F97kdSJmqkQtS0EOySFfkf
u/GbmMEuQ04ENJslJUMR1kio/rC4+IPOBZtTVU+tMZnTnO709SxhRumwFHlRZIDG
0XxkAEMhTn8UrQlSCQ6Cm/86/Dz/yWZjTVi9/uiyVYDc3sz0TuaNvCQnZs+5r93y
fzEbKL6b6TOICK6QsfPJl6bFz9/6IwqcR0HcixrsZWxvXINPDlZaE6YH3xM0nsNS
iEJMHguynE0R+ukKhzi0Np8zLlkDQpS824gvqgDSeussBQAtSoZLbIrQwqvEQCKC
TGuqvR/WgYT+mac2YFDg0ydbBs5LuhsWNeLsrxrNemU9hGjWsVoaVVUugzlDDS6a
X2iB0IGwKIL46JnX+B+sCglNXUKHEzxIGzFXqOpeicUMNInNpd4PZkSs7dx44lb5
jk8sGWF/t43Q2AOkhPpbV48V0K4pdkmplrEUFxVvFQv46YwgwOR7rdhpz9W2Kukp
kxfGYuTB/6jbrGT2A1jZww70UWs2YGnLm0vIJF5MHTzNkFjDGejlrUFgWFr2BIQe
qpxKgpzUyFwmT4FuLFeixURwge14atZ70oQlIC6POgBIh00QiSJHMjTKb2KSYcYZ
gs4Oxv/rznjmSS2owGOgTBUeG6BI4KhcdDvwaYbOaM5El8JDiEkGtG6HtAg67hKw
lTgrNqiJgc6oErc5jOurXvqsENxUSHO8jlyLeqKBcwWCqG8GvBB6fezb61MXGsLh
eSMBOU+B8sT+NTlSuysF9BDf8o50s7sZ4hD9zwsdrexgIP7In80P12etQbtaDza8
jABZWUl//LRkGjggoa3OgJTLdRCTbv+od8/q/XlBv7HzvkhTt8GOt6/dPqkXInTP
pGfR628KA/QWbylkTiJlaYVCaloUh3Vq0hNSKaPYIveB31uhsQVX8x4KZptoO/gr
5HweaF8oNLa50vf6mOEqqSPeHk4MZ0Wznv+mWgIBPXzzgCgOCoGt+CvRSt4u9tK+
L4JTrSk89o44R1DkJetcX1gRh3Ewb7wtRSM15iUAwcDuY6BqODQORmuaX5Z3XBuM
uHDpeWNzXvR/wbj/hYeBoAVmjMomHRcykERAqODj78jYCFJMAD/+duBL8HFmoqM+
ZdV/6LOiUtN2Hv09ColtXBK9E8ocffGDo1G3WvAzd37NAL7R31PjBDFsKwp6kJoa
9JlS7zEoB1+gm6gMf3QFCOwv0bxirs0NTnt18Y75SZ0VxUdIW+c/zRmv0wS4/PJ4
NMyQtMRIbyFSUfEpa1yCglC80lqrtrrbtipSQTkFZVGmSTnZjG8gdbiwXw+msvgL
5LlHiID0dL16c4mfgo0/wsbplyNFVMT+9i6gZfGBB/WreJXDM4XQHI3LrZdGbUic
0hHBup8bSu/o76wy+IonQUPMuolkZHmg8XhkDP3ZEpBLFJLFSzXAdGQZGME9pKy6
qNr1m/wqJ89/a+Jq1QNVoyNvHKSnaZzUOjnZRKzDInr2BViO/Xg958KTvT5nGSG7
YQKrzNMgCVxXV6MjUWC2xjgy1yyvB5qNX12XWF0bdT6Bl976mg3ziCmLFMv6WhDT
eLb+eAn0UDnIi3NYV6eR5yIuL3gbX7coTcCQcfgWk8d0RavR4JCrG3PBinmA0430
FsPp9BpqGcZlg/7gqXHZHe+V6BVt00xmangi+mszGgsPWSswrvkas3kek/OM0WWJ
X7YV+/v0MgBtHKBsp9jg2ahJn5dqrbyLXnYVREo9gG6dax3nZX9RRaNHjrA9WXi2
/unejp4KadOWUeRG/OyfXbFd2l1eVUGcIQtlESzpnbgGP+w2+STkR1ro43V8LPl/
y3JhMEZdR13Vy/jmji4X9Aj8SG394Ls4van1yEq37BawIAUUQ95Y4VmOm5M/+n3y
KH6J7P7w2WVkGD3Sr3ocJzYJj+d8keoZz03XXNzZIpQjhFpcIcECc+Qm33K+wt0N
+r3zVskHPq3Usza+AgRjwPEYb0Axn/B+LS80jw+cTZhAKriXpkyBZHkBehXX9Xr5
0TDjJhuQ5xbngZP/jRugw9Z5z27wqKY5FuLGGtJWD7f5avGWcjX/9NUmM9+QrtJq
SwAiVTM8VnRbw+Ip8lkh3/Jh6+8PX5rw2wEB+kp9O0bTq5DSkBnKZTxTVu2VO+VJ
BsquPBk/kK2YlYyjx7SWVW+fEncISjf4QjfiKwY+RVUj4XxQyIbjalflFv7/GiVx
ZiVq+IpP1G8v3QUy790nZrJe0DO/IjdOa4hmx6uUs2qpzl2f5VFeQi5FsbZZFHZ4
A0+hmNdqs2bf8VYH93zpswz1eYLCv0KLgYZG91uCkh/XubLLJTMyIXb0FfTj1aWW
dfQzeDBhgILgDPcpAIbPGAXPkExWfW+ZBA7Cg60fQaAhJn1QSGFi3GQRXAkS1asT
uxIAiZ0y44Weh04MfrnQJ+PK/0yb6vdCrn6kuHIfObJ1vtnNb5z2Ufxl+7DElqCj
6I90JEnIx05sjUXa0Nv/vfggY+Gp+R+VKQZUil3zfyJdn7LtFK/JsNDtZ3cz2PcL
xU1h75FLbp1OjM9WCgLtk1kXMTaAG/icGZwzsAsoQMECWoqKeCbbxTI/RQFBFXnh
kSiUaecJA8Hi5QSOQiJ8DsukXuXJcNkzBqIDb5D98zMBFJ6VtLCxMSWALMNp9tU7
7wGY9yqM57Uj81bqvJLZpEujr7cFFdEOqR0OngLu7gjhUz3qFfilfoDUDYozDtrV
8qk+byY/QVdGBqh/nxcWj0TQyLZWD1/gCyv34xrHdtVcPbbHlyoRGtaVFQryEa+J
jNADYMwXCXeoVzZhmvH0OL2nPLf/w6fetIVGR4WpLKEZ2YYBDPQWTfdMhk9lmQpv
EX7edx15JTv7l634PE5kwTJL9GS9MjMaXnzJRkNtknNh/UBiIdcUgzPJK3yDTsQm
b/ECISjPMva/X3MHBOLZF0YeLf9bvKou2cIo30R/sYVlIuzdC1lRppOjbQeLZ9wN
aJVguF3CVU6dBd3CGsVfYOddrfdIuDPpSigihjpEVxFIqDeaime6hqFUotgr+aPy
bVEgmmG4Npi2oalhbms1dGUYg3rOoAODshB55Bdn6yXX8R+jL09JRtcBpqgMl+os
E8IJK3LYhhSOa6i746K7DKkh1ucVFEN0uA+vNDrCdfV2OJDerC441iMBEiANyRan
2apGTUubOEc/0tE+T9ReasNXUYtj5xQyDGqoTTNcbp8PbvmStp/Q6oHnBxX6d1Rl
zInKjjWk0mIyvdFpk56MZBiuDHwm1eNX1htBVdlJQUn1HrA6bFe3aMdNETEIQdMZ
DqSSHGvbZVqVEChnrkRtUGi4sOtQmLUQVtZjol6hkk50BP3ceBcmZ/1OCLnX8KIP
rF9Z/hwKAe0wii1iQARQhqB6EDMeuHzyk7ewfvmoQYSaWp4iLyv+k0sHm7DxlCLU
sPDX7L5Zda5QrW0EWoAjdiuvxp4PBhbMPW6FAHzuFNNXU5npPrDkelQrhbN5H4ag
jxt3FVSrsu1O7EWC0Y8d6IeZRmCQcUtwuJ/0iSIogB/OunsmK5vNb5G0mIXZc9/Z
NBtg8OrM1j0e2Yyv2JCEX7qrX/ZLPs0noaK1Lu36wMxN6uuK18EyZB5R+VZUfTTY
lUmmNkgB1x27zngBP8ctU1brg4vO/12SuHev7tH5R8oIf44nbDbKm63DFi8BnDy6
cCqynMeRvPeoxLDi1WNRJgpFHZPCRsMBVVaXMM9lGozIdx9b3M3dQXykZx+Sf86e
OWbBPAc915WD/syUYQcdR9YF1QLwYNJnSMCdnHG+LS09XyCVYnXYON0wCrxrA3vr
Qw4yfKMU6O33aNfwvMm0sowCBkIXFNAL/JRkBSkofIee1UVW8ZLUWk6UwdDN2+ft
v2+9jjON35UierrkbeqWrqtJwpf1xwNiRajY6RnhENfS955MNMDOMTKs7kgC5iTt
VDSluEarMUScE5UGzViWDVHOxdB58Xs3DuPl/FS9ZuKmaoZT1jeW7eKWY4keqqul
e8/0niPg+xTUg7I/H3y/wy+4GtGsawz4FDfGdVuopE73BMLjlGySX9P3tG6Z7jTi
nJXVXJYsXOXA/nJ3jSIqrHOsNXov5WX8Dlj1hMG+6LAu9XXMqE+zy4ioPoxC5gxr
0pXQx8JAaYek8Wm+7Wbdc6NgDnCE9h0QFIseOe/eXoAbfToN55aN6/1hKf3gFH5m
7aO1ZrA/fP+qhD3MU/Jxcvu9bv++S4FxfZLho3oDXG7wme7OplOBxqZlMWTr4g5w
yPv+j2uvMCoPi++tnbg3zA4rzWuayvFpUkB/B4tD9yz3hUQ28kdPic+uCaPodN8E
Sn+Zl4oCY5NCwrcMdm7/+y1ct0ldWbjmgcokkhrXNZNBdMYC97QeT7ymezJIcg+U
vL0vkJlUBp8kGRvb1r1cWQVmqlJYOXT/nP5q7enblcXQYLHMi8YXab/skY9kLR+a
Jq8eHXOY+nirM23eP+DmU4l1fvkCzalxBcHOQGpchb34Ow+fWXK0Usm3fQy2Fy8h
geJeoiqB7+LKMoi76wY1BC54NdGB1vGoJT2MhRv5aEJIF0lVw1AC0Soj6PdSrZgw
BGmdjo68AQde8raqP5FOd5WS7SE4ZoaDZWdGozMS29g94hwXW+yIUl+Vwu5KCZi0
uETM503Jf23yQkKsvp3GbrxKoOevlaqdhDJ92PBV7+ksh1Qr1/HH+kHEcQzMvHoF
dIXzwz43lBjSbbhMBRqjceBsI6Ds50BMPN6G31cNHZcvNV0Wib+mD7fN+/fReX4p
BxsJcNZdgSLzujqv/EpicI0s1BR6AdGuzlN5oOT4Hm/K4xm/OjUxqCzZSajeNv+2
84skhJgQymhdexj240GpwV09mjxOCXm2U4CHmeRH9YOqrYvTdEie+FSA1XB3N36P
W/gQYSM9Gp9LT9W/sQn6IchsNcb8Aw/bRqBvnYVQyJl7xUld5HX1QgRe/Ys2qUVE
5E8d7JlL16oV9SYk7h4WmYIrq0Uw4NRWcvK12X0DgpA8CnwqGtyxVZsuJKzZFRbs
KKIy4MdahmJcAnikajroALlLI461u2m0eQ0dabeJbIQwKceSN4rhIH8Qgrs8LHou
fjnHVnEDw5p/T89kumaCTtTCq0JvqOn6ebQ/0ehGc3tM5PagBbMX08PFSlsCv3/O
uCb7ZFhuLUzPeCWvkRBGuF86WQNlRHEolXxdHB6ySONkW0CHRl/2ZgECPymCDB1A
eLovIWElk4XhBwvgEcwBXKDBOEPo5Flbuf01rVPkpDgoaqOXL04/Wd9gqgeL7EM2
biNPWS90et9+Xa0yRXefMIqi7aiM7PeXq37wRzgdgUKhwONpgmUIig1ZEt6tnc2q
GrpgKjffvFnKWBTloaVz3nJHHfiijxCAFjvXOd3d1zGlkxHs+6RqC9m9CfzkYSHr
4Roi7LTmiLjLecJwBau/ux5zFDxnpd1wEc5fIYdeyWUAzGkh4ym6BBAcoRpdesjH
Ozz4xjdVjkwjUpMGVrd4s3BZnN6LSirOkbIoZ2hPbBfo2OBrPJhLenAwLKSC4Y/I
zoDWr+dSn9AtZWSOQIIMUbWDrgK8ivP3wWq35IlR4hy3E+WRACnDIZsRlQAi9xpW
qnGvHI52i1f0i5E2gpF/4FHPlajzeXquiyciifXQzhX5URPmoK4pSOG7In9xL8xb
G07Cgrs3/TU5kqOIjuZvzVFMEG8Qo9i2dzbPRKefGxBrmRrqLlQjRvk7/GlW7Dsz
E3CLJnflkYjbHTXXGQh5b253YK2dmM+Lx+qw8LS+wFd8YxyJ9F9S9AHN19isT8ZJ
R7akjVxaqMtFqe/99ngfbVzdFjSZSJPdt71S8nyjFs7W0toTqYdcBjT/ki9S6K2Z
/TaYXwlgLRRxnUPjH1JgRBiZZqwgml4vimig8mY6r+naLW50Zyfsb76mYa0ES/Np
qTxtU27yYHXsCql4HPULJs8baMNcM6wMHRZE3lJZng7bk2h6tPygqrGDLMCAZg+G
bAG/uKM21RIB5rbtu64i1YXupvPeP7sCxB5QIwzS/W3NFhkySPEwCqYiVVBq1oGg
kTVJD11LdP2lRvEwwOTgdWQfrADnuJ5irwGD5+mHz/VbORr4h0CcMQYWbjEgACS+
h5tDJ4lPc4EN8L6tNrJ8BnEMXSK63tI7ObG+3TcRqe5sdxPeOwRR+khahjrx6TaX
We52X31J1ErPpW9SIMPLMoR56qUghnwHDq4tDHsKDZzgGCMluhrm54p9H1nNkPq+
PdSAwFw4Detgul+QXMN2jaFydoN3+YnfMSY8Tjs0b6RKCQI0yl5rMY3A56B5NCzB
13Pm5W1XXtV8TNDVls7gYRTRDFbfQGg1gtCWDlKha7Ucdc9H6GL3wZFPtaYmlrcb
IrVkiHwqX1EPcTfdir5JX3egRuqB0qus24OJhbMpmkL3ycpVLN+VHnM2R1pfGUKn
ACW2CUBvPs0XTxUrGf69+bZHi/ctNRB4fQtixmBlo6nqjcYyCKY27P+I9F3yEf0M
1hrOrSxBMHf6nDBr22eZBadRnTqWWLPb2yfXWa1xeKTK9O8FpBkAha1QHpC+aEci
EnKGXJ+7osLM/6xdayBDhgoQY7PBON+VIVV62pqf3p2TiTBDmQV4rDEhzVQV1DOQ
e+O9bsmDffOquh+ZdIfVbxgoJ63aGU1K8Q+j5E2VBRGu1HzrzqnnUUwiXXWfyyUF
WUb/1dISU7S+9UBwXsV7SKRdmVVPlyN/hjO1GQ3SR8EVgOJcXKy3L8QlnEhfl1Pg
x1KYrK5GqRXW3KbRhmzs+Z9AmCVrbPSrq4jIy6TWTxMsz/8gzc43TJcAzb/NFRdY
JJCTd1WzzBghDxbxpPbT4Nn16PuDf71v6QeK+sw/k9/g+yPurCvtsd5XUU/9DTSk
6YYFu6HK7IRoBOG4LYv6KprInEmRP2XLIPYcOmSMOPDn1Db3bdnGensrlRnbv/Em
V4Egw3kosfrIqmbbDrPD19FcnpfU6q9t+JIdGpEO+0+dvHgjW/f+8fmfbYJW8vQK
F9zJKvThP2tSgAwwUbbpbt9NDblITNZ4CHax6skXs0ZyygcTUfHSycp+7fKC3trR
CXuk1m8+CcdLBZatKncoEvGpFoZ333WTmyd2GBKr80uHJIYPbFEBTRIkukh5xvjm
N61Hx+CzfW4MzT2Z3CGCaq2aZoQQ7y8cf7LQfZ029PY3Z1FTUagCn/tGfgShrZis
nk86PJe0EcRrWzRPU5Lqa2bP1QZ4X1YUDYT5X++nk7tFg3z2sVwWD1aQ1kfdcw2N
n0lpiN0nf1CS/NOoeAYSmBB+Q9CsEnpJojTkev8Th5BKOy614k2eL0d86jrfZ49l
fWK91NB1KPw+HZuFjPwTG+Wo/3vBk81vRfyu/mVbV1kOfIhJoPTy6cziMprg8fy3
Cr0+ecZF3cZs0OvVWaEEkC5RPWlNyRgmLeQGaMWfJzp5IkLJrX9avu3ANQhmY6jY
+ujJKtqf3UgvHDVzTzt2sAY0zjIleg445QdyonFcszOaKgOARA5teoQBL6KKLIns
X3tWihVESbxz0SCucnyvsVgwjYUXRAaonyk2QQDm05nAI4wxPWAU1HGLb2Q52Y8o
8ckcMyYnOxxzU0TpG/fNAFfyTR9aUPqyHSpbp3naDN/N+dEoKctoDgUqqV2xj6P+
4Vqftn31DRyEpMoZRSAlUj6sIbdDdpLSIF09Ie9XLcA6jwudyq5HDoxoT7zERz2b
+kp5LHwBXs4lMEqT7uPVScfKIqrtLfIOhkplsxVtHqYbXuBpG5SUj3XrxBp5IeJD
GdysgKk1itJG2smvFe4w+nsVhgLIwUH5WkxuXjhlDF8vc/XRgWOOGJUjjCjMkxJO
HEAUNhbqMwdiNa6L5OGO5zeZtTh+H/0MDkfYX11zb1XJoJlMVCYsBeGAk7PUfaAk
VW9uI4BwfQWuc6pQRHUirIYWdoH29TzUMRDnTLfkkRurzLLsmtHYJjglEU8dHd5i
XKKFPq7AxYnw7wiw5hgTA/VDVfXqBpKIajeqN1kq3DtqxvuWL4JwmGruj78UHym4
G83g+sS49gJS/UeDgWpfCXJK+dHiyt0x2I/wkGUCe/4QksTSk+o/i05UM3ZWaZkz
+9+MLXjqxg5sxODC9+CJKYSocMqvVu1I+EC5wKhelH6diCQUPJ1xeR7n1QdIzb40
RPvbqI5LnsCRa3VbK2H6/LhbqT97F3pFJ0MfbfMLizzZmhRyEZ9VpsCNmW8gc9cH
8PjRjUgHgc19h2AVSH2qlnlY4BDrYTBblxUMlYKz6qwZNL/WJMAi0gZLDq4vfhWv
cXA7i76oabnPhxuZsOsvgmXvX7R42rmi43q/FdVY6F1zpqed7waz4MyLJCfJosaA
vuWCFYbSNfDNAvKqJtILZMCgZ+7E3NLi4mcZ/6yA9wZE5AodoTitAt/6TvJGGJMy
KC8BHPu7jTQ3R3fbfjw5KLhTm4GcZ0sL/OUEoituR+K5DPnf4LAfLHVw1kA1sb0u
/6MBMjZfQbwiVLVv7OLlNa6PKjYJz/7tX76IunFwWLzOVLNtdW0OWdgoWXmV0Wsg
r0kVj8SVoRnYZKzn9DeZe+Ojetf3Uv41u/0Zb7qYxR1J+ZNj6QScbEVnJ4GPpMKb
rQWKmbTViHgJ6x9CXbK7qh4nOW0tj/9/zma2nHyvzR/v/dxRtg3NbOknWisT0pkq
uVJQ8IdPNoA/pebmYS9mt8Zq46yn10krBsa2f7nulGBH8SchZnYZ5lgPkk6oF4cX
/lOoo4fnCAjtdCcLp+jS2jrhJ+hj0aMoQczIT7XhJWXog8BdVnPYbVkv0b+Gggdi
28CqlZwIj9txyQgUpCZ9b/n15KqVG93XfA/l7mOlmo9BPvBaul6+9cOGcda2po3t
K6KGLqUCJiEwXAMGVLEAV+9zJeHLGdNkQfnW3CkJ09cMSTyo7j/sPdMrXjoroMis
GSah2fNrjWG0GhPGylbbA3Rmwurg+IVSS0y+uJr1I4GqAL2fHw6nr6WejeGzZJnH
NPdDwMy+vLXZQ6XUxE+xwy8cuJCpincCNqCIHpYcTPqf9/vOJWI1FrKOK3T+QmgY
XoJ4HsoLZZ4v4ScggmLL2M/xOzkk6mRjpaH0A8UN5Usew1U2wAeMu55StJfGujBU
56pk3xIAgWDJtcHS161lyC6clEQLG9S9pHlr+wVAp29rWS7nIFjbyUqrvJF4/ugC
I/WYEZwbX+vstfTT3PuiqehaufxUcz02Fuzzo7yWscmNURYgq/OCwsNSlMGfNG6M
rt89L5SdPBPTLFyrYzmQHiV/K5Fn4dpOwmru0iQtuCL7xVXsSVZeFoslBNOjPscM
LBEQp/L+4n82Cag+XISvtSEDtMu4YfEN+MXsCNDavRhDlz4gzmCW9PdNIQXGsxZi
JUtqfYr9k33I7UoC/L/q9ZSpL0UrbTPtQEjcJTUedpxHVGF++qleMf2csbGr7SaJ
lnbKPPVJwLf++Tm81ddCsuvLyXQqZNMJlXCW4wEk8rxp/YYFIedtdpxlJV8OvLTd
IL9XHuBc5wdKJa8QXTTtSwzIBrpHkSLN+YvWIi023y820nXVzzPx/9qifzV/oW7f
SteySJMEU18vLxmomNcLQmoPAu1HJ89v50xbexG2Y5jeIdtMW/90pMxna4OxBHbz
MrPpiqdYVfB+r+q0Zdk7KHdD7uJJ17cRBpEgl+0QHxGNzY001wXo7nrxMUuU6aaL
eiOn/SrURsYRHxu320ezD+0WOJgApv7xL1WrBqH3olNZBuoL0ovFNGtO0/pfj0U+
NEHpkkbKcwV08jH4epm77Sj3rymdKZTrV1yIvkd4jpSb7+fpItLF5RYH6LAHXg5m
DPVR5EkokGtV3G/WPsLRd5SJbLtiZWGDRlaOqXIEsRo5s8ppYEPx+iJnjQjOiAYi
MPmQGgb8WpmxWNvGNBEfP7ERhJxOANcIEBEbF6rZTE4gmZ2cqYld+iC0SFTOpy09
WH9GERTCL4Ke1BgFIelsVwinLxoRn9kOMItiVnD4LpwTXRUSzy+3k3L2zhVXSSrC
qszeo4ZBxCTvD9v2vbd1/TUa6iOR38mlE6tuvZcXPAtalDK82RYD2xdvbgGXUypF
Ta3uOyCxd7wxxucrfcbe1E17I5P6hMdTY7JAFCoaVGIz8kaKv7lNa2O7Gawz9w/u
N4ykVQw4lago7Q1/ffXJimJXzPP8S6ddxfALqpe6eHTZ4Kp3hIiLv2mVw4/2NDjV
0tMjDDdrw3RzJS9slFXNcmhdk1bntg/vw/QS4rzv92urWrpJ8OnOJ9AByj/0n/td
RyWsaSLWyZDWYzaeZeCt9Ce3oX1BdeCcAtAvpa34wnS4hUHBf3lKTaI/3H7sXsNt
/F/iESyxNyFrPqHxecHx2rAk+RCZ9R8+0ACtQH6R0FTE/LrpMtGb877Tyq/fWqBk
6JukhXFwCtVXCCKik8cAjoYNfVx5v1lsXpSPtxyntpSbZwwmMZOfMkoWpW4vAp2g
vFYpZNCuhH1P/9A6UusCfAterXbl9i60k7zdbpHu7OBUD2y4CGC9ixk3MedPVbBl
m/QmcbSUkhYkNGfdwVQ8VzvuECtg1UAsXh7nZeZLRRQQTiZe/59JSvqZMpyorw35
ZBQ0FwrzyII+iy2X3cepS4Di/eFTu7TkEe9z2FzGQjoTDk47W6c/TuRI/KArxheo
dwUvmTq08kkN7+WTN0t7/lznMQyOro2LV6+2S8IhYXmFaUxkxL7SQmjU7HliFGPY
v/zmHfkFNzwtET6oCjaySrSVb1Kmrj6Nl9pnERwqDFvuvRV685gEyiZDG0yvYUk7
II72DwV8CV5LAvs99pCJufZ4yvDXfEQG7hjC2CpKz5QSkUgvCu7rpUd55Vvc88/l
Vir1ZT5+D4lBo23Wl1NNfO0WTNZrOUtf7FtE08+psObUnMo3fkCbYKmHgotfz5su
Xmcn+Vozv3YMumu6YSZ+mAon4ZldD1rBQr+KfmcPoP76wih+SP7XDpsYJCnvYMUg
rLgUqB7gR7YPKZcOYwDxG/bYlIME222GSW6r37LBCGuQpYJ6u7jVsxsKdSXdNO3v
QFByp5NibbDmg2q5O9TTfoeQYr5XreFKds+TPFUufXW5ZT7UkQBPaDasyZQmJL8g
/x7N1A7Q5VTkKSjBVzVHGRyXPCLyyOJd5swRp8SYPcukDgdgbB4Ro57vzWNooq6i
dDae/vStK8S+kO8RtzWb6fsSEt2/1X8yQmfH98DU6izN8WOpzoA12pQ8Wl8rvfvK
s2wwtpC10OJlBtD02LVG1NZbedFK4n3mDfvCszEyS8Jc5s/tLAbdbdJ2bSXIEkJ5
2gsVkWNrF1B+oRVItd85VioWlgX8klwQItvVmrMlQJQah4annuIPp8/7QMacoz/G
1en0YQgciOYIjN9tyqx+n3eYhiZvJieSnbwoFV5Dc+IVQkilaK4T3KEi+57J/9Hn
x0x8DmgF+ll6TG7CwpfdnJosQip0/0B0kVFrdn0BY/3Oy1hBc5kZ4HrTABykRbG0
Ik8o4ti1Q8HPFaYk+eq/QDd4pJ9+6H0wJLtzirOP2ehxx7UnReEAiXuyGkw/kl89
VK9kMpCT5Z3odzXgoNzzmwBncUqEY1hcnkiA1y6PgXYZ9wvnEi07xAlgQEDMUN2M
2mkt8bJ1T8+RCOM+DLpUOqcfb32plADht3iZ/PJ4VnJG221viWAubDAuKZQO/+Lw
fyrRS3X6GSguef71ke0F14OUJXNxD2LK7yKBEkiPGAW6e5ndJvalLc/U6akVwT2o
767vVxROi0g/45WloTRQ+VHmY/LrD8LhtFuJ+s8Jxb+C22qtihGu5cZ4wdq48XxK
+GEQ7Yk68LhARgpWyeWkj4IvpTJjlr7lKZr/EQ4v6ML6CrFaTVp7dwOPFyGYMkgr
a9sCFsBYpvqpKS/csuedZ5Yd2Zw3jg6x0xPKqAPKviOKhpfs+Et+AGwm9K76UXgC
UnCTnmhsMkXCe/wNXgu4MuyHO4nSUtIgcZu7Sbm0mtJiaXzYwzKbAzzQt86B7jcc
XnkorJFWqCPjW/rQOfyBdFBlMKDC9dHTl1ZIoFgtqKYRNDycMjw5OLok2/quAM4S
X6hWUbc6R1AidGYFv35KpPVXyJMRyczaOWpi6rCEaX84mxP/1yesXpsZezRykdbU
XWlBBXVIQ7SoB6qqbWp7ue+puWE+YFayPPG30kLfBoa2vGhLNyjlCBotJVjVBrgz
FIketnGCb7zHhD6124McWtFZ9wuS4ACXFABN/pSJHXRuzIH1Vi12izkriBAiQ0uA
v8hgumjZqFiP6ORNU77ywx88L+qe33BbiIkKOXR7V46PVtUTLmBXTQkYJqjUdGNT
+DTvfPdyQpvxDnTrbqsanEgM2gWl0HKJCUpuXXBmGESjfeXlQj4bspCV8OusMbbs
oa3JW9GsQi698WXjvzd2CqD+M+U3k/kNHst8Ci5+qkpn+9M0+VPNP0EDS6kXebLs
l+rkW6HRgnJFvLcEn6nNVKIiMN59wJgtSHbD7Z+Sbx7MA4yUUjeaBPnvrlBMbwcV
EI+RtKKWI5qBlBWgs6L2/sUtsDJK4ReOGtseDxjj2UPgxa3VzF3nEFTKH0zAkKW2
JF6F1+IE5woyaanh0ZRV8fJeQyF5WQH/m1jO/xBtVEVulCe+JGaDY6QKzfRTPVHd
Mx+VuQSQOOCxbkPORPHUkPSVGwSHP/v5CKT2iNMTe0T/1DPv4WE3LqD124/2ouqO
xHJtcvintR/JiVpYjq00c6vXHcYFR9k/bieNhLgv6emXNZ7K7oBEsrPvxSJn1cQg
QIxTqsf0ZBAkkkihXSaVSmaDtM9pV/QxDOwNtndwnzRsh5RYOt6V3N6cJfqn65Ak
Z7S9YYCD6jfTL4CejCLlAKQWLqlCbpJWDI9pI7rrYLwW21deqvfoyvUETquEf0Xi
b7sRikZdJ48nFB95EsKQQhmIjtTvStuGG7yn9JPd0DUfMRKSSQ7mlae2SMBrqqrz
GaX4gm3nd5bpeEkNOs7wc7kCm7ssNHIGTeI0w3rD22I2OaNd5L/qGZnK1yARGo+R
wTVIVxpgf6FCAV0P5EzuE+ox0JgjkqtWQJCxx6GVVivxokT6sBcRPDLyvinwUIVT
GsF7YrhW3Pdkzdj/ySIfsn+GQcKNNPs1YXnDMjq9MIHVDuGF7DX7iZU1ACvAXD+z
i2LYKOPq0tcBDd+kN1CXkKG3IWVo0H+Ayy9S57fT34dhBzJ535R7Ysz5JCHSDMfY
V9xfK0YldMApEwQTmMUlQGqRY2KWS7Vab+Jr8cA3dQuWHSkYOiRR6stNxK4W4MCl
BJA8rnbpSY3803tJMYQgq0CP1F+AMl4ttPTlreNPDSLbgK8i0Ba7Cd8lIVrTUzf9
VJgkgYeN/c7Vh6I6EzPr7463kj/DeiUU8rcGx4jF5PU0JkOio5Qgkv3fy7o28yBL
wguLjOHuGTnhxGBSIc4Cdd9Qw1x4ZWH6V4T0CZsGESdk7TH7836spMM97ussvBY7
IfLnqWcCTTDZKaSefdojF6Ik/Ollr2A8Arivlvb9k88YWpVu+Ul9p4lUWmXc8evq
Zu4A5iStrJh1wxnFwCIsjacop8PzXBFxRLbnmmADhAXEDllLSHJdl5Wk5Jsb6ytQ
YjcE/iYNkw2qj8i2gCtsC3HkRvoQLtREYEl2XclapbngD+m2pnASsY2p/ONkTkLa
2xGGBWQOROmh85dDhthrR/BObnNOaaMnORu8tK2SjLZNqxi8JGVOOs6+d6FAV0tF
56u42YMB03T0/8ii8TzsB45CHpuY2iq2RVYVnUTne8SqT5YRo0ES0Rj66OdLbWjL
Kf71cq0F69RkUnMZ5y7NB4xCLPBEEBgmTjvsA2ZK5Kv/ghOKEqyontaFlNrOihST
Yl/DivXoLWSD39Z5TFgWi+pyIX4SFcuYYR9qT8Fzu3EEV20TAHXJ94jkMNLUvO0Z
ZNtJVZ/BWCGsPX9+9UZUfqBZTb78/rr7tFnzns7uLtjWOgwu2fYJKQ0S6yAHP2xM
8PO8s1kTCHOZrV3epcH+zWZnSHCaIFpM91Dg+50k1WprCbm5bCYMNIdgRsoRweoT
YaZW2jD68HcAw1QjY0Wu7+Ad+RsaNtjZ+IUF94ci3/WjrFGnt44SYqBrtNnj2Ocv
4IQuZ72rZYwEqWdsGbVxzql9CncYOP6lgKPhvwcbzfmNaxxy3QU3CC68bQFWrURT
o8Mr2kCPfkHeXGyl9NBMG98i372JtwfnoxC0ZePhl/WLNtzw/bYlUv9WHTzHERuj
suLD83OftjfD8GdvLjRmWuX9+paYwoZ4ePBiDKyeaACRX7Ss12q8jTL4A3eFytI+
4By8HeXnhPaVe36HzyV7t4+zUupYLESPpgceYbwTUoeW0joDMxjsuOoTSM16ZrFv
uRiXYcp+R7FSAUA9DWpDLkVVTfPmWCuOWmDtSg6gOt01x333qS2OIRDfA/yfxvKS
GCsUddKb9Yv2BMbLVjdfsdiynyeIsYmAGNNyGWJJwsxyTskgFN5z07sZzrzIYhzP
15mYL4Y1LqaLuw4GimTzhdmWkWs3Hoi1MmJTAcnbYzc4jFQQ/nZfRG2b6sqbUgBL
oOVB7YU2yKmKC4HNbxp/MGXw69sgsIzz/chph7Dp7kTZvZH4AhSo+EJ9zjBs0xHh
FKQPFkDz1Q0nrhc932Hd55Rp/qKNLtkToYjNWPpaM/uPoUBFPIhIBROY//sAgxra
`protect end_protected