`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
ddtXksX2+yylW5zu6QL2Lhnb2d1sD00763mmSITNX595NcHTEkwn0zB1Dry37fOW
FufOhVzEJp80NC5qZ/+F0Vk7Ik02dIR0elf3clrjeJRK85K4e3Hoo4xn7YbFUIms
l/8VZSb14+JVGURjfswrIyCUotIzlzVYZ6gzoZwDXIi5gQIBf/gI+KxNXPaKV+PQ
Ufys/12rjO6aI/pPlqSm0hCvftmBcnezN2hk1UeXgOIuKZnogjOsf0iJVX2aOOWE
6pD/psybjbnsNB6kH5uFTA5frkzIzkzl5d9+YDm9OyC+k84E83I/7/j+rk4L2dah
QJOvksSIzN867/4Qt8qYTQ==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="MvBXkzurAa5VTw+1JJ70nePUfoQXBvZOku/SMmg4TwQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
oRtzZL4VJ4iwysPsC8SXYCzXS8Fw2gtZTOskLcDV+1B9Nzn1zTyNtlo6lNICRmmK
ZRVu2BmCc2G+fmzynYlNTnSa7C0Cuel6FYpxCBlOuk3OF2tzAmLAuDyOH3Z1Yjzk
a0aHuoCdIRKv7BrZCdALt03JeUmXKPdOmIlkVGFl8yw=
`protect rights_digest_method = "sha256"
`protect end_toolblock="Jn9CQpRhJt4rnzZPRk+dOpzAubz7omckX1MrFd4p81o="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 6272 )
`protect data_block
gD6l00tciPUa6pDNTk/+t0OO0nC/UTtBwLB41d4inuAUA3i/ALrNyoJVcBnAmEQW
ptbcNp5fxEUJjnOxnedyZEuEBxWRieZFQnkRdF269oOHX+LJHt+ekFVvkumsIFZ+
nsR76eq7yYPVyNncKLyUPa1CO956Y+W3rkSxl36/bNW3EG2A7EHfklgFfXLln1L8
yilIm4CoA1qDDlqslAZgNfyaauagxHAqn+fzgtdREj/pGlTVPy2vlPW5WtGn8WbC
uDzDl4DU4b9zPhcf3tLvTOgCIQEK689x8fyBlMUEPnZfwMnWk60zDSoqZU9Vz6kU
GJaNYn6wSTMPDq2UOMsd498wSdyE02g44EEQRMyG0wHZBD3Xspa8/YBiqO323MQ6
LUhujL6shXMzU8y3yImMDjytPrYHoF8Wooi80sAPzQCiTlCu0RCGIC0w8lV4oUmq
fe87Jvfp9Wn2aRuGMBhIqrgcaBn/8HQ0Avr2S8J5xhaYym2rzmt8WfOIAPavGZFr
eI+Jvc499nRfz+06y5Y5xne79csCKMgsLl6SMOGP12wVWtJdbBTu0cMbS822RfnO
Vtq5lugqlDcTTGEKjIadyVZvEFy2TW4gLoatKVl6LnQ6Yri97QDx7Cjuw3bcfX2P
T9AVkQ10gvobqp5ZzDOE3RraaqGhAx+rrF0a2mjiyPheHe9HYtMLWAmgw/wmtLLH
4+QiMxV4iq7T4V5whgQ1XwDpTdkir/a0Q+imHjQcFAEROa6PXlKBxzXS0Pk2mgGb
YL9fqm26LH5rd/Syd2v5Zun/fw1q0oJbQQ4GFGkNnIoTcKmfQeICY+qCKE3V6ibI
aCReG6EWkRUzyMJGfCN4/hOeY4I25F2oC4S7zNKNtimTwTceQMA6JBAiKhgkEuqx
eGC1zJYifQmbZMBEm7bv+2ZRIN58F/GdeK2doVDL23L5OHOXdoECSwk6LKdj45hH
JZ5dtO+aTXocW7qCPXVOdWJ3jK9o8B0oFu/x2/0tP7ihCUCBQ0kKrf44oM3XAnOQ
0iPfx04pL/rgbVF5Et14eVRUDHg0/gaBuXl1Lf8UJ83keEmz7jg/Tm434vRRSgKg
gw2wE2Hw6xaCa3Xxh1BRGz2xpJj9/dmKKI1qm2XyikihbWKpCQos0vEkbXR37fO2
vzbUU3h5Nsgcbg+s5unIZl9E5xJ31yDJPhkiWmaFZKSa5n+E18lcLoUf8oZejaO0
d28oyRF5rKmq1D2VyrGzfU/JNmOkj0Y+sTZ7Qg/k5LuisaJUhmLR/qLCUspuoBR9
cq6qQK1UqTpdBxbAm0cG7FQlb6K0eXGPHVDIbJGabIPww0ExqUqpC69bDUegskya
50Ov126osVI8IU7qxcf2Qtb49toizMu0vPIROVHxBjTsWkgINBUJtbvCBLBzvmYK
YfbMMPPbuLjTWqgQNVq7LKlNz4/YspMTByBFxDvkf85jKDak2DNETtBhI18K9QNZ
vPlDjN58vkFVOxCszgSDESasln+pE3LlI1pzKCe2Cn9ZiAbhdhYoOTSYRFWMuGjA
/ieDo6WrfouR0jcW2mqqij49EGmagKj+VA2NLmLkCyX0R3w2DVFDCmc21m0GT/oO
VGHSOF0bcfp2PYW/A+hcYwnroDl4s78MoYXi9upoenDnNc4aDtNQUKX4zo+7qs11
KVaGz7Ma6jGM3AlAzBKhEGg3OWcjpD9wzTO6ba6k34GH4kXdPBwzI5ZdOdv0yUyj
B6jFRr5hIxwEhUhhOxtr/iBdK/Uwl9jtznIKuOnuvmMOgbJ8xaScDHq8t6v6Kt8A
cqe3dfwqbP4q2lknqrbhELMHsIlPri/c5T+kRA/ykUvaRQp7rw4EHF8wKDklSYFb
GjC+mwi/DnRRNcXbLqckTojHJ365qOZwnfJnl5NdsUdP9pRxBgOeQa0C5X5hdB8T
e9DtWxCl/qD218vhwxuyrBxi1re/vKVGEB8g/wWd6BVyUVMmFTmNz3CZq0FT2u1H
CWqVh8kRvnTxPS9x4IYHWyToyehy8YQ1Jv+Nyju2Y7NrO07Z+nF6WBLwZ32t2bzw
0lFEvVx2nkjK/fk9OQ2egnt/PxBURo3QkYD3JJ5QGjI5ZohblbA88F6WP8XJR+QT
8hnv//WIKWkTCXoGCFxMQdEvgPiP20ShRL05J+hodWyKgIAaaOKSHxvshWPfHFTX
6vuq7K4P1d7D2LB23MFEdOJ9Tcrdweoi25qGhjc4MnxvcPFjfqWccHYVAOWKn6++
xpjidsepqfLjQ1IIJMG9c/KuH3jdRx0NqdRHzrG3c53Ga+W7jYlV2GiisFiKp1LZ
ajgyhc578PuRB4WTfHuYwo/8/YAliU76c5Uy4OVgqLmOpAB7OjCRrQFIhrZiu96N
Dpt6fDWLOH/0eqetDxS23EBVKF/NyhdniU7pbS0aR0S/lJ2diQGOuWsWkQLDp4tH
/w3SdoVh6JvDOnscDP7ZI+UJD4YfrZ3ZYVxl5jC/u0M9bqPCPxwAo5E95iJC9/6T
68+d+JKqvAlNAtDKHoXgk7DhPa2IftirGDg5AfGK6djal0QrGBCLH9q9B/8KtirI
KOORj098RuTTcz7Jz1eHmLnfq97V9ucUXfic+I1hCSPH5EoYHSBJolSavxj+6pWX
nBDc9L12FG979XgHkEjPQFAd0dhg0I/qxt71Z2bRkDeGwnGqcO136KhZ5eArMkIb
1e5OvZqrb99fLRQmeqN928Eql1+4Sdl/aDQyIfFhPK55G9YJ8AJlJqYaqMSY/O5M
DzYIO9rdDAb0gQd/BLokOStGCeBS/R156stgL9VJOaLj8NU3QmEDzNlhv8MlnAlH
ujMNBGDYNffNiikyIQn6FmTZM40EF4y6/ASyfVs8CsDOd5UmlZwe0CXUYdgLmFv5
V2jYAmneqcYytK4RrduJm0QSc1g0YSWTSW3FSAqI0mihAhhSmiHAMk6BHr82aP07
KxVSMUcu8CUK1HSECjHrjz29H1Nt3WC+8ho2V6lS8IxFE7akPI1M78XnnCefw1Fe
u2I65GpexDRezD95dzxm1++j4IUtAxO9C6LTP1Uy5v4eTmXw78+j2WuNL1mKi0xv
wcNC3ztHV0yjhQt2LMQCNTN0+CfWahb/oFq71xhIGRfQLvI5Uk2/b0lzWSVjloub
ekScPDt2oyN5V+lDiAWmLX2tFvivGT+H2yWQe7cVkESNkS1W4JCK44IFBi8+fPap
U9smrvwtYxuy3V5ZpNRi6ScT0ISWE2t0fGpAO+XRJJJROMIanuXuFMdl3gHcWaWZ
ZRYCCpTWjTYNHP7hDs4sm8Vnv7OBerqVvA+2nx7ZUEaxaN8AGiVlo8Kx8Pr9IRxC
/ggIx8DNP51cLia2iqFpymapINaRFHRNirbKjLlkccMDE7kXyvhTvIkepCc8DT8v
r2Kpz11li8f4XZlx84tk0/DtKDvOc07tXk31EkCA1UsUkDu8Zb9p7hiFriLcQnCC
4hMb/RWmtl2iz/7ldDNyv1MZ1kCXfsgK/Hm23ofiW9DkAdOIT3F/cnZ4cLab+OpP
+hc3nc7Ax2OvL205fEeEqXd2yeB6dp7eECdY53JpGT5rLLB+C6lLnb0DGfxjuM/f
/b7H27xZ8HYrQvupDreeFHkyGL0thG7zCjVxehyZCHAp1pmrIX3P8V6vw6KoMxwl
62zqAfiACp7JLkhJT4PFWDW6fxompJ1ihPUwcxkMcju5KmgtPy6Gu8lvZHKKto9t
mGaYM/MCaSMVgcys/Yd9nZLxXPxCRp8s2/Ak0ght0OEL/pgUs51Lwc4Z36JHJh5P
arUkkV+yNrttHntsyYCNcVeXa6yITsQBwNcXcIvnLAWP9FCEHigAQLfCAeId9YOz
SeD3wWPbKvurnpIKEtrA4dlmbQVR7j2llXSo+UCXzhPceh9HIJyPubOfuwa7uXpn
wdgHBCqSd6UkTj3s9+AqeJTHU7/lAXT4TOWZU+Oh828A2c3aRN+9IrBIo/VMvcBf
eW6gC7Na2T4EZlCCwjUCDfeVMQgKNAizC89n7An2BeZrGkBLIPYrhPMrUtURhhYY
Iwt6G5i3d+xb7K/Y2N8Zt7N8i6ie8EhtxXv2NOl7RMO4pHANC3zoxp6OKpYp7kLR
k71oddgSi0Gu/HMoegy803qZIVPD082hEWN6xfmRO8VNGXG8nElxH/IABU5+46RE
EdaX19YexFaml2hKvq+Qh2Fx886n92UyjnC6vlbGb+DOBTGmS+3D1JbiTpcwM/18
oLWxKF+dHRXMar6sKxH9AlaloGyxw6VHWZ8DU38Ro3k5d7oUUF1KFZWcmmJ5XHAn
T2d6YRQra+goC6+gl4U1kCOdtyf5aCEf6ttHp99MKasWceBI5LnecsKBET93qJqD
4orXmNSff9pqc3jn1dzA8Rb9aZsN5mEdRfWeOPzY+d7vNRFb0YOIDXAQ8FKHYXGn
FpewKBD4HR+Ex+qSy9jJyJU03qJ3ackkDb0tiqA5pQL8xqV74fJSzuFxKj7PR+6+
641zq1STsFriSjxl54mpd1r18Qpz7qBrvN9VbAJjKM52PMCcLvk0Ip2n5yDmQfo8
kEBgZrEkNtfgcXVFA2ANXrJkVV8Ak5jhBzbg6Em8X1v6TlaQpJQd4fj2hwvcvv3R
+1Bwr7inJL9ZPBcyl/8nTcvACz7gQO9b4OIw3b/YUZ++afqbY5cnxdnJVwGqe1du
WPH5oMK6iNKI807cL1R0nNElLjFyWHpMlERU+aJhZNkcJEE8Wk15gwOe2FJy5+iI
pEwU3Y0qkBFrl2nm9e/vgSQEf/cbhvfRLmwFt5jwL3Zwbvqoj7sDAAm6vfkhLswZ
m2fMwfhCauO+Ftlt4NZVUQ7DqRvBg+pbGC2OKEWYq0py/0u6hpS5AXYPwCUVrjy1
OfAP1gljzMmmofbo3HSxbcOrPEDJHu2APWBgcHAum8E6iJTqfH+H7iVBVaq5Sxyf
SL5XqVMO6m9YWRkVurZjze2lZQkWSCL1+dptj/nMHHY5y8vhIDGNZCqehT3bBqpg
pk1gLsAOZhKsN2OEry17W+Z761AQ2FLOpPo2m+zCo5N2+uD1ZrN+Lj7qMsaU1c/k
Ce5RnWxgye/uHD9wqsvdT5WKP7AOyIW0nJdpOj7vOGQKvqab8l/FjDoscA2mYu32
Ess7v1RATwXK2tf9UzVDOWU3DzL/nsnlUns0HRPCeZJy4kVHhT5JHkByi7ooKa6B
/QjJ1Pxwqp6I9WKR+sekifCG9D9le8rBowKBXdD5IxmouRHB9RZ0u59ZLMpR0GV2
ivmp8BJd54VI34JS0NRLcq7vKJIJIYr8SEBxd6en44Q3+xMZ2IQK/Ail4pBzVphi
6xWZY4cHK9lrJmzLWcowi92tJWAXchzXpdaXwGc8epxZP6Q9/yprB9OtcgCJDhH+
s44LOGOpslW4SjX0HaFm3PG3lDhsE/GhAV34bUdDceXiMBAOEV4sSRZiMUmS5l9h
YS8FdElRCygo7lYBtLyDyHpIHQQ4quK8X2jEQwi46xWnsWVpk6NK/75RWnPSnVGa
AW3lfQih9yZ/xdvxrjr/UZMwoMzffgWmajDhX2CdLUjXoKdwT5JuZQBAQzn8mSux
nq0lxXASWmtkshTF5irAxomxNApeBnRdrxRqbQm1PWw60GtqSRapCrZTEpAxsT3w
yYgsoFXNWoV6qFPja3kZ0RE0lydGqcm8v3Q8uQm0rVr2nCv9tSucJuCYFNy83VJw
ybwrjpQyOugezW52ES7+6tli5fyiEDt/4BWT1vq3jZ2MmSsDVJ12gT+VGRmQ3msY
NvUwq17X1ubpBWoZCaGwek5HiHtyU0k1Peh5fOm/lqHn1gCqng5RHFSGwWs8slI1
W0ZUBcB/DqoMdkVIFFljm4zUJZjBT7q4p0bNqL5UDjfDh7GeOj1IMtk7Mj5GtVqU
Kg3PfupCzG9l9r5pSs0p/4m5mFBc0xLVmQlg11gz8q5vSz8r6R1lqVY3aUlsCQgl
W8KXH0TEU1tip7WJdT20uhKZymyn0/xxPP5YCMXCE39rgyjdThp84KxElc1v3hKO
KrP9bKi8i0QZ+G5VyPbXwRfls0dM8WL5KUAeJgNMKJN3pXQigHsQP7ZxhtUgJM8Y
TdqZIwNg64hRExy4ablLqSJ4P9jgANbewZhDEFSVOHaTz8doj1KFlz3Y3jKP9wyB
kE1sFfyN+KZMYgYYBsRrj8DAyD/5JiiqOTnpn4VUkRhKSFNACJG0XJ94i3i4vzBC
8jHV3T4dEBvGv7rzPSpbnr/r1dqKfl5ptrYQ+/hlaJ5OBaMEmTwBLIKZ4aAgGfqm
GrEDBgVVWgWg04kM1CPVofZnuMqnQ1t59790JvsDyenxUYaMriUmGo5jJlFVsbBl
ZKb0jVXQPKyTIxZNBVITxPAoVSOLDtitX2QOAV6350nQg+6Ah4+2c4HdsnzoXztY
MJComvj7KNRWwWfI9Nsm+AptaQ6QSrz5cEykPQruj2Zz0Ct04mNmjZ+TOMDFpi14
1bB8lW3D0XpGlzyqydnZa9tUsz2YfFVeW+L254LXvrIg0GKaL3nPrfkUmb8aa8Jx
4uKeL0i32DkESgLBc7FVGDnIVlw+XJdD3cHfiSp2VcAYiu6vFzOhv73iLwQ5Dvpf
n5xGkMvZkD92vbAH7C+l9H9y2/LC0KTkT90OVPvS19od5gcw1x66RsePMW/O7DO8
hjIqB528Q6Fl2qkPCVwFQycrAPeL6SPe9zKSbISG/Iihw2XZf/0FKFaJUIYqoUKw
RyXLDSWQwTiGOWDKyipOJERPLBFASc9UsZp4xD66rGP6auMx8wGtqaGIkjmwVPLj
jEstVHp/lA0JNSrNUste0TiNMwbwVQhNLwOMoPU9UtoWH5cjT+OyNKllK5uAsmKp
iKHEVp57K7BPC1kpqEWI+Vl77TIlQBR7rVdB30OnWCh2HIs2zY8A99xMkyjcYD2C
royLOmjeDCt20CAgbW8zgEIZg6j/8H36sdAviLB2+QA29KRNqNIM/4rJTWIlFHZ2
ImivDzEaPytjNpmlL7zDg12Or5Q8EincELObSCPAV8Xd79i7v1aOW939A18Qvfga
dNcZzahg+tDLKcw9Cah01q3mm/fbQ05PCwrIlwDfSL0cG+pspav8PVQ6xJObZNvi
MrfJZ9OWMP8ovA1WGHC7n4EhVcDGxHPAQ/eoLPQ6rgwx+EcV3Z8A+KZRZW1gdCQU
6gnMN4z5vkKfqNTRSzTEgernzCheDCz9Ryar/NjWkon3tPxmClb7UVYbhEUaRSSm
JColZCoJ11QCh47K+V9TQpnQpg8esiqBrvF+uDN4qFL5zo9c/s3Xdpq1KyZnqNH3
r/Ja9HaqzA74TtGCnP/rZKcnfM6d5atUODeNbI89af8yFrAQ9AD5pva7VNba+oUY
GVX5RWLJ+P7tpl/51yrhKfQvUiBySqHFm21v1SQpXmIy3YkZnv4o44zcys6ZtHfG
pR4xpaWfRn+U970N7tXmt+kW3Kl5tFfH+g6Sm7lPPtKJbBpdAKy/aO5jxRL/y0Vt
ExoaOj+PhtDT9GsqwNErBm7EXrtA8HoGmXjiVBg0oStEw9ycGOJ4ZIl0AVf3EU77
blDVgBHEREJvVyx2FnjsqL6rmNGDfzsvi7yOEFM4nC8Wfuumd9pAUFcbd7GeH5L4
TbK8StmtUMkRNHNzFEJ419bhphLiwsZNkdvoea+ji67lWJFcAnJBZw0UYPdIGsfA
JDW+W4KvaZ2HyEQR1GWsPY4sXP7HRxBawn0ilitSEtELxqPahtKNMYQ6p2AvZ4kA
ofaV1GtNIQ+9nyooThR+RltQSP+q2gptWf/Wmj+TmpoZTmq0uhnZZOa3SfZDrRkx
XgZ/qcVnN3I3vG2P1WypmMaUUf1/2mb2fkihMk6Izm8X0dZSivcymIN6u3TV+T2j
3PEa0VbGUAqxP38NgP3R+uhlg310MoT4xYQLdDBGC4WhzQjiXeeU+fqaOqrRRbPr
Tph9OcdC7LOaSgiwIu5JfCLC/RzW8oB76hiNXBY06WfbiapFUxJZF3Glpg8xKHfW
/GKUOnx8uCa6AE61WHWxhggdnCFufVNAplhOMJiUta8xrGAhyNM5wc1CzQ4A3e87
U1IDmqqYCFnpixyvYEZww6ZSK1nVDa76rZkTmOaGFs2SPNMKRiAW0HSm0CVQvFlV
6OEbrGV482CX0YK04LT7o2nfbVhRQ4S4fvfeb+j3vEw96BGeFSiiAXpgC0sOzWdC
OqC51rTXpha9ev/0HZ8t4smUYQforu3o2dPIcoRW7PTdY2oXlY9zM00nqeaqygRA
z5Xk/OH03pUOGOYoDVlD/+s6VBpYnEqOCfvIdVtMzkQq/IG0OIwtbuCMlUM6m/Ec
u890yPRUDbsHLLlvG82Ac/Xd/txDEgfO3oVWVp74ZU8=
`protect end_protected