`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
ddtXksX2+yylW5zu6QL2Lhnb2d1sD00763mmSITNX595NcHTEkwn0zB1Dry37fOW
FufOhVzEJp80NC5qZ/+F0Vk7Ik02dIR0elf3clrjeJRK85K4e3Hoo4xn7YbFUIms
l/8VZSb14+JVGURjfswrIyCUotIzlzVYZ6gzoZwDXIi5gQIBf/gI+KxNXPaKV+PQ
Ufys/12rjO6aI/pPlqSm0hCvftmBcnezN2hk1UeXgOIuKZnogjOsf0iJVX2aOOWE
6pD/psybjbnsNB6kH5uFTA5frkzIzkzl5d9+YDm9OyC+k84E83I/7/j+rk4L2dah
QJOvksSIzN867/4Qt8qYTQ==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="MvBXkzurAa5VTw+1JJ70nePUfoQXBvZOku/SMmg4TwQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
oRtzZL4VJ4iwysPsC8SXYCzXS8Fw2gtZTOskLcDV+1B9Nzn1zTyNtlo6lNICRmmK
ZRVu2BmCc2G+fmzynYlNTnSa7C0Cuel6FYpxCBlOuk3OF2tzAmLAuDyOH3Z1Yjzk
a0aHuoCdIRKv7BrZCdALt03JeUmXKPdOmIlkVGFl8yw=
`protect rights_digest_method = "sha256"
`protect end_toolblock="Jn9CQpRhJt4rnzZPRk+dOpzAubz7omckX1MrFd4p81o="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 4672 )
`protect data_block
gD6l00tciPUa6pDNTk/+t0OO0nC/UTtBwLB41d4inuAUA3i/ALrNyoJVcBnAmEQW
ptbcNp5fxEUJjnOxnedyZEuEBxWRieZFQnkRdF269oOLzSg7Y4Q64FfThjx1IrSR
5NYepOwSZkGcwTHnbXRYVjBA/Ncc6tx4QiDxYwTd6qdM3E1n+9s+UnUfAVlYKLwl
QS++LcQEhC6rZ2bx+E/mkdhtsTrkOwUv704Aejkf/pdJp/R85mobzQHl+5Cz93kz
R68maJsc6Um7TDoPKldERYUPQ7JeMcnv0uIqohi4C4bTtv8em03yTF/3QTjhjJWf
g43YY+pDN8JsLk71CUOdgm3PZz6rFzgfrgx3D3HSPGjxDzugvHLxzYl6L6swDX8n
BglO2Q/t6F143QiR2ND3iYE1aqOadZkoti2yVE20czxNoBha7yhKh0IeFWnEBz0a
BM0hG41VgnuAwbvGfR5xjG2xJzHy+OKwoCnWUudbp3bfGnSbwgWIrhmp51Pzd37+
3yjAHiixc9NlTqOVFzvd684wq68qDXzmBgCxHrOOTC7YhbKqw4WJ5nXsn65JxSPb
5INpJo1pxE7DPEY5FRSktmpS+UTkMy46P58m0RMP7yeSRbajI7RAbhwPQ8BRElm7
s4C9DuqB6fmjc/4mKsTL9rk1uLwdfFpYlv/ZIA6uKXuRX6x013k2IkSZKNUn+VLs
waMliRclu4F3rYhYa7QV95auRfkmfLkbXwXAHXIlU4CT2lRBfkCPb1SGxF6r8xkA
m7lqU5rNjby6B1L8W3ws5pUvlWN/K3kz0xoW8tzunJSvxno14ttqp1gkLQ6zebCn
k8VrG1pYhAHm3Ogteng3fvt2Kd1x++dNfnu+ZQ17NlOlCoq7jTCuL+4IXlllS86c
yGoVquhfkuUDZd+CMi7YmFcL9wzGju+Q8OZV/w2JTDwy9H76uPVgr3iqAADfuZlv
iCQABCrhXyH+ZyCWZ+icwNuhgx++o5qTLVxr90SSVELDPM9WcvaRT9P/+u/4VuHq
/6sCGBLIilZnXaX8+ou4I+dUhMkrzDLU+C1u+9BE7+odzvHTgp4yyRv31ajRPwQQ
ijG+6eX8dKQqy2QsYHtDAEknbVS7V/QloIGPg27h8SnS64mKZ/cLiYHz/phJ0p1D
/edc+/Yt2Pfb1Fc6iXKiv6pj1j5TmNzN/7+tGEiRfQ85PFMChRfQ6bzNSn9TlxSp
836ihn+qSku9FJnmPUQF0TZ0QSSSOt5TgE9WxETWkoHxygooEDgXe4wXkTyj0hcW
QQskkLn5N8t/NimhX/nyyIMIAlpBBcotsE7BOxHAuABP4zgHcsL1TiTQq8y5ckJY
YbIZgT8bEP2bs4d26EmhXKYMzgSsqLyyAbP9O/Vddg+mO9pCUjbglhRm+J5lpDLR
cyVTGiptvQM0U7G/bDbFzV62GdSL20xy0SmUTCM9TO5FcBo9bSveviudI7V8puLl
/OXn1NueGZJeCpOxubJNv8FhBwCmDG/9qotLKb+/mu2xeJ8TLkGe4Vvvr/QT2Dbh
NDStaBONqCMj1V0EJ8el/wQppcYiyseyOKft0IhVtbpN42MXJiFIu00btnzCuVbX
DRVEDobvgDvA6jWyYShYBZyiLt5Pb0DHGsqTp6/wDxQfZu3n1iTFRhaQD2EZec78
DPKQuh+7FDLSpTkv7eICIQURGgfdxIi2+akGlqXlrChsPtAts2aYQ9ruoSjTXBJ1
/oRio6ICC6h/TWkIQiZGvGR405pvODAMz1etJcOSfjLd/7N7MzEwvVCcmoKsMzF1
PaILHh0+nmU2dksxAoSGf9+6ZtIBj85fJ0pE7wO4cOzMvXmM0rvv8FpYcrZy4NvK
qY28AEQRqdBWBiwvcnxts9JWmm0nZxWhd3aL1dXxsAhjR0AoyNOyil2g+8vOqntS
wcfp+BVNdduzxpF/r5AgHbV6zhYGU3l448zkTvMMNU2sAIDPRwLcA7MK1JKF+Vni
E45SUA7kyul0BXOoUpIa7keAm3Zu2Oq8X062wpaii8d5vOWZnoTRnxZtLNUQxrDn
ewu4Ijp9PGaCUJ4++bpc47PRvtBUL3d4rws+dwTqoXYNQWJYOGM3FXZtNw4bbavU
aaJUXAms/8i0hPEN6/T/lPWFuE2/WhX6FhPoNS2vFSVRL7xZle0z1FndKD0Io6mt
pjp4ChBDcpBXDqeQzOtZkthjXbJ83DpQNccxUOIn8M2zywUPpEpw+8kpGDTIaHjW
IwxjggMCkivyuaWxW39VrDogRzZKVDG8At3lObRQ6kApfcqClXv6exdnIESeKwdB
H+VbAZhpbYB7RVrF1NVm8d88V7y8i1aODpRqtKOhz/uZsDKK9pweK4UkTKVXM5yS
n51a3rnFPe2iClVsCYyWIdNUY+1QyM+XRE9q5y7OjQsKBuziyPVHbw0J+wKUvPM0
RbOAgLhvtOZjgKHEy/Q+u2sDI03JdNDDG5PLKZqCBMAkqiWe3/lJWilTUWi7A/k7
4a3fnrZJRBA7jD4bwMprryLADqF++rEQDvzGZqzclceX50h00cq9oXGaQ32rm/bS
q45TVdH7vdhXOZPVXiKnBhtkoILPHJ2PATLLAdkg5lENgPil/iWFGQdhcxr3dnTo
dPjdAU0gL/K2OEC5tY3s/yDgGPtAzM0yXVqeEfXcRHIUYqTpxuJ+JP5ZpvuwHbjM
JCrE/NFFpBEJrpL80Oe8LoZ1FhzNyD40EWfOFiFBBBMO7ZjO6e0HyIoiikujFLUq
XZeDhAxdCjMUBS3Wy5MCzPcScNZgOp7F8WUMSa0nKBLXd3jx9FYNlsAvzJxBZdRf
MGDKxnQm63gAEzM3Cmi0tJuEGgZUTa8Lfpr0KgBLTmskXIvQ1MXbFVCbcTU7TQlN
knr1PNDiGKbZ8Kt72KO4PNLZIHnuJieB5CKGtRP4ckNTNtWCFJWnDNUENiR8HXfE
zTLqFjzyvghH952WHDfpjHeHOpm9S3jg++JaHYlfaVAtIFxVEzoZZ275a+Jo75be
GJKY/0JWGqKivIgwFn9C2M8f8GT7sNcUo67+gow+kIoJVvMtTbwYOdavK1sGmcsB
mU8uRSqGB2MyaFfrBJ/oW1OrbrsOaDVy22Wq03w5feBo+c96JZxdPhC9F1tbHWs0
dX+deWWrsA8omIDplOMbzci4Cw3VWKZHUVwfs21E3x0S4/KeDoLIr1+XbzqB+w1b
wYBfqyH56RFj8emH0/nCDYEeg9NDk7xlGbVAJwMS2ubmsdsXifeOSC7rz/X3lBbt
3Gd1IXVa4r3DSF6WCipWG+XCTiAKxPBRWfb9tjirmqwayxU6SVB4PqrVu9E1oIjJ
EzLZp9eYjt2BP7F/QlF1lfcp8IlqN0X2gJI9B64owjtEkXhhyZtMmeVg1pwKGVg2
Mhh+hN9jQzvvsx6Oiz6zigk0hBvWo9gZS2zahov53gkefK3ZTPZj/lXzrJqHndKt
q1z9Phu/uKQRVTkL3eKNA3r5yfvvGDNet/E3zlYUdKn3NCNLCjk5pIMh1FBRRbQW
PhpzYaZrOEzviGy+R2HuHOpz0lPosB88ZKEb9a9HB81JyD4IAx44ukyV1LIzmC3d
INMMjdw3WJtcPK6AWxO2ZrggCNMufMxzD5Lxs4AsQTM53g9GOE47AFvN/lfGIrtn
HQdWQd2zk3TTrxx5hb4OOx5HtQbboBb8giLMh3BQ6ncAIDfLY1vlp907sIPaj/bB
LqA6VEND3gPo4WR3s9JZ7mixZNEk1lSDNlkOTnj+Hbd7T3ElREjj5LLr4E0RKEvD
/MjUwGD4lo6KxTK3iVZbl03T1AOH6umfbWwxD4GuoDAtc8nEQK8PEa7IPSFJ9tOM
439dIEA1QtP7xlj9HCGnbBOQiIunzMDdfngseGQhw6G6Pogc48aJ3zpxhSO1Df8U
zZZA2iPf8IKc1WmO9Pzl9tmD72PS/oCdmzXOd+68MBF5t5sgYBRCMzYB0Mpue7yd
hAtZv7WK39eCWx2wCT5wxp9OkIiqtgbDFQKyZ4kw43udnRm0MYS0wluzWa4y8+oH
CsuvyHlQ+5G9sdDzXtPoY9i/Vql9e6ia9UXO63d/+J0h/vNrXWRRE0aebSsy6Y9v
lmI6Xp5efxQJHwHO7SIVugGs38YE6FCF0swhQD+UYdRsqZ4nWe4QV0xNuqsx6pgK
3D3CaXjH6fT70B4ECph4IiV6Iq9HN7/1424CjDv2DpbZw3c+5XsXhTec9RMXpVMm
129LLNAH//3XB+2TrG7cCRcB3hzqRKbiNrKbrOA+DeiUiKUkKOxrP6sPLyHMAPDO
JuBPcVPLuUCK62QJ6kXWB4fsqsViAW2rtJL2qguHx/v9eT4cHIfPcpfN6GIL6fM8
rC9JO2BB1QHEdXaou/WsSFQhiZu0mRjqvMUSNBLxH0eeQApM3BT2qvGemv30Hzv2
YOQ+oxybG4YWTKOn3ZcSmOxZpHXX1PMbj6tugOmbfsEJXTbp3gLr4MPyYzitn4FY
ofFlZjaVLOsPkeJITmRLKVaEdpEWK7KqvqA2VYwhs6Ba1p+kfbvRIAPiFvdYSl98
l7OBdsROf0BseRCL1sSY43gXtCTHyeO/NaaBHii/t4QmKr3uyNFA6I0pH3Pel+Sg
G7LwZsgMFu+XJCL/O2I9RBtNhTajHa441iXD4Wj4kGx6A6z+GhcA8tgx3eBY2qQN
eUtFvwuhiV1N7kaNcLNOlcYjdU1lx5KSMYWJLUSkWCgS6IB+Gi0j6GuzQUjgKuxk
pFx5yH8OT6c+nacs4EhR2dB72K3pYo6QFHZ5Bv6DAUdQPAISouwM1i1SW13DS4QZ
t/obWvGlkd+2DuM5jV8cgqEE+HwGt7THk6xN581a2WjBNttTjyGqmN1VZ5VBMT8y
s+uATGkFg7QH+bAuv2mb8Kjvp1cr3uH5Yn4syBA+XWcELenL3PQ53YFuZ/yA9QS2
Us4sLtyPqxi1X/UaAfwNd/+dYGCwS1tgYuhUXH/8j9cnFuP9dB+E3tNhCC+SBsWv
zz/HBoYvULctVTnuOIoDsB1bZ8lZDaSq23VnonntRUWZDyc1kvGsGXNUw+fCU48e
0r0ZulVOzzXyHXLF5pH5PVeVbyKq8iLyicbMdtucVouQkfmRnqL5sF7BXABA4jjV
0nwq9yTacjEr8XyWnJ+8T8KbwoWzozAQNt0WLHTYGZ9r5x0Y1SdrAXoiqcfOFXLT
j3SrEhxPSNumScb7uXUfwEj2hb+uJQk0yu02rmP43seJbMu2Ay3Ksd53XMXxFQi2
mYx4l9ncAl4ib4bEeSzs4p4FFX+zORtl1VW30MMf9vYyWKPgVI7toGr8L8F4kTtK
7x1SAmlW3VGMM00jsYYRL8OqyVOaA14X2YPeSP+GrNPKGdVAzDsgvuGKda5xyCSP
UsTgIjjUTkDuh8Vc5kFmzmkAYDNG5e+dQ3Liq5cyUSPdmG3bwQ+vopvxCEeRGbf5
1bn0ouhO1O1K9np88k0A/mKDgspBDzZ3GkyCIAmjGuWvp1a/48Abd/bU3tOgRccp
cN4/VtZJH+PuCKPhE9cFPv4TZNEF7+pDMrjDaaCUuc1rVB+LhK7rXqbJSgWND0CM
yEXBwTVUiSFZSC2lO/umV0EBwIwoVYJqMsUGWa6DE+fYLRs3RS7M7nhRtM/c9F+v
iPxE+o4fOFBSB1momvFbt7CFLFK+i4zCYtj5WIHvRU041psUhn0xRyOhWudsYLJW
IqA8wYS9XaFo/M2O8EQd4qD9GmfuViNzwVh4keJTBS1rqCMMq+K1Ul19ca4M8wb+
9CwWh61G6KnuoxdgNRvwcLWDByHGlnt/2Yh7cP5tcJ7kffSlxa4+QZi4qXKNPKYj
tG4A5isXGPuqNgwPzA2vS9ydWBVbpwPQ94T176wJ7Acz6Zm5WSF44ZVuM8wAdU0y
LWNdqsbRH9wsS+i88a+gxnOXUpWICo6GnaSb9Q+06knTL2kC5FsYVTS/l9wkZRoH
bE4pOsDVG/19JD4lQ5flBB4L+sAlZkrfuanBh7sS6OwohcwfoIC62RlL0lqYOiXJ
Zb9q+2UCMFzHpt4ezp8gyNvmbFS1yxQRsvM5hBFMFkuDM7QHOHs6VcS1sc8+5o7e
IvOFned5IMLsn2lIDmBNLmEHDvswRFfI+1hchjFQl3RBSBbrbFrVWLUUlIB06Gb+
CA4+C/8hPIedCLn6rr1uHhXKVH5DINENQXE6NnM0x+6hB3zyw4qAtQqqUAkZx6T9
rXP8yTgSjuhBS32MMY5nrg==
`protect end_protected