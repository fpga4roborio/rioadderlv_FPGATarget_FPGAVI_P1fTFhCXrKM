`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
ddtXksX2+yylW5zu6QL2Lhnb2d1sD00763mmSITNX595NcHTEkwn0zB1Dry37fOW
FufOhVzEJp80NC5qZ/+F0Vk7Ik02dIR0elf3clrjeJRK85K4e3Hoo4xn7YbFUIms
l/8VZSb14+JVGURjfswrIyCUotIzlzVYZ6gzoZwDXIi5gQIBf/gI+KxNXPaKV+PQ
Ufys/12rjO6aI/pPlqSm0hCvftmBcnezN2hk1UeXgOIuKZnogjOsf0iJVX2aOOWE
6pD/psybjbnsNB6kH5uFTA5frkzIzkzl5d9+YDm9OyC+k84E83I/7/j+rk4L2dah
QJOvksSIzN867/4Qt8qYTQ==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="MvBXkzurAa5VTw+1JJ70nePUfoQXBvZOku/SMmg4TwQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
oRtzZL4VJ4iwysPsC8SXYCzXS8Fw2gtZTOskLcDV+1B9Nzn1zTyNtlo6lNICRmmK
ZRVu2BmCc2G+fmzynYlNTnSa7C0Cuel6FYpxCBlOuk3OF2tzAmLAuDyOH3Z1Yjzk
a0aHuoCdIRKv7BrZCdALt03JeUmXKPdOmIlkVGFl8yw=
`protect rights_digest_method = "sha256"
`protect end_toolblock="Jn9CQpRhJt4rnzZPRk+dOpzAubz7omckX1MrFd4p81o="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 8544 )
`protect data_block
gD6l00tciPUa6pDNTk/+t0OO0nC/UTtBwLB41d4inuAUA3i/ALrNyoJVcBnAmEQW
ptbcNp5fxEUJjnOxnedyZEuEBxWRieZFQnkRdF269oOVj8mimwnGch9jLKSFvLpe
pvGFLk3sgNSM2k0bSZ1D5LZb6QEyE0KYEenJtZ4SxGNJXG4KR+XBXOy+9eKSYA4N
EPXJFXe+4yvZsZy5vR75tn0MOa04R1bD2T8DCvI0c9TRy2xTrzqV1bPT0YOXnvQ0
TcoTAUJT5YkxTDNJq5AKRWqET2AUDfOZugVvcC0VzsmLRnx3VAmd0HCJRbDhTDny
CdREqB51kopO4FVo9bseZ2uIRoOOvOQhhAtO4SOICRlYImwrvsjxR4f9lPNXNddr
2zWmFtvf6EIC9ftDm6DDLNxhW3jInDdH1hH+q7ZslCDA7caR3NGTTcPqNWr9Ht6w
wczSomfBNreWtyTqL1+gZ0R+f5ESsmf7Jta8IG2P+dm2ooJz+5HkZALtx5OieWBY
l3Wt4/SaldpFhKXFG/wjO8cR1PeZsXGLwqCaRNNdGD7R/7QC+JOUA+jzPVo+gkCm
8ZPqhXB5prG989lTPdxOEh5SGdArUE5QfRV/GstnPdwAiuV0SlACL7cjyXSLINfJ
qm0HSekbpzbsRZT6LbAMD8bUljN3nN366EDB9VImp90aWX9oHXL2XkSb2MmsmXP3
zQITfkRSt5RPrOhnLhAMfjh4DJ5sAi+r6xyjvzjnio5Y7V0mDwG9rs2rcO76BonW
JkhRAcGnPu7ljDbvZBwsnGrwAUnF2vx4hYQveAVzfdVRzw3V9+o0phl6soOGT6UF
usv6Flyc6Uu6QvlXiWe0SsZ5qQ+EU1yMYvrWJEmzH4SWil+F8+YoJ29pAr8WBgDh
LCB8fQ+cGTeQeI7bW4KHfWUhFEeZ2Hr1NqBkG7e0F8jVn/clDFetosvjPxW/0c96
kHPShcWID2gYPvAc9bbQl9JcDSEb6gt19YMCOF970OPe/2vVReniab3we4OsVk1g
GSX9I5JZmHK2CdxLk5CHI/E2rhtZwJ9NLhL4G1AT+Su8QoPVj7z+77N/0dsnHSns
sNWBbRVbHVMPMLDKrmzU9AteEOm1nONN5jJOX5p1eOHCW0R3YxQKxPiztDLeGCTL
Hk7QeSitdjUSgz31SWUd5ar+oI6f9t9hl0Ot3AKL/E1un5gGdOVbowV06LAvDR+L
4FffLAib8qB6e2PwSBaBgpVmPbHwdZ+FrYQzvu+6CLVRJvqW8Q5IZoAV0Fn3lqpX
qZoiEwd7SwW6HHQiDRAVCPiOik640DvoP3VjkPUsOyoBJp/msAngXXZriEu7T5le
ZqcSX+XF4/Drau7zJoPaFBgFj0N+cjpUV6+69U2QV7pAOwLEH6HwVY0J3tZ6DLkL
boczPNnoAO6RWbRRmO7uKumYBYy4BeW8cb4xLXfTI3CEO2fzBO4+/2nMHq2kIuwv
jnQLDZKGwFnEe9eNWlMv3Rlk/HGS9lEZfFKrQnnsHmDYVUSp99HAdbTz64DSDVO6
VCiSN2hl6sPmEcusHgS/4wg4yo4lw4L3/xdXfwaoouyqA4E7k1Rfm93/LIjzkIpU
giUw9m+1qMhrSpV+1yDTEFDNjTYlavRdVSsNQ2OdUiecZllMMiobSxeGyUbyXBLo
udErxy6Tmo506qWhk/2D7ibMnFePM9JUHio48VJYf0YsZK7dgHXSWJkG1YyTwEX9
824Xkx5caHGUqfkynFiXrzpBerZ31Q+8tEEthgnfY/FJkofpNe0JH17vU0dq4Bge
isiFZfYaf1ghR0Qod1MwRSGE43KWtbTQ4HnVMxXHxWfhtIMqD0w5H4BmTwiHYRrI
eLXMGdH7EbKAaV7ekCzzJ2geagoa+5o0gz+YZWg8f38fUAWyc7HN3b7vynYoQYUW
m//F9qCgfmyA5ydvI5lilX8bfDzz/j2SjUl1EL77oqTn4041/K5ikuGGSJeHWw9t
TaptdT/wnuM23HIvtBVhNnG0XSf3mXeQlp6iaMp5HROLiWg+p55JxZwC6NWQAfrp
0nbKrANUBU+ba7T3YLWqiiUQggv6MFAAvhxJqvvEjRpTjWJPqb3QyyL7WSA+fqzQ
5ad56ZdD9usBsOes8Mn+WgFcnLul7bhm8eMzzmYpz+ukfLagqhq/ocF9hoSSSE6k
bo+BVRqcZgEFld6zlTUOX2O8EkMSoprKKgr++lyqrRmNyXOdd6nesFC10bhwihg0
FUeqXLRWcxz5n9uRJ9hU73GJztsLShd+BHC6+4AEfEYyBlt8gdNoSyGZ6pwT+3z2
f23NvbAkvHW5LAvcq/mG1uAkki/SjztAw5qoRfNVFKl8bUoTe8BmaQZln4p06fSY
tFbU6qIVnlC2+D59xh+m/l/P7XrMlguIfg7AqJ3g4QxtPk3V59M+ZwzM3UU1n+3b
CQ8ngHKr0N2UulN3A8EDFiSMeS/Z4uxqVjiTwHLTF43VC7/tgnlgvl6jR8Z343HF
kjI0MXjX4aHRBXCAt8ZS2/gpMcyKNc3g6UBXQeg0HTjIjhS8p7yfsXs4Cx/Mxn8S
0v3zWujHgSF4EvshnouKolwvdU3Q8w7Jo7lzheAnAXlZN1GJQPIC9EK9JAua6yP1
cA2g7OJ/vAt1vBuhxzfvC+/4oppuSpkidR6NnzHiLSsxCFt+yo9TN4lq+yFjWT/h
mGb/n8YUhuGrCmbmqlLa94g+daRTyLRhVa2v3NCGUE7stPQPbhQLCeI30nJqBQY6
QINL1v1DEWg21HKbOVeHo7b2qNQ0T287ggY4qMZHUFLDUTEe8eRDpFydqm4CNULU
f9a0aNyhze7G1coJq6u+bKSMWmXWwKQxpyFLDn8zpFP8scNUyTnppHGPOlsRv/F8
IdafFWn5AC7V5BSNDSuv3BHAH0yNp4IqweRud/JdLmQWo+/fcEjDBOmRwL0ryHZ/
r0PpjMkomQuuvFYPICwYyp74dI6oiX3LWL/s1yyEmJ6qYFFdOrDmyXVI5Z+jiNhz
Mp0giKKVBDEnMLIIYIoqs/YVqoQ9uFlMtTQFSAtYAzK7hooTL+ZDTB2hJljwKS8I
PiG6ycSEZV6tWV845DrqDYTH5LcUUfF8vRCJQExSIRf/b2U71Qr61iLDcKcTvyOP
wJgunr7OvIUk5ntvqgrdoMDTSZRWPEfv24RbmI3KQU6CtsbpGmOKrQvO+JzbAZN+
ublwgwbBC9t08dRtTfMnC/8S9WJSrziXsX2e63nmn15odjjW6lA08B60MlynGLOC
h38WFWtN018GWM/PU/w3NS5snLXfh/dQLZN89yUEM9zA4NQXy8OJIgUQCYMl2/2l
CzWmED06YJkPt96bxxLEUFJ+qfl9nItMlamYr9+7cArXy7gBfuM8tt5WF74jsayS
XqHkgvtqy/c/qJSo/q0uXzJwt1k/7aQpiqs0EItp3XiWjrLMDyCU46qVpBcbAl6C
ccEylCCp6mvzotNNriZr15m0jAz5w2B0hK217SyzEp6UiyOe8gtJOxWLd9aopCsn
nyFElK/s8PeXmrfIR8NQ2iozjy/POGzJOB1vn+ExQ/TTymZq8Y8Sfg6vGjmEArsu
c+yb65hL3TRdhRruqFd+GrTmOcCZS149+fUIu9qGVhm7lmkZG1z2HAeTvLEgkLZq
tOcSFGw1NlMTYncmQIbu33e/E9EQXJn1cSRcnA6aZu/2nkrKOWQjdbA2ODj9M7eV
5b/r3R1bi+cGDJNjKGPcE6hYnBMfM2MWqycRKYnrOWOhCEdocfOGN5+1gDTBByOG
ofOKyOISrbRe11T6LMJ7EKR0PsVdeJFt5DDUuP3UXFd0z2TkLfS4cXKddid5TZOV
+jLpbinOs1RZcy1aEe9x7e6UpnEQbTTwIQZzxNNJWZpbkjZpl4QZ651utADjW57v
kiGznusCZK/9H2pBcRie/+doqn0/Uz2es5tBbmDSs5uSI9gl3kck1qh8iPxaIMgF
rJ7gJZIbV9twa+lmtYlbVzBQPIXyOKr0U+D229j1YlvZNgOkQ2Bm2f/R9gLp2NmD
uN8616vvgCUczPm//s+KWrn7ZFgkm9trJiUKXT+FH6Pq4D/BBSJnahFD+EUG79rl
D1GWnt3xhEYpgwFyBAEvoOAzWjdCzz9mSqjgFacIAlJWAS5ppdHIXi4qnE1wBtWM
edcV+ewQe2p0kGsdSuzLF/DuPj/tA74mJ1ttaZCoHyJ5FaDUeAf79NxRV+0TPWS3
DCu8hiPXDWFN93Yar3J/HxWV00MOg4wxAxfwWJGjv55NaGSGm6pQPT25zmhMqBWT
4zsAOK7RIlnE32YckBXCuBR22JDukrmHyhntUKgwYHVSPDZB/QgqE3HsSZYcfKc3
Q+mF2rzVYN4TmG7FAl6k2d0yKWnTySsj5qLudhQbGWvFkeU61HQ1k6WBFhD5nqb0
uRA/nvdFaIh7OpkocS9no+tTIVwKm+hRPsc0pR7GEUylDWGx4EN6wipYmRTTfrTG
+QEhob/20ah3LJIh6c1MK2MSIlzmnVFnVP57YruGRfHovwQjcEwBDlvc65cev6el
KLfFmFE6TJ4TvHwIU3BKhPodcixPelAJquH9JzD7CCHBGXMse0PuwofcGPmcitPI
Wji0ryaP51J2YUDA1FvllImSy0tISCbhMo6DvcKiIXBrLARnUiTlWCtHLZ0oeUe6
CDp0PaaqkAPNLfmbIGESmKo4qvCgIKojMPH3qOl1lns1wOXdKor4Qv16xVdlfux1
BJdEXtcvt9qTU5OQAKQbqAP8B4rPz7TBV6ya6gpxPrfQC41wk+Au0QwuDOmxJ/q+
CKZ3TERHJh1A0M47yJiLoW6L/LtaSUcAAlDIRvosH/AA60a3a8l4J3482CkfB2HD
O3dAhDJNR+EoJY5shh3lRjfjOLoumCX8zy7Fl/rssInn+jegD1PAjWEnzITLcQxF
vTAFvrjMjf/HVtzHAAsnlwYsUi5Xo5U4rI+02zEg5xq+2AyAu3/xIF0xETGmEmqQ
qd8beolyJuiDK2XnOi9Kp95ESXFkOnbey/pngFZZMH9xZqeoKoFRRb6ggqvxUMQw
+mgv17LhIIu9ImjBFg9VE+bDhUVIcGRIEf0sRZtOCPhFYkfwXyS44T2ZlLu1AkBX
tw9na73JzH8EXU5XvI8sfW9R2Hh2H9JqqcNQg8AX1nodzil1xBA4Rm94bi2RVUBD
zXlMYg23+x0tC70Lk4deNVqB4KvQUqUHWMkRRpkkLvx+Mg7k3ex4f3zUIOd65xFf
21KeRcrHb9SPJsm4SK0awoXUQhDV+Y7nYTN68uvKTTSaY4rXLP4hdQeyYB7sx3t7
s8XbM+k5w5YlfFSc/SLhdSxIs38TBxkC+ZWlS1j/3FCFX07QcUzuEJlKgdIGBOwN
P9xX97lTVr3O4BoyEH8FPopo8vI/5B5gf89goXwW7pJ4SrBeNzI1VKFPenjk+mN/
NRfuAYEQsIuUvJi/tPCEsQfcGp0f9Z638RHeI9Ogp79GzpUSQVfEPRDHid10lYah
+cES9C3bp1Cfr7UTRk7Qrnf4Y3D6W8yH5YScXNUKUoGk1Le/yitvo7TiIE/VmBjM
BgUi4xp670qS/N8HUF817zcS3ywyIJzrQoHWs48+0a+yh80ebyBNusQvrPaEGStK
alnnpLo/xSqds35mYwX0sq23kSnq2frDngIft5Q30zGfQ8VK3ts4951Ti8xtMJbm
HIIJNLPZ5DzvOML/I2MCbEJemCPBC5uGYqAitJ9p4xo1wwdnb4fCBJ+ZeMp0+ByQ
ee8dwmF0dLyudF8dbIl5b/AzIEWz1zbWbNUfTj4naN+TOZEZTjaAqmO03Q+Sxs63
QY13OSPuHWEeum0ypUWFprYQH6sehdQQXtLRky+aEbNujxgVl7yVzGpGCPeltydj
DADImGQxvVKrbxV15GYh5tU7+2R2aHasmjEVEx7DMbItIMASiXcTY6MNKJWnhWNF
n+ovimof4SDwGSX6gKNK+8Jbcf+98j1w8g3G6kW3pyW2o0iCCFCbYjvDc142rs+y
NBL7ii+I0heQ9irc9eWUEUvqdEm2ui0mbWL2F5WJcUKrDkC8CD5I81SCkDI4rRe+
oPLbSLKQ4g0G42Gb+hyKqvdr7zNvEAvYLTZkSZfBgN6K2JoiKKcroqQZs3uvrFlg
pCnHd03qO2W1JWxT8+Qt4/OTY69jfnfwx0XJ+lhuJJ4/L7T35/yEmeib+TT7RN+P
Uaqo6lJzINt2ZiP3yQMkMwIfrayrMGEs2m0OJf55vm26p/558VMrLp/5+8a2juA1
Ohal4lf+2AQPwNXDkTLPr41Tth7BS3pukQ0TS8jg3ScuaqMcZ2RU39ZHCEaEUo2/
bYFhXWw/gURF3OgBIJzY0KJ+sohVV9IEK/C04O6gexbLlp4KLzZv2sIUI9dh42nj
aoqG1xusLw6xoMUaralvjFTAdtjQmOTOQHhc69zM3QtbMe+t8TO54EmP9jzydMzP
QuQNmvQfNr8CeTYIUB4SEIjB0WhQ5Hrn1BrJAq/shD2Pku6y4JhwxghzMhzt3lRO
ZtkNGb1XqUH6J3b1QUQbo8sYHgeSx8hC7EYwsaCNVNS1aWsrWYIOCITN/dwJfYPX
hF3QDZ5iwFphwsgQWe9SbZ2g5teE/bdqGcIrHDyL6VYcaASHydUFLLzKXQFqomqA
UhUbM4XvT4NbqKiDpaAJ4YRSi9yXspH8pMoJNirOZi2LW9ir7Rj+EsLSMt72PFgu
LFsO375Tt18TR8bvQazv9wa89iBhUP8EMAY6W2SHBBwvp4VCD2zgXMfNWVdcg3fk
p9h/CPos7/0eHKT2tvJ0OOEVgW/R35LyNaxEvztOFv3wPREaeL7mOIIG66URaBPa
wzDZ1bHJzPYdsjF3Rf8Jt3rWEl7K4A2PHpolOOlgZr9OLen6L3oQQpRifSP3F/L6
qkKtzhC2INTMTBthNlb6XtdQmyI7vlZWllMcjCsxF/f3sQK1PhMwk2a/XDrQA/gt
XNUyO85PtkzEg/JjXePZeY/6+5bzf+8vs7ocscjuz1FbJ6KRRDt16GpYIdz1KQw5
JGIiYhFy5nfPlmVOSxvv+PfB7XgQYN5l9laAMaHWw9KzBdLNactirHOiUZG1ESj7
/OA0OUN/Y5q/Kgonh10YELEgf6BW7N1JqEtSdrjDgEThKHcmDQb7+ktoxb6kQ/rD
KG4fmp7hFmWDDDPGKEGW9SpzRfJt27SsaOQjERpBRfsDDYxN4CVzCj1kOnFLq6r2
4y/77duXQK2gvTTUcufFzAy9H8ZWGx6bffn9y9N/dmvLNiqakbvXIzmdIzbn+6hI
sZ40lnkI+6cs87pYxXZFnBf+JkzE6wWq5Gvjsvz6Fu61fujhaLOzot6id9sy+8Pn
rIzYdkdqMS+IkV/SyWXzSv3j+neqfB+S+m9+svbxl2zubtdtvvPTPhsiD9gtx5/9
9aPmgkd+rCd5cAVXjh4+HwS58OYULzzwZTD6OSaHrUD0lhwbWUbB+bZcSCCFfQwg
TKqk140F1xxnspc3DHkfvFeR0Sx039GM9/eJncHw5CRVOw1LV4wppv7//Rs9u4dN
/+wO7oo33hOqC7dL0esrBQZNZVqLVPVMGAc+mVYgYV7uuoYnxsKg2wugdHHeWA6o
Lglu1Y6W8xNMUcG73pBQo9TP+iPD89MLwaQKJt3AIxukymM/uV/ov5VUVtmUgnLt
f4F0DBxNyAw4btKRGcK2hWXUxoVjyoK4Hf9hcxyjWKfr1vP5HnFl0kILjrAQMCwa
lDR51QWBQ2Inn0/FbAsVxuMy3A+ZFvYxngOOv+icXOWbo8VH+xINuwl0nEUzvFhW
TZLbjuMsqLAvcOFEsyuKUS2ax+lShn/fHtitbiu+AnCt2F5nDlCD1yFXwsAuq0U0
HF4UdSvnYpStViZPbIRaTNsMXVW8r2ID7vNgEIvXjQSjw3e1f6WDDQLP7cZ7xsuy
PKjZQkUPylkWiiXBQesliNMyJUmhaoMMvrjtUGnJ8UjZE8QP8yeJiKaq5hUZrO+U
e8fgAkln2CUhkNKk1ffZToTGMFFAgFe0H2cqr6xkrfoMZZhUwZA/GORScKlWpG+d
4TO28EdumxPSSV7w+DCijfHnPMWe2AuJuM/m9Rb2vvo8hsVIGdyeW1jLF23CxCUF
NTrxgoYQlLdNPoDOqEXklIGS8bnPhmrz6toWxHlNUhk9ZFYviXTvW3+gsgx1A7TO
c9M0zHvBw6CuZCtqnVL8EFUALCY/eRDZuimzjfurtdqSaCJ3evdIhktgS4CnYXaZ
XeX05FAZ+YdQeQKbB+HlotBbVaDiMT10px8PYFbkLyvjiUWuPgcU7l/+bp5c4NX7
Aa4p7uDo5Pd1f0UEJlmZu0/bGzgieDVojiE75NYF+ZGYuGsLZhMxk8pC7jkMk7ZI
/3JqdJN5WmexxVjShQjPe2EKwIFWaImX5BubCs3pwcTtQDpOiEZVjfOWnS5QWZAG
RObzQ96ZV9OGan/HbPIXKAEVwPApGxWE38noSgPc7VolPliTmdK9Fh7A5OWBkDGk
kW8uSeBkvLz76sF+iS8X6ZUciNd3ketDYK+SNSMZ1j4ubr2yx5Z+U5AXkSLLVSSK
WI08/9TX+WmYwNujLCOqBPelKFsqFW27Cl0WnQ8Jj1vnEabHU6GS2vKNmn83JLfw
bFL1xaPpOBZbfdg2eMPpMpV1f/9aKbv84dyafqbW+ybHyi7Vf8pzDol5IovhqBe8
5VAXBnsqGf5NrS1dLyeDF0cZGUab4WZ9XYthz7ZjchRgO1zq/S+AEgdEEvsOmSZG
U66voU6Dsn4iKq5jmzGLJPBZuRSAtfvJaDBhA+nUFEaAKqoKbsIAfAy8GuoG+yNq
eYiSe1WA7y0EzeVqcxy7nBocwgeykQ6+HYqmJ8mCV3ASvLOaCLVLEBSpxg2qKNG9
fK+gt2Nnbt1qXKTRJjfYhV1rBUc27IU/bR/a0VkgCKM4Z0jx7/cgLKbe9nTTzOMr
iXTdvPqYegH6EkazKPDKPjbBYxxlrm/tcUQm5UHLmUfbbyzO4RMdf4vBhZeo5o82
y7PzQ8DklhZgeprhkS7ZaQ7FQ7GVCtXlMXmO9ZpXCKsGD4GKABiVeDPZrZR0+h+P
rsL/eWSbiSXaCvHAQMW3f63XEa5notLY59rddaE0Zx9LOfJOpgyUIb81W+mI4+Kn
IDVuE41+gwhFyTpgYqg0TTZAvJLT2KZBour+i4Uag4IFprLfo+Gvs+z+tQth+ICA
zgUQgHTSHB1J2bfob8w/nH+mF6pRP27erk3r4/rvJjoB74sGuKTrSHBSU5iStFAY
YrSzQDLVoDimas54SFAyZ8CKhsZs3B2okcHFxvZZo2Tf5OnyIg0FWSkysg/8NlgX
OFTrBb1MyOksN4+c6K+JT02qXwbQSjDuolPR1khefkW6jg/cbydNmF5RDW7ue2yL
njOtuDl6JNDXhjV3CApTiKlAFLHbxCBaotRczPv5baq9gLK0sJGfPFHq62GrJQYo
JQHnRjf9ci3usP/XncgzhmE/mZ7ADeaVUBKMUpr/G6ETZatFddOmu7D9d/8PeA4y
P4qxCJj5SM05XK3ja81mD4wGNgNgYaJQLoKgDOnpRCdOdAufXqbMac3MPUHSNLzy
nNVKbrnzDBoW4OH20JWZIiAkU/7BIMmGz52WWxnrcb5JKjTPFLcMXt8v0A3kPoUB
BXOQB2pZ33rLwaz0I9f+W3R6UTKAgLc/QiWs/b8zmmwJfO/s1O+MQifXchj/1UUD
JiZhWUZeXucjAtlrltgkxepvtRb7wDKOjuKRkfequHLmadUaSTE4bxuaoklf94Kw
pxLye0c3+j7l0BtSTKnOuv1N5yDQeeuN8l43+8u2zI7QlYCzvxYB8NuPuXDAZwAs
mhWz81gzGurKR/iURP9kNo+Xbwcga38bf4GbMmZDUnPx/StxIvY6uT3pFO16bFyf
k4iE80CON9wERgd3SMbAgBEj9FgmgnnQYnniLvSvHnQV+KQeer/Zg0buyPL1XaGl
SnC9ijTHnLhr1vogO0kyUuHNH0RrqhukWvbDcmU1uLF6Raad3KL5lUKCvmFMj+M/
MoJZxEYkbvotAyfYMWIfRvjhgp0BhfTww9NEvxNcNXUpNXME3U9fuxKvQW2DFhsa
DyBabp+apjHkqvgFO3/Y4am3tqi5SopFH5tj1KyqNnOJin6LXY47wqBSwsEmLNnk
K+4/MtA2aza/kZi4ov0w0TR2N6CqrJ17xy7SnDNy3vkyMida8UdCRBcQpRJt8ypM
IomxefksZrLQtefSu2doMVZHSKBAzVLvCCs1ZFM+S+TEsnSU2O26cv+KWfBwpM3D
4y0Wl/GGzfPvlJlTwUy0q7gVnMX37sXaoQotCu2Sa2cGoJDnMEYTyI+hshgKwkUW
3SHKWrAVbep+MDDa261cGNY+FrsbVZONtSxn4C7XCS8biDm6jRoUtsC/pN8GVt6Q
QSY7WRXQw7lM801AGXCJJpm6cu3io7NiGf3Bcw21fHzyBfLkY1j387KQOIuDnr/i
UdmmaoJRais8v6wjuxj/5dI3yMzrArQHZIrgQ4oj/itvUJZbJCEbXTn4n88QKwL+
NV8ZS/S4VXpiWKMx0Eg9L+fjwlro/Sa2Ivf4D5pLYb5ZsTnxzyoiqBg6Zt9U7dVD
Za9kmDCSBRvJlkKXb80i2dp/4nFuzJiXNLiDZe6VRHgHPeSbsEp4DhTd074ZUGB/
7fSQAky5gE/q4rKs5CQUd1J2clZ+k0NoFHkol84Cih+Ruse1+nmTS02gD3eh+Mh2
aHN60lSp06ljs3/jqdPVHtBMN6YYfA075yN6yGWQOr2LxhtmVWHZiflH39sWe1oK
aYNMpD/ai4uZYF+KQCB5N0IPT7PhSYBFtSE6M/T2b+uvDz5IrbTvVZ9vgug0oywi
v6utCk9sKBVhOtiLk5Pz6U26Aj7CflzZ2wnOt0tdah4r0Gqv7VAJHukFK69e9O7F
VP/ktCxNEuoYuIe3HMXDUIjVflM8mHvm1PT6z6P+5c2A6nwH3jxoDyN84/vJDcyE
M9mbwBCm8sv30mu1tO1bJUtw0B8/t85VZ0Y6yBRpOkayTlkiJ1j+RkZobr7XKpY4
dpR+1SbC4kjX9EnlCYvd1SYqOWigK4ifq13h3ZKNt/sMyPETl/qrYQnzvnVlsclV
PdwHOwuWn1VjxagIQtLuIpiITTglzY4wBfYOiT5V8mrWFlhmSs7oiiO+wgkQWAQZ
BDfd6feITfXZ8trQMIUudVxzkSqDV+ANn6LWGMWZEkAMkIRBa+xtTNIs6aSMHNmB
bId/VgZFG6R3bvHPbl/9UPnMSjPOh/dPFnQEttucKW70NuHr+Bp664wlpyoLm6X+
qN2uXbdHiKZDsmxQEYqSk+8umXNJeY5cv/Kb5KI7lE821bTRcTSgXlP7G7wEfrxw
`protect end_protected