`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
ddtXksX2+yylW5zu6QL2Lhnb2d1sD00763mmSITNX595NcHTEkwn0zB1Dry37fOW
FufOhVzEJp80NC5qZ/+F0Vk7Ik02dIR0elf3clrjeJRK85K4e3Hoo4xn7YbFUIms
l/8VZSb14+JVGURjfswrIyCUotIzlzVYZ6gzoZwDXIi5gQIBf/gI+KxNXPaKV+PQ
Ufys/12rjO6aI/pPlqSm0hCvftmBcnezN2hk1UeXgOIuKZnogjOsf0iJVX2aOOWE
6pD/psybjbnsNB6kH5uFTA5frkzIzkzl5d9+YDm9OyC+k84E83I/7/j+rk4L2dah
QJOvksSIzN867/4Qt8qYTQ==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="MvBXkzurAa5VTw+1JJ70nePUfoQXBvZOku/SMmg4TwQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
oRtzZL4VJ4iwysPsC8SXYCzXS8Fw2gtZTOskLcDV+1B9Nzn1zTyNtlo6lNICRmmK
ZRVu2BmCc2G+fmzynYlNTnSa7C0Cuel6FYpxCBlOuk3OF2tzAmLAuDyOH3Z1Yjzk
a0aHuoCdIRKv7BrZCdALt03JeUmXKPdOmIlkVGFl8yw=
`protect rights_digest_method = "sha256"
`protect end_toolblock="Jn9CQpRhJt4rnzZPRk+dOpzAubz7omckX1MrFd4p81o="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 18224 )
`protect data_block
gD6l00tciPUa6pDNTk/+t0OO0nC/UTtBwLB41d4inuAUA3i/ALrNyoJVcBnAmEQW
ptbcNp5fxEUJjnOxnedyZEuEBxWRieZFQnkRdF269oMmPauSIg0aoDyPjFiNCWzs
bGZJVdc3NOEPIbWS8zu8xzcAjEM7Dg33cOfgj6LuDdGlQVYwPMt5BZVHPyqwkAud
4f69ajgfKv0ejfSvnxfJ51qEjpF3vCcqkZe4TemeuooJs4RBSIF78MW/kkP+AaWe
GgSU14rgILzTMqVbiRB7gPPRzPobgIwVqQiDDbY1SI87yZlo1siUv8JuqwLaneot
onCNIxS7RU1PPoDAxF+c/P6gij9P1KUW2gNYCLoskoS9woIcqzN+UeBrPGXEeHt8
ZY2EMKEOOjsids/fgIYNEFEQQvGFCrTRG+vu5hPnUPu85KfZoAIvj8iJjtsch87r
983ykJGBYglQkzMNuEmVjs6bioxFta7zKHcOfZnrDoRwnz5DEPQ5m+OeTYfdcxcQ
W5RqCCkH6l66UtoqA02iKG742eMIAfWAL0llvesHzGAPkZS09iFoEYKmLxcqBnbm
1uXkCODsuJBAjPd6psU0bQnMeZhrWDkS0VfQUnHu2yQRZqlNvTH6VHZmNi9s7i3f
Vf4z4S22rjowyL8/dPh7kBxZ2e9QKZOh0T2cLZe0f7r+7zFYpkZ2qCf+ICqq7cTN
pBF/7syqbsHGD1IN94Epgf6oPVMiKqwtxhBSGFPJyz3EK2fxvThpSKd/x0YLztsx
DE0QVy9BOP4hMx2nLqTgVJlu8by81+pe4rn7yu0Sc24UB/UW72hY17Jx2QzWf99Y
oHXAnFRjUiNcvNXnF61X+JQBABT6/TTuWi6X2M6BGQkhH16pxvXEJfReYh1dspJ4
uCNIaJbohVgfQZxyLSwmmhY5wK5vQrtuLqJew2VduTmmQT2g0h7ynC3mL22AabHM
181HM2Jxr4eokvuyNPP7GkZX10XtdfXHLPysXjPDlnee5lf8k/IMWHPLGMnls2pJ
3WbIfv2R9BmCmG5fNFnz1xyWdjb4H3MSJ7Qpr227wpPCAV0cUOVV3K2b4aXbd0oN
B2rTIgGPoe/BnVmX+c0uDo71LVT6bCINUhURB5Y1z0UD0849m8gyeNKS6CE5jiBC
805DM5pntQLiqoIsYbeHK0MRtMTW4GV7FM1d0OZ7dBiequfBM7Pd/WJaGAyYj2Nb
8O08EjfNUlY/3uQHYSphbpQUGH8zDRH6rXT2QUXDQGDf/mpfX496xHjR/sHKD01z
JhnRtNjzgHQR5CU4PsG+tdzV8Q0enTtwqP4k3u1vdy3J2XnItVUG1hhD1KRGFbNR
rOK5cxRXjlxc3eNMJV3H0XhGjijxIHwmIXlJyH7wrbGWFtsmFQTRWHI+BSyZv34m
UWa4ZiCz/QfvLiYlrhm2BjYJcT1i5QuMqb6ZDtNtZYiY9zetxQMc8QpIROZl9FI0
6x+VXACPtsvxG54NKYko/ep7GLY63A3sH5/x/kXvyD6Lzk99mCf9t5jUZCdrivyE
15dPNSQp2fCygyubqukVp8GHCvk4fRdY1SiduZE7U8ABNDY6AR6XWGE6hlXUJ60/
69EnLOS+IOrJ86Xrwo2lrv2BMUS/4G464/ISkAnVv4nLsRvSRCEzOIBYWG3LfagW
u5bt5W6Kv3+mtSRyJag4Wj+7GDO4Ohed+qMSw0dPdzdhOTIy8TFEHeLVIDmzQMfK
UIK6Fki20uilFzQoHKZMCBCB+Ypfmb+q18+2lQS22OgMVG4Fc9bixFd6LJFSakPh
1Sqv5WwHQQdjWyNKfjj2Po1a5jdiV19ZpN2pKCJw8/7/olw7f2Sjafda/1+RNdI9
7OgqH9mKsquQ7v0cBT91GCFg/ozMxAu6rKvpYAZGSQtyzjiW3EVEW5lRMRa6twUh
/GFpwK/rAqyQ5MlcqB40Hw3OO/fh6/wLpDwwgGkcLGIcDJaz5pK+W0ZdkAbHB4pS
imZ3d1WT+vzdO0AAl94lKAxcclg+tLxfw+0WNMirz2EaT8BVDACJ6mJonS8/wNvw
wu+EmNsiGHI396uL5nDhl18Rn+YM+N+ra3E6kIEkpn8B18TxU++XPdHaKTAsg/+t
cTLIJGJnrGaLaGGf+LBmHa5qxuIM3HznK5xgnJlnK5Ec7utl3kNZliPA+5Q9fBpb
5pOuB5yMC8S5wvCRIo5s0Qj4wI3cfhS+8TSna4jwcerdDWboj8R6gHcJf1xyk01Q
i2ce6BZkIbxWtZjKjTswTnvGEyOCQpt4uvH+1WzP3smCmUAnqArHFn2IeXqDmK4x
3xVChc7EgaQsqG1carLGB462FOTSBiD+p1I/09e2w8AAxBJfegk94NiAwWvCJEwi
69wl43NMn+1LhSV7XxvGAKD9rsOVSw8EMvpLDtpoDZTKhxR4xDokQqNaJbR29scp
jTA+njFxM2STyxapjb7f88INbifktebjaJoP9u7Tvtg5+EjIulTGqJhXDbF4ohBP
z032zaR4EU+nYDbWraMWfM2U0nVJuv1d7QALo74bql0EDHclsEEkTPN21Y8Wi2RT
9GSvJfR4d26+2X7PqLya9/LXRs8/pbtn2kQz08nclg8I18F0I569dBIskEKRbp7C
viJ3wEwd2YPwY9thbVE7uMM1QxNuYRUAj0L75Ro7y0bQ7PaHe/BH+vs85UY2HgyX
vAKo2yGqm5r8K8hBNki3Ni1Z3mliWZsd64y54th05QCxZU3Dfs8Y8soMOO7bvJwA
qyj2P8c5bwTIhBV9rM1JTaeBdTnuNulm6tcGZtWxyE16LohGnuxlsp06PrQybN9i
lte+wK9acLnJNqY9sVPABShUHi0VrU+LQMJmS0xUs1vvbxG+mKC3hYaLuF5Y6hV7
yBMtXAtJIdq98M5SjPbwxEzQnanOhN5vq1ewvV9JEudBJJWes3OcL73fWQYyQinb
lZkawm1TqzM2L+SNXcI6Kwh5lblM4sxTqOpngRk+cfgA7n+wqHZGLy6o4Xvyzxfq
/coVE9bbzb6NcbhRtDV3289ZPjYsHPmwnuOhG4GEk6aJVaV1TBV5W0mKGT0NKR1x
GG+5AV4AzuSKBSDad8B53K6gm79XVbk82wqC7HpmW967yxcRFNhvgc9X6O166GWS
CbWbqi1EvMc82hP0RQhS1ttfCl5Bnop0yg0t7P4Qshxi1ZhgDyiAopOFjg//Og17
rJtSJ3FvhaGRKuLfmownrFPAa9ELHZHFuI4S7x3kwm574kUhLL2v/jDPds/HtP41
wW8O29/Ph3NfY2pm1WpKqehQbhNaC2kZGJJfR/7Q9C1kRcfs7VXQLN2YNY4bIcln
fTCP6+naQ93cXrUQSe4oLXt4FyvPI0MmNmJ96kAaVo6XckAWPcHT8NcBQxk7URFZ
C/uZI+Icqz7k96d4Av5TEajI7ZMmgMAtGlLTqvZfDGVwH5OIwAiERDIlWDlqENDN
2965LzF5e6exghkBZW4vzPfj3JXzIw7ZqyOtGeS35BzRNoXNvsImw2pr4Rxvyj/P
dV8EreLCUpFuFyFE/XbYcjhPHqW3VOF1jsToFmJHHIzKwgQYVcqNNkD8uRkhKSJo
c8JDkS0gWkhFVg+CZWCW9ooMWIvEDK8OkjX/WDyEs8GsiBtqS2oLkSQAt7GGi6uA
1BOefhb3gUHihmRhbVfOEMfZPvS4HzmuJ+ns7gSFOc/EX6X93iurVDVMhzuL+OlK
r5nKVSmo6qWKNfAQ1bhxq/qB9yOfNRBcyjO+FCTjsCFxVo0WeYYXX4NhLUzONcE3
VHpM0TcaZT8IeJxBvNGtKBNKoTPYVwgBtuIbzOxGN2s03e9Rx2o0QcRRioI9xPn0
dRLYB6TotOKrtma/b+KGR5rgcShsKvCedDBTM11LLdenfFVgjnRFCcXS7Ju67cj4
eXRDY1aiZPjluuFsASBi9iLGAZrLeL3ihvq3IhvZ7XvGOgePx1gzJ/HCxxUYjlZW
u/+3BF4FagCtCY3EgzCiANtj6JTlyYuYvN3sZ8bomA+/SB1CSIfjqHvY/penPvgE
7kumUdCUioGhgYRO4brGHUjYBrr6B0dHnPnbor6/vwguPSka0KMw4dOuTvfF0gEb
YqByCm3B8y0tJPJMwEzQuC64noV6CPSMAv0UEylZppFH1oC03hQdLrhumC11zk43
aavm7sPhFkAzlesCKM7jbpmfqtERQ6w0I+RMSLF+31aVn24mlUXRkThlXUMi6ECt
wFuQ1xIxQUz/TKPezaHi61N+lxuBML+7J6jTpyl49/LyVl6c15Z9JuiK+avpnyec
ncX7pmdaWihXtixhLCa4cM4PUAMK/c/UKdejl72SMP/mODQLfbI3QLgys0x/tVIe
qbOg5pyZsLwDPHcUju06zoOQsGVa1EZqfDanpxL2QZc1wOBZTRZOTPoSUkvaIvIM
bfrnaVwTs+drWM6Hhj4HLx5UWEjOpGxOvjCvxNmElxQ3toSUOklQ2/lyc/UxgAks
f3OC6wcm0bCa3lAJH5spjgw6PM72ixg51UtBEF1UdwM2NOCeaGg9NGOk1IwMLw2w
FrprZzYkAxQhcWnK+7hXH7RSRSZ+aea3ZCnAKJivHwDHO0hbSb9d9jajMhQ3pVdc
QKzLgWwD0KL668ftESVR2KgVhsljJCR7uwJfjzQm1Yd94WMvBPAEHbcuuoBTcDLt
QpWwPJ34mYOaGEm1A4/m5AZk1bb+5MWtIpRegfWi5wkfk2z/nR4XFgD0cqCBlG4F
r7VIdYGHfxIePA9/hg7VvKDNGBwdfwwwXqASLo2tQv6baLEHR7g3YQwKHcqWciGk
9pmzQtmjHsXFOkNoHgx5g0AErr2YHSDhtRM/yA+LZF2VyRBNOeTwycrKIPnwshbV
vt0lcR9ZHgb61CTCIQmGWlVmUIT969/fBmysrw0Ewp8JWSDgyWOxIlr97dic/azf
U9B7cs2YQs1ZshXRpgXsIanRsvXPG1N00IBcKgpAJZ8gwAGZ7KCLp/cw2jvGfK4O
tM62D8/RchjAfB7WVVW/nbBSH41PkqGttJw5I2FgtxT+1O+zSJSdo9zukksyo8Yf
tjl7QxJBTDahzWyWPeD7HejCv5/dPw/C6J6hONUnVk55LYUo3+njm3FZF25mX1eq
ZVs2tViXfosJJ7o0TZ3xZ14mw8IpealjApcqpI5JtU2MhXYqzpOdJRrn0i8DeK5E
UNCZji+4s3g53mFhRWOm6tshWnnPXCtzX/CGQLd7V0sHgGPkemCaO/TVRGuqj64g
JZK8y+mbuR4n+xvsUir0pPWW9yam8N54+beE5x3WX+R0GB5GIyVJnmj1qjiFUQf3
aYK0wn8q12ssEZSBOdQxeLEKygoSnWObLvXhne8GJLnfL7p3cL8GzybdPK5UmzFF
MN02vRTbETcO+TnnWg4MfCCb30M+T4XzuNuowJtZdnEnrMUz/rYYPmxnVn5wWiLC
8sS7W6NBE8BWFgkHDgLhV2pkFEgHgCvU7BtlhVFeF21jZScqT/35JGex3Z/N2b46
s4jQsVK8aNk9+OVqndsjwLi51XxJ4Ami8v3e2gZCGk+k9pxB66eAKmNJ81b6XfL3
j7QFUlz+Kvz4XbkL5FcTHzJFcw2DEdVQyTE15Y8hIbT3e/SrBn/LxJjO4eIgX/7s
6YoWc2xURPfdFxd5XQmkF6rOUfqI+OUrXh9WTE3CPI4FXOo02ZTUtICYGdvIHaO7
PjE3J9NOR4v3VNGRs0sAEgV36hh+8vnLQH+LpsdvIxUwkWpMbuMtlbk9snnN+a6V
tUADkCh4nbwvsn9UJEAbStweLnzIBJdeVAiVfy44wc8ABJ9a/b1gQbXRFWnz0mvt
N/nzHjCznutiGXZd6PEEY0Rj9kw/AYKMDjY2JpFU2+JLcA3sIReFweAwi2/2n+a6
XoFEWLfNBxLVEWjnL3emWJZTulfPofcuKZZ9zdsyKOQRKhxC9H0aP1INRE2AdFLl
yL69j/Hy+2saaFcEsiN1SGKElOkAdgQN3vEjVW8aGH76d8vPrcJyfxBL52zl98yk
M1UZKJNNw2IPzjc93XOBNrZKtwjnVGwN2Qyr4/pjGKEhlvyJqIeA9KkvkmIGWLt9
P1BEQE3+v6kEubPrROqQx/pwq3MgMk/z41+Eqd41iF5GxnIinDz5ynczLdPkBPf9
2tQqqT63sEX4+tWc1V/YdVMwxPADLqWEDeAM9pGrl1HQHK8wqcoFm9uzNuhYL+ak
KoRoDVepO4IRBR/XLdUqIAJ311iFNFZXj5gqv4VViKXaIizwDCY5BqfgFO7GHz9A
4LnZIfEtuoen8lepcNttJoBBEICgfKoEv/IC9pXMGgVtMbQ4hEYc/4ioTZgLTiVb
sCXVPSyotzXA/4/wmmoBfLONG34fkAsJ73fE/+jPy2AXXUF45z1oIFAKCtX1/adz
gYcPynpYuBp8RYcMOJj31usYXXQGM8obnt1sU6y/QOQccNZnJo8zEewPZqKA4uGq
eNYbQso+4u8xeo3amnPi+OP2INE2lxL0DFxPDjHelspRvIXnAtY3sKIod7ugygK4
ccMwkL1kK6TcJYaIyTb4BOjExQW+Hs+/HiTiG2515BcFq0rvaN9XixH+I1MjdhXd
g7FUyXsFKdKy0Z2ETvJkRyHaf/HHVw0Jg9yQj1FT4Jazv48my5qWywyy1IB8B1nh
8qytrtH7iBE5HIgTthH7COCbGzAF/4k4Nn4U6yFS4C1O73lWyXtxCJTmr+8Yr2XF
9WBhOshSB/qBJsfIUNX3flyjijpDKvrQU2/OeQvjTNToEhJiwWmfVUJ6vspVf++t
fVtt4JbJaUIL3C4SjwLIzSb7CBIviCdZfEkt7r7Lun5Df7kVCvTdISlVPHUFWG3b
it6BZQuPWn0aY5A+jjrNaVBYWvmx1LfOtY4CaMT82zMV4sTovMMazJv9QBsSQ9cg
Os6pd5CBKO6FAGbURty3RcCl5f3/T1Pf5oLJx2gEYeCDAqROPhG4IP72N+Y2h6pt
uLSzX6XbSLFgDwGtKOB/mPMjDJj8sy8PxvdJLLDpwZHIylgMZX+rWQ7X1Hr2Zwct
rVAnGUt8CxiVB3bLsYqIuWVFKQpvRcvPZJ0vby39DZzLr5qdPkSoIh5O9XJP9fjG
sFKiM1WDkKMqRvpEhBrsUEHd712j1+04NVmnKA2UIfecaUbOHKOttbqsu9Amu5qk
phaMS8LopVytak60fto64q3s6TIU6sHxLL8gv+vkTAdj6LTj08N1rdT6XCO9n4cz
dYHeviEJf2b/7nR/5c3NEvV3SOlGtjGJFkrV+ACaj4zUI/kId1qzrm2v5etB0mYS
ann+FImscCBNR0NvhMUpZwemZXRPMytCiLDovZzQ2AozXOednfg0nIzJV1DUKhUg
/B1hMDKjNbI8vfmH2UWtZQh/rprcMwSAccgjZ6d/l3pztZWOlt6ihKr713Lmv/ct
6KLdVXWuzo1zkUWuxIIF0ki66ypTIf4QLxRDy//pxIWVhC4E5z9Yv6FaP3FLVqYi
8PlYbzPCMTi8huR87MtnqMKx9e6RRUNcCrLgrmDSKOHV16Zq7rlPDv4Zb2rb+lg6
fw65dSwT27CWLAn3/6YDPMGn2vXP7gKyaOwsVRfaulKZK+Rn9zvciif/3lD+R2t4
lRn6RxJNYTMHYASTRMp5RMxAessIpF96SHKbduyWKvq64r8jm6/cB6Ay6+Kj79Go
G790x4hqlPUq4HBpJg5tHyZ8KKqWJv1eRk4EgiGLtCiObwB8iUSWibEXou9Re4Gp
AACSaiDvOuQ1/NmiVG+Fu0jcOQqu32/scEXpt7575kkDfcHJRqtzEQ2ZqSwXXmBz
04pVJhPkJ4RzW9jQ9KtXShshNJ9DhLvuTlS8uTAlN+H48CkXJ4svJxfnAaGbxcfs
A5+iRoBH9lfnsjB4RZDeM0IoKUsG7BMMfYaji+d1gRUo9HTpnu3XWs9qxZIoZzeQ
ju5GvS5hU2ASHb0gIO9VvaaxxZCaDp7wWelKYexD5PuiKqPxNOQ1QXN8+M7GbrJy
F/B+vLYTzM0aqmA40hoktxgkxyb5xfF40pBOH0NRYGffnAhQX5GYMcyA9sKxfJDB
2tmQEY6dNrhNhXss3Av5KBMj7MW+BoV1uBdKpfyL3s3i0BpLvp5bg8KaM8V3lEzi
rydhtw/lOo1d3WqDUKFnhzLfvK89szTUI2PQS+VVxzK4IstFYm7YudoY3m2uTBXP
rMSl865bbwjbOAHak783Af7/pSL9NYR6m+VS3Q5ZfPAKfEo+QTsmn8Tb1mw2gkHc
h0GqnZXRzNtbWAjenShUQJoMKGnynSKcAAs+0+q2T7NfBqWKSXuUrohNGyp1F+OK
4yIwtDIYygXCVbQwfbz0BKNHngMOhvDK1eoe/2aGKqVP5kA3sP5N+ffeRGi+Umjw
qlFH1g8srn8+JUeYeuJ9hpo680rLQeHp1yzbs21GroiDFCgE+oSGpGxLh28JUqEy
DOPDZgGeJvwWaLAEWOAfvBchS7rMbiAuWO5FkpgZGWjRLq3ui3VSETqenOhmmeEr
yNYARnP005AP1/ssKZT4gRiH6VAtZaw7LH3BZbCguNwbVSnhsKssF8snX7oCoF2w
dzuVjTNkZAZU/AssZHKx6DufQL+IJ4oziYdUcTNsrMmcvqd6UJR6/kwdXI8Id1Rk
sqdbwox2dNWmLkG7J1R1K5MdENUUVoA5CARV4n3LczXc4OPNfx5+gOrLnEnvAm98
ntkbLw7bDRdHI0gzUfINiaZ6puTnIrTRgN6uvfvITWh7hQqu8Xs/4t1TV+9dJehc
Il02M5S67ejA2pKob1TSSC4w98oz5iWTdhMnPH0VRbjeolNgmCeSawmmybNPOoZk
v5ehha3wuufiaJgh6tr71lS6+pjB0ueynP2iQmgpS8m3COY3ld8iIBVw2Ud3HNoZ
SjpbrNuMzjU5jZW9O/po2dQqdM1Gp4QgqCF57TxeVv0oMaVYE5oMo9ROjsAUWfn3
GbmPlU28NEF+XuoVvEMxlXpgw0YiRhd8M/ZPa9hJJWG8+zRhkZR7PZPr1lUz75zY
Ncz/D07NWHirfcmbh/Ee6inPTjeQlP3arDD/MVFia6irxmf0vMx1ZiD0+drAczje
nBqNtoOPkvL5jhgCzvIDO2xMcArWkYdFERmNo2poL7gyU7UHpOF+IWSwrncRUNiU
vXYa5D8D/X3eAIOG2MzeUmpMhHVUXuZ7o8HWZaGPSKAOtnrNUZFU64e17vslGAoW
WvGIIaHYEEFw0rsLOplydnaKCUhmt/25j2ANMlFtjuJKB2NuxIaOcO+Rz7SwZqoZ
2lRolFDFzXpUQtaMDoeOQZy8eIxupbT8yjzYlaKCmuRpq3e+jkOd++aO3imaND9Q
8gjNa/Da6tXHjLHE6MVTKBjODrDloqqvzFDAkd/T6ft+wmIPVCxCi3i1awRy1bN2
eMCeT8BTtDR43Q2to96hxtm828nbyWGoZZXTQ2k6sGa+p3TC++ZWdwD2F7ccHk6L
irpVKZaiZBejiBY75RiQgVE51jqLgweAaFc3fbqM/+DmYnY5T49W2RuOEaF3oEzE
j5/m/m5vDvNKuDDq27qn/P3cNUTHZjuy4zGOHJPGZcJFqlWcc1lB1Zl0I1WQIgaA
GiPnjY4KPq+WpoHgMG59jbKipATyxMN47/Bszf9MxsQo+3Z2QLZYN5jcG4lUZzmn
qK2tGx9HlWwZ7PBMjtIZP01wOFbMiwA/O/7Ec53dPWNvZX5/nYtqxENYhuruB77q
EvW6gb4cIvswQ/bh7ZoCMoH7+GjqMkTykRbj3XGq4/6OSZIvGoAJY1KFy5oCOF00
wSFmvLX7uQC6a8MCTeTbBo6V1qrQsCh3fw1Wr65ldMBKbgm4FeXwfVbUAVYa216F
KC8cH7Ka762rLNvWA+rIjiWymbnGEC4yMGAZvzUrAGpFyiN2tWUw9y5Wxnvq/EKU
O6zuhTGH9n/ikhne6Wfb3Hhs9hGRx3a8drAVGcqlWyu2/ciabDwIZNZYGxdStZU9
rE/lXtpWcibqB6CDPtyRp143TmDEiWh9SqJJbhwkuWUFEuXwUlZ+LWVB74LKvJE5
fJ0eWLiSbTiqyJZnRR2tqHj30lFSSA6QFVSVJ80IBTJM2w6JynQh/HgIzwZIKPNp
oRx/JIIfgevfvCho/pPi65LM9ZU/+kzk7fN1DEiDLDP+5nSssahZjwNpvh6fH3d7
pk4nHlZLTwCSx2rsbOPh8qvpnq2DXelmGN0FT9Ibffv9+ZWHndmuwDJUpdYJ1E0j
QeM/8BZCKP5GcgwDHtViPW1n//SfmBtfxN9HMnLgTSCz6icim8gO9DGyEc5gIJj9
8ggAjHmJCuc1kgKXOyjAExiJw/x/R8tSf5ex+YLDl46Zbz5yiT3rjCYuJF/JFhYI
XfEMXSQYvENYQwz/tU0H9eRKwndVDhX5h54ruO0V16am51QGsmYqBIYs2EZWyMVt
rKZW2Lf4CJAgDL5dXZXvEEz7JNmDdSBMwWp0B5kro1zlFjIXCU5xw82530JE3U29
YyQoVUuN8F1C3VayEP37fR9dkjvTUMzxHqKSz2EXxp61KCiyMk1F62UNvhOiw8A4
PafmZ97n3qssnpA2WwjD1tkyckU3pmFc+3K734oSxXrQeI91Q+tAc4qj+hBbBE4C
pPHLQYzy3Zj84RqJkbAHPDhJ7nx1N1v9E/rMmFTMN0NpATMyIv6NsnIIfMWW7s4w
XXmCow5OCAkRq1cyW93+eETIuxADp48Bg/iZk3ty8IKIVI1HwpeRktCg9SCtYlJz
wwn56++NJPPJbH7+o98wDDFt8G5t8UQ7K3uZHcudwIFp1VfzphtUkPgJWxmzeomF
hjkXDo5/MG3VrHT9dft3uvNZE2VzDfeQSB9+/m39ZlHGg6tLIT+DM0i/SQbxOMSV
ugXg9hQXVSrbPtNhj3GIp5lQXS636chTMaEJDTFlgXV/w/OSaf0KFWugIWaytZXZ
JezqNqduppaexNitqUsFSaKqR9NdMHj4wrScFv9qn/qFs9VRWNZ7ibM9ctYN1IqR
z6qYIEYrPUFdRpKF+PVsOGQEZW9pG/6SXkS/6dzGKqP0AIyajKzkzBH6BubIVYGK
bp8eeyX7KORbN3FEOMo/XZPbR6i5C6JeJfnqqxDZ9aaoQK96VjddRjSTy7jzxj9C
tkGeLLjis0Em03voj3w21rSSspWPRrq+zC+RKnOd8MGldZ92fs9Mnvi4mR3GDBp5
g2TUA5KFllZf+k4RqNBsu3T8gEAH34O+H0mqLYO2jVydPQls2aAir4uTrGTYbEyD
uQzcROleJqjNUJ+DMkdkzJb/cBzKN816YkntxHSpGuQdirw9ZUBNruqwsZtW3oNa
NxuRlr+HnqPso2gNvLpqCE/p5AI3tkIwf1mgjqcjkUvsnU3N1CkUHmTtDCGn2ldL
1IduCBq2uihc6Fk+B1+Y+rGAGG2VcG6WbcBP3TFG9MptdxJbo5DKIiD0RIABRG4p
ZdQ0QZYMr2h9HmDc0pACwe4PHVowDydAaQc4v2cUGVoOJxw5JyTOVh87XSoWQb2r
go/WQQFvuqT4JOSj/ayKNt9EO1Ewb+zm+LwHrNOsmV/lVx4aL/FQPIfIw9aY0wg1
r4rOQ2ptGc1GDd37QJPuAUFE3+4jPQvIu4e3Gj8sjsmoR9ukyjSPWXH8wVfi3PPC
6sJZEPPyOmvBTEc5S0bKwP0SMpLu5rdqkZJoivsOF61scPz6blHxPX/hq5GraZhv
omSfaGAwAXg+4uTp5B6pY8NCX9G7TkcZwS/FGgoy8i0biOqQyUcP3GQLz99+feGf
LOfwcF4XJwaeNerrQotn9vM90yjOl1sglNRgo4qUe0odJWhTRo7jJEwY0DrhMxIB
RpbE4DUdxmYqVyr9TlIFsdMxe61u7lZrvyTapw0OMjCF+k49LV4a4m//ZVjiwGit
NZZlIdEyjHX/Sx8BW7gq7ytO4fbCB1CoQU19bbNOUps/bopH/p7OgCm+7i/PAv/R
a6wZNSxJCkD4Gn7SJcTVxk4urRArJEQFWCt+dRwXTvIGp9++rmim0xv85K6sWUXE
ikcE7Dg09EmMdSJIue50Lj5vCiW3Yc7Z5KY1TIzp+ujqWesyr2pNnAmBuyaI3FLm
8lGczWIAzzAFMdoweodJzKS2p3CZwfELkZhTPr6s1XlDkVXw6vtWWNo0icyI5kFE
2zbk9oKD99sHqscvRhE9qrABqiEHVmNszfu7mWgZMt+Ta2vO6ywhSWDBlvmdpslW
2+jozD+vCZLJkM1jBb4v/Fl9TZa8IcrTIGa+stOxwo1neOzVuW7x09GyYreKHbUg
wIdW39Gk8Taawk4WDn35O7DyzGgKlcCoTmvEnARwTYYwx8VuZ/dfv9iQEHiBrvW1
9KStaUMIYSVadLZEfQKip3MXpg7VymA9mmvsfdhIx4WnbbeEm3twUcT1RjITn1vT
HBeo7iF3c6YTt8oflUEk5p9CU0JcvoijjUbG2m9RvDhqYFlaqtVVUTSDsW2Isj+k
FzkpQS/U+tLMBxx7vdXUkxFbMFuTTVXJrgRwGB1G/9OZ9+FXf9mRPV1Pwadun6Re
WqAe+NQbIg9zBQnItCaPopZTZLD3T+rCNyHZQL+Y1ZAydhA6+rzDd8MLnB6uFLJ/
eE/8kwYkm6mvWEMVtORz42Wz9QcXUl5F2NYJSII4Nmoq100RCYoorCz7zThrpi77
YHhzGpQG6i/QNEODQXhMMyT/wau1gSgJw8bNyZmPep+FAQcxvmSM2cPqylVUhK7o
pJeyyMSgOSlySgzadda7nsak1YR+DtvTUXJx3UeBsTe/0q7NToeytKdrh04zrCu7
q6ZN1cFzxTd0CqxCKw2f5LZapFHeHwrFB4Mlwzmv1ZmYpYbsuAfQO7LDDJLp0+ED
79pAfLD9m+nAuPIdRINOcrd27Vzq/3aWt3i0KW78gcCm98NoQ447A1Gkhv83hrHF
/6pOLDHjEq39xz6JX81kdAbuQHqs6mbmwIsPnVOm/671t3+X5jUVzQaL9Cpu6P9P
whLDC2K1kXx4Rszkt2QSGHCex2WxRQQMSrSPz/4RebizLni7/EvD+HuLGbZ+ag1P
Y1IuSai1TX997NNfFdqbsqYvQIY4hOXB01ASI9uQ319SO0+QEy/Xa7d85FuNos8J
uwKbjgWt9hlnXc7G6CwUUly2VJem/BQcwINJkBqbGwX1QUVL1n62B5nWGatEXFQ5
wT959LzBmqcdEA+phrSK9/DWv7TrEu0NBunOrKF08g5a/3kgSpuV/LrQgWlOki+O
lUbSncmibQMddD9YWtwV0+YuMl5APr1nw70KLr7Ifgbr+tFIgDjwIonIKCh/By1j
66YvPwSziCeZ+y5WFRZecevIlQJnsEC/AkhDTwrOq0OAzRrvlsl+CuDa9q6ohkpM
KORQINwj20iq1hYIA00EB2QeNdY+Bfn/ZbwShp1Bg2lKgCsVuxQqX/uA0iNBlQma
MIPjRrwRHIwJGAMMgjarHpYuJI99ljd9yNKCBohX369cZC2ZAjjErOrdBdbM25Yf
r/95C0kTPttjAcB+D3xqWzOkay4nVaqFvvd9PuczDZRZrDJ55pb5qDd2nrfMx9jJ
NIawgRGb7FgV5N4YDxadfyh7Wk/iY3AF2aTt6Y7Nfe6DBWLrfjwXAIGX0pOPbMzb
rOKjCIsHkU9ojVfgWAm3B7+2wD1L5tGk15QiPE63zBp2/sfORblXztH0+pLSQBJg
0VzTPgrdJRLWfBWQHNJV2pBFZI/eEapZXK3bj6MS0k7KAZzBq2G/UB3n/Rj3klfN
Id+3rOoNUte3h3pJs2ewtOKlYrI6ciDip0GjRpAm6jS92DMFX11bqoPW8ZZ91gfw
OYGSiccJ7NtU33n1RM1oKnJ1REOU2ItPNHHc4HI13X/JHRdvHEh6XGD5hYhb2vqG
1I5B7YRkZnfiTItNncOCPRZNnKRJCJ/Zhv4ad4kuV7cd1lZUlxbzP+qWP2l5LYOj
egM2gTVULmoFIPs8rZhd01bbQPb0egCoPP4yyhWeZPQg1n/8BNSRBuPaL9qTXLvO
/vzrXWpFHHJDJ7YI7JU3TPd7NawiqgONB7rceGUUzaT4YG2b48H//9W+FO1MSqsR
JMFmzmn0FBxPKcA6dJGv8BRYLjQ3loBG1DXi7yMviGlmETJ+G//n3hc+1r9aTvX9
Fyfa45nvmKbdhStreb6uQLFtsLiJ+OJk+vrj3zhHaQuEGY/+CUhvBxMixYLJ3kcZ
ltqccDJj2yhF9sbRQ0r4iZlodPdJJE1+uUHu8z1coQsDRAPgJVP6zTDM7znz4mEW
wb9X4YukWzHVBDdVrH009ZnDDkvqUai7PTLVnEmQaH1f7HfTcwvrVULxp1ep9SFW
Xmi0l7TEPXpKY7/wkUL3D0fFP1bwyRSJFCVO/ZZQMgY45QUDcP99H1QpU2l4+7sK
II1a5PyMkkQ+wuXCrk9sj+mXN4Lp1TphS4vc7Fsuto/pXJcP5fthFR5RzlGnue0j
PuR3ODJySSJJrqLr7JYlVBReXmmpFZHvVJL+XWatWBlxk73dOBbTwGc4eFCXRuTQ
t00WEAsb60IeET54vNESCrwai/JSe7jCRLI7cZccpkfsvRKYZKwsCRNEEoUW+q+9
kL5tG3m2m3C/DfYC2QXTGBM8mSjYw3Mr3qthps84JkMavNzPMcgnkzYxj1aDtyMp
c8eFf2yZ1goxnYD73VLNQIh79Sy6qs8DnaQtHEHBulMrsoEx/GhTnoRs1GiJJ7+y
okw+Z/xZp3VvPUE8ydoQ1hJjyVgFwd+wSnLwiSSTQkZyqFgerTULqQgRMUCDgoXy
bUuffRYmrd/SXwq6NryD5n6OC4EE/4as4NGNXVM6FYLofNu9B/vBGvJ8uANdkGR/
CRMDXhN/PkJmC/bDeneuVEES98/XS9lp/iHv9j4HwYSxPeUABvVd4kk0UFZChgEV
ZrJBZ4IuhbqjysgTQHJoEcReNnGw97vAmJG0ZgYGSEfSHwJD/yAwEVSXA6Ffettu
8VCSCR//g0BuouHo7XnbKLM0Jn+UCXqSiJiknVYK3oNTkmo+7T5WVyB/Qg3FGNe0
XQP6ygKdvGIPVNiz5ktH3jeOkU/adVFHEnV2F7DqlsJyEQu4WYKh8MT5xxO2MJcH
1bHHnuat4fq97poXeNvfPJ1U6bhHZ4m+Vij2n/R5rQIEXTl/MhVQ/1grvCKSPsC2
bxO0TP+esjdlrqyF8QOYejli7qSGVHwRn6HP0h7uPSENrZ+yq0MdgZNDmMcSHdPP
vJxCxBD++/81K0OjbQoDF+ALm5upc3Oh6VLF6ueY2jROmePPbWhtHcw+PZ43Abnd
hBEZHTZolOScAb4//He/DFEoIUlSwiiTitkjx9s+AM9VItrLeA3ugUBx17K0J28q
fXnoDvGBvgcFmaZespjG+jI5+0OsJUlR2mSUwFKnqClfQkyR8yq2itBEbvzZEXjA
SRF5jF1Dj516SjeK4iKm8cWxPmmD2QLvYxhQ1O7xZqzDtAsGbVTd3vmttrcmEsZs
bhaphOooluJKMr60hirpGpH4iQONDMIKmkMVX1hh8WpVr8vOdpSpriJtkWCH/bLZ
Scbsww/jgy3CrNT0zsB/d5jA9Adnc2HYao+VQmqkThuePWOPAAfP7WVHy2rLtq2A
5cHYwgvI2Q1PI1oPgDeGjIMk2xG5fEgLD7BQy7b6Tf+/Tfc1IOXVq/5GAwrLmqXD
vuVL9VBfGqCs22KcgMyKEVeB9LiRR5/x6Gq1rb5LCWx17NbY721QOM5VuFzp49yL
L9KHwdluxp1bhUqksM0PAg0M6WLmEuAoZvimhjZfbY85mTTmIJmuN3YQjtU65L65
Y3Dxg5mLiiHpUgck0SELxOJP14vO6XDPbm1dcZP1NHlgsCYDVSbNMX+AToRQADK+
7toE0xDkGrR3p0dCrheENrNFVRtxuY11HrSkvKFeTfI3z+8hs6bfgitxDLqx1BzU
RD2CthKRAtThEXJ+Ag9WRq+UTHJaBp07xjMnNkBSGxQnCoYC4fqpElV7oNLzpdW0
ZczylDVc3vOSGXqkJDP4gIJumtl5w3pQgakL8aIE6Ex9LLvKQjWSvMGkJEacKI+f
1y228vgpfhTY8djsiFxsawOfd8uZh4hq5XxdLlF7Tt5vj3D0lG36z4ATAAB2/p9N
L2ljbAaqAeIoFCDH49Kvt8VgNM/OCi8oSpFP1qTvjqhH0wCFJLGU3PDqbRVoi+1z
f3ggWk7kWrHppths+77X1Z+kOrWodcliBKGJCxtk/+Naysrh//WmpXx3P3TQhVbZ
6vwnAhKJ4uqNZfySwVbV/ENqJhJ0PnrZuPnrKCiA4YguEEPu7se0PGKoMzyboziB
K3NMoEV79ZeIvg8K3jEZTB1fbqq0sE+9HZJjLAxuEKY5qNfHFwhfvazGKNhQVepj
ir4PN91pRwX/MOuXDUINml3FxswIgf0ljR2+PzJozdCtzfjKp78o5FCZYMqsnXHT
K0kHhxtzc0Ex9BkZrox0PFW/cQ+OFxICmRcyyepfcLsjD9EBuu5RTdD7uHOaXQfU
bD1pmsC5eoFsPYyOnUhix8DA/ghKNJQriwQwQu+Folr2E8NTosmu2V+hSXVwp6SZ
+/4oWtWhVyyYlBjB1kfy8P5iLcyQPToZPAIgMf65RHLs8pfjgXOt291cyfI3CxZ9
JMoprswMC+cywMy0atjOq1BDoHX2JdPABbNRNDV9EZweS3KjLd9P3U+wkOG85w0G
VzciCA9oQ1JwanVLAjnuprFHL/7F2AXJvrQn4dUhNINUYefIKdqvJmhkykmr2XfX
/ugHdJCFvz5N39nrki/ABDVEjadH3O7475lDGqGosmlJxCsA4md1FCmVod0y4pd0
VrwWfBsvf2UyMU25MKhyIBK8x4dVTL4kTlA5EA4ZflobCRASekZzcKO9Tu/oJ2VK
A+UADlANGczetdAmlOuthLd604I3ZOlLpLotirFi5zaaIzgXHuodRmFByWR9BMtx
0yHkZHbiJQHaz766US5SusT5Tbqhah7K7tRyLTL2dHEU+YmH3rey4wM6m4IqnFUl
10UMx+rjsFM4Ali/UkZ1+1Z1AcZxnvdwLqabvCOoY2UJR1KFE3npNaJ7YWF8RLcF
u3CHVRvmNs5CwUVSNwkVx45iNz38bb5/S271Jdw+CL/3Y0ZcpG96wtkTWm5oLrJv
2g+tmxlsUcn9ZEyyNSolKcmwpnVlQszssv2dOdQ10vbFuVj8tboMm/ogNbzq89Gf
Lh0q46B0vlAA5twor9T+EjSqsvm/hoBFQMFe8bFt8CctJzkNtd1bhdD2t9DzxMDC
xP0IoNNTdMLhd2d6xGpWTls3okS0DWek5MmrfM707cuSdyxyv+sEoqT1TqZaEyGU
skS0s9Ld0mah0RxvNtRt0HuEtRVF9Rbq59p6Y+ftMSaeh/OqCNn5VSya+ZYg9a6f
nzoUQ4Vm/uNXkxpBHk2NekF2aQEL8opJ99coe2biv3TFb/ZAgw7OaGghyUhlhWWN
wZxtDOaq0sJOeWs13qFB+AyzcCnr/fholIGRf+h4RDIdVDy1GdkkCIh3adLsYYhx
CkUnaHXR5lyV+y9NgNN0eoGgtGrpP9SprYqynDcSjx8Cvyaq2KLwPU3o71UCY0Q6
oHoW3qeZ2NRxp2xqVMk0L5bsNWKYPBHMF0XsEru3ebotRjWdqZI6eIgmE0c6N/XD
/AbpgK77Y/ZV6oOCDar7d1Tq/Ezq0DnkhitFNMyUTfNMfD1HkWH/pTTeVs9Qcf7c
POk7xYQ5TbWRD8FlRPtzQaYFvBxhv6SEJxfUkuMzRCj9druHGBTlg8VfxcO504iQ
jHK2dkNwS8AhA4FIQJAhh2LVSx0HpDcF25Qa+KIZYMl0tq7HxCyYuBOveUmLgmPU
xBnKMVKlTrrsWhVXejtXmr9CcOFksHGSQ1pNQNdY5XHPxhqXwpxCD7q18k90NdDE
8dfYnpf4lNVm2DjUgZFvhWQ0YVs3V1JXzdy20SOAZHRZ9kpeZMl245TznUijqXip
hHq6ChX2gJdzV2wUsLP3E2wNoNZsquf6xeSMVHwqX3BuPlnIQSLGbmRTXnHys/CE
07Q/1pwyY9X2lNil03g5wkJv/KhCO6Dnrk8LG/M+hx8TdVOuJK+NBT8KKULd0rx1
6rAQpoBfSDo51LLTf3Z1KKpR1mAH8dMD2g5El2nKgFrK6sq5mKx9QlEl1v7rqtAz
+Rt/+6+B9GhdXy2EEFyK0WpXiI8oq2Et0phYZN/L2hFRnhOu4Q/sAF3UC7JwRLlV
dYX+iDNZiRV6tWzTaweW4eLYzbgNIvr03vJa93+OeAJc+gvgfLFjZu7jlF/oII1g
HklCLaJ0impCQ1mXUfCkuzDZ2E7jYnIFsqMKoiWabrQbP+yLz7lrRh3xiY3tFIAJ
WwseaxbTIE9X+SvQKdGC4w/XU0kEho1EZtY2uchs5wNNUXzKhsJytqiu7Jn2wDcU
ev/CBYLYe2mvfJbWq5Fdfot2E87ArodTSdiu8xMvuVYiIX5uNgmp8uYU2RkGXiO0
NaCycFxe9+bJ9GyjddWtPHpfDYKYqhSvH2EIZ93LszrU4iDE05xIZlbSogIZ/RfL
yLzDV8CFkYhx/REQM0i+8Z+w/kFFK7zyf+tV3jST9xAx/CYJGyfz2ilrQ2Sk+iwL
oBA438z5seT+Xt2yQ/DhI4zlcxzRjCMmnyUYUvsYi7sjluP2TRFfy7hWRNpEAliu
JlCk/O7dAU+hxdbdJjgp6Qmu1uy3SiIAShZNoVcj1QItTZ4Oyuop083Fh4TFDaKa
h4o++fm9ZxCH5UZNHi0amTQMc4mpVoArcHmMIyqibgOnJOdVSG5F/g7af6CqMvf+
HdsdCM6/dScNWbd8xrEeWIqK5BKE1Sfl78Pj2wG114DbceMacRplucB57yKWGPe2
PannQRdztMRN8H7U2sihQ3dqZy2bjzixuv2HKphaY79/0xSiap/6K6Z6Ps9ZlYWt
M1rlvo73/z9FtiC2oj5eH6Lze06SRYJwNh++ZnSEKJl8mUN1wHvu7n23jaoYyH75
tPWvvRaVObm3w1FJ/kSZ/b17fCwSRUR6JOn4R2opozS3KmhudImI+DHOu21YzchT
VCsFsLHojc2iUNlnP3dYoqL9EZxt/WscKv2yYWYS+pEDqiNAmtaLwzX1zDVkoNLT
HwtwfQgFxY7xdcQSjIzy0cz+c+2JkOiL9g6bDWiGseLTTyAWXMk3YSaMIypx2Ngm
03U1zLbyTggzcIg6NGiPfsH22YL3q2lixT24T30NzPQc2BEUBHEow2qstTclA4L3
UmzTq1F13d12e1nHYFW3jOlvYClfp5GP9AL4BSvMwEpgUQxqhJiiF2RaYKRUAcBo
RW4y30k8yeEkP8NAZxmisucFqUnk+O2GofJGYvpCvuXbQMnmvXIF/5dqrmIf2RUb
KwHHodOVglf2ntqUpHO6zYS8a+lx8+MSrvhKQQaxKomDIM97cI9vXUCPz9s+KpUn
PcM33VelVEFM5DP2eIXW5YQO/Sox+sBqR/Z7aPpPRU5OfbVGMWcmWAbMMjUBjeMS
1+M2OmnGLiiCMP74XwRB2CWrAgMnlLAenqAOyxluKsNKDJlzDEBuWraY4SAvWj3K
bXxntdiq/+Xxf9bBvSYLSAlf26W9orACAjIZIHhOJY3GvOYs8xAsElDfTGx8a73O
KjB6s/Un2YzXgxoSfjJASu3Vze5UAA0ZpxPlpro0waatu7Oq6tUwzPanzkj8/RZ+
YuOhlLghzCLgmlKcVV3cp8aMnSzB9FrN2RhkZcFlu5xRHBKON9vyUwFVj66dcrIA
n7+9uoYUrgvx3/myHLF1uLUYqEElyLfv19pnnE6YIyzHgNEqr491+645oSFf9yKY
OxQSeR28WdEZ5JbOdlBzmMevZKc+mouxTrA4FMjgOIgU+PA2jObuU40hEgVhCKEY
XRwRiqXOLBhGq1XFW1i7N9ATuWthVYU5oXrE38DdqVCY+uvCZU3HzIHUI8m7fw3P
XCYREhXgpdehPh8u2zZuyYa5E5cRFqY6lUuuk+cQWnMYMkO4kcWK4SQSskX6p9uI
aPmMcQ+gwH5sCzsFWM/I9udK16iwNrJ+v+bMuqhuGCpT1GNkKNqEpnSwiV0UO/QW
HhvcjslQxqVI34ecCegl45zgUZfUIMgUGK7ezRbV2Ion7FXZUPtgyOf7FlPFFGAL
7aE5bGQ3MsXoqQ+arqCiOGDf2/K0q30Xe2oXrnc7RMgoG80ZQ6egDUY0vAxhQfpx
tnJw/T8sR6RiLDvUrxt1i4UgyxfrBDFlVjQoLXiXZbxunEUBdHb+Hyk3Os8j0+Ay
80B8tuhWkqDrj0fcInehiqNX2mumsyBvSp1WpzqRCWo++3S0oKiuZM+F0rSBHCIt
g582QyEni/qkkGe0CWbWvbSBxj5DqxNmk31ab4wIFmhFwF0EyPbwlNV9bxPKcEop
fny8UidaZGz6jA3vtl3MLDd9jyYe1NusTXAjRy2Ji8wSufKPnaU8F9B7TqUbI491
CdHfse5F494qUnXptJPlkYRZLnGgIVl6VCLsFJGkONaB6jnj13fQ7tj/UkGXbyJU
+07I+xYI/cdqrddWXPHNTcZ33uQWIqAjtu1oQLJNjAUxPJblyRugi+2lwN7E/D7N
u+DcYYd91HDtllj8YWRgHA51eyJcN2t6iNASkqWUhTiGyzzS4ZIwLmgnooN9oAgx
7X+kXWH8psrq2uQQeOT1QKA+WkYV+Zy4TBVZU2CFWWRclvkC6lcU3+jyqLtazd6b
SFIqmaRQLAL7zbzFWMYr5FmRfpd419ndlW1/z3hDSW3t1CI2z8MTvwYHLhwBDDMz
kRx1I4TBDtI0N6HiaOXRM8WUgHzddCCtv81YcEFyKoHXmgBsitOIx34bNUzZMye+
94LzlnCJ1d2w4f6gUVSREx5Tz8B11h/mmuDzCdmiNbtFTxn7k7S53cvXH9aGVLaL
+QmFBXcgD39Mp9acIGUCnVSHc6UCHA/Ch+bfYi5IiadXTGKxIA0I8sMiIljQ970h
1qZ0r1jrzp5X812rtTEO4qsVAhDY/8IwZ62E2HyZE2enDVRyY1bHoQw4VH34BB5S
vsWi65Mpnw/VNpZPoukFHrz6Bedx/kBMyR/ivDCnsxOMWxJBEDIZaNXgdnsl+D7Q
5TVUFBuPoqZM4j/6RLxXnGkYupKuYfu8AcvDdx4weMP83Lcq85hPBILPOvY0CbYo
XRgBmjkTqVFZmF9esvgmqyj1/hIzG7m8b4psaibmkSBMGiXnUkFvmB/CawdsWRYN
zzLE3x03YHEJyY8NQMAUzaP6KtImPLq2A4H8GspAnn2A3GHUZn09GmwcDkpNJsgL
qbJkYcnwenaS7HcgS9WWxoFkZid0z6vWSXRs0Q1/7qYe7MgiXkaNIAsVu9rcUp5Y
+BhZN3MBLk/pdQts5XE49F+WltLxtnaVAis6PvOfqqMiBJ4oH8jmk/JF4RZciso8
TSsuJ2UqTTnmNMT8UUZ2ATEtK7vH+tryP1jrKmVi+NUCmq/ggYAWUHAxOxp92CTR
24OZxu8NA6JUnyI4h6/EN6nnM2aSLg0st+9wDyKi1R+iYbBiOq59gyHt2BBCMT1L
h9dFGK6aT1nSISSIl3LVHFqOHhd9Er+igKHjoh76FZoDTC4Xty8Y3osM0P0A0P10
dCjh9hzeWbRh7/9rrzlnos+hM8mhnzOfAOpdm0w496PeBQb03gJ32dgy2/V/TNHo
tJpuyrl/exs9oxgQI2z9QHKYuZOFIZfie6JdQOYh129OyS1xsZXct80nwaR7wacg
HBATVA8Xiqur9FoeeL0jaQbycjde7Ig7yRQK1gnc4DqyYv4hFxJniqCg2Yo21Zpf
VgDkCyp/B4VNGoZFSmUsZMinCsgJlQNsFW8vaVHiIqYiHQPLdaL7gcYZWOrhjcVC
GS+Ui6msvN5hP6w+eu69wu1v3FNhLXGGfuhb+0K/Foa47f0A6KLR4gLlXxTXZDU3
GqvgSRpnQ5+AlO2fQWwJhOpKOTmm+BZBu33PfamGlRT0n2qxcrI3NPbaNNFF+i82
QLkwWk1Aufer3famyQjvGLv/A5iIZzL/0ZU6l1/rX1RG0xiPkgfghFxrlkuKyvoj
pGByczD7HKT81vAEp5c45UM6EBA/RMcY/RihW6eQSvecRTvtmrL8ryhHLqrk5qUx
YZrknb1IGKukZDO50Xvmn3BfUE7a+OLSraqK7s8ki/Kl+DFL5EZQgFsnmmYqOlHS
j+ffzNFa/NZ8owZstAEI5MAKFwNhyGQ5YHZZOHz0TVP5Ohgzhtd9/v7MdBQqmVhH
ud5TT3ZI3fVFm5wpyDinlLIyuhhG3YurBRIvDE0nJyIjq8Nf4cAr9qO6/ljS8BKc
76lFZE2GJFBdx8HljpfmlMbg9zq6CrB7/ngjHGEaFfz/8FfQnC95nPtXlETCmLKc
MGdEuzI7KU/qur43v/0ywpaInyQz/3PNL+4dDgDPpH0Jqm9eTUBgmXV/IgZJ65vy
wl1wFVsZSRwiErF4upfbnZINggKoQW+oM3nKjYOp5kw3cqnuyzMmTPfCCP/bQnC9
+yzzuLSnZJDwVXB1770Ngyj/cQFYIDAagsy4f0Xeb9Oy+mLbbng+GP7QC86STZ4o
fSIEF9WFOYRPf/CbrNp72KyCpyvA4pxoS/ahrUMngnhbf5nUl5S5+SYSuZlleu6c
RS1Wpx9etZwRO7YF63ZOrXDjZCCaD2NkEY6iZC4laNsK4JEwyjKPEjWso6QZ6V0O
B+/zV27LLl+V3UucgPj+Za/fgEJyC0sMErOCIjjRDOgb7MrWYndl9fhCyfXBJvhn
zM6iTBvCwrUzNogPjxEX79+Te+4PQIUcK0P4r+LHwA8EefIc9qYEqkJXVEmr9aPy
+dD49b9JMD/HKBhDrBCmNnIyGwqW3aHz19Ev65a5oHOrSPRC6R76WcQAtmEPsc3m
YwwcLkHrPTVlhtoQjWcGxQhRjtmj+u60gw2UYjsd4PwJyVyKVAHEG0q02mPerVaG
if/8cXkFLPJR+sVuoXlzYJiOtakl4pUAI/vsBijIdBKdV40CN6+WOZvK1Ohhk1VW
WxIF/3FdE5xBpl6Tm4Dd9LSjEwVeFUsbpsYaczb8D0H1jONXlTGiwjm6Nhvdlfu1
BT7Jhme/86m5M6DDtPF0umXMOyctKWSzcRyUGvNPWmVS+MT1fyr4+JELn/89qwBW
kTphw4vnyklYcinuudNJjIrU9+iez1ZrIjXkSFNJP28XzCFuIBmGrTZH191xeqek
KMe/XG61/49hcXHzPKk/Kvc6kF3/rJhmQ3rmUPzFKXp7d2nKBPZftkohDEc4YjZC
v88bAAU3SGvPOg8f7s9YAEXzTal6aDJjZYi7ENLcYW0sSNjfSlh3ur1oCJ9mCywk
Vt0Pqv8BiBtRLTgtjLd0rwJuw02rwC7Yx/VISAj9zpI8dSXP95I2farhr63BeTr1
N9lhpOjMWApDXlcE6jSzY4FFGigdk3ZTK3L4Ho1v0D5HLxtZWFM5wtJFgGXdm9s4
6Y98mFn1PPNyPAwpcrTvO0Z78Ds5MBKkH7o5hOO6f/P/Nor/Ez/N+2oglgnwSxtO
sVnCaAwRfBpZZ77hprciCQNI0WVru2biuRHIPaQhTXjTDLmnxpA/wl+HvrfbxmUx
bxT/whgvDKD9SoE4CGf4ZarpGCXag2XlLxEIGQd9ZraTwoESeVbwB/OLkeZrDIZu
Q4op7ljsV6yqlGmO2ZERsxrr5yEsrKGmswUYmT0OLw6xOlfr422hgcwcLflZeT6X
AgW1ZR/xbWrKs3403GkCoY2R8w1v/Hq7okaitEfZW2lxiXVaGfXrRy/sdlTWsAnj
/RiNmfLasY5Iw4HOP8wFktWbtJtFVThyvJi+B/Uy2ZeFSFCge6g6jfIhhLaiDq0Q
DeXRkxO/Z9/M552AvBGrtryiGkVpGF+Y9fCCFrxZk6+gJBgVfWujxgJ3zpvG4nU9
QXBRPUDY1woIBoUav7eIlaxoI/XRx80IpvX0cnoyt7ulGUiy7tE4H85oeV0bv/eI
EGege1GaSkA9gn4XiOCYToLjN6dhry6jIbQO3NJ/TTR+ta58za0dx8TITiVLyYbL
5+tEYbKxXT6jxCoYscJ+495leS6OW9sP8d9zo+6mK5T4fZhkT3Q3QMyCXV78zUbs
QfQ4Gy5t8HD94NQFOCmR1MhVwghE7mM1dH2E+ai+xbeuZgwPse7woS88aJIlHit+
LRbMSwE8LNtnonRDvPN4IH7lVIYrZjUVgadDDmcPnr/Z8kIhLePOkS5lQbXJHNyq
Zb2GfOcsap2LDmueQXBuaf3JfSMZVesRAWhT+HJHd3U=
`protect end_protected