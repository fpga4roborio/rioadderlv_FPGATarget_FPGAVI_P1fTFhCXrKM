`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
ddtXksX2+yylW5zu6QL2Lhnb2d1sD00763mmSITNX595NcHTEkwn0zB1Dry37fOW
FufOhVzEJp80NC5qZ/+F0Vk7Ik02dIR0elf3clrjeJRK85K4e3Hoo4xn7YbFUIms
l/8VZSb14+JVGURjfswrIyCUotIzlzVYZ6gzoZwDXIi5gQIBf/gI+KxNXPaKV+PQ
Ufys/12rjO6aI/pPlqSm0hCvftmBcnezN2hk1UeXgOIuKZnogjOsf0iJVX2aOOWE
6pD/psybjbnsNB6kH5uFTA5frkzIzkzl5d9+YDm9OyC+k84E83I/7/j+rk4L2dah
QJOvksSIzN867/4Qt8qYTQ==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="MvBXkzurAa5VTw+1JJ70nePUfoQXBvZOku/SMmg4TwQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
oRtzZL4VJ4iwysPsC8SXYCzXS8Fw2gtZTOskLcDV+1B9Nzn1zTyNtlo6lNICRmmK
ZRVu2BmCc2G+fmzynYlNTnSa7C0Cuel6FYpxCBlOuk3OF2tzAmLAuDyOH3Z1Yjzk
a0aHuoCdIRKv7BrZCdALt03JeUmXKPdOmIlkVGFl8yw=
`protect rights_digest_method = "sha256"
`protect end_toolblock="Jn9CQpRhJt4rnzZPRk+dOpzAubz7omckX1MrFd4p81o="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 20576 )
`protect data_block
gD6l00tciPUa6pDNTk/+t0OO0nC/UTtBwLB41d4inuAUA3i/ALrNyoJVcBnAmEQW
ptbcNp5fxEUJjnOxnedyZEuEBxWRieZFQnkRdF269oO1fdn3IMSlrBbkxq6xJqwm
D8rzfuOaU633gz6UDdydq/PIPVHyfO5gIzSlVp1cHXIy5Yig6bEzPTpX6RJ+2jx2
bMVAWoilelUJ4NF5DaglSCgyQLXPug5H4zjDG6ncHXqlVG/9njeyonmLfXSUe0Nh
YWLrJWdnGg2k0ma6ZiZH452CRDOXW465LFy2ySweOVRyyKDVDN8cEXg/vCjEmaBW
Rg71PGgoaXdKZEQ6qfgQ5yUMZypGYkJhjiwEhGfM16ZyIeEUAqJ4E/PWMMst80Bc
BkNwTe3wxsAsMF7r64DQBtAVCGSHdHYgEK7M6LvepVb7yM7BDUOZaX1tX2q7ig94
oDCsyM4IxXKGk1N5gWXkBaeDbKNcmVNaqjh6zhV8blh3G1cVpZ8aiOq21FW2sDIj
lFqsqdXguWlcSYYC4X20adUjHg1CBucwu8PfNaBA5tkEyeJu6WWYt6/l8Rbd5YcG
mOwQ4cpezpMxMmZAZb3E+Un25EccigEVTxvhsGi8gIsNUJPvM8z8uo/f8iwjhbpf
+dBKE/rrnv65NaIdk8l07YdogJ7m+6jIxFk/msKJrtGVTds7oV/Peu7BW39LUTtO
vacHGrjbyIMMuj7W97kQ6bOzXJf18OIHrLAYRrKzjJu3EIOX4PZh0qV3vXQVrN59
6gvli/GS9bUogxVyEXQky8fS5u258yMgKlcf/G/dSXBGWqP5SciIeCNedX1oKw5o
DM76GQBNFaLSH5z6UoYsotRRJJDFCy1JzLx054PGDb8Q1JImyPRK2ULkdWqKp1pm
hR133qbN1GKGxK/eRmUDXPT2VTDWv3qJh4jpJOIDsk2vgXRI4AHKLwih+YLikQ+s
P7qfxPBL1FaneZbCwO9gpYfSVCX/gR8ZFk5O0+5Jtr83CoINa/arHc7LTK4z9248
/2PCuBW8oZqX9rydMVxRDdydr06y8rMAoXUkmt23hGsz/0Yh0812jJfbPZ4PQqdB
7MrY8UBztifMIkJu/aZ6GEuDCN+YpgJb0JqrN6JTaFNuIMpZz1HomNrxfSzdhVBp
24FIe1E6VUWKkr8TOOoDRB8g5jSKiMQba0CMFrk3sXepw8HneNpzmTqjulD5Ortp
ebO+4KVyYW5k9hesgVngP1W/5gGRYi6AfZb3u9idyXTX40eiYylw1B4tUX6o3k41
zg/A1PJpPk59ojyEQowH5ILZ+Xo8+aChqs2ksgi7i5F6gDkkUDKboQKD6Tah1pN7
JD1/wANDSOUdcLdmM1+Wd60bZKvXCqo5BI5qA0ixzlvvLr6JAvT19ENxf3xylCdQ
9KdSxvtgSmbsGu9FEUPjHkoO5bNrKRh/skfEL3bkjsCbAjTuOTTYk3B2ZbU2IBkg
UlNRlDiMEoMm9X8aJtbYw2DINk5h7F4D9cmQucEqck1/ObOO4OvW6nK55+M9BeXy
yuRk0iyz9GSBDUfCMw07lA1wflEn4iR04pyD8hearrLisyaR35wFAt/tZQ1KeQnT
RzzV7guzqAl9tyH/X1/NaBXLHLlkr3xi1vuRmvGuwN5Et6BgUIhl1ou4EVTo8JbV
K6d7jofLXHjiifqNspCY86HvalCr/ZBQaZZxr5erQzW8kBW+Th3BhRzdnL7OTCkL
6vizkO89simkXzfQ4tDK0ERs1fKVusYJYEysjY+UDmzDnuT69M+A2T5E5U/6E+Fp
nXa6V55rxoAfbIyQISLITqAWYI5IkcGL84fPDJCSKmAyoJgO7gQzk2g9UC5w7TUo
0xUZZpszPwAx3Ay3ypFRoiF+qhi1RzIEO6zCBL6NBvnBThBMEXGxQl88oLAorTll
IYYWyyHDSSIjW4GyNR3k8SbjDXQDnGGs3dO85aJjfrLxu2vQ4iTOq8iBhVSZW4UR
JBgIFrKvuR7bAGqSSWjawziwVglQJItUNfjQ43CC7y8EARABGDRX2oVDcV4d/TWR
k3qBPjWs+HS4G+9AiCvXKg3jGVKWF6dK/9Q4RrWbassTdF9UfIUq5s2L0z1UNVR8
7XE4SqB2v9RP1OBsRd56tFnpwgccrmyEl59zbZ7m1foNaUQOfm5b+qygX4DQohxX
B7uO4zqk1lTNlEOpTdy+Und/8gdjSYSyHOEHHJCJYApS9yBTBvnA+cn9SU1k1aKb
VY8LYow/thqc3W3S2aKTS8KDLQtvkvXTl7up7GUDdlKpbC9VqFa1zX4iwT+wzGNG
6WpyVugKhLXD2vWAqfqlxZW71x+kRzkD8L7oAKNA7blFNVb44KgG/0qmN6US3QhD
0nAxQZ+3j//0QddPhSKwKy8+a2k1a4wyT2jHaYWWiMylEnPlhilguqE7jHl+Jwb3
QUy821c2py4Vupvfwpj/cpo4vsaT5yBKZI9cwOurqIsxAMATnB6pocgblkUOn/7N
y3taixmSm05+gCeOXgzf1/hYJpjnEuBQGXmdME95VJ3EGEH/y0rIRWXeHxOuTbI5
Y8YHBe5IYRK5+GQ8vcCc8tv2CM2G9/8i14Tu7sFs7W2liDbYgM+8i7mJysRk0hMm
EMbQx4xcWCPdoBWlGCkFyEfaUobLR5MGwf29QNTPdhr3c6VQ38E4EhB4sbUBBteV
miuPtj124fDqzwkFkt+q+EiQ1xNZiUCuZp8h1AJy1N9HvmFzms66J/wBIPnJhfmK
28iW/ShbG99BbZaPqyW5HJa63cdw2Otsnnw20ZBUs4d2/j7Nc/CyV1+MhaZg52T+
S4/fFonv2HhYwMPfHqUEyUkG/W2sqeUy8T1t/1s4NyHYOmyClTeNOiB2Vc5rqogC
m62faSizKtGhz01GKJ4UguFQocPwmIzanyivPMLTkZVEGRYqGnDZNxiWL/ocWjyE
ZDq9vie6gxzc6LvNG/flJmIhma5szRNv8w01GDd0FYBh3MU+wlgxMJ0wkTkMl0gy
f2rEcVDSE1aYQMZPrtsv+odArN6W5jvZNSvcuuRTapevDvfdQBIMCu1d0z9hTmAC
l4lZlCQjlx+RFErEl+bMu2FqU2XCopcCvcLIKxx2KWjKuySZpruK5uu4rwE1JLQr
H/SRkgNsA5n/BTqUGZTsg2mS97BOuwhM7TDK40BNhqIWO/d1PpSjIzkyn1+h/B+c
ZereeEPgv6YaMnE1gnIbe1sb5URV6x+uMOfSrFko/qoPPBfg3j94mfRM+iaiI1W0
Y4yxhfX+WJKdU1TqS/rjSLk5ZRzGTFeEBibM/PRTiXyLHVeZ+aGseZhYeSxlYwfB
daxwmmA2atsbrrTd0qwsIAYjHKEIcxwAI6QjLMj4UAX+wqoNk/doG/X5B9BSONCl
Ixq3pnr50cOotnA5jnIG/mGEE6UcjohjZVKiFB6XfNNClxQWAV1OvNZtZfUsBF2n
P6nPrZZBkDdl9Rmk7tVToFxenEHWwAeVDEmclMSx8UtKAwQMnx95I4gKy9ZedA73
02WmrwAtB2aqa47cU0jjPEI3npbOZzhNSnSy0VQzcOT76QSBtWgWO1q7SPRffPgV
gsnZWmhLgFHaikD/MdPql4+JKQAO3SKySatijieOJzgMJDcK6R+55SEuJseE+Xm4
XDqY/Pmq84ZdbRIGTbiK0EqRQWc+h8B64YaOn1tLzUa5F+NwcrLGmTBVGEzWe49S
d4saP5JqRvYh+CBrEqlTdvmTe/er9rbcp/u3h6PfT1I3kguWiL+bRJeJahF3bMFQ
9RTRjI8K5yt8E7/D+SoB/K8HykZEr5dO0DtWJw+B9ECTTftPYesP6tkz6TsY3JJV
bkfY8JvTdBKI4awNvkkkeXiVkIi1FuuSxOw7XfNHB8PsjL3S9wiaVIRgvLw1Fype
5w87pEJIPUPnHix/B3ve1sDZDLotRqH8N/WMHLaqlKZQclkqGj3549PX8wv/Awgj
hFGMyKph91hHnTKMyGmuRGGTZ+Rr3jxwYWC8oO5GpoD2KupemaE0h222nsfiEt+V
7lqb/JL9/yEurEKXjIJ/7o/rCbmORGXbjevIbPS3t6ekoWMIKV962fMfKcHPCQbj
hp+N8SL3d3kGQMyYJDB7pFt4hd6XXdvveVNaYoB+gfxq2W79F6sQLz1y0bBkEQxC
ypbmNTIxRolQSsRhTKqEanRfunZC9iR6o1hY9Rk2EPgt7dNyevIphZG9d8iavh41
ffJrezI/OlEAyJqd0MT2+U4DrMqxhBn6dmSfD0fYeQTskOLCTpti/AL5X2G09xA4
0YIQf9UZzqc/x5CEtquCh0xXCjo6mShTjYD+D6gdSV1ZSGYsFMViC9G8SvLj0pro
d7Dml8qZU70UdGk1WO5wl3pKHtXMN/iH6fnP0IaIGpwBWRrg+do7CA2SGTEBahpM
lO0/ZAdHlm0NEdkejtbGlwUAaaNvy0LNsgEhcHjegocGOCWpGW0O+owA84n6Swva
CoIMLTOfqjvVV2ZB7K+C/1yHGFCzh7snsLZJGj5iqi7XGoyE8EEKcqHcOEJawjYv
MQzAmLcuiuN05/HfNZ9FQSFweDiNiCZDzghU2m3XNM9MF0xeV40NYTHI2PwWOmRv
0tSIK0b2KplqzjNZS21INclH0PhMFssTlU3pHm82cRnjFZ7kGpGbgQXpKvIaRQdH
QsBX47s6SMwvNLu8RLzXT2OyquSBinuW5cj8XmLpmDQSk9tp3Nj26Mf48tfIEmr1
sCcQ7Ci0ZJPVu/bgNMlEykNENlAGncEIn7Oug0Schbkj1/iGYnXHflZfBUvvUPhj
3u0uCyH4AQqksWRxUndZNq/koPd/6qZS3U+6uc9Z2G33vC4NJs9S+VoojHz7Nenz
0Du2FOwo5sZ/wz5vGR7gFZQXQ8Y7PJVnbAGwWj5zyVgxqtP3Cmiu7DL6DyCCb3AR
UZQ1WTo+JKJnICYQxmapAihI7l2OfzSgvkMhqE33LHNrnYB5j1ksuPUDH5FFsagZ
BGVhanwsZ4XVPJ1fyWeDKGyNpczt46ZSF3cZmDqksC4rKwyykTHZ5/OhE6isXHnP
cZys8fuIhVVvCNczQPTJaxvnkboDjUJf5rLA+gxQgNQ76HVwQW3WJrsVcprDoThp
Bzq1xbzwjRPzGnMg1s2WmNVQZb5xKvvMe/JccuPTY2SI8LXlXTB4ujM4AXc/duL9
NojxUMeUuLiM3NEBI4sHomxhZhHDL6rmtIWf6dsEiA2de936BbyWgwp3NTteSAoM
OaL+FvijUYn/2ayZ34t9fMdh/3Q2FadiaJFG9uXNVbpJkR0Se+I587h+oFtazlJW
Qxh8QUgtbR3N6SACjdU9A0djHCJ7PKOMOfL9uH/w3/t55WxYUdThFVvD3SKlitVH
xMDGniUm8v4BWn/y26jrPpYkeG5pydCN2zEoKnwrju+eDXQX7DuMSB+imVgOLsKR
zvtTgr17/JKMhNaPVHRiw6JQpe+xGmMr30IirnQpFEG2j83iM8ALBnLT2nbh0wRv
UtMzn4qxKHvCxmHZZOFmiY49X6EyKzOhi29CcRxQXbyf6F/sDauSGbdl66CW2yn0
Jtbtnz9liG6DA6iOXmmQbAG/xGoA0kGLgPvRjSpvoYPYsyRwCGHXjquDuNbBAKKu
0U2dGUl2hZgGaGUZV8tYbn42GYRAXwgmdFHCQq1MYA7pAXCfLmC/v6j2Byxtsrtc
WoQQuqg2qL3G60cvgibkqIptdUnp+mQvu3STYk5LsWnZq27CAo6fM+BkH2ZrNpeO
UEWeUG6/axRDOBZhJvH46jSUmOGE9bKQGbsejYUSfRKiaMVUovsEQIk7mZROnI6k
jAhjVXzhfIfBmuGvm2qEWVsjJ6dZ/UW2mcUWmAYdBCsqqvN2lFPTkenPBvZIDXbp
n1fRN8Z4dGAs1C8fL9GAZ+WIvXlWB7p5IOlykjpZW3GYMlqcMlYQWst19Nbw1JMk
rvjxqfH2GV7LeYpegGxaOV30gvVz4YuOmlebyeg6eBuS5wybfP9JH5VIdtrFN3lS
lq47yDz6bCrTvZv4XM95RYgzWSD9ReU5vp+AnDfqR36PaPUg0AzS2OFtujoqG0Au
XTkfidHZsfTt0YlPf8bvFbkKSudeyGT8JDXmDAVLsHMFSv0meRdxrg16rCUZrjI/
CLYGtw6mdL7aQRQ16aQxBen8zQbtahLqPH0Qq4EJnG3NVWc9cCnJs2BWKEFWHAPt
1JhJyF8py46ZvYAhCZEqITAKYVK+2bQzhLHprmwhqjy0JjC6BK5zGmLTsb0AZI8s
XdX0a78uK0PkQ3VQLWuiIADws+K1/GHM5jaanWWDbPWkOo5Q1yuvONZ4549+QtDF
mB1r2ffy+sTlED83Aht9qyVBmnzFNon/NKiJuU+AlCbk4g5nkJsFQivdNHBQDQ6L
Mm2QCTNzVIO90pCbv9JTS4/3UHr4FBH5DuvjUYWRkH8VrWr3iTv/O12C+RiXlvU5
mSR+NeBKJU3cCiLM0eWRy+A42X+jRkx7vuNa8cUPzsb7F5D7QZFZz3YoQgKiED1W
qKALSyNfuP2kgbaWUwaF/wLKO5pMZuFGuqA0EZWQLr5+JJmDOOrBlzIRMvl35Yc8
3et2G7E0GE5BPa4AQ1/N9MJPd3y83B8rZNaeXG/Id9r1sAGFV2HAFQ9OWLtwQpOU
LvGBS8j6b7hxKZRWSbAzFTuU1UqiybSKfXOe9c5WbEXPUVZKrgoaQCLoWRGcGyFY
KRsOsh/cRuLckD3L9tA8A5qm8aLELij7SomAbxkFG6rNYUcGK1K9VPpO6oCV53XG
FVuYez6DvKwg6PcUw04icNvUq7ZYUbFumIjQLD4e4c+PWFbx0/npbC+Fz4eju3my
JKiYRaW1fCWvDUIDC4Kb7/q0Udn0W38BQKEVFlzW/1RmAfj+CAeXcU160/oM6DQ/
Kwj4/Zz5InMJbiCfCx4u0hhUpoX2mYdunzJ4Fxy7v1QcoPtX55LVymPHCeqB8y7H
l6FhMV6qn3SKwVFQXE2l85cgzdyVZl8Rb3JDQRj49LuUHBUkXdN81JTh+WPM3XdL
mQ6oJO2M+FdzeQLMZC+dyDGUy9kcER1/cUcLR+BL5bydvGeEcvh6ZvA5a7XZqnNE
44MAHyMe2+R++P5yOELBBD4mMZcXuxLNnSi2VBBkTkrnZtUngoLUYhtZKAXdeu9X
9/5Y2ROcjG1aZQKwr/j0/2tLRkO0WkZ5ekmnU0PickFNa4YF+mTppZ1tadZWj85I
bno+nfB8VfNJbzggh6XKOfZ/0gl5SKl3FjByPp4oMf6qISWM+KR5SqXDgWxL1JsH
bdNkRZBvrPncnmrZ0HlNEYpB5EZvHmPIysBAwtT9/8uh3R+t7COZrK3if702zy1q
l7BhMouoBjaPByPairDY7yjkgt6ajZ3sqWKS6ZwGiRShpTEpEm29TDq1Sz/pXZi/
ysUSSInxu38n6E5uay7OHEVZBlQGufJoGMYya0PNv+PJMCNStej7MftrS4jcj6Kp
cXZhURZcsR6MtoyPe2/suosAXM8GgBp8PSlafaSXVODQXvPKwR1CMCP55htAJbZX
m1yPjlqBNt/HekwRxRVcr5bqPBoMbBPOSdkNeLLZ0DLHioOXqeJSce2RP7rQTNf5
9pvFByR/UsSqwAU/yTIbOMr0IZ4fqN1tfsoHPHUldNPqDR22PEd7JvieYI9nkBDm
66GyIWD+RhPfPFUgFiMk0IW3K8mpnJrw6L35ioVReXnQcyPTun9B/S3ce00PChOL
I5swO2oNzldRcgV7enlR1k8IL1KSkSEg/ZzrYg44+SCDcQQPVKX6FJBZyf1nXnHl
b3yOiRc+Ei5XVtw7UiRN/7EC0DZEN41LYD/aHqjCS8diW1R9062t0RuSV0T/7Oup
LFrjOgGbvpB1WD8bUUEdm/jq21lzbKDzXcl8BSO1W9L/8HKuggYEGD2evqYYkR2R
yLswhNIvxVSUwPEcmnnby/rHmqfbHOUrpo9mUQuOVK9rOA8cXG/2sOB76LZsEBD0
8nmiVLodgF81HzIfjVoEoVsXwhTFcV//MKLpKccgcIFzrFllmsNig9iL6xl5991Z
oErz4v4J1W/luk9u+af2yhhmJFZiQrj1FYrWi5I3icL9F+N39gkPZmLefBAtAU21
zX2HdEQfXuHEansWA8sdIm4SWiLFhAxzpkMLDLV1O3qrXwMZNk78Q0UrEbfSdEFB
9cDhef2DfiDx0t7wrZi+h1m/6aYQamagsd8BMCbrdc3Sunr/3gtgcYwcuznpg1aa
HQ89LJ0WX0/SEXomK6G3IN5yF1ozn25cEHG/bwSHR4sCr5bvqhJtNTQ86G1uV1RP
9yyDtxClv7YcLspp8p8R5d4JifaA1WQLCHhHXSkIaelWL8jOjAbGUsVUf0mTrYWU
IFHs8z15XJqLySKXHt6Rk8MRGLeLgqjVzeD29UtmM/nOvWoIDY1gwXi+lFwYAYen
sbstXJAS/jf5MG/u2PizCAH4/ICPz+F/+XLvbDsWQ2cwi/4z7U4X+XmX2wyq/FMg
3uQrDADuv1FXrqyvm4tTgLs/WqpYVe1U1OFgiTknfjs8cLm2LKHf2E4htZkAb7NN
qqdV4no/OH6+i7/1YaSGZZFEAV++97I3CauJXfWM1gNiy/CZcTsRK+GE652XL8gr
7JBO1fwik5XRUMNvfO/B9/cW9320nBXbuqy9BnJe0WVTqmz+nsHL3Z2cqbcGudbq
FDHG8DlRgNNqwGSa3/maA7teE/86v/8VShROTNFAxnsexcsiafmvWJe56Pwkn5KI
7zF1NImdG3ATrGBLR/qyI8/XinvGeHPpkCmKEkOhtO7BOJAYZpyIkfeeIsUz5sCG
iLE3k6VkKR2VwxKtp7pJlP6Vg0xiPqfqAIbRKCWokoNStLKXu3M1mpSBx9W0ddFh
u7t8obJASxH/sIMNNkMdqvbo/iUy9V7QhkKozPLlpEWx5pNoRxx/jNYt3qgKggAi
WImPy2I/rTAeQlbiwpeVP1rsmMtYlYuAiNMBcKxqr8fFOb9Olg3X/QCGNkLlOAoI
kHN+h9Gp21iTp3eHI9MNgf5At56zB47ZW8074IkfhuT5DmzUSHlIudxQ3o93Wgqk
oxjHiy/B2s83TK2MpJVH2ga25ICa7BO5OWJm5Qzeek7uUGgjoJhuX6ekN8TyCi5K
BndDVuB/pqeRKOse3jAk7vuT2kOMkRpCx4yIUn2IrtpbEwtZQNDL5NJIexUuyDSf
qt80XEi2gtvdTyFMrh5e37Kj5szJeYmw5ZqGGvIeAb7yNcravlt93+ZdSXSawxGb
gLoZ1iW/VglSNcMm/+SRV7SaIr3Du6BZA4gpX6iipRRqboEMod8+wODslkvfMqny
9oj5ZrdnWQPpfrR5S5koO1PEuaVfIX/2oA8lf5iXQIfFMUKKFW0Ej2d5HiTVYIGn
NRbi9GDS64Mtq0WatT5vLwvv3vAWOi5d5+XQj5Oq8f4erV5aU03QFg7/U3vaefsa
FO2TdDZV+T1YFg5vyU8aRUnGnD0m1G/lDcllEoXjHhqhlLx3y5azTlZ4pVxRu1Y6
HnSr/AGtu5u9pHD8OGWpWGoVBzqyfILTxX0/hEVhOKHQoYKT4bVSsdKNHU6PEcDQ
kczMdlq+pxxmPilbmFbsnHsxik75SgjJuAro4fs4m+MA7G15hsLxus0jeEwBpntc
yybCOeinGJc/V0kjBFZkLagyRDbcMGRw06lJYRhSCj912sdofUNiXPpQ7up02wPF
tV012mudCrFbjX1umTTdYTfziV1MyxSo8r8YIymv6T9OEBcWoPBxU2GXZunuUZ35
qV3yrSs5eMO/27viAbt0ElHo/fYtdEW0PhpKr/3dHjd3pYfJGNcRQBv7DaHrXmi/
/TkjR5pgkwz9JIh96QgBWp1UBR486/2l1EbsXvcjqWhx2YLpfaMd9o50aeKaCUYy
RwSUb/8lZkl4tqZlv6dNRORsFZP+kpb65gcIUkH4GjSb7yF/qJ/oAbamNKnDnFlD
LrupTJBL/D994FpFYZoJRBKkJSiCVGP9x3EDYMU3CuJDIq/3aPtSbid8H8UL0OCq
AiNR/aw6KVPhLM3b0NdGf2GORtFSXHc8NEzwpOVG+G8lg3zpCxRwXfEi6QTGt1lh
y+VnUVFdmTsyMq3s4hcsIyihPqSL4RZQhZwgjdwRK7Wqx/zem4JzQ7k0oX9j4jqp
A9BvFxud0gpdPHlYA6ajshqnrApjOgEJgKd2SuvxUUXaeCSihZUFSu4hXvutMmsu
o2/TPctMR76TiPgfEmOuQ2gqtgwywtLfPsdtBkXN1tf0Jbk6iNt0x6ZIYSszN5R/
qBc6gGbBr1Hb372CmADgXGMKCF+VRrRgEL/I0l5jENATmIusB8/VdH1OImXbVnqd
FWqhP/xFJYYJvF8HOj3mfMexz/KAuU3/TPwruy3/ak0Kcs2iXhU176MGgcTrVYaJ
RH9h1bCfJxjwstdrJ4v/04wd7Axk4cW6/0OOntyB6ne1oNWp2ex7cnVPzgrmcAex
2gX96ERrPsHTYkzU42wDaQCtZmAqlhjHkTJ5N8+/h7y8kVngQzMFpfehDUhk/9mv
sI6XchfjfE3Oz0XPyz5R3OYH50fBJ223TSi1SDwdVarzjbgzaj7jpoVruthG2yaa
teNme18rwD2bjNvZZdJUPJhQm8N9343sYrAsNemDaz0uP15hEvfYVzjD0uwMsIGR
QgISIBPJaWba3AGb1ntrqlZjy/rcMtZNWegsXGJQD39z52PRlZQ2CJFo2RucVGIc
bdCw3af89K7GR0CVG1j3svBUlhBNf5KKw+CtYsKiuNL8EacGhysM8FbuPDawsQqR
1q0en7xipJ/OgVoDgAuIxV9CCnJuQqC6td+QI2Vm0SDZgicsFL6O9JD5hEN5S29C
x6A3ydBWqacXUloRiBR0mnTygoo1H6KpaZkaFo7h7RhziAP7e0SpwbYiO1DhzKQ0
x6lwZBiXPt83x4ECc93Bktq2Rf45gcEE+A6+lsaMbrkKiLZK4R4oCW1cLKHDyUva
vrcpsxHNKUJ6P2zU2TpgSMCtEgc+IYXKSJtymKXh9nm2a76/Jo3of86YuLc7306j
eB54fbW7T2sFbZxayNVBjHBy5x9wLwqIg7koiSpOJvbgvYo4qaruPvZ4NDPV8BsK
m4qa5AQ+4YHh7vNjHpNOrttgTtjRD5eP2uS1y91DRbNhKPJKpSn05HIEEuS3pro9
qtWbFsOAaK4sZlKLGasogtQ0VJzpwGl/d/YHGx/I7743uw5iFKjJ8EZVhyc5XL+9
YfCNV1ulxTJyeTsseRgkURa45S6Z4swMq0+iwDAJEDqk134QemgSqFlMa/scVBK/
Bc9bIP2JBXLoGZLegwuIGVg5LSxb/dYgO/saqj4q1ClbDkldhF52KGVpgo9Bq21y
U3g3jCsnBJ6hPTaof7kHQ5MkbcQ69AiGaOxSicrrsMBVsHmbWRaErunRTfMuk0cd
+glFMo8VOgJf7R2vd6jkDJFfbhjLNPLfVsOZr7qrxBfxZhlKEZwZmEwg9/4cxycm
cUU2KwU+db6gejMOzqq5QJ2u/zxxKgOYKxvQrj+H2bN9YLrlgqFPVbhZGY0xPZFb
68dSNVrGBQAScQRRY+5eqfNW4cXuOGIVOVsK4FKX0Mx8C4d6f33JgALdJv/H/SgT
mSxNt4MUZD4VH23NhvOfoTsIv1YSqp7ko9IdDCE6PBIQBTt6F13+13/S1+hw2ABH
mkLOxgNQAB0BEXN7gGADfYspHoJ6F+oru5DAbVxl6aOjBsRG1/7rc1NZFkIHKg3U
RFpc2VMsBzyr3RB95cdrgecQO2qZkKurvOGenqNxWBhp0cqUo98guxLR5SPI/9+9
FDOwhVJiTdC/a7MzWwpdc4+NugF4Y8qFFtcmpp3GKl6VdlUjj5ff9nFsYgRdnFWr
ExaLELY8RT1Hy6Pra+wCFH+cYtPEOc+ffhJkpjOxsi4iVXaFQLpCbpXMwEsV0ICp
88/PDqykow/xrwIR6su+1IcB/QJrFl6ZmXwn1SVywbAha444x/7+872va4zldzt7
1BtSgIuyOTpJnHG/F+9rrr3XlSjNfrphZ/B5Jl8et+eObgThcXWv25/nYZMfzLhN
mcc2D174pXDJvp9HKX9St7VmwwYuvGafl/zM4Y8tBwyG8Mbg4r/N28x1C3vAMhZJ
fIsskCVTBpF/P0dd+HR+KoLdUWkEuIem55GdpT2GuiW0HnXbkUqTLgInC32G5iMi
AYObROzoELN8nujPTeN5OpTkdte1S/zvjnhLm9FW/JRtzVPCXf/BM9cAqAQCTh7p
UCxpU84br/EG7ywTTixaMId0x7+W9+XvW2jVV8DkwzopJIa7O9H1M82O1CiBS4ab
0U7MzrLGg/DkeK3mAXumTU8ZazO2T7QNXtio8QQZOZhTZ665TtyxhqI3B615jdRe
WS8FnBEBx1ekhmFKv3V5oxF/tD1HuMeBui1T144ozerdT+17a96AXpc+O5pNLHpi
WeGk7qa77mFwLjESJGdfm5aQGQMHnCpdiGfkykk1Z2LyGMfRXz5NkmJdeN8/rlke
xUPpb3XWurRtcC2RxTucx9BQyvIQ/pnWS4Lmtd3QcePmWIWYyqo7NgRxFaJLDHNJ
6v5tNRK3WMTdR2PwnpCq+qqVmzlT/TBwsJ2cZ1jEsoXMFDTdkcjlEZPzkCs27WLr
B7yTvrsVW5LEV2hj5rwE+VyC84uSY0ym4PTK0txOf/0sV1JrdG3dMvzCSa5leOYV
+NL3CncATxQu92n1VNE/I/buEmiRrrV3d8FjLSeiZCkbcQoKCGbBE+mhpJL5g47t
S13yWoAyw/IuUv+ZIsTqiW4ARj7VZImUlKPO9V0r7bJjXRFDQN9uAXmoYJFKvBYb
prhjUvigi5v+AiKgMSf3L44Z2eJ7TdiQnpHSqp4dHZM9aZT+f4FavB8duNNlmkVK
kSZryK7zOniEHkswPjMgr7AaiiRwL+kLgG9wmSfzaUzchYlkv/p975tS3t+Uuqj7
INRZjbQnlxdGbdUF6xrqEyAUpS8TjvohJlEbSfT0k1d4WUd0JEWmnshbcO1Xpica
D0OqLK6KMrhDmMuJf0lfSvSflvizL8b4prMqIWHqNX1GOxS0ccAXhtwQh56txVzE
1ZLqrOXzKIi1JVlGWBHHEoLoD+MInOL/NulH7xafHzqxyd7CWaligodFfxjP8dxN
CMXCwgUSvDBxNfoM/y0WPte9AAMMK5bG2PYE+vDDeEoJ5ysdWGSCkS4ylM/yl/9M
FOs47f0uUUf448sDc32TN7HegNzfUpiaoYSDBvNfRuqV+k4e1/G5kjswnTdbvjju
9t54H5gdlcxvPMAm1Lf5TdUI19DgpVdIi/MzusD1oFxRDVPpabLaS+tyK/BBoAsS
I2I2wIl4LQnL0Uwr3nXeuCPPeUZTE4Xo434+PI5zJfBthlIBAGtoOshQEWh95M/Q
76Wa/s4rYg4Rj1fPygEm4p1IrE/hr9w2abl29pLut3koMe4Z71PCpPoGzv1RusVi
TswIgRPZYv+fa/g/PJ2U14BcUsn/SRlZ8qXblrYtoz5y0TRNMKVkNtHloXs0DyeO
ZQ+4TCNL394lSJl3199p8dGlnFx8WQCmRzdABJKZBoozbvaX1dLsPmfxs5ITf1WC
xK7EeMTGiD1SvBWX8BdUlO7kMfXdV+c0i3im42ZMY46e2ObQMj1glo2HaPjqpnMS
5NU7tgdq8u7VZuxpT+d/aDLRj8RLlEpGcZINGuUxhEaVCUJXUo9on6c3SuFd1+Kl
ov7UsWba88IdKqAPuv4rPW+wh3iMvfW5kL54LI0te03l1l/NhuOgYdGDKzhoYw0f
uqHtgE5//n9s+L18+LtAaSHLfqAulGfA7PyDzXCt6ff6KAoFxEbS37tSbqKFNKjO
WMgqiFoR7ZTlag1svpEV68GRlz96nnl2CKEAvxwDh2d6sVpXh/CYZjFXIRZ56cCe
PLh2F3QvbFDJGNnjlM3wdu++j87KEy/5/4iFmbjfvgaxA8wAs9nAeUtLo7WSFOU6
nTWKe4b3sDeoYYFj8ZGVihR2sgB5Smk/nmSBuydv0w9JQTo89hOa4x3YtswF/0+n
MMltxibeg2kD9gWvUcRkWfSP6z6C+SWFjXfDetmWGh+elB0cDDeJT0RnZWpuTFkT
Ozyb5UQt5VCP8WKrUpBdP6NfPSmaLDYIBD/ayx8OvSRzhuAva32f4ck1tsXyfCfQ
hcIAV5TtV/gHWxrFJeK/JYX4Z2wyX5MS7F4BZ4IZQdjyJhaRofXnThHzKxmBpaAe
0y/pcqGWnkDX3NRfFWwnQEFkw5/7bkytSIaoHaS5D2kTH361Ro/IucaVD2yc0S/Q
oSdwXoX4b+pY+DsAoaRqkVJnh+cMtc0hoZIhsXzqhK4v/IRXNdsESfjiKoPzXXuB
CKz6X5afmr2wx8o+gleAb48/eAZPkrTaRaMai4fodCVO+dtjp4nJxwCLizQg4iCK
YDN7MOgF8JY6iDTcFSu5QaUe4rgx9SjcOEWxGwDPIMIXnMz1acL87jSctoqgJW6y
A1IbJ+QKfbkAqW587LIHqhFwYcqQdkHzkIYluMnoYLRroxwkIgZRwTSIzvj5vSv4
WdWIi7Mgp/3GkS/0hDtUkTbPtUuKyuh1xqGBwytwOahu3izB6vfPqIfgeKVkBZ1b
TCta+ZT2idYmHSwkWwx5fYRFKP8BuiPcUMhmVBAgd45SMMOqAh0oE4AAqFQjJwHn
JAEgtP99iKW/O+Youg1F5HDd18aGy844rpoE4uamgF5mVczGzs+6ybFBhCLV7+rx
UzatHisuu3CEFwHyVD/2d0QcOx7yTfZUoNzfAk1tAL+sW3Gt1UU5hGk6OZuu6mTA
sw602KTuW5YzzBj9jUCVrA8cajIqGZmLoAsPSOsXJNjHWGgtVRSQEbgrQaYtXVMy
smo2rKf+AXy/ycBzO684Fh002oX76zJ4AXcfQR0soC4SpHCvhPcNKd8Ri22K2HwO
M+WF7pQux6ziYynIn2jW3vbfd1JqD/U5SSZZygmEMenE4yvA/SiLU06xJ4lyMAwu
dnqam0fdCU0yzVKXwwdwq9niIE/xzWyEfHA/TjSgmq7FMVYLbfFjAoAaY3KLGw1K
+vdfocsXJySIvyVdNUOIvNXEZwLK7qC1FCH7yTBKxx3vSRDJ4C0gFI+9pgtYPZw2
bjzDu2kAq5Q8ZtQqh+VDpkQlzc1Zu8eSB7lMV2gQAy+Gj/VAZhx8JskFbP/qKv8k
bu4b7pycn3jk9Ar7Ly/clkzs3pcfCzCF3WGX6SZPVifV9zOkIeRP2ply8rxSFggy
yU8qQ/39fg8ictdZ0nZXDy+6LM34LCeh3k9aeQx14vFbaOwXFaGWHE5vCQd+jUgp
NbVLvlvgxOZh+ZjZE4C7DmrMIyA0myYCI+M3GxZthkO4dSE4j0u/SDfSKDSYUyan
Sg8ucdY8pS1fjGaiZOmFRVbXYEBAhytbLnuYDaw6izqgZ3JSOStyNn05HspoUmt2
xgcNLjNVXVl4A8Rj93ZSGMRn4hse6l/t1E+7rYmorUp6LPpoWkBp9SQoA4E+5bZi
60S2/N57e4SpmnQT42KU5wgmLV6jTis4xieeqDD7T4vCyaT3jSsP7o0lSpf3xRBO
pOPp2+WUa1rHYQq74HeVLSePXlLwAmQI29LbciEqSU6leLTURVH9AzhwAvA8ZzSf
C3U9zXufAWWjSDo90p6yKWn+2uRmwFnkFnol2g+nbuhuAWikVDRErGksjIQS2d8a
g3wZDAHnbg0RajVM0ALbhV9dcPgMs+kUWRarkKoORloVwxJ0OO87j1BJoskeGioZ
eIz5GZESiNUphJNDbYj4+gY9CcN31yhyf6duQlOfqKPY8M1RDc6Td/wfDM8VM4x8
3sKHJsFcDDMTWPl4cNeTF5TnajteUEJ798Mo+Wa19Uuqc1P5TZQR8cvAsD3ikEGP
WXXANXiszRDHwyPswI7Lp931iMTCsS2WuQqCCt8lKLl6y3UFerPlORm99Mz9NChS
ZA3d2JrPszRYFBtnp/UW5LAPGOCpWJKKYAZnuIMDO37V8DiR022LbR+xk4DtSiaY
5duejI/vhwv2R5pJOjwVtuhiguxE0x/InjA0MuPnzBrBAPPeq89wd/R7tMK5GwKX
zH6A/M6iLXyTeYg/3uOyJj5Umh3EhxR1z14+0TBxP4ty1LBTmZItrWxbSDNSGspC
E/ONIXYsrDDKhxD7h8jOfskyH0u/5TVOq3slW9C2M4XU+R5Ju5uTbQ1ndZY+fQHf
Z5lLp58/vJBEv8RNkzRn3pxEsD9Nd7j3xtntCTKK0FBfs+UDy5WgkCRzq6QEcfwh
KUdgT2KAK4AI/oGD+BogXxyC83wR+9hEDoPByfchWfIcteF1NNRvcB9zwPEjpIAj
PWhIRhQChKmaK0MQ2FXy3hVLTiuqb4we3URL8f5kDrSdueHdEqex5iGq7QV+yZr+
6Q20mYPyN1/0ir5vyOeb7NafyYYDq7hwBwCn9/PjoT7xgY5/g0B5PD93aOV8J+pf
fBQPFR2K8lXNxlpm1imDXOu5DJkWH9Dvx4qKsG/2GbNKlMTw/OpDBV5SuP242vRP
8rn8eucxasyKueOtHCSiJsXH1N1CQ5tkM58ELEeo5rJt7dDjCGuL8zWMvx7nKC2t
psPYs+MaV9aI5Mjfbq7qVEqUPshrLevY1B8/vAhSHUcqOtDNi/zA+I2SWW18Sdux
5T2Y+Z5M/QjBaCNpyYocWrkZvUK9v5M4w2sfnjvbp/RWVdntd9lZA1y6EXs0b5T9
XAa2sA6HRGq5zYmeN7f8bQLMQTwaizzpZLzOmPJOgYYXGq50xW1Uctg6t3nVcNgx
3oTeX2ti0Cy4PAXMB31tnOE/x5Uc6AdLJH89NHu6nf8GhuVsGmmR5gj0sddCiJOa
c4gcmnn+2mWqb39LdJqXfGQuGSblKQEjuNn6iFVUklkFO02b7OrBO74PfLnRE/Yr
2T+Ecnusfx5KWH/n1rNdvk8bQWTkroITN2WsSdnPcjJ/jmbtmjVxMXXPKvpe6wJ4
daIopMoD8O5oPDww18DZ5hc/4mWTk00nHbXUhv0vOF4vhP/O9Txb1ZPTA4ieOu+B
IsUhJigIUPT18lsbrZZhF8AjaWNhiA2K/ctTdU44RSxVOLMf+098MODMeNLHm6td
EFG+vj2ktzoxyIbvRdVVhHOsD6DinDazjRV7FoMy8gLGOlwbNWjbr1pDVnWAf3dK
p8nGi4/VBXn60YxqqrZJv2N6fA+X7zDlaKQm/C4NVKYfoModavZjwrzmLMNZLqKG
9HirCId+Oz9DBIt1AotH2gJkM22PbIMtKfmAoT9cu6lzIZdRETrLe/PNHVb4T93D
LLoxZ4M/ZYn+Qx9/pl/7BcfdqXJCrYdAzA7AZLa3eI/QFwWI6Ta3S+uNncuEzQvk
rlHEMLftkQFjlFI/LJ+1rurZG3irHOOZCVqKRjFAkx8L3Emy6/SKJpfX5YPAk5/p
1BDApoEBN8PtPUyYfPaLcRm5d50r+PoXE5U7+svaLJoNWV67SpTKmtiqF40xHygX
aym7DGmC4+nX4+fskyL93kzlMi1FlDOBnRNNYRW3uMd/wT/dZK8dgsm+GmMXO8NT
KjOZvQ0/VPGN5gsAl8BSE5p0ySPcLqDpbjaIbGhbK8hO506s6lQDorkOYuJ0MsJZ
L8PECNEiIBqYUnOunN0bCy6dptOyGDZfwrPj1wUzz7pJS/htBhx7iSurGSYG+g0o
ojc0OnrvvviC3hMeEicWU3TBeOCJI1yzkJIQyeb1NXET00TT9PWMNPkLRCDPHFlP
vLOuxpAGJPrQBYX86r7BqbXsSzkcm8wsTUI4fihZMnN+OP/pIjjAMP00Gw7K3b7s
2rjK51/D+w3nxE2fjC/JV57ypBSlTR5xf+aRzrTUmcq3rdwLEOk1wDH4JrEedi/N
ZAHbpYaWisaVDI/tKVEpY7tR2HH2pw2M8X3ROoler/u6SZyG+39cMOu6lTQ9zCVK
ZqTujhK5OC1dtObPlkzy5pPFAu7RrOfh9oOWTvMnjl19ewtPpH760Rvqa98o5/5B
o8KwUX16KtoNJgS7REp9n0haCeiY4JpBfpctW+0/PXLqu6CVrPUxhK9/DY14lXJb
+CJJtH48N6HAewt7nCMsnPwQP1jR04F8tQdrtkL3XXTF0ZFneNwrgVkgPxmyjTbj
hkZTdAJG3E8CC8gI3ljvsBtZR0Scvq9haVKF7+aUP8jzlf5mc6MQhGNpmIyZDxbg
Pd+uPbvdw88B/vKA61wucLORzEXpATbKHfpTssK//sAJ9o2J5UddXb2KpLdVlANQ
qW+czvrZc7FNoWzIi3KFtcbBWxX6upBtIEYyP3nbaWvREjHU8Z6mwXpNUgK8686E
WO9PnGnbDuVjw/Ioib0Rl37OaVpbQaznbDsa+x9OCOnAGES7puQmpS34p6XJbmXy
e6Irb+MF3vEf7D0W+WkijGN9IjU/+qyx8iCYQh8bJdXSyiw9ahPyrokxnoDDC8uU
IAutQ67EFrSj55MvgHpBG+ulsMYztJf+Updn7Kw9bJzlxtMODrmqsQp90OL9aEeY
it0IXn/QuJZuYUn0NG1JORhQ8rjbJsS28m91mIU2aGVeCHw66cw+xu8NNza21hxp
0CBCxX0ife1qC/kn4dSMxgaeuyea4JC2f8YKdL7G1dRX3NYO1KTLhpHMlDnDY4RL
IkmqV3+DE2VyYNiAY8KpsakEP9rm1+XPVs8tQ0w0DIk9dlyGzmexvJ7plhN/72jY
ASBGfYP5TiYae2CwL7qzrGx8WpTCH03mKhJ5HEArOGes5lZHxx5NU5Q4EYG/FjYN
0kgf7iZBH2wsMYSKsA+FO1Au/Xs+gVLdH046xKBvy7/wzbvr9lbFEEGiWklq96nB
mlzFCE3OWPZtSegZYxOwcjpVJ/l3F1bBWdkloMIBvEfkzIjubWs13V+7DBVdXwyW
TA/mcTEmNyNBCIIxwmOX/klBgRVs1i7QzEFktOZG3USXfqGVVuVWbP+sU293shJG
OlW7wyRn6K23C5nFykAp3OvbYBxGXRz58IFMtFefnQISiIjA0WbnWdX5Tifw3rn7
+/MeVPKT+bvTCfPVdjC37Fu8NsMgvhQ4ORfbRlUGRfStItX+HZuWUZdYa4Vf9dlu
SiSpJEaCKC9bFIUfPkPAwTgA3hZqGeKB1WI9SzQWLSA92yhFbiN6py+oCunK8/P4
dqsWz6XfxFfN6TWM94sWjDnsC6LfuIvY8XNFn2Z5bCY2fOzjG1/DtMvBKdEees9B
bJeCkNXdaKcA2O9Vf7S12iN+p5V2kdj39AR7B4qWtxNXPtxg1Z7AnCTNL5qrWdBV
fW/3RZTRUPzYfnOr+oGDkvgg2ZmJfQ5BA6PH/fAGCPalbU+Crs9PGt98/oPBqBkv
HbxVtURh0o+xHr81voMD++z/zAVBgdxSyq6yHeCUVPHv4e5NqfF8oJgZXaU6T8O4
qZgYWAtVoJPy7GZdBceL9+oZ0cw1wlwHyuu74ccW2ISbFAnG8KQhBejG2sWVoxAF
+H0aab+9efeL7+r0n+brJpfVWZRVe5VIBSL58QlYBVMpY0zDmOZM1+YgvgaedIHZ
62oJrd1AeMlWXGdmaaJuFVJnff+mCKv21t/YTYbHQ3Xm+GSY7W6I8IM4pQh7mgKI
3X5CHrNLGg0mAv0rOkfsR9GoHU2t4WuKb2W4JAx5y/HKHfm4K0KRF01wWGjzIfvR
Zl1cD8p+MLbk01Tcy6tPzM9tHXHjllWcNbaPqiqXKX3qtKDqtLxtH+gI1hc4pgL0
aaJ6qB5NpCaX36fAUVplZG0hc4GdTnrpfPq1MA35Cy6Bf7cfwpoh4wpSAVC1cmmw
DLdNUrlhAmErZx8tCumvUwRKUIIbLckx1v/QeAkRs5Z8QnSx+z3InT/Y5WSlKzAa
3Br8XP8TWurOPd08gOq+7mY6kRY+TmoCoVUOa1Anelvh6XwSihCuFpK7hqWG49pd
klaZqPqr5NduwPrqRN3w5KRkBC45izzqwbL+sXhAcvRqvN7ohWwCVGiF92EX7L1I
aW/G9PJC/3Z3aO0b7QP/SiR+IGlGsxAjcbqtMYC91KO76RKrT8VLArAwNDueQCIs
JgABTglL+wku4T9jmncLymzSJy5kFFNg/ZBVS/zlDYfc8Kv1orb6A6ytpj1chwLt
NlQ580KrNbKVMzHXjUrwE9fnXU4GkzhsDFuaeJuX47ITEJNfRo+gMxu3DMazfvT6
QiparqW5a+sPxoT2xcw7oix+1yEau4mzucdzwq1S7k57fVK/R3qilAO7Nxa96zjk
AOVaG7V+BZt8knUi3kyOOSmGXDVgeoz+oSGxf7FJyW3ygJxnmtzd0fvIjsgd/xU6
D7q1jwNKc2AYYF++NIK5xaineO0/DkdsT/XI54WyMEoFg+noUBoxc8GzUIr1XBN8
8QDk+DzOUHDNiK+ht7hlu7Ei/bGlBg3HNWmXi7d3oBePp3FFC2oC9ekINj9chBiD
HqFc7mtoBUPB+glrkbHZ9+3ONKz5e3DQbQP80NdSUAYNwsrEoRbAMo6pXSw320P+
wTi9k3djBGXOT2brrXx3LyQ/Lp0ETJWhkK5tXfipKAWO+ZQ/w4qrCVdr3wV08eOM
MGZy7Czkz8PjHBQuvc9mJDchN/EWymhwGw4BctSCMreLv6GJfus00+SZL9bHmhEg
221di2j2uOC+A4EfMQvjE0Zj1cm+WtZgJjq04cbAO0ZSp7jqnOTlJHUqFtcD9BHz
LTyXT3MtDjiFmK9o5/4DlNHUTumYUttdRjVV8nYYuBlgOix38ithVyxXZG/4oW18
0ZkqD7FUwltslAy8how9sajBjqzwbNlGd1dHFooFd3UCvrQf4gFIK9wCR1H1Z4+v
ZTAuDljqVxrlrIZNqbaZuwMOSg7jePx5fUJ1Xwamazbla91p/zw3Qg/mCjnlvneV
7ugxUZ2ADFulZLy/lzSciuRJpRXACPhHteUfT9HyXK9+ia5K4CcRxYnFIEd3mBeZ
cYIg5vSmGWvKFHzpJZ6v7DHiRDMPTgwfN5p6Qhmb0e/jWZvGeH1bMwYjFVrrdmq2
UgQ51CvGlX0+zlCyCdJguGKjq4irUAFAVwesbpwVIyyBdxGMCtpnpBL7fKY0AzC8
/cqcV7eap+SVpH3ixvXXq9RHdREII/E4NF31iQynPQmmcVgB35WrVG6VlB63R6F3
yDPtvKTwquarv7nWeNYERX9btmpD7RuNOOCmfC5po1uK7TOl4Ho8wbmv5o4KK2nt
dj6TZqvU9Dp5GLf/dHS0Dw7MSQgqzawhGDveObBwBVNfouRsgevyLnZuruJxhEn8
s2qnIUKFh9tYqqtGGShYd7Mz3Z/C0cDkRaE71ZLez+rdEHVQHR8cXg5Jqs862JZW
waXv5pt4AxAjU3R5+OQMgn5cn4SmEsTFUwCNA6dDzV5QYcSq9C/bLZ2XKsUCEK+H
7CjioJ4dZj5+ulEnW6mbatnzC3t2dK5I6zRc8PcaDB5PoOL5xCFxhOQaxqYXdBtR
atnIyqQJ8qtWShQ5g3w9rys+uPqAdZExKLEQBPHUksiAcqGU/JD02fWYiEoZxezG
TwrG8xb+61Sb85eJBO8WP8A1OFCVmCqJ6NpTvXctn8d0O6G3+KeqstE+IJAwDiT7
TEiSicNn/WMYcVpeU2wUy4noYoK9V9YiCxxzsEgjvOBoW9eXaQwbYfQMhmic8RyJ
StwGcmGSvVXgB6+YlYCtojBpk4RLO/1Kgenkj4lhwJ3YmJONOXny+/mOb7qtibKg
/RKhiE7MPkkdRqFQHE7t523BFrpiv4cbXHKIMjQ+3aQoW7q8u29jeieZuG4UYGY8
bV4D6wysA2D/eB681LT4md+0Q5YjllS3nxD2r+EX13SdBzctdnchM17fjBkTd9ig
0XFlp130lWDxOK4LtVDVQIn8WoAUAm5eoORzHhGJVTTas5ud9SZKRoMWGRBJRrpI
JszhIK9sm+kmOZDJvAMr0/6WrkZrap6OAAmck2a07iiStHal9VL6xS4azcYCuwMf
JJjRY9M+uFRxeLjgl6wieumszJ9qThFl6oAH2NVFB8fwCejsFggJiLMTqJxoyetB
vsrykLN8M0OBhyOGpxp9CMjsQzOGU0oicDPxS7tch8mEZIptTfVCLWCO1TAUJiJX
9HPV3tTrhtPh15nUnrnEYCPsu8X9P/oPgXCyN3r4euPJ25GGxkJuzTyDvgnVXFLu
yFy8z9E8IMHGPukUza8Sb4AeF8vM11kNNsIs0ON5ZitCdtpfWcQg6C+KbN0SGSHR
G0wGb/OcY//LUyRB+wu/OGtzQu55O8k4iLZoDe4RkqgelQmqO+mO5uoo83t53XuB
lBj5nVks3cczLhzWqRj7snwiAOU1TeKKrlo4ZgMaRikHsFAly7Hm2vRl10lyQv6V
kZcMn3kKgs2fADuCauWYJVUuqFBPrfh7yAR4w5IyUg+yZV1HoJwzS5bxcfgmTo+N
cJaJIMq6BcWlXcUWM57ws06DlyuKrd6jCFhWFlvh52xPDBFtrcqkR+S5A+WyVt61
GommV+8ERbBDMd1dGjTLMMkFOWFTXt26+T5R2ZHDvv+QgCbUCtPxugE7vwaWGCwL
5ezqh2JfRQO39SnEdEZH2ZRJnPoLGClc5An694kOH4KOt/vYdNTf1TiZCSR17hmT
+KDpQVf1ublSfZvEk+QhK3pFfCE7+S9bLjseuNfHy6+jGVwLkdkvdbMrJM8P6exd
98a0GvR75hot+pOiCwDkwCNMYSFBLFjuLbu+yG+pXN36q4TnJXIl96fuKsFLewy2
K5xHRFeWt0DQ9ZjOGHyRWGH2h9A0rhpdwjhq4Ax+Vq8lW/Wr6z0bnsalnbIau6G7
4lw0FLveY8XKMJWdGx46P/lSJ1ak8TRykxC+TS9knYNL9HV94fPyxEh+PaaDuzfB
76ejJOPZ9GuWfyRwTJyPYjQbpbAxgB9t7DnIvVlLMpin4RSWWSY/h0zbuM1Kk9P+
Cx3TvwLCcbHD7fU5THbue0x4l8/GPOwqrfW76DxrTC3HYFoaLoa+K0DoLwFRosCc
c52lrk3mRqtgmzwPnm4jqERtlW4Hc7Z6eBsPzpP5lDP9EtRm4xHeQnsR6D2G1wYG
t932uaOqIihnOvkUjyZkO15H/KZdQFXtyrrph33CD5vaXCPgvoQl7qkzdEQiwOAP
P3i/HIxYGixy0JGBpnX4jmN+tjY8oZNqmvo2tO5oXQtvNIlqzxdJHbV8m23YYu0g
bDWc9Zv2ApIWZ/+6OrgN6uBl8GiWAkMSJsgb2Suqh+6Z3o/hjZDUuS8HTIZv0coY
GjVU1nWIig0fl9XGMo8agMIFCaTcsrS642FVdNFmseweTpeaz4kuQy/18VbRJBu1
Wu+TFK1NokLxPdCJfwiVCBQWc7C86/LYLb1YHZhHfAY+z5XUoXhz2jrG3Qh2bvcM
QaLRjK+LoWl1idW61pRCwMGyLMy56ZjJHFBK+rEJ/p5aYU5Y0Soog4HedR7Lz+5M
WND0/eISqN5koV5W51KoSPzZhx4D6cxo3VLN36y6aIbcZH4N3V+bR4O2hUo0Q3Ga
eHhzBWiuzJg8FMMayxS6MrelCIq1J9CZzB30fPo3RHWNOobvKbJWhGzS39HTvock
clDvK3dyOvvojwO6TFDzXbUyTenMcH8Hkql4i7qmiWpHbPCZp1tS8wOOUUl/LLIb
JfUnbF9mcvZCwPo+hJT3mQF7Rv+aZeKPzvtki7VSoS+jsVNU2WUwwYiTEKLsYJEo
VxMHVrVSl5/w3MCfHL9KKyWlP65RmZjwSnk74Uwlza8ZmEEgsuyOe69cAYXTOrkB
lsqBQ0v15T0mEhiPUHNfmjZNwB2rdWVH1nU/0rUTPeaaYPQ/uAlDw4SsVW0Q+cp5
AcaHVIyzDd+7ckabW3AdVG+zA4AUCixIPfImaKeGdh84q0bdOiYVWqccSadoffUw
YHvIw02KT9vXLJsWnutJFpReQPOQuXgx/0Glm6g08UtI9l3PGgCEwlXV96tI9XUq
jyujjLpZxDnJm/QTi9sm+JHxQ6T1nY90StcKZeXsC65JqIV0jW+KMKRdYV4aNDj4
BmxUJejwRd/aoFITVbFPnwAfMcfW1rHXN7E9z/oshDaJnwPooVwl80zaq06S0YAH
WQDmwyEDZ70sg52kzkgUZPivAjG12+sqwvwKQvAWfPTumsB6Ldu2neDTzgyzo6VZ
pnxwxhGtJFCT6yCk3dg8fHtZQ9gsOjR7KrjN8Q3HG5otbAI4p5uOfOGH1EPX2Dq8
ZLXqtClclqQx1tASuePJt3pJU36AGJ4ZceZj3QalrUK87WUIPdhKFhA6Fshe/+K9
5qjwUgne1eNsp+VUBcHEHAdVJs4JXPNgFXiWFRIy1ilyN1gRd76/s4tV4W3dDDXN
1B9lzgdsuDu0wLJvsarMbPIejD94SRHB+disDwMAry3SaBPKIfWrVCjdq7HOcAcn
siS6tkI92xRywRyd3PZMMMB29lih5QZlkWcQ8qYHY45evryEeCx8FD7kqf199BIQ
g6u4LUcKV/0MhhBPd8KvYZIvECNZbT9z4rU3x8g2I5pwcA1KwDHM8BJ3FDY8Lq+F
E6WrbKlvHcmtSximhdSgvTzZtqp8UVvlW8CdtePibt+V+P6OVO8PwCpK1Ly0DxKQ
zzxzc5NRNzM1vZDRRMLXapeK+k8Q8Mz1tKh3qixD9mBS4tXQHUl97XcJydvH1rMr
bEZiY/uk9MkAyCpg+S8sROtwHDCXw5onsv14r24xl2Lk8LzOEDJrw1g/Wsk+Uo2W
UI5fBMemHQ5KIiWu7j0z/ORVRLeU1gAX3uSnsKwnbsPqoXTAFRPPXTEN86C2WpP4
ghAnr5eRf6/CdUmTebjuT2pVYbWb8ZZtcBjBOYqVDmARQ3n0koJd487W5w1fXDHH
9dpka79lg9Ff1L7Y6XK+zHqfT3hQhmN3cBUfq18b/PNVz2kPin00FMkFUd2Z/Ub+
wB5VQJG/LLT05UbwZUif6DR4GZt2N5PG5Jor/VFIw4OCwil5NUA4FSIAdLTZTQZB
fcGhJq6bfKiPwOab2mMbuwC8By7eygJgwq7Q+cEFWBbgaC0afmwIzJ1qyBJY92DG
OPK37HU0cyitDKu1ILmEJw7N9329+r2+C2uFF3BJnQ4upnNQb2bLwRGmDt6OtWKZ
AWZWNGS2A/3VfU8CaskqPkBxquDlfm2d5BRbj75EaYby/RGMelJ4Lpery1hyF6d7
pzG3eg0GohLgGiGXMrxGTHUD0SFPKu9b7nSUaaLEhswqNXYNy6xQ3E4HvORvG9HA
L/DQn/EVpU1RGRXWXVDAmCqFSWaxlTM9+dN8qjz7MHfV2gpovPmEO+FrY3qWOi/0
KMe58s7YChkUZDuPMNkoVC+9hNrwOZnwYykY9omsP/w6ic95rRoCSte6JQTh0qoj
m5dXICYEA6tO+lsgJBqFBYv7kSq+90Avwute6wuQmC9zN2ZGasAvLQqTNLKjXYe1
g3hTWY2RQs1u6T4MAvvPI4umHI3z+W8tUOBnppCjFLx8hnOYcQ/hdwupyXFKf7E8
/eyHlqcJD2oueB9LpMON0LSS/b/I30BKL2Xv3iHcZjXyabHZa2uBmmAtjWuINidZ
zT/zsB/2+nS/0nf+WfzcB/EjC3Bh6pBsvCkD5h9pFBPkVrglLUNCDwzMu4zOGqS5
rdtE9cttSNKBNdxYHHDvdzgesvBlfj2YXZF4UjjWGn+wQIbn3PWtDsxS24qqr37x
wTiWfK0/gQ/CfMYPJcEyef5KZm8kNC9//yGxwK5f8A+lKOCpLRBiYANRCRoxLyXw
lSJg/DhSbkbWpyxRoCsSG7+uGju2jqwrAy625TfYXQCB1w1z40aVdY8ngzcoBpxZ
733GtofwJK7Qn/DhkwAOBnjedC4aX6au9897dp2+s39yPPWjy6sMS48rDQ47vGvl
eTUgkJO82G3xULpV5Dmn6e4spwUNG6IbemPvkuxQhzChOd0N6GCDzw/AIgHF8gxP
tqpdOv2DGcET9Gbce/A0fLoNS6pD9FvDh4ehrcsusS0J2ZSe358jr0TZhmELI6//
x2I6wE8Yfpf9Ii2kS9NiPJZIydQL0WgnwENvNZtoqa90nJrlO5TlRrAq0BiVEp5+
2Nn/RDn1JXYtoKMQFLlb/kldxEpgBreFXYKaPV1lu6AobXOsJZ8hUoxBDvNB/n50
lZXhzoEzmhnWYEzsTIE93yg5iWTZtRaRKdjoFzmGf8Bp06BlOs5ADGt35aY+pAFo
th/ZS+3Gm9ZT6T/n8Il/KiUn9Gr5RgKSLGifaS3sSuUNduLL0FVy9jXDZV+2F9i+
tTWG08twA5j4aYYkxruutI2CB4Lz5DALod/keFsLFAw4xuIXnLvHa8k8baW/RYSA
6CT5VyJGA3duy0/+BDPlv9HIsMiXDvWYJ0cTX5KTyI8mk4aGUwwzg8KIJvnIjf1z
ClF8jRcyjI+1RLLVlDagEnMXNqJYvqn+nGWjhAD5XznYTroTG2CC7fb6kT8AMtPQ
aDg13hPqQdL/JEbIx/SxP//Y4GuYj9qK5cqOOqycFdQO62ebavbcsCrKETsAjPZV
Rpw4ljgIn7OkwXZkWgAhcBAMvT2FSqMtgrDGYmDqhhUrMJWg4vR0F/ETwv6zqlFC
xb4VzL8+ARszRYLceDjfHkgku1dVQnQrGlYBXhx6NhipA3ODbV4CXCF/bEM0DdBb
sgxvh51IPASUDtfNnoAKzK8MCFKWFD/LEzbnCbzOqFkMNqWuKCMo7WaV0STnoAAE
0MG7nsk9PZFWQzDxn+CZ0AZ86paSW+3M1l32e+S5Jz5772lQ7ZSIpKtHtr1ix8co
hygGahBX3ykwoe3zDyKGIm1Izr/3kkt2cvbavYi0FNy2Jtq7Fj7zW3xOSSL3Q5To
fIQx4ktg/4ZE6YlZjrzBmVOVtrk8W8HRNWgDTsPovPQdezpT7qbzFNi5DaNsroTO
w8rHNcHlthATASAm2FIKywypMqOKdE4HBytsKgFq8cpKUfXfXjXF56ceCe5rbN3Z
uYk97F6FruWjOLLMc73Y+5KezociihYLjeEuG5HQVNWBtn3PLARkgyutsCGH/LnH
hcr5fDjSRg+hzT6PQhDTS6DO98UNvjkOoLY53697fkMW3Y5vSNiKGdlH3AtBQ9yL
sxTgZ6KB7/gXCwJP8W1fLV1UZxXeVVg+kY4uy7wDWINURrO+QHVAGEM6d8tCtHO2
rzQB17RXCpGxWVqRI4w5Bcx7mijp6vDYSRhBsdg9g1lyD4jzGaiVs6X82yArIqrp
6j4Zus9MmL3QcyUbbR/bZh1JAJs1GntAUp2qPBwfpn6l7M12s/OfdP95YN648R+h
uA+5NhPdkWCrywOA737szRGVWgkF/hcIp/SAmzSgjXQ+21vL7a8GxGMqnXHh8RKU
Oamb3PUPvm4cV97ygyYSwWWtEXWLLew8n0KlHdx0XjY=
`protect end_protected