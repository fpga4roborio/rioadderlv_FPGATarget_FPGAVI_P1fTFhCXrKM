`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
ddtXksX2+yylW5zu6QL2Lhnb2d1sD00763mmSITNX595NcHTEkwn0zB1Dry37fOW
FufOhVzEJp80NC5qZ/+F0Vk7Ik02dIR0elf3clrjeJRK85K4e3Hoo4xn7YbFUIms
l/8VZSb14+JVGURjfswrIyCUotIzlzVYZ6gzoZwDXIi5gQIBf/gI+KxNXPaKV+PQ
Ufys/12rjO6aI/pPlqSm0hCvftmBcnezN2hk1UeXgOIuKZnogjOsf0iJVX2aOOWE
6pD/psybjbnsNB6kH5uFTA5frkzIzkzl5d9+YDm9OyC+k84E83I/7/j+rk4L2dah
QJOvksSIzN867/4Qt8qYTQ==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="MvBXkzurAa5VTw+1JJ70nePUfoQXBvZOku/SMmg4TwQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
oRtzZL4VJ4iwysPsC8SXYCzXS8Fw2gtZTOskLcDV+1B9Nzn1zTyNtlo6lNICRmmK
ZRVu2BmCc2G+fmzynYlNTnSa7C0Cuel6FYpxCBlOuk3OF2tzAmLAuDyOH3Z1Yjzk
a0aHuoCdIRKv7BrZCdALt03JeUmXKPdOmIlkVGFl8yw=
`protect rights_digest_method = "sha256"
`protect end_toolblock="Jn9CQpRhJt4rnzZPRk+dOpzAubz7omckX1MrFd4p81o="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 9824 )
`protect data_block
gD6l00tciPUa6pDNTk/+tzLxvdHE2s3DQL3/JqqujQBC/Ei+vcAB8wM3doqg5vTg
mdfn9XB1bLOis2CVSfu295W2DNwHfMSTc/8BhCDRnTlLIX0UCJs9Za0+LoM0rMrV
T7EjVWppbP+Em6PkVKCwlmIQ7JKaifJ+Y+kjw9HCGboYo5074hY+K/CBbfsBQY86
AyoN0MKhsIx+eViNgnWjA1/Mz4yWLcxRJz8yyt3iik6/zz9TcvWJRm4oNO2t8hU8
j7dfof0kYAUGIuD1eEPQRp7s4z6fTcYxpfX0qfRMB6ZaBpPlUJbJySB+FtYGsNjr
AhHPegCoMoBKzQRgtGFcoGbMreJigEGuLSLah7iN+jDEEfZNeiKQ52L8jJ3nK8z5
t+hNPHzaKjmAJppqGN71E4l7GJINKxHY+5YLVuwcZrwXvkvdT5qAFCq43ayCXZUh
m71/46wgcoVpc61JBX3GXKcE11SaGZho1MQ7viAwxTsGaT+/H8qUUbZuXUL6OFR5
Zz1LEI6+Kw6ynDDmFOzMfCqy1W2ngprQzEUOrWv5zmnV36bMwr73JUN/1fVBSi9V
AWVZEuVeQzyiglkCq9Acla2TkTosQYNui6sAFGnG5pUSREiMvctLZFMUDLSRyIxy
EOv4NvKBbxw4B1gFGnl7IXK4el/if9GdOAG8idmAU9kWRyQw9uVmJJauAr3SBZcU
MJdljs0SF4CZY07mU4McIFbRswD+zPHKVKZhpgfQqHlTRVQjWJ9ujgh1jD/C/GCm
o9wI9Xr9ULFqGtS2ZufXg2XjCj4fqViuimVWWP3Amn83ZpPge+klMrVlqm5c8SDe
LS4hrNPMRo0nvDkL+8Y6H/gO6TfxgP1fipz6O+HRok4TnlEXzaysF4vNifpSnfm4
6E6g+E5m00C8ac4klr3vQ/JT+SEUQ4zJ70l1i0QUdcTSWvfOv+4Ji5X5AxKH8sRM
rW/vCfHtutYZWE45WTFdNVARqJHaS6pMsF/DSy0dCzyiRUTzCHo6/BmOB3XWi1P8
Y66w13UmAwSjwBSre46Tp2IVA8l0yq9OiXi5N26qFXKlXduhkVvuvKI5eH0nf6Lz
WBHbL0I7Qre8nzaLhp9oNFSv2Ndzua5Spd2p8l7LQIcuZW4xM430QFRrL3QypUch
4NtiPlAf9/VCQr0tSStlS2uQcbjSKO+0HWzyyOxmpRQUdXqAz5hobdtpVlDoa221
m/v/bsUq3JildUgi4M7E4viCsgs76ZhbcICDLVsVNfcduy2nXdzN4RRbiPZYYshO
j1GME9TZsw7G6NWcT98/XcO1x38xJO2qMUDK83UV629FHGHzdie4tXMBeUKgvHY4
F5Pj/qIN1DZ4bUvNosJjZkLW/s9DXqel2EN8OxMv6ht2D+Ikzok7yGyJKf0a1VAR
9Gul5HY30icNXyCMm2xSdtXZkLo1X7/DxxIaSnL42uO9vlIrUYPbuXhjZy8GMoQc
PW0yinGm15/2/e/YlKrx90QxY/oPcFA5GeF/ZbaTHIjHY8gemI5FCv2GjuAIS0Kb
Ty0VfeAirvzM08osrdtA6j5z1JfJPQllFfCXfxiackYOQBBol6QtwWB/mvwRPDwn
npodDMpE3x6IK7YJ8omh7YsqoyKnO8EftVeZvNpReXYakqpYXpoiKbzzsGWI1Jto
MQp/UbEUhcdbpuEd0/vhcn/tDwRpl1Ms5pzpXxQ6BYgtC/szJIK0x3BER+RzQZ+J
XSiCKBZUvlQcVlZqEmMmSSfKvvJA+N97tSYZYhuOw0DFz0J9YwwAZYsLLxR3CEuz
Mh0JlKLNSo9LZJNxK5UJXWUFbPTvCGlRK1JD0MPRS2O4Sa+lp1BDHZmoRSiyzGpM
QnqnsV6pXcV0IvLKgCQ/Qxtc5KghOr93iRLFjDL2K088wQr9l/LMwb8JBw4y8Oiz
Ws+y2QEisGIMDPU9m/Bo3C/XEGvRKrrRZhFi7YIX777mqQFm/qcpmH0ZS1CT1RjN
Pyk2CnT2744v4B7k5bIf3f88Wx4HQrM1CSqlBy/9OIuSQ3O1a6brlVFLlxLQC1id
Kw3dc+lSQ53iMdnv4QboNIP/ohu9b8NhzWrbO95JC6WowSH+n6BvAzAhczIQXuI+
flp/vXnw5nhxEcubGObqoxaDXTE2ZHseXC/BPmFVVv8bwFJz7EyuyMKGb7nGHZWO
xXdEONYNzYPd34/DNjL+V12FIxj2tBf5YuDIfZ1TnoOPvnkdTPxd8OSyCYZrfOHB
/hb0YKkNPOkKYMHppljwqXqOMbHxpAnQNSaeXZ7bxiAYt7A0NGjWB2hw5G9Dydpd
fQ8WUJ4Ihjrzthq0EDdBQJoljZAdcXYBLkRWMPH0tSjOhd+qGtMlmS2SYoOMKoO+
ZxLYukQhXmm+SgF/+cXuKy8HU2jWsqkMI5Wx8GvAnTIluTdXI8mv3poIeG9SilPE
A13uyIbrxD91i1LC9HToqXNVlXUFT+uIiSBWFCnHTWh1DFaUgwFo95y1CL0khvDz
/tz83lzhhOLHyrQJtdjg14fl9TK2r3cYYBRWwYruOL86uZHbrYzS0AdI9YJPWS69
zUFMJxNAFbURc8mdX7uDtz9Blv8+TCJQz5PT4LZHltTwU7bE1YrnuPeaPLFl9X+B
7kZOsAzp/YVye/frQYDAAdG8z5xz0aRONuC/ADVDrjFYKxF90eL9uT8Z6F7nbk9N
NyVrxxd46rpfVW40YDTui8jvBt4GvaI7ZOXv9GiyNNrLtUySdOeXnniHtoVHhVak
XAtAw1biLPWozEqB6B7jSkM6N7ZjtCZ11+X1maIlnVXhcDv4IDG3pd05xnJtvqe9
2bX0SkN/ZEIJvNjpTmwpCWVWX9IM9X38Z4oy94qwHywzL/0V4YsCySXSzFKVbj0S
Apy0PZhDbhKaxKZsB394Qc5ouBKrfWXKjnX6D9xDrt4rLB+yt224NbaHAI+Um46Y
VdAP2F7j4VwaL1u3R6iRRqcGPRD29gzM+8gg3XEHQbxp1BxBunVW19rTg+FcVEi6
C3lrHrzBzSYuh56BNE1r5MNYbyoPfS2eas4PcnojTUp7o6DG1O98+io82U+epNTd
Y7BmQlRkTLfGOAp8a7j1TDfiJSSyTNFSZnLkuSCHdnoMaDeOz5eq2ESRgFLqZcuB
WrXCraZrsar5W/HVlTXPE8jtlhjyX+KA7cEy3IlmYNB//JvyBQCU8R4qw74H8NpP
YizDj69ZRegfHTKL2C7SwSO8VQDr2L5Fohe3+zRepBpwhDm06aSQtzPfd51oNRQo
amt9ADVeQKPP0MlVL+5QjL2y/97RSg68ZHaeEKQ4eGTCJInU0RuxbSUlh5Q6YacJ
63M8hm1l3cmqJWJ30FUqYtRP79EEZJUkyzWDvXrAE0ePMuTNUfe4tqYoy9vnxRWo
vVzH5u34ahx80aFNls1Cb7xQVM9Cb9loGvgOWeBOUuxzFwu8sOB7p4ZIuaZgObo/
nFAKfmPYF+1gB4AUuXlD9CBRUcD3ZMNUJs98qRyrnMahV0zS5OPyTqP/QIkSFomb
cmbPibMXT1n5zQJpCthngM9S27gLbnix8lBxPOnybdrqJcdqvVFVpeVXkCE6aOdt
MiM4N/yiKDW/jnyHte6VVQe0riWsC9Vj7F9LK9q9nduVrecw5emmnDnCCa/7CiER
RYMObjRs3YFToxDoWUk4DDymCBGnyT43ur/3YD04PiatqMtbLFi+d5CDoYKtbg2F
Aoo99Xmu05PEQEPFnaX8Kc8jPBT6Z1HNmQHQM9W4NbIMpKokmKZuHzec8bCzFg4F
WJ/wtQ2GVklUx1Q0S6H8+GIxgS5DNp2jid1TUvzDmUMD1PjbwoO3aOlc1b5p1uLU
wv0k6wheGTxWvl/4VaOSNubqrPnlInie2oUqit3EOua031Q1sRibYUOy2fmjE4QF
EiDiPi+9Unnq41tBO+3CMycDWdflPG3/fYN9CfcEHQUG+nKweIntSheWIlSSSyQM
zd+flC4Hi5uxU7cAj4kcmjszhbf6RijCuuazgfizg0PZ5ExCgTOz6TrVZ8ated5k
UJ57PtOh1T/Kac8XGwCnWW7E+rf2TUmLRNIP8iCkBexfo8RIBiCFy+Mb6B28jr4Q
Z7LoLGT2ZoOCctjVIA2/gGSuYCmCWliGUPbL8EnwjEz3lJKZsn6tOQBcIve2p5LD
zDdHTlp6NEdpFjv7A0ou3/uz9WeVqwcOI8vParyK9jqqwdo1xRjs2s6PFLFHaZWa
zfmE8xpx5Xajowad4pbLTZDzswDVQh2DVdJ5ujlKBJ2eCKkMtfOClVwKfU3NOcYr
4NNRdnvS+7vQOPPvsqPWOknXaUnaNj9Cf1mYqSQdwnu24/aY+B7Jn0JsA/8YkYva
4kFfPdL3KnkYd2bEyU1l1qm0jPt3KA3qV4+cFoe/FYOSdBti7b4VSAkK4VYUDQhf
rLnMo93UsO6b0tW0wDZgdvbYB4UV/VdZooSypBpWs+iUuwI+KP3SqkWqdyrc+qGx
hktRZBD+S4mpiXfDLYD9U0FVLrIvTSY694GLa7XnUMvkDFwXW/5AxG+brsO0XCkB
xO2dt7DFRGZK23iu8X1zKWvz/7vhI+lPcMj25EHVJl7il4VG9UtrO7ivRvWykXux
NTPisx31Vps8ZUqQRely4hRFL+5hAavjFxXpBsyfgYIx+DuGOCJXmKbKUIky8rjl
8iK8+Et9zi++c5RCW6Ouf48t3dD6rVneswggSWVkgVsZ39r7Azvi/OAk1pf57Tug
v5RzRVAePgnkCTeA8DXj2uJ1R6GfYCM1UBIzHq2ANOKVRJ0OQ+rU6KqpSYnDdvSU
9S59D1RHdavmxKDCZQQqB6T3eMH26XuzTPxlS6f+EiaUjlep4sxn/I6YiEEIhh6G
yLVLUGD3mV+rv6w/SoBrydACWno6yPo/l33dAI/SBnXESL0usyLSfJdhKySZk1Cj
JR4GNV7Ecapt/qIzCMGFCJm1RH2XPBvpMT3S6zlQYvS7MtCAZAynAjjpMdL0qzzn
A8gTq+nlid9wTVEQHFN4/2IPDpLxYvRfTBNAhkEq/00WNDVCWc6niyMycFBBbwyk
rWdtR6JiZ1wNwkzjEjajXjgcn7y6c73OgEFcp9wb5IqlU+s+8lPLCI8oaMiFVg2E
pL41yMTwZobhw3bqbdPKLWyztEm9gAiBsOAaqAhs/RmG2hg4i0DcmZdLGM9SaqGo
nUF8Cqc7uEnMO4uZBbEQlLasespmLh11k6085+JPQsZtyVVCPRSIS+XQIx0Pq99N
To+l3T8Lvu8HrZ0AEKknVZ1eWpKgo2F71W+GU8+3XYx2EpYGRTPju2+0JlzJ66rH
qTmTEE/BBAnFergzDo2nKLZ06yCbSHUKaUEVO/wP6JuxfGW/ZyYzEYHxYXjK5401
lxbpXV5MGD5fdWxfvvSjTQoK9pBfRCC1s1KwMt9Bp+Bqx6rekq8fCWEYo973ft/E
we5dlUI3/6dUDhQUhJEchi7vqfdf3ueOfaXQ3PfEYhekX/qqePJZXGcZ/tCy5/vY
6ua23ZtSD3DxvNcdc2t8TEtQaDEZubVplgw5bVNwZSnGzIawfX+3dWFRskz9tWUC
De4dM6LOnOFXNtyFsBq8zJUGQhMAKnD/DciUGMfBmUaYIJyvX8PQHzO2FJ1By0rj
Uki09/o6p3+cSoS8cOLqRb37wne+b+rvr56Dzqqs3WaH887fpNZkopQdILR9Kl8l
OLX0rECuqkNkwIx8XlaY4gYbm81Rk7267HLl3v7X1VrdSya8nIkpBKcE0V09Et95
hGcO4Rs0kjW5ZbYykj9htWt5v7yNfEE4CO8V3GwlseUOGtvegYrjTyeuax1hPPoC
Se3QB3PsTpBwY/wOGyp5f6dcIp8rbk/X/qKAAjKUxjceNeMwUyMFv5WKRG6B7rQB
TOKp2WhYQB/J4v3IeMD5UGGDVixJmT+XpSVa4z6M1BSrCPFUTkqFAw1os5CRaCC2
FJdRegHXTtJbO2FI5m60FO7KOscChuMv/euRPNH4ygrhjILNvA8ODQ+TLEU+ARdH
fucX4jlFm/5IulvbrG57xM9r+4pS03DkpxWMViJ+Zueqpw/f65G+xysfoHVsUU2l
YY8tImZqKr0QCnQbMcUi33HM41pFTi0aipkfItdHSxx1RX7YszxkDe7J9JPYpr0L
T8Jx83RK/doSiVZss26eTu5d5eLJVxl59qpfQl7xBZYSx7uAnetOzTExEu8LVj/v
uPN+joHYsKBN0M8NRQ7EfUyIm524X/SjhdL6riNxfap6IVi354WK4jEdRtMo89PO
Hip84E+NUKB8gTPljXuTxPDhq0PfS4+LKwuMZFGDG9/L0RGPyxGbzTM+armY2Eyh
jGzuwOtiYI65EbCideOj3Hag5HxxsjiEu3Uy5xwGy7IUtnencDzOMVc0QL6xRCUu
HtFw80+xs7jTfekGOlo9z6Q3UDeHLOoshVH7FOqUBxhDjRJFda/BKmY8MfXMdivn
DZNiAP4bubbSOS1tzs9MTMaFThnahuJkTXeqsmfqOMNLOOTyoxsgNwByQvhbAAm2
Kn7JTiiTanyNLokTQ0yaPHWXey2bCtW0LnpCyGtnm8o+G2MDywRel7yFqS8r1y1u
cenqs9UBZszp2upEz9PGOIbIO1gKIjAEIZY1ITlHUQARt/1rZLbEI3TI3hqqfKJV
d5A9kbYKdY8vcD3kW6UUbqg9UMjbjHuAy6CZM5sPsOCDpoUVYCDxYUBXhutjUCNP
GnVLNR5Zt0/pa1apgC29RphQ0XUo8x+lreJvnLfy1XCM8UCGVTFGLjrHvQm/FudL
jsqaZXmKeQKmBiTFG5quwcG0hZyhT+r5BlLJ4V/7yOn+sccTGPFUDtOvrnYpWgh5
llMWCpTyirBQgMEFUOLOo00ROc1lWudx3BFIxuFzxKzaE6BzQ6c+gzD3BUhHROzN
M61S+Md4w1ziEYJxLbpdLkmXCyq2bs6l59ZXZf1nmDm+a3BfXEK/xP5rcPtSEHii
WFn8+xfjoBZ72mr+FvRYoG4UAWguhOP6LrMFYUiDjl9erZ8yaNnyGjDzY+K2nTwk
dy2aouoiMFzFxQ2h7yuq7jFfYmqVzCeIhaiUkukQsUyrdmp0NJuO9rtYghD9fg0s
f3LyfDVn8fiSMm6f8oeug6oxH8gwpnZ6zJ1WA9jMTEWdlp61Q4ns4X8/chqaQWXm
DvNURQsiojQht93Uve0Q3IPQMdyqnZ+R82C87oo3u8fJHZmKxaPEQ1YATLc0dVG1
AyRXIgfvlRBmxPjhOi/ovFyT3QrRq8+wM05hkTZQTvjFjuVH6PMVZ870rbwDErcG
xnrTcIRd70cGkTYRT/a+TbDr7o3PAh+3IKInU/BfE3qbU/1MUz8dsPLmk57o92TV
98ZfSNymlMhMwa7xQcz84Xq6XD0I39KdNgFtN1p0lWcpLh/rrlUNADhAv0LjMYsS
G1TcrHiB3e5G92b9FUjsVzMYFwfyrKhyuWHBrT53jt/6XdItwHRbhgGC4Y9tf3XQ
MZRHLoLYEGMC/vkLa+YUsiacwVgsAwT8H0Tk7xecFMCC93rDXap45HakWxAfVkGv
DUBCXd4ifaAGmsf8vI9gjL4oILvOvxEG5dSY8U+mFncg0rM3C82rwMJ7ucBCJFA2
aibr5liEuyoA190Ob/ezMeWm1t3U2IVfu84//j2hMdFEADRod1Y8ZjFQgclfPHM1
zxP4kQcwzjM5moGxcyUIVy6FvksB3HA2mN+uPw2V9Z/jd1WAI59rLFV+XKvj94Q6
BgxbvVfk/bEfXsALgW+KKzJmIcY/uEZZH0R/WJ//tuCsffSkckEjNevIbWR2lx7f
pX1iAsVzubF/wfU8J9OK28jtZXHrpUYKo9ozVs9kU7kxNB/EVqusRB4CxkuJiPQu
IwBVEMbfKBLN6EKFs/sR7WHSrR9vcMHkSF+PWBSjw4bMYo3e2uu+E+Mb2fhS8w1A
PQgCk7Oz/VXVLOFBw4ldxAelXTejbhwgRa0sBtqjU8p0eX+h+Put74vnuwi99BXb
VxzDWeE26KsgIlfT/YliXgmCNsinSCDx9I+G+3ENU9QdAgj4hseQkDw1KxYG+sfT
VMGqZJpuIguUHqYik55ZFXKBIiDinGVZLaWVXTP1woKDbrkIHY8o+DHN9OjE8USm
ABlfe11U67cJ3pV19vygm9D6lbDWKbqeBM2R+MlA8hhyvQwRwYsKHmUrmCAXOvOu
I2NU73x4XYG97E4pl3Jc5JraaoFJtxL5rjz8dRGhz4UXOHAFa5P0y2IalPZlZPqY
ETrkSdWNlKgjH7aHeRG44WAap+90N62woVH972rmXtlGVmqnP/i3YJKyd5LGPia8
VSIFZDGXVClVkuLQfhM0X888gwR3OKeinLhhqV94JyiDJfgH7frV7HwQ5KCWSPf5
3l2ATL7zQsNnxr4Th+f8rLxTAtlvojyXPvLDg2hdCROuE7dZZmD0YZ2hbLmegi8Y
pZpUITfgItvH59xcehWHJsyYrkXWzcTPBw822vfGL8AMbzS89635gHOmFzvRNgyi
GCnxr7lyeINFcvmPSNqm9layUU+y5HUoQA28l5vYGf/PYp8TGbjRWRREehsIU/oC
LMsb326QCXQAu8oS322asglYBP/HQV44mCm7NJnunGM77OJM3P52wSsKjyIy5N/9
NUF+m24/SbfKEd3HovdLMvzY3cOtr0HKIailfssv//dQ8iELfIn+9Hq149V4qDyD
4E1xoPz03ixdyP3+Qm7WN6QO3gQ6Zcm7PRc7QMDTgWmkAz5SjfCffdVr7CEjLE8a
Sk0JhkOnt3AfFk/aviINhTm/dbDbcL0qz8zbykzNOmy+Ar5gv/KaJ1MpzTCw1Kvp
Y48bO+xE0UQQ+58Ae9Jzs378b3r+fWMk27moA5j4JGjK/ZMMG0scpmv4cILB0Bog
HFBdHmhbT5L5+AAOOV8uytakxh3+7a8ajLSQqqj95+1U2MpxdlozC+R7qcBGx1N5
BJxeAOc7YIjHhkPpyF7AOB8yN5DN2APasFey7embv36sgMsf0r/JDeCoqJE/f2jP
xMm2HCC0fmrVCi16H/GjGxOrKcDriPYnZDFluVf7yHrkEf7289hYSmdGCVVqNYq7
h/I6GINVZ+1+vbuUIMU792wDtdLG1aq1J6/LWSoCHiMKEs6E4HXL6EIDjvjNDXhZ
szGJ15eBI9WDlFiU9zOR4Fv3rKnn1RCqEqnbAzsUDeWdvJ8u2bXIoBBb9H/x1kld
z0SEMhOhgD9D3+lG+aDHo74dPx+O/nJUqxk7XweG+rugj770Ns8B8Dz/C6kzU1x3
vY35ly2yGwaT904Q4jnR4F9U4+nwRGX87BkYftcVuaamAQoMS5fBo2psFhXxBC0C
w/IDq5LXKVB4qjlqI8JsUFDtnz7VmSeB/2ij7FtUZdtPXS3/S0AUyYpkd5PtZwWD
Y8o7RZX0+KFPlLz/9Y3SmC4o++tia4JzvaZ5kT89xA3ZwSM91m7MfoOiL/0OE1sV
Hk39W/Tvd6OFaLd1lc2qUaRB/NziDcPVTvYH504kiWyAJ5hnuBOvMR9T7ulfbfgo
lP9sdw+fY0I3AFPHpFLo23xZ1RAZyEgREGtvJeCZufylDOyfUfjwi5y/a0+oNURb
bWTPdkRCy/r3algWyZX8nEDung6BbKjQMj/Tx6tPS68xA1BInm0J37ugYc3Y3qTu
ittvP2Lk/S5O0QGEpJr5BeWkypTVyIug0OJq2ncoaBTUxziTjpWH7HNUwRXe1zWg
VXfVJ+dMwpmegP+aVwC4tFY5GS5dTpKF5YjN9H3kkuhv4v92UQz9/GLoilnyfvsY
UUifw5JEM2VY8g8ZlleN9HSIfahrI7f5bEJyMWeVZ1qUpnqglYWLFjuXQCHclkm/
BUl6USiZIhJGSKtpdXLeeq1nPHL5R7++flV0mDffVNVy0opD3FeYkMISJYPTIz4F
PQa0Gwl6Rgb3vfJD5Ix0hKICR9xe4lMJjZBV+6HIQc2LuwFmv+TQsCeK45Gx9zR4
JIDhjtvQHYXwQ5GMrm0Ce3jyrgQUvyaiuZEqlaAWyjvUOInPB6GzLDGzols3EZSj
jhu3jghVz0kvZdYfVBaS77Qwdg2cNKfooxSeiMSy/IAxCH54TPclJhp0YSlKLMJy
oUu5ZCOxCkbxFivwZ+YivhPhk1CN9IO0MBOVs3GRvTigHkdTAAbrB2Tzefs/RO2O
o98NPva5h7p2Q11tR7jNRLcnLyzILnooXtjTWHcbFQExq7ZHmttbFzgbaFa7smR5
DixoUQOmdKuKLFv6bJ5Ug7KaffP2SH6hBY7t4J+VPEKBPejAHEoUnG2M0e40ldPP
s3Mx+9wdM6Tx55n2fTfo0/iQZvq3o2BW4IROXEn9Q8rzQMFoMS27oxrKQs6/kR8y
J7B3QwI40nsWvPzAcxyJwtYVyPuc3fPuMzCo8T/13UevHkyFzcHXoBbb+rmqBedm
WMTb3VPawECv3HWmTUMGKuDlK/n04F/wESyovi3bVJm+0tToojk5Euw9MkxK11jN
PytdapLNZbyweOqwcOCvw03NQWK2b4gWfun5Ye9EfTsmBbfh1ISe7TeDA8Ez3R+D
bWmyhbnUWpJ8qUOcf+nXSdIznduEJkSWpvSfsKJrSWQIjHHKe3zyBPoNMGjAknKv
6eIYXbWmQWUZMq+dWfx3CSh7bAIcP941Zrsfb/RNX3tWmEwNLBe5Mh4R47vZYtoC
RnF7CvH79wO5mL5MP/vFOr6MQcbX3JA6/V4iA12W9Ge8gYTpbx13PEnlmFQ3d6xD
LIlBFyWh5fMNXG8qpbvcC8qP+MjYYq2QqLtdcACQXPn9AoJ39O+nkPW3dgqOlcsd
tWBPoguAGh7Ml2hj8+8iqB8ojFt//ASc8HdhOrEvdKRFqCqa80MgpUGHtMCliC7t
Wk3fCcaEvesLYv7fzR4lwTbCyzaxKI/z+Ts5a3oCk2FYp5gGCJfhGxlT+p4OVpQQ
eY3PnxSYbgN6/q/1ih6dTYcu3shpmXNsKGtt1/RLVh2Y4tE0E6wyUZ+AalwSXSE0
/g95UE2S1l9hTD0jM3lPtUyk8sYK8TDmYc3LUWRkFIYdbMnJLdpptP7tfzcf0x0x
ma7GHCydB/Qjce0lgWszLhs9KLtpBRvGFvLASbACvo+WVFB2uj4MZjadeHJmwHf8
z1EX1klkbJV9xZCKfyq/Y4t/v3MbIq7ksPGujuKX4YALMAYkfbkWkQCCX8C7d1f5
RAK0JdpF0UrfpAdeA2bSmBoQABC5TcgH2ewUiI0hqH6a9dbTugXnjZYFBTDG+fMQ
v7bfP0DdN5J+IjQI7WVCVET2tOefWOQUOLmiEeuiXgqthMp+Y3dcLM8aqu88q8TM
pQBvmcR3yDwYL/9DJtelIfK2rdgjudpZFei7zOGIEcEKKk/2/EjzdNYu+lrVTW9V
OG51Zp9u9HR5c7ohs4c+eLc6GcSm4ZFjU4vB6RaPhTg+a5CHzseRRLEuTbQv9pUl
CiIj9De+UdslgffwEgDxdgSd7HW9dXVm4ZQExByx0ga0cW4CnDQau6zWh9aURapL
GuA0VxaikCY1/PCVnbmNDoXknMFAaoYjNNoWq4NSHq+icrQDXq9UlyI22F7kndqX
Hx1vFRqnUSXx0xalz0FdRsR+oXLaOIY8jzQJpVbppObSBTayn7KPU5qbl70nRJGT
ojOzkCSQU/Yiz2TtBhq0vmfOy3hwvl3Vx3F/zgtEDVioQNhfu0+tz4kzVZf2nQ9P
/Ku0SJmitX81678zaHM/hw5U3JLM130o2Jyi3/k75aqWVgFEXFP76Pfm75xz3ugb
qAndHiGRl/7QJHFKki961k8kEvXFHzZ3Xvon2BMvZLpMzMjoAc6q7lUs13VNr2Ao
m7OlccvEyJSmY6IZq26+NaHxGguHRr2+7LnZCzwJIzfJkWQ2IcgU3OVxb2hhb2DA
Fm7nu/ueCf/O6Z+a8lryifwEeQcSUK9RIZjQ7Hal3DENU3asO24IWS/x1EUYliGB
E4HwCQPf4AYa0awKMzy1eW8In18wx47mNIHbn7oxvGHVucMZLGut4ztbnYkKu6f1
Q9IM+vUpq6vvYuc+LwEw0EKI9/Rd+2GEmrXALJJBpcHyvdJqCWYaJVkApeBYn5oe
BK8o5LTd1w+VbKwV1HCDAohLK44WbqPtBzMGQ9D98ozRPSo57STOxiyWsz9UjtZf
svXeY0prbjO0/1WC6a4zC7aylew5UkwQ7XTuz+qQ5kBucx91gAbkaygWmN7eSVPq
eWwXS9HgZbRDVasqDAMaoYrxJQJ5ahpcfqNTmHr9hK2r4CktK1GFoP7WJII3l/xr
A2znE7jizt+F9a8l0uaHeVjUGSjWzvxWz+hH+3pbllCLdF5kn/CzPWcWTzd0ZoZO
2dAZFVXXouEfisRfXjos978b/fdJ5zgQMfXMnm6IJKP1xwa8WmUsgOWKAMDwhZDF
r5eLfVbDUPgF1lPFzvuZtd6HMcXR3BdmAJwsIDkvKZk2EgZdDM7v+EZcHezDd1Yd
65x6CO4nK9+PJWSqGsYaovnCEUnldoDicQXplFCrExgJKpu2kUJ5KDOiYxFznD5l
5MOf+7MNCAWnaDRUT1eMAf+CMjLLuCOnldbp1fGgm0IfQ75WMo3HaChYH/3uA4BL
Z03dKCq/Hfy395jHnsrK01zwoxrHkl9lgBuaC8xII0MMkjaX2BWcDEQ9L3QDiWjG
UrW6BxPN+AvZaQuml8Ii3ayONqZ7RY+XH2RrF9UU1pPviTcSdr8ozXxeMSi3g3J/
vKxKMtiSwL3hWY7nl0Vh6KIXxEp5D/v+9kDfkNHti4acot8MW/uOQcw9NxLUuo14
IuX5k0aReb5FZO+UC2zUFksbrjWaHv2UWdovG9xOEgyLPVrs3j17Az3ogin+j7iZ
Sn9/Hwn4bzug569is+W6LPHKHx8Zoz2+Bd5A5FUIe5bLAldm4z7mCbm7bIiNh7z8
P09sKiXBrakqlcMRMlTOdQHs7LZiIQZVcQuNZHrVUrsrRsRj8IT6OFX2vRti4OE4
FlYB+pGxqSYRXAow9+SewJGMzAMb12CFBsWDdq46g/+Phmw5qToWvjGDv/mJ7xti
7JWE3/YNcsS810WDV4TesSOeviv6g/12nDZICZtcdsE=
`protect end_protected