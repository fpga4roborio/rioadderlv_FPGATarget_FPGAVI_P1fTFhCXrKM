`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
ddtXksX2+yylW5zu6QL2Lhnb2d1sD00763mmSITNX595NcHTEkwn0zB1Dry37fOW
FufOhVzEJp80NC5qZ/+F0Vk7Ik02dIR0elf3clrjeJRK85K4e3Hoo4xn7YbFUIms
l/8VZSb14+JVGURjfswrIyCUotIzlzVYZ6gzoZwDXIi5gQIBf/gI+KxNXPaKV+PQ
Ufys/12rjO6aI/pPlqSm0hCvftmBcnezN2hk1UeXgOIuKZnogjOsf0iJVX2aOOWE
6pD/psybjbnsNB6kH5uFTA5frkzIzkzl5d9+YDm9OyC+k84E83I/7/j+rk4L2dah
QJOvksSIzN867/4Qt8qYTQ==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="MvBXkzurAa5VTw+1JJ70nePUfoQXBvZOku/SMmg4TwQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
oRtzZL4VJ4iwysPsC8SXYCzXS8Fw2gtZTOskLcDV+1B9Nzn1zTyNtlo6lNICRmmK
ZRVu2BmCc2G+fmzynYlNTnSa7C0Cuel6FYpxCBlOuk3OF2tzAmLAuDyOH3Z1Yjzk
a0aHuoCdIRKv7BrZCdALt03JeUmXKPdOmIlkVGFl8yw=
`protect rights_digest_method = "sha256"
`protect end_toolblock="Jn9CQpRhJt4rnzZPRk+dOpzAubz7omckX1MrFd4p81o="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 3792 )
`protect data_block
gD6l00tciPUa6pDNTk/+t0OO0nC/UTtBwLB41d4inuAUA3i/ALrNyoJVcBnAmEQW
ptbcNp5fxEUJjnOxnedyZEuEBxWRieZFQnkRdF269oM8eXOHcKycjkKP85lWa0yg
5fVYgHv56yDuHMiicHqL1PEDfcbT3bsqbDEX4UypFURuGdwcCUUoZ31DINDaFzii
OmfcD7ZLLk8PnAsVDCTxyjbJg6tFRDpwXu5BfKDsi7EKBARPTgwS84myrucy5Dpg
vtUZyzA2FdBTvn9N3OPkR9dAMMsKgLgkAQRD3rezzV6w+U4Z3c448CdiyRutw13R
zbBu2pE3RJah/LbO3mK148BrZE3wDf6RceHMJ9h0UVl8RgPp9ICRtWkIf6ZOgWwh
f6osi8gP1KoOfbz1A0O+V7S4TXklcnrQNaLlfXTQzJXkh+7BxrTsxVZP4h+8n7a7
EjcEkbXPQAXzV6i/GoOpywoHyvSS62G3w7F3lrh8EV3UCAd5KR8mm2D92r0uUv6+
fcTOnyvNOpfxtxxAicSe4JdN1yjVR90Q3qlJnyWIbGkMDOMbO+iYDHxVN7yB0n7V
Aam93GIrpT8SguiL3v2t3QsjYwApbl3rWQmmZoBb2rI/lYWW0Z6muDvUIPiQTBtH
0BiiVRTD1usH4vlE4NIED7xuB7JoHpzYmn7Qfhv3g/pG2ldLwJWpEDZ/aiIeAJM8
J1BzhJnXiOGgHNmEHGn4WZUoZR2dTr5jbglPEhe6iEebvE4a85KM4OWAzz37UYsj
INEOjr7p6SOtmsZdwibea/ohbr79Kcj94CWcx5q56NprbuCLI0/h2gcCpbcMzF5t
l/S5c+Igg2ZJfUUOFz9nWJ53tf5mRwWjyu46P1PiCrE/n8a3AwP3mM2L46SbsyvL
N4BPcxKuD472I3PSuubf5BX505ANHCBHwrBniwGKFo8OqvkS212v1p7RAryUhvPk
sujUlTYg19Gg/PyzhwT/0k1Ex4RqReeaRib4cSkf2h7XzM3ySOEEMun6gDXnUNa5
yJdy0iwu8aQBjO6F+vDfJgTsm8z7E9CKFZezCcQpVPIOKXJDQwXf5YIu0sj/7M1d
FZR09lDq/WLiX5b52h3OyNHL5EGpJtlLVoUtShmU36IjfgotIev9S9z4D4+zrXfK
DORtHFA7c14dQiBSm66PEh+nTbwjjxlgHDXmHkIX18PEU8Rwg8fEavzv9IrghDUR
GNbjGYaPq37gsWJW4k2+5cGU9MLFsPT5WgL80prELiAU8tTIwae74zWI6xpArTKV
ccgLmosouzcvD293fSPF41jmpbIeuwMXLj/CuFcCHdUHbqJBE2uCFPgKYJZGsM43
3pKrtuZKV3joCs/pRJ0nw8/QUm3Fop0uzOE0EJ8CfMGjAhUKAoQy0d/+41L3MEbJ
1lXJJTJE8/iiM1L7yXxMTm2h2fix0Zjfqx9NG4U476/a8LEmSjr1yGAGml/tUPE0
Kxtpcebf05fExQppNH2AgqJ9+H/pa+cQdvgfa2egUgjSbSwVBpPeLv5eO14IUhPN
uA05R18g292c5C2GrQHI9L9gteYA9QEIO4DetS9eQBto3047nwa90NsLeeFh4s+2
HWu2WHTLRJ5xEztCn8hQEXuTe23r7mlSxTBLvXf7isE9alp40th9XP958mdvhQ/N
DHUalQyrfTCjPUeq+TjF5pbLCXUNLm4ycv35pzB4OtG+iDDCnzyGGU4JjrmdE+TV
lfm9mTdO1Y9wyzZD258gN1QsXKTIjVrQu8RK5KxgQWWdwvMCEVL/caHtgZCwQh7P
LrXE+dbg7X3KigJNeAfw3LSUF29htkkx9wu/Jl0/8rxLPUXI93WxNPMm/an0XsMS
w+UmeDP3XT5wWs6JgaWXKLrF4Z7uLUPJniPDbWqQLIhZGmyOHxe+sfyULv6Jz4MX
Regi1JIVtAWQ9FhQXFbhIaMKaQUNnseQkO1k6O5lNk6ZP3RxHEwvYlU2UFRLTZN3
D1+N7yIlX5P9L02VN//yh2pXHQO1hZ8jiSDTNnFog+mmIPuXG8SUOyMFkZUZjC6/
KX3v6Pgl136Pl8DFe4q2MKDG0ITMT0HXbYggnRpFL+1++IstV7KEdUY1ArWScpeK
3as31BX6N9b/igvmAfHe78if92rds9r8pZ8eli1g27jQuYXIauBJWYB7sM7v5kyL
ZyHhUSbqkvxkLcgA+k/t5bq5NC+1NfkeuqqphuV3ZNg32NQcoavzAkri9NuRKNoH
b1O/TKRdDSwEuWHQUVZVAnz7f/AWK+UJEJKtjosWM2Essvi3VFNdHcBHpeVKHEma
hBrtL353J3a9C74FexUaw8dx171FdcFEm4vFEIXdWcapLnsw6pQWlRLG8X32+MHc
kTkJTR62k79N44ZbahbdaBMl9XQEcJR2B3KTgprc7BJbZImUE8Xq6+neyTJY12rj
bu4SZ6ACGA2Kh5XkVV1hJyaYXg5TqNH3v34mpaVaJcMnz4YbC9PlzJqqZgd8Y0LX
j0eC2PeKehr4LqKPXQzZVYVQJupr/KuvQfYc/y5eXXnyk/cJdor9DKWsnButUUSd
nWzI0IsJT0Rpg1FbdKJIc7Mr3cC7y553PTM3T0xbxyyKHocs4YnKX1CE+ByvYVzW
tgph4srUbtMCS+XwtVw5wvEb1OagXivRPSiHphFAnRbpMeXcHmFltokhwtNnQFkf
VZ8cfHTI9Q4M+HIBKo/c5Qgpr+0zm1b4FsgkiMchtBOXQqJy9TpThfh3UQ+Hypbx
iXNVaCqrzkznFc+lQ4R+uOQxD9IDgTpFGLtoxFDuAjVFsjfjYQ5Pla9VZJ/Xd/Zo
RAllEy2CZZBvSe+TOPFF/vdx8R7ZhBdkpbAoWePfk01kR/rOIGY97oRuWYbPZT4v
VfqcsqHwtgMTbeq4gJlTVnkhO/F4T/Eke27J1vXRmtz+9WS8hrX2Ue+Q8M9m5qh0
9XNiFyGlxwyMpqs9dEJGDfjd0iwFZ3ACwJutTPzYfUUqY+SzU4ECHICgUoiWtK0d
E+sEA+EvKoVq6nubJTC/+L2YoD0C364i9RXHWn7Lw8FfQcKFlZ7AyOZtyM6hP7n8
UAOYFtqaBm2CqSGXgn7RDmTNDHtdRCnfqDtTb6TS5WdQUpvsURZtkjUn4CzHNnJb
9GOE5yIIUmN2Uk4PU80x1KJKjug2fzTwowMXtePpCN7tdo/7DMmsqTZ41op9cp3N
RzXZo944B6kGGOb2L8hKwOXPZHN6wessmsfMC8m8S7KVCS5ZyQvFKPEh8Zo3eoeG
7ilZltpM+yVCimG2BmRvbYDyaIhYZI4NNrD/Ui8r6euORBqu6bJffQJi8j47N740
r4mnxc1jvvjHUJ7MHBOXSKIGnyxTT+37R8D44G04kop9/qT29Bqi5dPKrr6bbVSY
9wavtZPJsc7Zt4OcB02jsMAjmlMNfEXTF4ndIzuzERAUOWkMlI8ON+WRBogDEL0d
BfJjBifXiwemlVYwPGPxRXgg7EoBdvlvWEEECpX1d4k73Z+n4UELqvcOl0InZBda
7N4zyZCXmrHWWCjsPNdkX/285L7qIN7Etp0bwLWe1tsrPWMVx7EpRt0qHMjUxL+9
MrgUSafw3NG0+u6Tdaexk225ow4h1AvXzzPBFbZm3EewQnHePgwMA7i3lznKIMGY
6ewnLsfjzPvdmPayT29EILXpCPRHeuBm/f6YI9b33KtSRFn/PAkqYSMUdfiNsFck
2UssBftKafxlSYptw9s74DWHlDNqEIFldx08mZ4tCTW6BgigK7eZBj/L6skSqMmA
SU3P2yG1vCl3+j7JBR1WY81GM1GqArKsSAGOukFLtDJtonsakpmLG9s67D0g+5X4
LGe+NnKw35TN+97KMe/u1Sf7+ROhBDKqPUkfuyv+bTtYZlIWh1AuSu5LyHyu2o/7
U2b4hZb30xit8uiOgVqSWXw4v5ZomGtb+wy9uUZoTQFzB0YLn9X5iPETXMhUzYDQ
zEoCK7+oDsIAQTbXyQ5DYY+hM6bfWa4VgmE735Soprj0ajaGbW8EDvWBNubZL76K
S0Mps77reBLSeq5Tv1dGmTgyQchVxhqIa4CIfjZUjPK/YBHbuwsEEKr4DnO/7mf1
SDOrbp3mLAZ5brhayBCI2SddDfAVtzbXnLPWXgl6KhwKrrMmlEhdRZqwDRsgJI0u
wd2eqOVN3xI9HaTjXAoZAmVbVnuF1gFhgGNUcorXCyqY+dSIhztiqVVWM4pwwJQp
GKugDx/ArOZIJJju0WMxf4gMB0azDTPpw01fC+voYEwuvflRXZmGyIlLbvamqNPm
DFzJzmqwxU6wEjP+j4/6W23K9mezGs+adrDQq+vZwCzLnphaM8+saYS9WLpRipAl
UTorIWHkhdSQeaXlmefIjI3ekoA5l6SfctkygfuPuAbjAsNlsNSq8tuPi/yjLcTy
mvw2VBAwJzh5Vb+Gz8XXOBsXUq8/JygSat5FH+4u63qWbl/XRmATW5P9wzGRi2nt
XZGyKqeXd4AT/o7yAlKMNWj6NS+ldMT38uY8Tot/gT3KaARU0QbnLcXTahbI9pIg
o5kp+4JGw3NAUy/YfQfnEPtiCq2xxsNUjo6Ojd65xn7/8XdFZyBuOp5Vykl86E8+
vrNCNAMvnCe8awn23SvqriX5UZ8DJeZCbLeVtDq29syWudsc06wp76vsjRJyZjQT
u3yEQnD6aDABr51o3E0BZ8H/AbZX+x1yyL+483afuN6NE+O1IsKKcbK1xcxTKPrH
7ooMi0BqpDXB//RV/c9ZgmcG8KJ72cvfHbCrVd7eH279UobgN9hTKygat5On9Gvc
/DeJxJGOSSkuSS+jJuUEqeJTUZEU9oddr2FASjYM375TSwrmZMdc1ZEJJa4q/IEe
bz/yjKJ+zR4kDfwaoV4pKXzt28vbC5idYr3GhsMDP5ol+7I9LZaSauJfiwr+dZ2u
aG9qSFFsSZlwV3XylqFV5lCxxLPfFtvsTz81oiD0UX6OF8KUjzxP31nP5hvjUnii
LxmRC9VgEMDnyfxacWikOzJTrNSrYd6w5oNonfJQcWKehvqeSEz8Zv/BvFFypxua
`protect end_protected