`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
ddtXksX2+yylW5zu6QL2Lhnb2d1sD00763mmSITNX595NcHTEkwn0zB1Dry37fOW
FufOhVzEJp80NC5qZ/+F0Vk7Ik02dIR0elf3clrjeJRK85K4e3Hoo4xn7YbFUIms
l/8VZSb14+JVGURjfswrIyCUotIzlzVYZ6gzoZwDXIi5gQIBf/gI+KxNXPaKV+PQ
Ufys/12rjO6aI/pPlqSm0hCvftmBcnezN2hk1UeXgOIuKZnogjOsf0iJVX2aOOWE
6pD/psybjbnsNB6kH5uFTA5frkzIzkzl5d9+YDm9OyC+k84E83I/7/j+rk4L2dah
QJOvksSIzN867/4Qt8qYTQ==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="MvBXkzurAa5VTw+1JJ70nePUfoQXBvZOku/SMmg4TwQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
oRtzZL4VJ4iwysPsC8SXYCzXS8Fw2gtZTOskLcDV+1B9Nzn1zTyNtlo6lNICRmmK
ZRVu2BmCc2G+fmzynYlNTnSa7C0Cuel6FYpxCBlOuk3OF2tzAmLAuDyOH3Z1Yjzk
a0aHuoCdIRKv7BrZCdALt03JeUmXKPdOmIlkVGFl8yw=
`protect rights_digest_method = "sha256"
`protect end_toolblock="Jn9CQpRhJt4rnzZPRk+dOpzAubz7omckX1MrFd4p81o="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 4352 )
`protect data_block
gD6l00tciPUa6pDNTk/+tzLxvdHE2s3DQL3/JqqujQBC/Ei+vcAB8wM3doqg5vTg
mdfn9XB1bLOis2CVSfu295W2DNwHfMSTc/8BhCDRnTlLIX0UCJs9Za0+LoM0rMrV
T7EjVWppbP+Em6PkVKCwlmIQ7JKaifJ+Y+kjw9HCGboYo5074hY+K/CBbfsBQY86
AyoN0MKhsIx+eViNgnWjA4oHW4fXc57/W2kQuu3jllT3zitThKnfTp20tdWMl+3Y
I1Tc1KerQR/SRc19dkw15G7RrCyHBV6CFgpcZsr1ucZ4SraSWHADCApG6qn/thIx
1CdEyOjZVNOnq0udnBdQptj6pj+xCYbagjq9KiR7r7YCyOnoGJDI6cZnnrkYPQY7
pBu2/K183dCYKALIeCJLJQQBH4P7IvjUQEg1oMKqyagbR+g52zkMwmFONxU3V9Qm
E/D0O1HVQW47iXivREGxwjcGVWlK1A6a1dthAxzKJYdczDqJO2LX/KZFSeBcLsDa
yr/HEwheBx2jIYtebjTC8jZcjhMBiKK+ReFE9WfCNhQdXS2OTHu5MxAvc6K+VISs
Hpe1JKkvrgHbT6+jh/ICjvrdKSh/43GzTXHNiB4vpGaifEwVHUHaqVzNGZKvPNkU
X3wplbB3v1ugavTmZcfFVkDYXpOAYhDZ5DtwRqHMHQAsEVMb7F8unCnxRQ16OKiV
xxXS+GxI+f5UuTPvDuw8GqQlk3I1h8p6E57Kfig0mBFLav0VVScxsYwQ7u+U1tEU
ZePfZ2Gz4wXlZ6DSwQahMhf0ye999BnYfSndNy40mLopdSrUloEFomzfb/aanXuV
dya/9WuETxq0GYVLsTeMKvaXaMNdfc3resLzE1QZ2/1yf5fIr8/lqhQrZyb9CsmQ
gJGbD3+7e6TfuPqof6PhYjGq1UVcIkKLMx6QSlyldhL92VzSygfQtYN79KXNyXgI
9uiV9Yw4mKax2jWqHrPHkcCdaEmWXU0WDUR8kl3QM5THVO11bPVtcjWhaEwFEr69
LvOuW1bOBaFPzjm7YcFw8qF0Q3En6EHPNxg6T/IdvuHCsaK56cKU05rGScSrjuE0
TBsTlWxjXE1B6JNUkmj2VmI+ZVYfYne4w6z3gpsw8/LItzKf2yejm3LE0TqEMl0a
GmvjIHfqH8fUPzFxi/0kyT+UCrli+JUjxeld3qQIs6nAic4R4utseaLsHIxf1ZPq
Txe9t1WAmByRYrFNsAw57tm4WvXw+FqstKEtD4zZk/II4i/+E7DiIVJ4SoBlyuyf
Qhgs3hRDEhaPfkmm39l4Zp2cJiqMi2qBhhKN/rD0u842geaNiStaakz3Olncd40A
VCH91fF6IDCGPvg5/mJjbBhj6343Cfzbsqvba8DCQ20g5vS9aAidkB7PwHyfXGFt
ML4k3RIVZRS/zmyJyNbL8NSo39jkmuv8yLY1WSVEm2e0sywHIfMrhCwlHMPHFe3K
E0r0In8mct4FqXBYN3r/5XuD/yYK3CvTLjHzjMkkllJfDaSr9cvEmWKLHRHCDtVa
ehzdKlObVp71jSfAM4PGHRH/T9VUzruBa88SSjwZQF86vaN+PgU/mpTOpA0ug0Oj
LjwfEOPPhMSZyRZ7oKkQWvmvcz8C06AO+lo+ZcvrdlBDsLok/cLfRfiz/fC8T+qj
z9CW56/qiH7ARDplsLit0s0HyZNK/hVjMNcFIbg2ZKSAPZLqWKBMPXIkx+n7tTKj
Y2oljx7P46QMXUNP5V2XHNfNOZT0uTYfj1bT8ccSX09faGE30JHVD4mljdYCyDjt
bNE+z2OeLnQE7/XC53/zhqI0vnXv/o9U2Ng8WXtdnRA2FKxaawiEqQg8ihoO8Y7W
CafVHoaBuLL/khvLmbmHGol0tm6R67yOE6SeUl5759HhpPQJE8gCFdMdBvymQuzc
WT/gBIystuIbMPW0WN7eNmnY0nQ6bmyqzXLzJSS60u+to9FI/nf9nOf+JCLs0eBy
iYfgy7pF9gIwG3DWyaVe8oniv3JlGYgE3cNq7+OBPw02gWoSFPXM3s88psBcxzcc
lgrPsibdEYvDZ6xq2mfvkzcpA0+q8WZ2+9zlqW18aaH/eNAhLYnkr/bkde+7FIvA
9zloeRRZS5+fctdbY0VokzS+RvR+Y69ymkNGMcmoGI58qiW8BUuZ5Yb/Ud9uZ4Ja
RybduZvSCZ0fmgayimC+JLiXykj1CHHMBYMA1+iDIhELE8wcTSA6tI+CSjYdcTga
5pQuTa75YonShPLVzMticrDOx5J3da3FPhAzx+bHKEZRlgaXW9asLX87f6TYKeg4
5a5PUmRXhEFJf8C0X0q/vKqnPXYovURusezUAW+fUukyi8KiUoxsqqlQQ6prL605
DfEUkBpmd3a2NpshZFlzK7e8Hou7O7l6kwken6rf522mwWb8FxIpF20Gtq0ZVmTD
hIMxoBPc8klt6hv6S2I6Nq05WtFpaCWjUQHI/iVfo+o7a033KIGzMH9qlAzcnohP
WuoG54Hkhbp3y8oVOQfQwJgNaCQYyBMNO3EHlCDXfgi00t0wxqc0n7eDpWPItP4z
RvjbUecycoE/yRqy+OxfL4/mAV0MYKSbvDVN/S1HhqtWLJYFIlo3UcEOAebbRamz
nm82QHw2stdHv2oXfNyu/MVs9vk2YLQ7/E5Mmr6x+93STej2R3L916hB6Esxz8V9
124bm8+ifVMEV5QDz9AMfHn6fvkj6xaziI4q5OOYinobT6Dz3wZKJd8ejQIScaL2
Ol99mKGYY1A7dn2b0B7eqsavXcWryQ1DnKP6ePkSbEQDTzsDZW+eMvxcTXpmG9el
CdHtdy4HYwLDO/9rOhOgFehEznqScyXLCjJ/t+vFhDTeFC9DOXZt4TiXAdmW6jl2
o+pHgFKrQON5LJWufkzYnB2MNXDluLzYWPdHgPnIVOPCsBsqEEKlFF04dy0f0PpF
PWM4Wk1DQnUWNJiiMEKeru9H+QplpKEjrW1bKHyWoRSKRYbEhsilX7ndfh+Ogo2q
XoGSygVDVtErnQD8R7USdWR7lCcCJ+GCWkuv6pE09v7KdtInpe9hPCY9zhzl1Uyu
X317B6xIxzL+H16BRj4AZTaeIkjChBo3ONBY/5dAXZ++F2eHLvVRWuQVQpthL6NN
hKmlHLG4xIrrZUJLi0XCCWWybL/DAfJNCnPcD5skM9Q3VqpPOHpM6eNygFVvmQJ2
NUhS5tSMaj7YxemQT58dUXTHo//za+pLl2TF5zuIUIZvo+0WPNlr9ZDz5MJ2ii+8
mM9vd3VaJ2Ur8u1j2ucuGnw8tnsz1edpWNSzyqt3eOzEDlLZz4dD4ysOl2Wi1LMQ
apd2YqLZowfN8HfRUVLt4TPFwYY40BnlcHAdZZo74v66ukjR9+gxy4GgYV+8WSko
og1oFlLtVLOiqmWh5ciDm1Ff41U4Jp8lfWWtFc9kjyOm0KVaIbKY8n7lV/TPU/9A
ttn6lDubfKrS6xxOZ/RJhLKCnTSAn5DohgLQa+2rKzvPyoQQlRRWb2+0SRMjiesp
nQcEh01WkxxxIXmU0ekomVh13aSDj0sH+5qlLE3nNtjUu7GMzzMOt1/LPaZbfJ1E
0C6vl5EshFuE+SdYx5r+7QwUtlm1pptd31S6rL0riayiPxp1YZHIWoi7xcMdjE/j
WYyIXLTQGapGSkgiWYWxKamnhkNDp8PPPckIH7Dsi8FGKjP+oSQdEZe1Nqx6gFgC
NbIzbryegYDWERwusuSWc6WG158fxkX1HwRwITBPWqKBX7sUaXD7CelHzAHBM/9M
dJLvCLJq/moh1L1usoBQF3KKwDx5AHJjzAn6hi2zcpRzOwwcZ8cr3sYE/xnpTB8E
jImqYnn6eegcm3huga3klI86RKPmn+vN6z9Y3JwkcLSjV2aMQPRmDRyyzNqFMD5z
7qo/bxCs4IB4G7WUvzgvo4TBQQXHRve+Tvc4K2xq8leG0hIy7pGtgmShlHmuraXe
DHCks/4j3e5FE+Rp3jitJdjpiyArtkRKDxD4K9sCZ16o7/JCnmLAyQ7999zm8s+5
Ow7DePzm2nysadQaM9wPXl1i0QrHm0P7lp+FdSf/4pc0Yo8jfw8uZ5/2wpEd6Izv
o2FkK0ZXYW9KCSUdI+0Gthdt8mQfv5RvgFKBg0SITaaXe3IAk/eiEqoDRGDRf9fI
Aqs1fxj0aW/6ANCqdVjQc26iqmKuW04N5VQdl5nSj1w5mCLjD1CvZ24Jkx9N04e0
1kmj+y/BG82jQCCm/451E/zoleUtflvEqtfqBgcwdzq5vcU8wExtgD624xQS8ROD
v0u/cEofr941j1JSX0mqQh+U0F8jZX9LIPWGtopWN8yV/1KPbq5G4xPwOx77MyoW
yl88liHKlaZwMzd9MuqnCUAMXH9HVE97ciE33DcEoqXB063HEwXZuRC37NIgauo5
OfVpUw8gFMknMV5YZ0od2THKTPcL7o0U7kHvn6R/WhiKyrxKrcG2nGTKAMoo4qlv
WQJQhy3GGhbfZtg+zvqI1ja1dr2OSSTRg0H/cEROZaTfT+0D2njAcUoHJkcgoav7
yM6eI57+Ll+/zDgaENCFUiCr9uq/qfNuR8HPINoE+dNED6un7r1ejLOT4MOMbjui
NttHuBv2e0wUR2Ucyy3ubpvO1k0ZPf7zO4RaRGyCG1jIYbFROhF/+g9diCVR1QYd
NyV1Ia0UQJte0ILvq6MVAhxJ03DqJiRqRpqrxc9PGye2LXqVlMk/+DjnEUPxR/uX
MIYCNg1J++BpTpAkS02DBgEPyEz9UIaDUSP61ULuR1/Dy3+4uRhz35nc2QzMrPta
zbj+VosFgOWmxtHCAtp8pHZn9WHAnMrsKiUT0YN0vhQRxbK0d1GcgyUAgXBMJAJU
IKUcCKbtniGP5RBHieKYcEKSywzwLtwrPrXsOtqKsWeR8v5nIBCXd3k/Gkhnw3wX
+IUDyD7u3nJ5yhkbyEiUnTvnXJPgXeVSzQfZVwBOW9POEcHN2K0Q8y0K57hAObKV
qmaZMeVw1h2U98cMUfRsSycM6wwacwwqX9hyWD8vFRHAy67YXW19JriBH3IXyIfK
YU6CQw9MofxuFwyajBlnoJCpcrDewJR9dVR3EdHTKK4O7aNekkECKpdeiQfQbukW
qtZmKaea/S6OkvQvkysya6V6zHE1D3DiWf7YzmkjBNPAkM0jQb3HCx6atbHvm5SC
Epk5qytrpxObZ9hR2BGVbZI//XmHEQNoLKhhE4ZxvwXbECmm1sWR62PdeayjMh55
c7CSCEtIjP6Db2eRA0aFEL/+MQxmhougoNZhaM5nNO2XYvsJXouz5v6z4B8pg3If
XEqkYZIxkE50lugklIqCqdYWMBdHu4VOLfhR2Qv3rdHh9SHonSxne1srnKcxyBkX
/4aQku4Ea6+CiQIcy6KessNtBlUshyXm3c1FzL15N0LBTD4PX1PLYwitwKOeC6uv
OeiSxaUTnkq2C879bmXwKYu9DlCbJundzCDAjZlRtxvI0kfTqoAXA4b6ZdQRszh0
FwZ8HhVg9mtzKNRG49o1vYHDCjUYFVRWDA88BoKTuLIUztEhCmXXfRHFDrtrgNRj
qyPrAkJugHn+EYfCu9OzR5jWaYala853AhDOnCk4YaTyKOT10czZvZl4G+o6X7QB
0IMY1YhjKcU0Eay3hU/0dI4SD2nOdo/tT5SuDI43/e8jzJQ2aFpxHtnOA51tF74n
uhz9/c4SI6e5qX8nnMKvYGTndRIYmffHLni1Atb/dXo00Yhxby18UQGTjhxXZcKT
N8qPCCKmG22mUSbe3rJA9een9CNnyaM6VziJXzNx1Us=
`protect end_protected