`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
ddtXksX2+yylW5zu6QL2Lhnb2d1sD00763mmSITNX595NcHTEkwn0zB1Dry37fOW
FufOhVzEJp80NC5qZ/+F0Vk7Ik02dIR0elf3clrjeJRK85K4e3Hoo4xn7YbFUIms
l/8VZSb14+JVGURjfswrIyCUotIzlzVYZ6gzoZwDXIi5gQIBf/gI+KxNXPaKV+PQ
Ufys/12rjO6aI/pPlqSm0hCvftmBcnezN2hk1UeXgOIuKZnogjOsf0iJVX2aOOWE
6pD/psybjbnsNB6kH5uFTA5frkzIzkzl5d9+YDm9OyC+k84E83I/7/j+rk4L2dah
QJOvksSIzN867/4Qt8qYTQ==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="MvBXkzurAa5VTw+1JJ70nePUfoQXBvZOku/SMmg4TwQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
oRtzZL4VJ4iwysPsC8SXYCzXS8Fw2gtZTOskLcDV+1B9Nzn1zTyNtlo6lNICRmmK
ZRVu2BmCc2G+fmzynYlNTnSa7C0Cuel6FYpxCBlOuk3OF2tzAmLAuDyOH3Z1Yjzk
a0aHuoCdIRKv7BrZCdALt03JeUmXKPdOmIlkVGFl8yw=
`protect rights_digest_method = "sha256"
`protect end_toolblock="Jn9CQpRhJt4rnzZPRk+dOpzAubz7omckX1MrFd4p81o="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 17632 )
`protect data_block
gD6l00tciPUa6pDNTk/+t0OO0nC/UTtBwLB41d4inuAUA3i/ALrNyoJVcBnAmEQW
ptbcNp5fxEUJjnOxnedyZEuEBxWRieZFQnkRdF269oPUdBParg+87IzqdHaKxl2n
dr/qOosfc1UCFiwPtg2/anKbINNtu8Ap0+QFi9EApo0uEJBjvpJGpwaahZs+kd+B
jpVBF5GGWM1/YNLTgtYwsTc5Va45amfjFqpznVsVI8vlo0WpkhxJDCStnV98X/zl
U//jCAN/OZXViOMONHJRsfKIXiaueEI0evS49Hal133muu2/4sWwCaPqXdbqiQBP
FfTw3d7PsFc0Spx7+eXmkc/N9RLhjEqofcixSePkcChX3JAWUjIRzHEEtg8y3395
rgWHFiVN0AvJ18/EvvY96FLnn7F7OKwVY7rNcY0ktlesr8Mgz97UYqeadkfpPtIj
JXpGBBfNdjBr3VH3O54j8CY0luuittmkpS/dqmY6Sv1xxw9xP1LzGqguau+1gVAh
iCTdfBrUMFsDBiWjVvc1/K17z/hKiqUt5Lf0vND2OLCmymigYVwOBGnwsr5/dRCs
fsNP6R4O9i3fe2t6Lm/7fQQ53XgbGEWK4oEtvOvlRgl4DpbvMF5gX/hOGV7lYz2x
yHJpxZy1bqLntUFEOrgKVaFvVG7mXqlQCPrJiZFM1lOAF+r+9PrtQx0QUpxtk6aL
N3xybFhuQF5kwnHyp4YBGo3o/Duef2g+ElSA/aqItIGRxCCkK3Wa/+B/amPC5U8P
DuMG+ug2/sg50yeDBrGvcKV0wsmrM6mrqZRKBFF9jzMELREwtXOo2pYxBRwAyK5B
NgE4pMwOMZdl+r92BbmKZN/XKb8PbT30Gzf23REiE7wPhgOVa310Mp+AZSaO0Luq
a/gOJhHZ1r6FU9fVk71Qm3gvgMoq/ekRti5g8zXccEIZ2Pn1pkrPo+8yPHZhdqwf
CFY7CVMhchrIT3vaS35w+6z1ForgLFukJcOBLOpejdXYiJGNBlUcdbnx3o1UI/ii
US33c7o0GZ9vXiPrlVxuhoiof8Kz7HGDOowYJK0g8Sv/y3TRVTF3aYhkdlIP/qk4
/mWdLnwP+RqlpGvXXY4KM55roHpGQk3bQVdSbFsS2045bi7lZil7FHvVkD0mMrgB
LgIf/GxO79+1rhJYimjWfc9tA0JVgDv9lNLdON/bLhTMkK/aIwoHW8jL4kG23wr4
aNXG49BD/4MfX5bTt+CromE07FXTDFdl9twWI7LJd3JtWxezyMVU7SzBrzrWQPHo
SF786JJQS56uGC3ZOa8VNS36oesto/ni2Lz6vQ2i/HceRpUk8K5IaqABAo6XCcL7
e1ga/r4MnMFSVxixl/lzlKbuVV5bFk/EEbOdO2olmEUG0s4ORjaFLfvg3yfiIzVs
AX9cK5WLtAdeq7jwkS5+Fsha8e2+8e0RPWDQKcLYQIEFJKlCAG3vr3EaGFezvR7b
Oac/pmP8vpBwAN5JO7Y0WJTPCT4D9CDKWkTAmegTF2O7O8PurufYcbmOCbJb4VBz
dWebQvgCci61VmrX1BEQJn1Zkr47krKhVDWb1wUKjnguMm8NIMHkrf5NJCh8SaLi
oXxGe35t0WRM9vTk4ib++v6lT2dZEdLQPJHbFOAbN04X6F+7qBQN9+pUQAVC/+wl
ceDc9168T1JKvtccXulE7ufyjx4Ge9d1VcBaC/NPXmC12tvWWbnKfv63urevc98C
JRNidyrjKP/2AAUbASkDlfgam2EnevDkrJnJwBMMrhTjYdIsHRequWwKZUu8k1bF
0z/xDjO/k6xRdSmZze2lIrdPfrmqN57VcG/g5iJZsV/KXZ/ybF/O5HyxaR9bTmnM
Ax5eZgiVF3aZ/0D9+VyR0WiA4q9g7BFfASetNxy0qmLg4qNXRU3At3vwq+iYkgrv
6N5aN6/WiZxYMwQV3UKeTS3POqzhnOM07fxS3kX7PzZSLaRQwEPJ7ew2neVs2QSd
io6N54SSSED2XDHjiitWh5WSOQ2eCBMokvxJNrkm/elZtveo50XN8rjUSgiihXTg
ASHHc3kXEK4PD8kcmcm3U5FctDtXf/cMP9QxYAB58DRvkj5I/+3w2Zlp8pN/lFHh
PSEE2GPmDdnFiNy4ZXV0pLQ6xkWhDDnmL56F6soFRtkcAu5K422KwoPUQBFinTpD
ZSL1ptGejE5ptMQNDHDgGSrQoAMNqaEhIMJ3JS2Zi4WO/jvs6uKcDu1Oz/lf3jAJ
Wlmt4weag+MOZ/EroAlbUES2qvzKN6lXOzR4tYeGr8RDOsJ8uvBTx8/2OBseuNCo
syMtDfCz8nMmFbVgf5Eaciy/gDWq81yFJZlaLc6dANVPhtxobsTDX9A9DW64WbFY
c/p3HHVzYWeGwTdBYUcWUWNhDdVpWQpGYUm0RJLABebwjF0wURS+WYvOeZ9MsdVz
6mo1xh1dxN0rROxVJ1dC6q33HkOr5GxiuDnzAV7iGpcTzQzs/tsNLeSG5yhYQlCS
k/yCELMEx9DBclkOz1Jn/NyswSC5rBQRegfFh4UCH71moWgrjxHGh4Zpsf7OqlgP
opt8fZAlmmL/JPta1Qq5j3EfkRAQ67QQrYmEasB54/cIArk9ebvy1Gg7I4eAoRLj
MaUs4EjM80mvzpvzL93ugn9ebsKiUVeAwwGHwqM0qX9ED2UcHqJWagYoxbNBEbpa
WOunDGcAkfOG+kC4xF70YmUwH+CYJU/uvnba2vQFeu0wEtvQjPojxzNy098IcGyg
AuTKlfh07FFolKzEdH4FlAAWLsBlLCQt4F6Bntt0ef2ar0QI7j/srlbsAFGoTTwb
eRFJLJ1HTiDEdMtxgbHUT+DKqtiQ4q1cwG+dh6hFYVv8CHGuycUTbxqXOjcZrDZN
yosFyfOhHcql02B9cmhMYTTbwCoKC9F5ioa1eZk9659vbsBkP3IepyGskxZu0qti
dE8OfWcWU/OuOqlsQ8sQSUzGjxbMerqMUkC/4ccYEgSAzoFRUeBhQh/zcW6GlMrH
TYPhSY2PayX3ouVxiXEU9RlgBn3yJCZh8rGBI7RXyGyOb8hNTmBQVPwARvrYCA1W
FvXOQi+esqYlHqydjiTQ7AV5hqVwbLncIQnzFcQVQcuB6tVcu0zAHHwem2luzRcr
Pv0KlBIrppPYFSaAoRXENsu7fpn9wLBWoQxOepDQmoCXLveRHCF+M6Tjll5MtwxR
RncWTqIfHUFNjKKlSglwZHQAgkbsftHMstOUkU0QowsDH0GcI8x1OHRUSByKvBsm
SpjsJ5d16z2HFI2PGX76B3H33S3YSgTyB5sFVpdhjxXlwuqc6Lo1s8tBrUmN3ptr
jH4Ucr0ESpRF8YPjkdOspz7unl2z0TOgpDSSIs8tkbWipd3Mm3g1aD5kDeL8B8vR
+NuibiFB4GdRYkuBKJMSvlnPQyq6H9YU3IC8zTNn5cBIFdA9z7/+1vnLSfRqPyYt
D0RQmJUkPiP1HJHQMqLapFJBEoGHe6kM7I6pSt0xOFEuqV7tIAK3fQaXytlA3Lus
lOr6DCma29bRG/g3xov8pFKqPUfrNro6IbABnih/um37BpbtRXBZHhLau6rcLG2n
CX2ZJOqjp8KQ/1qTnICxIdhqKJjzVU1tyA7yWLZf//UApmP7vtPwHEsbdnjSvZ8X
YG2aA03PxsOYYliB/7/UFZ1s0XdvjHqYdJl+divraHn0XtDzb8kC02Ed6xrdBvVz
+5OdLPL4S/WEhaPgW2GzPKym3BRTU1Ec/9StQYn5uMRkyL9Y7zoGLC2jcYjnqPwP
dNQk98YM28VZ0duW5Wg0wOSL1rx9+YthanOJTrOLE+QkvrNdOOtFMJATewkvvTZP
PhO19cgHi4IVCaGmLMEvtYpDFl3DOM08ateCSKI3UGOwkq+F965N1n6NRWBBUmyx
PAaPdBlBNThzUERbvFDnaNJFPjOQdgYW0rbmrRcMZ3HnECkrckbgSj9w5ldoFgof
9Fai7I7/laPmH08Pf+2FTc61PXchlV/elchjjxYkmIPD1BfmZFAswk/nj8aq/KlG
+MtFlCWN9AvDKJPcYs3oyorkaC2+ZFg6NmcT4nhU2zb9tgCH0X98GKh6odH/RY+7
alPlQnxXtk6y4W+vHxDqH+NPmDfTIH85PLhcoVyfCKvCnZIx9B9fkZf0/p1Z/j53
tYzjy7FAlDYRhc6HGCYYPiYDNyNpowdFnNfBvUc+AlSMHqazANx4gkC1Cm3QE1qC
wV/2lYjLyqVXrrkg7VXPICKG66J+fT769cVJ6rRKVj0pEDldIO5igAegZoQeiOTi
ggz7Fh2Zgdk7zHf96xpA0ViZaJj8JnALDW1c1jZog7o+YGuMuFFkoy3/rtiydlwM
XkKF+9exemnFNu9wFqBhwcQAf7433Eo9PrnfejCXJRCsNiQ+ZjX0infZZyLdXaTc
ZKXQ0YebO1AZgnl8X8KciKUFg2oyC7OzaAXbdPJh0ZHBIEaUQhpabDLOV4OltjTH
kSYqJj+H2UJt4EtyDDPavA30ZcwKCL3cMI9tBpak0w1xQegplViHZo2dHIhlUB55
EL290rV7mdP6dgHh6+f7xmYKKEK4YhzHMgSCjyqcFrtYMXo4m0sl6M87wBMldCM/
p3ujpZSn870or0IWKrPNsrzXskTt3wEsI7iq2Z7thlQ8LG2+CEOSC5JgkrqXkr10
NfPgnUh6NyNEVZHOurjx3aQmlZ3bbW94Ub4ZB9apaFL/N5IpcxVgYZejVCZoku+E
CCgMB1pbXD+yAyAgdrSMLVYnRMNN+BKdC1tkyLkjqyqnJsoUfrmHsoWxYF7n1rqz
BZfzPwsqGuo/61QgKdpLMhfSgNHzKd4RWQ9tlqbOTJIe794+JqXwW29P5PV4T120
EcD31KuWGWain8ozPZjPD0mUUJNVwVxCKbNic0JssfAuvbMRcqZrZbWgqFZOHHlf
ZQxnQLnuJXJnQKSoInWl23hvRmOLQz8D/49ODaJOnf4rvpeYcXVuGA4UCa4Z+dGQ
TufItABApXxQ5VR7qWgjS5jlLfcqh/G9z3Xkcs+RpYC2k6jcD2Bdv2aWG9yFI2Gm
v10XkHo1khiif+tT6RMmcn0relMnQ9ls3G+9ATeH0D1M7RAT8XkhexCpM+VHbbY3
eQCovd1deTfYx8+xHJ2hANxaTr6fmlbxEXrT+P0L3kkFC0lSf9iYVC/VlOYPzpZr
d3za3mbmHlLJGHNm3YT3jtd3hZxjxEENXwc97PNZqbQj6myLX8qekGYUYCiEQ6NM
g6LPL3hJ7O1aRrd7x37Wqwdp9MClGAvTRWxSgkVqsAc93AUsnLc6QoTowJ/o1Dwo
MNKfanH2vtTldrI4RVOjYg91nr8eQAvCtgtTCmaV/JGQKfEDaovZQQGuPTxbFpFs
+9YGzY7xNqvZJRcR0goLCv7h736GMVyE93QmOMyuvfevCRpkyoBS4NAL96ytwMj5
asaPbbM+O+qAhJYMpOUFWykDou+U0Ct+olPLwg/xMV0UQw7F5TFuXDF3KcAujUaz
iP5/8feaVCJULSxMrfim/a8c3GG3mrJdmEZR13TshEzvjsmawCA6tq3CjQ9T5xTv
IZ67cnr0dgsw8CS+3yIxT3BTtN+eX0Pes1aLeWLC6ygxedtKlhnCX0EDuTubxkt6
zf6THoUl5/s1LxY9wwK01Y25DhMwtcXRbJgewW3AQ4DsYSua3VrjxxVsMprXJN3O
hI4Ruc+4Ky6JSWxuQA2i1mF4CV0P062XKI7cSx0aR5bsq9pNyDjg2r13lgZKAJDu
zWfOc5wMwxXEYY8nrSeGu2pEYonPXk7T5BunCjdqSLMm1uc8IPLiFVUoTU8m0Lr7
+YWQ+Pvcw0J9dxTkm0RWdFvAznnFBZ80ZXMR49jIYmat9KkEujF/NkIacMGB6IeL
fFrjmxXHAvPnNA9KQnbXtn0jPIVYrtvJEiIM4XftT1J5HqAEatIE1IVsPvKK3bBj
GlS44KOLkrvcCey7ZEL9pXMXIvsj3aixFTqpFS7JnfZAq4zKTq/jAdQlwFOyHHwk
j5m7PP3rjcVOlBmCvtmfcrjOwiKuri81oyHchVkFEV2QX14E3QO+jMZHUgfOQOJX
q8WMygTCsJSqNznpqRXLfYQFnHVVKav0EE/UEqVyGOb2FuaGTW/ws1gBfO4DkRk5
W8Ck+2C8/4DdlT9bt8cViwtYJuv08gIkFflayaaRgaI1FqsGCA8GE3vm71rLjpM4
fMGBkmDNM+KmvWL0LeeIIhoj5gCxBBMScZNHbqSLs7LE+eYqge3X5Yho7mgGp+69
mbVf2pIt2YnARNuC9W7sZsk+8U2xuaNlr6U9BqTaGZp4r75YF0TNI6c0FL7la+VU
ooQAQt2wcXCr1d908OOd7ju1Rd+EA8lahXVRerAC6FEL6jet093V8bH991+bSVbr
BsglCvEZBGHSHJZ0qK3heKhu1G6f6a8KBRGujzJaSiOLQczScaNpfGAqvLVrORKH
c0IsMXYCjJ4Jq80FgxeQsI5dSwGIK0cN0Gr81V9aElOwCg2peHnGsUtF0280v5AX
Dy49EGXtyG52d13t9g9YmYOBK/mdgr/odtFO19JxnAGvMuYr+R4KF95Hvu+/OR8i
kHQpKbz5Stg3TxczpDCVdmlYkdWED+9ATWjk7eElZbWa7TrZhhAn1Tu21oD/pVt1
eTFmgr4UZuSwgj/9QlMy6IC53Ql5CtAAor95xwYqfocQwlxngOlo5YK1BHnPUG7v
guoAVkjVmxmFRkWHvEJ+XpsnnJuztJRMgxLGe86piu0Gh4H6uB82SFCNGt6Setya
l4iS01XlCDeRQVLKmG0T6jkPEkRMTm3ehcZAnZGcEtHXrn6KcMqQGn/rszNcXoiS
IE36DztTqfkwUsa6hgKRwK0VfsmPwladJ/SuVN6Fa94aogW1tvHRwPEgGkl8Um2y
bTKah8F9owIeIrnWBV4++jF91pQjLowFwX+SRuO54JcxhdtTskVnYCI5BUURQGqD
YagjwP/AZWHoB7eLy6segndGjDkINshOMBWVAiwyVsUtAiahIutovSW28gqfCKq5
7f6IWTEmVKMzWYAqZH19WLcOFqnww2ce+9hU1pDOYFrwXUiXEjdRcTdBcPuX9FWF
ZtuHBjHY+fFZpapyX3Sf2b5kO0Firzh41RKl7I13NbaeXzpHubP6ATThGUw7yKFG
UCYHp22Tk6hFSRsHqT/GdUu4UJh528iUcDaPShd6rnFewrOEj8eqDG34XPrYtzlB
PNJyMg13Sq6vXutqj66n8ol8jlEdGq+SzyAg7pKr8qChSpSxVZvnS3tTFWmoIQcl
V/0acuaJHgoYFAt1qvL3h9ygF12PSpts/yEsr3C5PRyFnRD+H95KBftJMKe5vW+2
dOOAy1gB5fV3bk70HhMw3UQ4PdDqn3HZoxu5m1XvSIKY+5vgfUQHMBNhsr1Qr3DO
ypFaGKIaBGiQ8UqrvanUWCkOPmERjdX+R3fVqik77znkXshtSZVAE8JWWhbOZ7pH
+1et843o5o9+m1/L19nvIAS2x6fuTGigL3YF7hA03VN/8YWEqdtOKuIJuf6fCbES
SFOMjYTZMwIazkIW/NFou3AN6P7NgL0HAkUDO+MKdLP/8fPhAFMS3W2b0gb1XSwT
A6KseOCzpje1g86CcX2RN+zpXSb9BFBcQFxnTivY50dCUjPWKH6KWHcsgtnO1u4h
Mb7fOa2y1Lm8YyukUlZdP2prCDJrhDagBvKMCU30vkMU41waX15Fa1Yop3pQbpk2
g4T4XhlKobCZxA/IcfBglEUml61BF9LplvqY4GYejMyjUOprkHs8bGHVZdJ1O1UE
+MyZ+5XqfTq7xeHkAx90HhkdP4qURS8mfrI7+mQ5WKO0G+piaypIukeO35JPYqy+
sOvqH7LcnDXM32c1bXmlMDUsMGKQse8C5HUrRzaw7MQMscoKmR07hbuWoN5kE55C
Zy3ClBsQQfz2njeYxTONZT7bGMrgVzrPpCIoP7+zPfE/fZLc9mxGQi/O41ThJOfn
YIZGbSQpX2Yb8iZ8AsiwMGdyEGLSNBItDj9ZE/jpw/HyFkbsFyZTeYrRQmlr3uVg
zjrHCTZtEgpx5w6MsZiRdCmVVX5Zh5MupcKi0udJBmJTZvRm8fCYuxXf3iN3vV7q
di2op0ZPcD89Fk4PFrlrsUXnax3zpGN6XLl8qZRN1oLHMoVg2N9/OHshpMi36O9c
pawkImQqzrB+3UZWqnUMPcdg+USiiKEkbqqL/8MqY6Qz687//kdNhJ9zngovXah3
468nj0yo7s+DVPppRpwEsgYE7CnA2rf4ZGH/CqLmlD8seuRR2EYejEqVO7Ll1LZY
igomR/cgcCMS0SOKCVYp45okkDIQvm3dkjebPm7XCvKiDRiAzrYz0BplWjT9e+Zh
TYd+QVPRVqfhYkRYFpNq0B+E8JBQk1P3EMQusymGdOMMZ9VOdhAG2od3B7HISUzH
TSYXUgBPNscg0ByyQdjNyfmda+w/yFVmw3W8kU5rRsEjyZJKClB2yK29v7ot5N7t
YNO1KdBqrWMmWUm6e9q5xNY6Uab+64Hyhm5QcYR3bJlGTJ3Z9maQDLBZfQfMJFeH
5vd97PIDwVi9FQvdGP+uIW7o58zmMLpMrNOft4hts14G0/NBQeVMmBfy2oVEomt2
Y6GrViGJQfco6+6OHssju/dpRAHPtiuALmuggUGHNRvCoFxYFTrQ3nh4nLYpfLIi
joDIlk27jYlUHkzz8k0S2a+3ffEDffOAjf9DRta3L/UIB3ZioL7/dX8GQqDbYjdf
EkGh2HtRnuJZwwZ6FsbaZhwxCf74TVsEJMtpdqEpuVyDLn1YPhp39qtvWQzZs8yI
Siu1NcyvVIs+2sLhLM20V4QaOO13c8mBSB92PPYDHTbV+lKitVI1kBLxFXjB1Hta
M6K7Cw9UEqX9sx4YS5TY0yF5LPRc/0Ju6OVdAPJ3xsScmXRnz7yUxFczlcTrjQs7
alBOj+sWuV5eqg2PdKAxaz96R5xhpIh72Nzl3lF1VjnNlQTmWhaliEQgeFERfjy3
KJzwPn0AcVW8kTuFZM9kDLCHEC2WMODMPnnuavl/vKfI9+O1rwFdCdUY40hblWmc
f6NsBLcZvUIsU5nOhSUfazvJJSFdABEYUpy4ezwVIYE1S/LsoSRp2N2EfX5tf31G
GJ9BKLXFlVD6ypLPssQZw76XeihFrVwC4THGnlu8xvH96Q7gWHHjVLCEucVKrts1
3DoeR+8WfOxmRplXuCVPz9ozPQZ+xYxqg7vqF9YmaFn/SboVO22YPNVWBmg3Br3u
Lkz6vkougWx41lvgSdSxg48NuSCvSH4DTVUXhw47y4+GtN5/eqZH8b8L3gyO44Uu
aqEw1WIChSqXvE84k5+nUm6U1KCxp7ppAbXEX2GuH5c2ejPiaF5UQZakRHIZhfVW
3qlsTczU4h70Lis2KvGXFvCKnKlo8ITvMnZyGEvX2+u02xSsjbx3z7nKs1rfXKNC
b8Wv/yMesOjkH9sV+Clb/xohZUKUHlpXEym3N10aXCkC3jqTRMa1iyahhrKMj7Qb
bZt2Kem7/bP8+Yoyy0kYEcmHRX2z+3qFEL7njmqJCSc9V2nCtUg8QZxvnEUNdXHM
G1HFIHz55M5B5r2qhK5qVONL7/EJd2vRZciYWkMUIViN+sOWJUJpr8n2CY4ywUSA
mfnpxZ5IOAP50O/RD3thjH8rlVKV8dAnUJfXRxfS2qg0l1Omzq2wSFtIqQVg/3I5
6jNPcAyMWDdssPpMDgSlJhQheWVfM0d41TJYYIjdHqxmQo/Dl7b096xlCblI0fHb
3FHGvfwMHr55qNlfm+w0gKcGWXjgIplcaSJRyrdLBIw3OV+038jW+dxl8P94VM57
vKdopcB0UH7C39qSVEUmEeORABCgSKkOSo306YlWtQKfHAtOwqhYaHq3McfWsovV
7z+4orxcw/mMreAZDm92yoZLhckK7gAZecG0ZC+b2okLbohAfUdhIvk0SGab2jLm
Dtxd+r7S/w8p5VYc+TpE1+RULjTElDyFOfKYhDeCkOfPjbm86oEYJ+V8xZmAVp/k
aLNhAiRAaAEvjxfHBRjXISLsRNvM6PUc6vXnDK8rqrzbrGLqBcMl4xr+ADLcUSIT
5KVD35g2eBfCko2hwuCgb7Qm7U0SJJP/sKWxnOvWAbTVaM2Y5f7LakOFYFtqkIO+
OeYgL9MQ1OOsHl+KCvdFPZTQlL3wT+kupcU9HUqJEgspRRPtJkYrfOFDn5fUiEPi
Nmy8i8MJDJhRfYGAWQev+qvHvPlY1Zew5YelkARmG+49qUdtBmhAPpgxGhbfRO4S
c+7CE8XzrP45sj/kq0p5/6qhTXcEhKRtSX788kj2Hl//q5WHqOIep52dpMFf0ARz
TulziPRjjLzyk4Oaar48+CseEi8Y2u01o7y39H+4KlW5GSuiP81Ux3RHkhcowp62
7pLC+4cB3u+nq0JnSwYY0aGBXEYu5i+0j7PZoTLb63AYL81aI+d1xsjLhinutbcG
oi5uvtz+pgnNVrvVAJnOk27My98sVjHttQB42zTiC6pf2gvh4+J/5P3M1WBo5fv0
tqKpFbd5zNDRNyYA6lBWAhlH5VpWE23QNQdridef9HGXgugUEJqgKYEL1yxlpbQ9
o6UeR8eJT5vMdWJ+j3R0uscMEGXEUm2elq7aEPoGFuvzZp9xjbOzqCR0BLyx73B0
78O/VoQg9pWYVyErYgJtZN5UHUBacxzacKkDD6ppKYkmSlnEsL4VZQ6DqiO5W7oB
50oBxUJWCDlnvxY3HiIbm76XOF/o4nHx89w4yfwIxcdE862tQy6Qe0vECepEKqc7
r3RNuPL6Tsv1ArUj+O5fARbGx0u12sz5jd/fUaNHeSgjQVi+oWiOFOcnKVRnrl8X
Ft59x7W5qBpCy5Q4VEdNjbZNYH4o7Fco0P0jWceQX5SyiLwKWGQfuYILe2lDwbaE
wlf9qOvBEy0+GqKHZQz77sr2KThU43Ui4JicgLm7/euMCgi9ZVLhSrj6LOhseax+
ok4oQHutljKHegvZ8d6FWY8UhSS1N1r3+AgU2vNid2BA+LzEex1zqFv3t2mcIQ4/
3t8dLUJPNSc/EgOTW+n4BmS0HPX0cIgY+eF/BMP8lMbN4bmbFMIMVwPj2loWd7KD
uFLwS//wa+2YdsLywA+XwFohZBSBpjYZnrRkSX4nfQ8ynBG+NVqKsOemtO0ipMCR
+C+O7U3U3ORQ3tU7qDpcWTAN0zvLzvdEAadxYi6lNICVyk/tC1ePqqgVzaW5dbsF
hK/K7il6Zu/i0LrUdxIuzgwAqlbRcTfEFnGvdyDwXj2elJLQIKfpY2rN67aQiegw
nuAJvFHBprnr8QusnYhBMVN1YKrOf3DZtjG1xxcORmyOLWg+kcutHERbvh/W1EnJ
LagNwqHC3y+VISck/tiNTjFJTlyTyeKkZjmVWdMp7/qDXKi2dghUGosREGYOpdPK
Eqm25z59VMxwod24grvzArfSKeYLnbbJJgBtlgVucZzeoc88b2ivtecgxwQ9iq+B
XeEIgalK6740TyLy9hi47054NYAbTUgt5yvefDX9aSe/fMFzIGL89AjwG4ZZ1mR6
LqqvNgoHLwQrKljgcjxmhacVHV3FttKOcNgULNXIBHQuYeWbq96XJv+U6Y4MMsFN
8sByLjiIGNFLP+itu0qqchEQGS/uVG9qMVhRAMOct/0cOpR/P3QGl6IyeoV+hVV3
lzkLTGRFWM8e4RK74e37eDbTCXGbPjZv7T36Fe7TOAD+Z/TKeE91q+oAFNLh95rj
rQK32HElIePBubJA9yhHp5Iwm9eF840wu8YzNs6/Ba/M9lIPfQBB+eyaJrweg+6n
9/Mi9epmziCr2TLmdUbKH03klFu/N67DKFulsD8RGBHo78HnEF4l3lImO3Cnglsn
4MW5Ugubd827H8OCX8P7vXgwtz8UBZOSkyuXC3ESIrwhEQzR5R2a0GDTqzAJUCjQ
ygD10B/eJBfiNW2Qm7r+GJs4xMaAVwWNJRFg6ba8Zb+avLUlhzvMITZYASI2R7MD
Wxgasng07vrfvqa/20VFqMtWzEsUx0P+ItyfQm1XVSm2YBdHubuGyBO2N65sZLA2
zGElwiNwNo5n77nYL/895ywnM2e2aBmWjRRe+P0PvD+VMANqYyvysXzsHqgiWNZK
i5rBUNJLuUlhaAI2JPlKDOHJIZXQB5OApNGQf4CfaBMetphDPn2zJqWkvFbvUoIp
t1i9InkHiBkczMobX+E91QwwoKa80EtlO9a1HfRE/j2Wq0sQ7hKnGfXfs1+KTTRp
dLRLSe0c4CuLoYldkA7QoKd+TedoLUgJDEJHXGJWFEl+r9G+vgkx3FMvbr+Fpzdh
210rmvhqUPxPqge64jElVl3PVAa57bOrNps7T/BqR4OHrUrPDGPZukFfZdpi74Db
sMNghfoi5u13N4VU8shP3RZXUMSYc8zVKodiGqJnqXc6kV4SMDa1ffuZhDk3OsnR
QvwRBWNA1NGtmAZ0Tm3eaKrowli03wQx+I9kNLbFZxR5CYMNb6KChur9TTwoKVx1
ZW+ajFcmYMSwdk7vv0n2gNMIYRF+Csn5infmkGWQFlv4bvJb4SRqFhbklyNLlmxt
JBlnXeVtZsL6WcunK3BFFeU6Qb1i0hVEnS84UV1LVx4JHyA3o4PX6uUiXgKQHvxt
6kBTIx92iLE0Sn0WlssVr9Te9dVjCDyDeeJTl+nsT0mCS09pfiZ5KEzHuARxHsvb
3cbF2bXGGb30HqE/wVTDiJGPuZcCeXkIZLe3ApWzCC9nh9w89rfP0IsaCMFW7CJP
KZsh7aVBrNO0vkIWYm2HHwnfySOPjV0jYzQ3X/0clyD3cJJOu2pa5o5ZdyOoIVz3
hl9ubftT+67Nj+Bp/t9IN7H/+LWj5+zL4Yr5hSV39QsZEXFjRhHeQQoYdRlKrpDy
PaMXNPo/SPu0jD9jP/AhssjGF2f7pE7yoqp8wNhngOCDXF4nVVCIuZ6S0cf4MsSC
9K1MIyHtqX8xI+kuyw6Dj7TcVXcJ/um51MK4GNRuPDEKj+M1SBmJU4yTinbVai9q
NQYAWXEq7X//4eprKDWE3d9qsODRZuLoQNzL96X2Q93xCqSfg8s9U/mIw3ozs/l6
BKazhbqzi2A5OurgG+LNG5GCd0B4mL+uxcBgYbBzISHpIUjtb5bQrmETLr8UK4Wq
pK+p+xv8qa7BBrASsX9ydvYUtlXYNMSo+fYL/wdHx4U04TFsdyVijhyqPlH6MoKK
FI3rejj4AqriJDGqaysatjdWoXN9Q/GLOpZzMv1Ge2MHf+ttFG7+NAk1A1EkMS02
L89hiyobeY8ct9mXk7F6jVUeMtXSs19s3XDJbV0OFZT6MzhoPqAJAyrY1tSfuOTx
Ga6NlNNytF1i7vOe74245Rp27JQAu7iwlU7EF4DnCxHBy8wlFDBID8hwnNsShNG3
cPWuWE9Sog3qxcEV5ZE1BLBOLkXuFR9CgEUfszefKKTnE8+o0k9bQWm6yyJ/Tuxh
md08DT8L0slqi3gxGGryblv8JZAfnh68r90Be8qATH/VuQO6ODhN5R4lx3k5mr7N
2SoBABTffKFu14B25S/SUFB55m0+RRKgo2iAsM1rwff8UqRgEllt7knRRCbBR04q
j8D3CsTJQfurpkrazFTMX93KOl1HxCHfjR/3zhWK5ffIeBscNoCaaixcm1z0oyjB
BGqzn95vV/Os7T72v5scw8uTh4g+G3DizUhtCz09i4R4dmIFYfZE1UMcNQQgTq7P
DJiWk3LlJzMulTmkYIYUxBJkRvlzv0hIRaGugGEVnmum9ucP78SNcP8H8iZsn019
AJmAmsxGC5FWU/ES85Su2tmaP3ZlYeLS2fkmNS8chsSaxzaj8RFNtdk2DTkSueFu
Fu6J2ravgHNbDFg/huCVSmoZgcAcECZULdcFlauU7Gfj3IKtIDc+LII2DnvyTJhQ
b6yUn27dpyR3GWGb2nIhbIh1Sp1nD9HtXFEWIR9E7V6cqBMgb/CdBd0OjTy8k8L1
6EpjtAMOcs+7XckKMThUaL+c0kYRz591+Tl3TESUXdbRO0/LZbTqtu9GPdMlv+o9
FgqKUVDidrGqubG4KBZH5+rFWFkg97tT1pf28YQ2NEhS30IUEP38n2rygmTX6bdm
UD6vyaY8+VhPSt5i/F9GVvb3YULOrpfzCXRppNCKi5ey/ltHf0Eb7fDK+jjioqSb
+E6xShcjoiy8jYPnGnJPUprV1RaeeRz4KelgWFFMYcP2MEhdlo+IH8uUGDOrieAq
hV1vkneSuPsRMoTlri7KvlRSp2ZSZstM1NLtl4f96OLWh7KlgVr+Nvs+LthUIn5f
8JjnoZ3BhxQcVZJfoUa5QsJDiFnFi8VMAXwh+OfCf+5+DtudKvy05ciIN9Zkg6SV
fgSaCRlF757sPT2mCpQCCaLNE1vLZmivIbCa4oozSfe/kp0ACjdKDBlw3o+inr++
QUyKJsM88NQzIzVBC8SU3UvZwQVhM4R0+8xrXkR/OYsSQSzSaeJ0YfXMMHekGxN2
dahJI58KUtsxq8JGWi5b0rqq4FXTk8s1PbzL8LsDeTNSH6klGbfsLtyyN6Px9yq3
taAbTEcfScx1uDfy3H+nMzppfC+kcPCtTAVY0kHM9lLSZic7exdyKuu1W++S0KrL
oZenKFGocYtmO6GVwa6AiGdgzNt/kH8wX+5rK5D5+vvkcsJ1nx5cVKGaCqLZDseA
elPVB+LYPm3psqaJNNtJnB4c2RUsybqSvqxqc5vOm2Iw6oB9BGf8tpWJdBfdeGfX
eeDWoqSbyOo45Jss9Coo+dgzkQsdVMxGCzzEMIeb3Rmkxbx8nXfXINFAe1GeyYmB
liafqWLBrRD/ZJw2BKSD4sYJoWGJ3O8ip2k1lleLyiZ7YHrHZ/gp68RWs22zJ3Y7
xQrd8FPtqOtgpBR/2ebcnENlAOuYmXh/+OgxkVA8Y5IQWjSruXA8PF05gdHSZg2+
9rkQRl20rA+boTVe1RmG8mnBJX5mdOCFWTF7eGx7ylM/xoFWwQM+A9M6Oxe7Kbyt
nHWQwG6F0sPfkC4ki62paZDY08HYLrI59w/oukV5d682zvCYcCaXXLZYQ6hueF4e
RMMg9tGJFfLMaynlkQv+APNcuBl2OjCK1fVDidvBOQrfa90jw7Qmn/cr977ahD54
7nnSO4FFD+g24GvxTkqhcUR07nzjN9HnaOcwD7h9Z7LJs/jwTIlRBHc+PelJwnl4
VteB63wYM1ocAD2VzcLR8I/3nIqMDV24QZKG6IiWVf+Jo9OjMo7hKdpLDHw3/w9C
iWgfn9RdECPRhR5YdwLlBih5rMQg766ju1hnqFnZ1i2FhEdiqpu/5BWbT3CJ672p
9iJ89DIZAgo4V0UhUX9Sqll5mYZeME/1Nw/AEDGhcWlcfgQ/uwGIjr11ByFrYU4u
abX5dY8Wv/wraObLeF8ME1RIB3rcUVHaurD1qUPWKn8D4y1Mnqq4+6cerHic29oo
KuQuQ84ps/ezUWiwpVN6IFP+2oiQYLL2h0zR98mhrQfavI1+4ieGA+hMStUi63Pz
ivYiitxvX7EZOfANUG2Hde0svf1fm29YyN7G1ZZXsotClQDAT5Cdkt0qvjWNtTRw
X5kbyw0jPpnf0M/+VKatGtwUoORkwJY7qRIuWQJZhuQCFun/0qXbUCrMtM6w0QW6
hMcGtEf3TBEBHdfYvE1gAALOtPrQ7EuYnsyYHynduyeUFV8p6e3fdKWPfd7Fy8AA
cl/vNZoMWJzHaF0xbN6zoqBP93HGtCLMjcrNC35me7CiRbB07+Pq405iz0rRcVAj
OpzPekoxmKvv9ClICoN586eNMNas6S7tqBHVRMkajpTPDoXSpWfGo0wffnt1BDPz
XYG0acwhcC+ylMRyQQWwV8P/ykaPMESmflS8BDzEM7ifCWwMZCDFXYOU5AAuMYk9
dO5foMVEah/ngtykSib1y3sOKy4zc8xcQrrZyO8zPz8Q5NJxi3Oc41qY+BU5Kh4o
pcyNF7WR6qkVNXggWgpt2y7gkN2eNBb2pfGXlcQJj1HcUbm4b+yNy7WCK027tUzp
CvalFEyosGrfX4sRD7iCFFRQ/XbxpKAknsPeAA2lTF0hN7wDMTrg6r4WrcRenNUb
SgfFz6h9fExuaDX482XqNQEZrBkcXM3NsBgq8wevtKznaEzBH9yd7rClWK6undkI
arvt8e8ivwfSRgQSkgKn+rh4F5s5qwvuMg/idGP5L1skZoAGkvHmhITIVO8SdBgZ
OhEWqvoYE+fDxkqW439g1CbEcsYBV0BAYdAaERF9UzMJ8Ph7RwGKEuzi2fduk1lA
HgLAaFXDguyPvdqlst0J76z6RLpnkYp3pugkRROQtKILNHs3pZVQVeIe++2vmV9x
GCd/tP4tcsdt5RpFXvwXzNyAb6qDGsPYN8eFxG9aDL8J4knm0VCyCswvLOhtxyJt
Ywrvb6009hr8g7K6C4pXmLY0itY2B8nYiqNcvN0sgyjY2ktv6bGPy8IvH31f6tFg
CPKm1DAsWTNOGMzsLg++K1KgS55HkIUJYNMGL44bYQvsZokUgr+/wpp0as9lrrNU
Q3WeI4cff6duod8KRpmT1v/EHVMWCmo+ULqXdaKgHj2gD1c9Be7jFzIaMUA09qO/
m3Ox6vZ6tNQtIBJxCbL4Z6ypeKTmUe9pNnqDje6Lys5zIRJCQ/ji4q9aKDM6GmtL
OYb5tdkMYnM/PKXAXZtWKtRa/Tw01r+aw6YaJtKOM80DWEOu+GLOWFqanZfVZAPn
BDvBeKkFk6oex/rw2I7rQYo9YNsEi3u9DjYo07oxoz17hG/yAZ2QLHGmYKSfmVke
9ZrVcXZi6HqIZcHglhS1HoedP09C5CS6vt4Gcg/WwfSXObuB5r9lmEX9ccs83y6h
1ZrhYXV4y9m6swW1ABLmjq9IxEDiMIMcRCkOJoECR+vyFCUVlXy+UCxGPwmH53Kr
UsDln8ykLwrYQcNNZqZgHlz9oeZISBfRg/1+1a4F46FlLrZh9UfgHX+5gftJ+Tjj
06LpV70UjhRIpRZKDJfaM0A/SBkCLS85EADUVgsitEQibkVOnt1bTf5Bld/VVZ40
ZmM2EYSIL1Mq8auUGx/j0rTGQ73lIyHnTkHoEz53/TZTqwGL4xyP7ujGLn38AAsJ
EqYFX33/qK1YXKKQWdO9Mxq/JZ9QQaCgF1VDD18cq/ku2SMBHRzaP+bGN/g+15A3
RASiPtjt0rUW1hzPngAI0r5Xyqiqc3N16oPzM6ZqMoiXpM8Yq1h+wInQFUpFUGq8
PbDzA3Mf0wRVEGQp/64zMFkwA6VC2/5RZXnkw71N33pTil1F2RHzCu4Cklk4oQza
wK3QLcT54F43wl1glJLS5yJ1aUJ30RP9DSozgThoJ0vb5zEB/fewyfMRKCTi5naj
30z1JpXR02OyX0DsY4hETqmmEhtTGrvn5+l5QOlSqo9tHAXZUHdMrA7VtTV/EDlp
n0e3uX1QJ7RsBV3Bb2fDOdFmA9TN3/zJ8x/91ZPePy4Viyf0b8c6RBIC68A0o+Oj
MhGq+vuIeTY9CtJksGMZv7ncclsJla5zpe5Yto05bm5QWyU7n4W+67/JxC3yYRRl
Q9fSkeOH/WZFiCewTDFGUOTDPmPithgSyt0/Xm+c5S91w7vkAMqZ6ecT846zfyiM
Fv+GtQEq+xCnzlVvwCcoqQL+sI3TTjzqb+90vliOpZENZZAP7rWus+kL5P8TJLUn
j1wA4IIdJ8dpjMoPyPxsuVrOaBlG7HQRUQ+90QLetapDwNPa07srRW5rL82+HEjM
iJD6g1owSth7yvT3Q94erfn/wmOecyTdxx0/fvYxvjfTNVmjAS6Ge0lUB9sg5K0s
P5xybHp591/hsrIV8Eijr4FbQwojFRVcXquAZdmDkT96gm6sKtgpGfJt8CvGBmqH
qySStBZB90o/HeD+8qxDaV9rzn79OW3CjciNSxlilGZad/hxVy4QWr7cWrKht/YR
F/71+RIzIz8nLSAxkc/SyDUYPH6WnFDeLwQpgcGw5ps0dUuumjUoVducwwPt7RQv
9HU+4OquP3AXzD7Vav1J3kToUHl5lgkxrdOA34XGpJhXrCcKNYTCo3fslp64kMGl
UJ7KfBvsgE6g0rVC98j/OpsQwNaiC2hJwpXa4iXSATtOj+OBihCC9VPcK/MiKEMm
HZP3TkQqcAzoIWug7Eylt86siTVZzdP1yPqchv4BnJ8dHYe/JCx7NGbuC5PgENID
Oa+p5MExqEGWmTYIYMeNqFfHUwewn3cQahK2/6HcaBNZJuTraOeN6xTn+4dRlCds
+rxbbkm73DAWbwds2vkmquF8bjg1hDacdSaE8Ma/E6whTWacy+So1TiBkojTjFEf
lnvdabH6raUWVSJmP0Sbehup6IoDm6lmBBYMPwzmSGvInhlF/z5uh6xzKVJTIf+R
X7pUnw0/27tzhubfDWj/+fH1oLHmBSlJZGya9+KA5w1yCFJ8dE2St33w2R/1Ms0K
OfsCUSOw0nM+Y2CPXCVKIfUkRTV9Ans/VUTthoSI6pmE1kp8cN7kuDpov1MEooxW
Pks7TtaAs+5YFnqx0MXLAm9/VbNSp4kRxgGYPszIDEFUI1CtA/k65FxxyjXc1/N5
k5NHQn7/siYZX8mN8yvsWhDWAVjopMlA8ulIMwV7XBT92holywq+k355/LkxZ2EU
RIqmn1txQfVjFPAigXXdAeWJa7PO9eiq+PP0B+incIL6Cx9eyo2yBc0Y7b6e9Kse
WJZpgbzSCG0L/Q81q9DAjFCy270yiOkX/M7UcvXxScvaHqpwVDSqtcpqF8n3nAII
fhmJyRA5rmOdiBCvqhf7CHbTf4uHprcn6VQ6/Rd6LhJpMBe5GNuTRqgiwnUt8Rq3
MrBOUyYyLxASYXTm69tMftLh5isId691GGe68eUECR5K57aIrhp9rwFFYNTwvpsF
YRa4aup5lBHwgK4awrArmuku46BYK+sV/bylZoM9XJDtful8cRzz5KESqjVwB2c0
POj6r7oy8hdvWO0S7LBlsVCE5rsdGoOitOj29RG38OQgaGPwPz+otCCNKoX/sKVf
sMEM1Zez/OOaJEEU4uouLZeXKroN2q7qcIFEmQiUSK+dMq41tNfvdgCXC5MCCnXz
TV1f3R2qJV4z8/YmqZ9NOXZSeCy6eMIHarp61GE7cK2MBQjSbWlPjwaAY1dFyt/+
ewRZ2bKZhPKpfIGucq6MM7uukiuZV5utLEd4bK1R05tYWa4X2d3Rb+YvtBnaSrRr
q8p0Yyl5bWunG4UkI+WLljSFE2y92jqWnCbiJOtodmq6hySdsf8jmFUwUQbmhyx5
CPlKyYsU+43SYtzeXYQwOM135gWtFeVGlAe4wclBjx6zP8YqaYdl2MXu0V19qiCH
M2hNcRmzFcpqDvxxFODvNS4WZuyCjS9LWvvj5I36dbfWYku+Crj5f2SDSfvmH4eY
9zoOsu1MZ/rqst7tiJavjTBtrmiQDxg7CdSx4Rc/3MmjXWegcaBFx25rbKzVqAUT
lYM2/MpdwrGmG9obc/5BT4MMCN88fh9O+kFXBET0kj/2hoyT5FnSKPXkBoktT5mt
1vgyq5LOm6TYA1Eb6xah6OuV3Csi9weix5ILuCBr+TYm27lz8X/3jdypILXFSMxr
wDyGV54FtJ6XzZSOOhnDcFD9XfxMDjCa4TC0v9ygjDMrE+xyPqY8eDNN2Uvxjdzq
WIT2/A+rknBHbc7Ytchn6lfgS6eThrH0y7a0ga7008WcrA+LZvYGLs/OE8MK49X2
09MdmdowLsfKlQ5R0XcqjVee7mV0ARFF6VqYjLnY/5kD+HRoAcwMhuA6kVWfvYZ6
W5hCyUHBdqbqlIyDMoUyHvUOIPcukYlglHw/ZbeWsWHqoP/BlQ1SWjq49PLd3apw
gryL5IjVxnM13FfZu1fd6mNjngWjuyi+CjqfX+gV76P66xWitst1w27DV6sNuu8k
OsJ93qdvtOgYgKq42L8EnUXrQm1pEkRiJgIlePqtBX2b+S142DONb87yqEH3PIaB
ZdmLTRHdwsYMhorhX2n0FgHEEW/XQ+yfQ7BoN8dQAgtrY+NGVoOecDyz2hsxRNm2
BxDlVV8bsU7heGVvKtZEThUAAholHALgHqeVof7KTZqO5JOOkfi0gIW4+soQcnp6
ZdZ/ARIC08B4VTorpTEiSTseANJzt9+XKCsGRKC2lpKqXuaUo8YmWuCQ61PnhGYq
PcS97Hl9UxRMrXiZOpA/0t88O43CZD3wwLqcW2qQutOH1y8qWT5GfT8Jjx0V2kZ6
3tfnTmwPMuyL2H4nnarxqthQkRW0iSQWE/R2qUdk2ofvvTgwjZslpckDrd/fF+Fb
37vZOxn+2FhH0TbcAU3CAUG8Vj3JfOdk2kKVQ4XTZH3l3qFghUh263WGAwzT/EiM
TrCc5SI2ZivZyAwOSubwqvtDLquQq07lwlEo74zlB5A9ljijqxUIuEcglBpStotG
NtB5ALTx7jf7KtsHqfDn8HDXQ+MxXRxpa0yAxSKNabxYlNKNT6tk6YjCEN99z1Qb
f4/WfCJyfYEPTpCJYOPPjHimeyan5xAu9WqoOUNe/jQetoh1WBDwGaK2+KtV8wL7
m4xxHK1yBKQoYGxuOVTygOvSLPVFYM3GZh1rtlSEajTFAa5ijH1g9uwS3rxIYaI1
FXgtT+IB+wA6hFavgCXqTSIXK1UQ5R7kEx9JpbHmobFMKSwgTnrTLuSEoB67iXJo
iPdwh9WJLvteQHrYslw6tY9HBxbNwj0a+O8gnuvJE7eqgE8zJ9dpfHoqMq5wsxPK
/OFPlG04EG4s7LDNfJyFazBw8UZjfJf/E1BQL1vNvIOEnBSrxvqkQFQ4PPMcP5Wb
v9LhoeKjTIsG2iLS91FwYzER++6O6CQQIAd3zibz8iaKC03h0Bw4XJpGdthNRBgl
raRDjt9cgYkovVCHFg8utxgBdViY4rQotqcWozx08n5cfflTU1hZN/bHXAB/xfCQ
K9fhO17RRiAy+Vodg551ApsHJdoSFQ6Ikf4Ik1j95LnXoulx7GteWgEWLQ4Vmfg8
N+pkH0HiURWvv6CR8sfSmhb3xhxezC8Y4+2md//C7Py42Rh9m86UUuBrkNalRNSR
2HAj/ZxwxCsp9viqq8uxg/+XBZx1bRSWoXXr3D/dvArrvPle82sJxK1fFHTVgqdj
mAPAIC0X7XQTknL78jvFt8UGtcRsdNvNxheXHNxVbM9EvT/LndFks6sTYCTc5/pr
jQhkSmuEN43D+VspERbi/TYreOxOld1LWBCs3wq6wX3nFximZOs+n6pLU/XprCP7
our4azJdCWvAqU2mPHgfIQFCHEbk4412itcyZo4xv86Axvzp3aXPHTAXOxT825Fc
9LM7+wSwKoogpCdxUS2JnbzyLbTwmy4/HNiL9mW7QU+b2brFY8OS0pvljlp4ekv4
nHgsXK0ToIKBNN3XTxmJkYBfqUmlFEf8wg8QnPf4wD8zBBJsuh7oN5Ibyk5BR1ST
Nw08NiyCxziFPhofCffZUVCRL3G8hoJpNw+yi79c4hHZ+QzpQrvCTGtEycFqihho
wSmsb2XJCVdz3rby1fC3bo/WK576THYWDEidYxZnEGdqEerf6FUqbJQD0to9G46+
dxfjS2nYVguLyPOIlgkPV0FNoVYnsnrUN+hP8oNE/6MR/cV9KCDmwk9kirEx6xfw
plySddJtpIepJKO6B6bPor53oPzsfx/OVbcr8hyPnzviBugTOHdNep3YL/VqVDmR
QE1K7yizfO7NOi8XhQKRKv8gl2H/OrJgGuwiIJ94a+aOAJsn9544h/keys+BVY38
k+j2ItZguzcw/u2XbNstCcpTK2ywwPA6KV39UAUOzSbPJA8NxtiIo/Q1Jzc+n0/I
Gjzsm42M+12NQfu4o1jnptjOvxCPEMQeqHR8Rd9weXQ/nYMHlnVIN5HNNUpVIZC6
lQi4LHfrSdqIbHBqoC8yut9c0sZ93EZiyH1Q22jeU+yGLVLa/9GKSiKO5c406ZoT
NCgj4SGcm9/XnPz9c+efGN8LO5cljY4z9Is8N8GYUeNSfb0lDlNi4EYsy+B9vy1L
n9z29hGUigiDXpYxnFZfUNgvBegdVI3wMSsBCh3DHQMDYbsJg61HvSVncJbB2sBz
oLBUS8udK2W4DjMs+vYH8umx9JX4vpOHbgvJmic2+TlgdKqaQprPyeIo1gs1kjNM
dprlJ8X9Ed9JOcQsJJFniDIS7jZU+4J7ds/uoSABSPET4Rj9K+0iiVVEwC1BQFaW
V8L14XAX1mwnG0Xw/q0YNKhVIJFfXEQiSDXorVslM8PxlORTYwErufcR6iCYHftc
Lc0KnPWcnfO3YQpnzEUZuU91A50zZj4DLSYLfRleku3wCHVYRCRxZUG35ifXtAKn
osR3TeRaN3N9GHHCw9Mduq5Z9YRMf6LTHzXDalRBsgd297Ak1B84qlp36d2jVug/
Rx1UMr1vgvi3Ym0OQTa8dr2JjIw9sNsOFJRgVwYm+d+SzWACNNnvtkRkNreOcBF6
grGHcIdoHkAIsIhEXz1Fq+uT96I0eqoivXcLXP9lJKIw5Bgj5sMmTeYUTlFMFb0N
L/YyDkcnBwR7YWgPhtS2PjeFdpSv5FmIrs1ykdGrSU0y8r7rbhBNTVYxAe474d6F
rYXDxdULdCmyKt+jkueTgESOVKnGRzXcBQThwsnILU9CiVstQbvPfFKg6Ni/6657
IdmkGwx0AxY6HXHKrirFjxLJDsXFHKUIoUNZK75Uwpmb4/hXXp+hBS5+Lr92ZpkG
0lCtCCKeZBdtTW1LQ2cH6pdt+0vR0H3SAmu+ROzWoz/vNQGdhOkEAzETHNaHjI8i
VsvFYm2DWnk66Dc+Zoupv8wxvDipNPY/76alsNw6JPjpoMN9s9aAaaecviN3/2CR
wMXfK6oAZNZiAKOlHuvQy/O6khRNmx3J17U4dS0OP5iiuRCQdOtHmipxXNW2sQGa
owG3Wo7tF3h934u2rBfHo1xxJl3UqYe/kRuHYAKR8kXit8gstxJSZyaFQuv3dIgq
lEGAibJVe9huQXPWO/rZYFnYC784lc7wofGnX/GzzCJ8tTGykyIsnTa3k28sgA+n
Luj+fCpS4eSyXj9AFmKFr/+wpCWwSge293II805eSLYewm4pDjACf+OwA+Lt7w/c
zDvv/JFephrXs6yb2w9DLQltrc0NklJTE40vjXZs3c07qxd2FMRgBhNtu2DTOEEr
b9rkUl141uz5T/j9sZO+qfNLk/DyV38uNfXD/9up84i/yLnsK9wwcwJB9dcnZS6W
aK1V1RzCbmpX2PtABVeusRQbzPoUbxEa5V07UeGyEzWtLYwJ5oC4uEfd15oQT7mg
XjW/5FiOjjAORjFJBzhgZIdx+d7KJCyj6SAbRsBGUHD3SWMfqDiuU/GJHB9NSW/M
sMq0I805xjdWo7zDm6OCv+0s/gX/ChPt3H5WANNVhwbLhecgbzEIRE7X1JBGM7mY
yh6eDEaOl4g/tEaPFNjOeg==
`protect end_protected