`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
ddtXksX2+yylW5zu6QL2Lhnb2d1sD00763mmSITNX595NcHTEkwn0zB1Dry37fOW
FufOhVzEJp80NC5qZ/+F0Vk7Ik02dIR0elf3clrjeJRK85K4e3Hoo4xn7YbFUIms
l/8VZSb14+JVGURjfswrIyCUotIzlzVYZ6gzoZwDXIi5gQIBf/gI+KxNXPaKV+PQ
Ufys/12rjO6aI/pPlqSm0hCvftmBcnezN2hk1UeXgOIuKZnogjOsf0iJVX2aOOWE
6pD/psybjbnsNB6kH5uFTA5frkzIzkzl5d9+YDm9OyC+k84E83I/7/j+rk4L2dah
QJOvksSIzN867/4Qt8qYTQ==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="MvBXkzurAa5VTw+1JJ70nePUfoQXBvZOku/SMmg4TwQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
oRtzZL4VJ4iwysPsC8SXYCzXS8Fw2gtZTOskLcDV+1B9Nzn1zTyNtlo6lNICRmmK
ZRVu2BmCc2G+fmzynYlNTnSa7C0Cuel6FYpxCBlOuk3OF2tzAmLAuDyOH3Z1Yjzk
a0aHuoCdIRKv7BrZCdALt03JeUmXKPdOmIlkVGFl8yw=
`protect rights_digest_method = "sha256"
`protect end_toolblock="Jn9CQpRhJt4rnzZPRk+dOpzAubz7omckX1MrFd4p81o="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 4128 )
`protect data_block
gD6l00tciPUa6pDNTk/+t0OO0nC/UTtBwLB41d4inuAUA3i/ALrNyoJVcBnAmEQW
ptbcNp5fxEUJjnOxnedyZEuEBxWRieZFQnkRdF269oM6TvXiIjcYTqyz2GO462ZH
m2uXuGm5N4ExnG3uINDVkkXopPu/22bIpECJdTvl8h4Kh1snWRMPfgegeJXvrG0+
9tWsdt+seAzyFZeP9Og2TVQ8fdfiKjU7mL/RkQSUpkGiI9Z+cVwZ0lHTGqX+nXZE
3vIP+A2qEUrlVv94xEwKpieGkfPElohaYIapCJkXF+rLeInn9/Ue/m6lOQS33Awx
QOSXQrapqjeUkfKK3WgW9dXzeKOiogZ62KpNMb7nv0rG5vGrS4y/PWA8bkgdfKnh
Asc5qvLCWjcO1T11nvfXwiLEzWkOZY31zxfbalwDg6hJ54TKW3/kyQyDnfopt6wW
ToVcYJ1O3S8t4NWi4hmMYvUHL68p7omsXQ9cRTV2+I2pQ235uBHvuraPQqwXKUlv
PqYKht45CMGcX8JwsmfEk/5Qh4jOxNq0mfGP+xujG/cr+UG+fGY6y6uartp/bjFq
vlURNM6jLNRMhyNbN9600ytI30XpJ5Ll2lZtXwKjz7ryOYqL9BMLMuoGlnYo6uJW
+v/bQNpp34PP4ij+ElMjulCsjZsVxpl1FhOcix73uarpMaxExV5jgpCmrdCTHxUT
376oWDqiH1C/m2LV2hoZDSWs2yuQmST+z07u57R2a402tAnayGSWsy/F3ecfPG/8
MFfbQYi6WOLULZh7OTb0OSpH1e+h8w7BGfLE3ZVqKf4E6st7DhU2JejZkrO5l7Tr
yKYjbU12k71FA9ODWn6TwQXkgeMO4CN92E+PsR1/XzCTskhMxM08mp5xMJaYNa+k
TTw1xiEuYQ9rifn5BhNVpSBXdD7UQHKtZ3d6JDCwvpFFMdqgxcWOynNqLdlPzCZP
9zwDHloSbw52vX/qu2mj6H+DPIsJrHVcEgpqTreZhI/7FQnOd88nESdz2J/e8gI3
8F3j5J6UDleQNF6nz+Pc0kdktwxZb2AFM9SGhnl5eqi4NWuNMCWf6wtocjwNGhbM
S7pNaN4n+Q9GdC6uuvd1+BNoHXEaBVuA/Ykk5emLR7PBvHuq4H5W7/Oe7ZsfQA+k
PWBvh7nP3XGB5eOCT32DVRrofZ3o/i6sAIL0aP4XUrikhozKNPIN1UY9oSXx4CR6
FSHqKwC8+a++fxKn4SYiHXlqAHW48S+1u1svuNcjs1Xp86/GtCrDxOE0ufTSiX13
ukK7WYFLdryKCUy4t+8J5ppTHqzIpzCuvN/JSBqDgEQEgPnnqR9Z2fjHbGy6KhVR
Xg6Z4nqczNyItxHh7R22TWGNy/QKDJ+TnYX2hknsBEUP9FXQe6Ssf6OaH9xth+PV
GDNq87tXNNyKScruqak3ML/wUnAZNsrPzWjZa5Aic9Jjc7W1iD+t3LX+NQ8cC6J+
LDo9OXnuxhirUHBUSqQeeVZf+nz+mUVWPnOLSdZwzZ7gRX731D64qXofgMs6nOg9
/OukFqU20ufs4juu6nwznGpjsQb1Ji2xA+1LLIC8nIqJxiPoRtEWK6rd7t3aR5gF
7VC5FZkbWUszI4ZSlqgCYfhrB5gA8Us71KG7HNFGH3jDwsyqM08ICMBkOxRMevbR
H0jKDDGfFTo/FwQYWMSkRqGZac8333jLgKLGFZN5L3F2nU98mKSKXGH1vxQq8lle
NTF0BkJhWHfagmVavbbJzBrUC8GaIjS9fT6zL8cKOZQRzUy6YOji309gG5wh/NmI
1vfqIbws/0fRVWYb0NP2r9AQ+YcHBPBN1sksyd80UPr1Uhxvsy8sc21t0rbizEoA
zCdx3ScgWG/bi1Ewd8FJVOjv6+Mo75F2LMjI81kVQjGW0jiN0NDHHqQqWQZzdumS
hrB+rrNnFd6BfCl5kIxFgu2wNVZCQ6pMd5iA+ui5P47mvLXdsa0HFG8UCfaVqRt5
Y+8bHbzqvXEIv5KjjotGS/41YR2f0pEKFXHN3/gDHGbP/YWLYFPdS0YV55nxXN35
YgIp3XrIo6AzSRNhacEKe1i7x69n4iVLSWyVZwKKWORmVfL5R35GZ7pudGcHvVpy
40CLISKrvZUPxoVocUli3YaCGhwvecNIjBJDa/oO3W8Xk7/s2I7ptaEKnJV9/Sr2
O9AHVII2CplHzonJRJ6vgUCdodX2k2nuzcR9T8kezm/xxRTDrjZr5xAlca+BoOFc
dnXQsdy81FYQJzYZxppyyyK8op4v9oXjPy1FJGqJ+GWJGADnaiMH7bh6k0HBheNC
H0DbHxqrrrbge/xgpJOQ70lAQHFREDlGxlkfWfqtMq6TlpUOIzV2OX4k+kkR97UO
2tflWa+/pkRoTjL+O8WP4dRNFcrTJsnSm7l+7BTOvgJRpcP20NvBx8inDqeuMKE7
2L12QG+UbaCQYv81F3J7euNSe0/iuhS6v3NfG4o23DCB099Zy49ueD8iZ2jJEwi3
Dh2A/MS4WTahkkj08867GHujhhAP7Gg00avdXEvwOjDcNdoSKXaNEUY02uRWEaTA
kdATH99T5hXvp6GUU+B6psrSO0jFacN0uoW0WEWVA8bMB9Kn0dpOSC2DOl2gVlRx
O18FL20e57LjUrrbb8bv2SFasRKA/UHnYZbtfioBzPRtIGpfMN2K/RpjEX5IN1kE
CDmznfUR66qpoRV3pttLKBJGgKD6vk+hTmYP6+znmFNgVnAVhLnxXCrrS1uWapz/
dG1g4DSF/hlXRhQo7kIfVN/deGph/BgRdVvPEMmsf78yNXySH4YLpxHBR88qxFD0
BnqLkpOEngunLs6PY03FrCfSnXChjmWs77iEJ+L5wHDqjRYAqxh3GngpcZxrAwKa
/unVYSweXKY0BzSc2oqNyBBWzHayEHJWh0g2m8jiRMSizqvGOe8rMmTLZenWN1TA
Vd68NjRsGKIw4t+S4+SyJRfs/HSFM2cPxpBjnmlo684t5TBwGMrqDZ6LpeNt/ibv
zip53KxMySvFAgIw/OMuSA4lpkJ/fWTS+G/VisjHQ2GTgcDVsRuDxmZ8coiV8CtB
wFB9w1+9qiBaKTDc0iR1KM6iSpBIpnrwSI8wqzNADHANqPjN7Ql2iMSS6c1uTizi
LisrGHn+VXqGl1SECXyuXKLSt/8ewdyrhOQXIZlWt8mMFvyOV3fx6kPC+f6BOggC
U6iR4A95jW+xV1tCZwr80/EjhvOLhKuGus7kw1/cXvk1h3SMelCoetBFmT6pWcBu
PDvTqjgfQYPxOb69PZ7q9RH2oHpmkhx2ZEhStjM9enFBhN6sf6Xs3TbPARUPiHZF
tuOzZzghHJ5nOUAx9BJ+OXd9U9x3gMeI/n6ytohWzn+o8rTgkn4nKv8soV7iLT1m
oqaKxrHU6gKzby8P6mpZUR3kj4UQMBqarAJonwYz0KbdVXqQHIqeV7DfVvQFEU2c
6VXg6/E4ab6WbedYI5P0alu0eplKImgw82ZftcQC1Pnh36X50dcr+V/09XiUY9Kw
AlQNcRYZQzdy9ydZ2rtU8aak3qxhvkFWngIffqXfQROpeNPZjE3Kc9nLv0shBHMO
gp8wToJVXjF67TQ8ti1nk44S2DAIRA1Kq+1A5ydWJ+4eR8ZC2/A07heAuMp57KZB
NjLXtPZlSF4WhynLdqTqK3Lt3nuzQvLHPRYCumK4yVfNKc5iJZAX/N7k4NEju9Cl
14Zi3g8pfgOK3k5+auTbqvzrfhRyqGetfBF3gRuHfws2HVp+zWsLsTg7vHIC6rgN
y0qPS/ucm/YYe0VveZ/h4+rWxQUC6ettkBMAA+L9eH9ErDHqm2YmSG3m8kAnXAGm
g7Y4fUgv1pxeqHamnllv8N3GHlVYlmIgokHXv3WsLqPfEXs05/vZ+R/LDwOQHT9Q
EbBOLlQ4Yza+SqJHYpXiZcxewRYJ1RZtaYVjF93AJuiO/Xb1DmPpalg05f7cDN1M
eeAGJ3eJTdKNZ2EI2X4qQkfTgTW/wMo1Oz9++fwnu5jNkfymxQjDvPswEj0rKt0V
+zGSRjXtGn32qlnsBuFakPfHWfiHHZCAZqRqyXEe+m4LL+rnUa7MchNMD4+v+VkN
PgJFb76jyoIRYldvbc6MIifW68Zn8YZaGGIqEwxY7adWFRAv3+1S4t18VONE8tDd
4O84nqTLlDq0ZdTWekN9NmzayUB4uWYVYVUYYh4QgBc+Wxv+d9A1zOf46QGMFgha
adOGPBa7bJFRoaaf+3Y132AjaQdk4v94+rD8Mb9QH11Npr7rdO3oRG8/6m9maKU7
XVvf0a8zwR8aZVGx05xVPlUz6JDNZtB/t6vNBYTOPa4wezqcGLcO1OvU/6ztcvcW
JH1Bm1QgZ86S//QSQLkBeAFmt6wUGsq4nt55/7ZMnm0Ot0E3ksWBlmyVpnbfNziK
9UEzfiimmikpw14q0sPyprsGdznY2N47fP68CjF/0rROStkWtqRpxc6AvSTbkfpV
PMhIUa+g9xfPTM43uEKOyCjNlunC+9VSWskEs5wNM+P2sIqg2OOGw5VuryDFvvEH
g+gvUBceMWc24wccdGJGDofGOaOuMKyMLZrD5Ghk4XUoomi5CZREwrEHWJeH/t/w
vXIzN7nTowq5AlAZJugFP3ryR7Y/p3vNYkeFyyDB/JEHT6clmB5dVW/4WP9qt1vT
fvLgfimkSzT33sD/mHSXs/wbPGbRDZXcUJC16zr0By8w8LWO84e+7EsG3YguqNWz
i2ePvw/P0ao5n4qDDHNQNJxIPf5u0dh8WXqwPPo/B0IkgoxvmBS4Z46YiSvNA7lW
4RY++hRNAuwyTq+69HQViNwP+7xjYODchTkT1k/fke6ZujxhfyTVx3uzNuoo6OdM
98dmEjEx2LlO81ltCTvxohZ7KWhyv3NAxXMg9r6t217Fb6MEPTV+bBtWzTbRSDXg
t2o6LN/YPHV3fWgXUHMQ0Z522hHr9cpopidL2UUq9FUHcxszr33mn7OQ/GouIWgj
PwCj0w9RJpaIR5MyqlDptxUvhliK66MV3N0LrjQcdv35um38xBBOgK93JNTPdUo7
PI0lUarN6/ROsgCzld6Aq0l57hT6UaB9/Dl+61UbBs9blJh5M748qrj2E2fGqmH/
IoPSthYYldnBaw+aunkglIhjMuOc2tLbVdFPXVgOYARdV3YUCGZV+pik8Ka7s2h7
b6aL5CcVn85BF295STWaPsqgb4teFWRnApM1vFfkoepdpWEZVxA4KweEnBQyCLwF
cLuGB6tW4d6HJg65Wam3zE4x9sYGJf3FmNbe2hcJSEizlacFo6P9AL/zXylbBpSx
/JyEXAyebAVCOgbGlj7fYWgdoT71fOAGvjIxUFji1rxeUe+uaQXTfTAsWZIlXyY+
lF55W0pzwg3UIRJsc0lrdtZaTR33u/oSkC03caZLHXScQjy9ayciCu2G4JkPeKQa
2sVVgoQkyayivmd3sQZ4kYd19H0cR3TZFr8p00Nmb4HwO4c+uJZmD3Z3bQFkaY52
`protect end_protected