`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
ddtXksX2+yylW5zu6QL2Lhnb2d1sD00763mmSITNX595NcHTEkwn0zB1Dry37fOW
FufOhVzEJp80NC5qZ/+F0Vk7Ik02dIR0elf3clrjeJRK85K4e3Hoo4xn7YbFUIms
l/8VZSb14+JVGURjfswrIyCUotIzlzVYZ6gzoZwDXIi5gQIBf/gI+KxNXPaKV+PQ
Ufys/12rjO6aI/pPlqSm0hCvftmBcnezN2hk1UeXgOIuKZnogjOsf0iJVX2aOOWE
6pD/psybjbnsNB6kH5uFTA5frkzIzkzl5d9+YDm9OyC+k84E83I/7/j+rk4L2dah
QJOvksSIzN867/4Qt8qYTQ==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="MvBXkzurAa5VTw+1JJ70nePUfoQXBvZOku/SMmg4TwQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
oRtzZL4VJ4iwysPsC8SXYCzXS8Fw2gtZTOskLcDV+1B9Nzn1zTyNtlo6lNICRmmK
ZRVu2BmCc2G+fmzynYlNTnSa7C0Cuel6FYpxCBlOuk3OF2tzAmLAuDyOH3Z1Yjzk
a0aHuoCdIRKv7BrZCdALt03JeUmXKPdOmIlkVGFl8yw=
`protect rights_digest_method = "sha256"
`protect end_toolblock="Jn9CQpRhJt4rnzZPRk+dOpzAubz7omckX1MrFd4p81o="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 62320 )
`protect data_block
gD6l00tciPUa6pDNTk/+t0OO0nC/UTtBwLB41d4inuAUA3i/ALrNyoJVcBnAmEQW
ptbcNp5fxEUJjnOxnedyZEuEBxWRieZFQnkRdF269oPt1p2a3NMrBvKpNtsUQb92
yRE5YKhtm6cAvU1bZFqtKkV4yEDT/gCTGyXgTEhaGXRsP9oX1esR5NrnQSXM7PWv
uaLbg8gnARjocdAVW+YPMg8JZCONw2JatNYnj8TqlYpdF++iNycuYcoKhOYXlrYL
w9FRzyWuZiIy0m7LY1L/8bIL20k34HyqO53iNNFB034oIxIK8v71hdWE/OgpxNPW
/eHhCBSpkmyGq+/S583XxCszWs1hICLFvjDqiGmZtfwxgq1nv95247ENnyqGh7DT
VxAq+pacn4mVPYtgNCf2yBRTslfcbjkWWgpPcbPAOC/kOJgw0D45X7PyExOd+9ta
ZfxerzrBsBM8HkfKSQfkrs3D5/HLZacBU7OBnVbvYTK3bn4hG4zO2rO7XMST8DqT
6/SEP3MuxP5mi3JavSb2TwbfnNquzuI+LXtndKwtYjqMWTSTLtmaanRDK5Rdr73L
Bb6Z9OxXEIig638gFndeT7gGqG1nOUaYigs95jWTszc+r6aHODQKA8H6/54Pogc1
lmwC+5H7CKsERyGrFWrVkxo+0GyA+MVDoJKnIloOsYRzaunzWCbSKMacu2AicaQV
rqxfE7exyElbbOg4UCP7A6JAghVWR577IQPH2qZqjXUNuG9Q6mAaPGertEb5KNU/
TRCn9abp8phOQzBqYK4C8Xet+lL5WkWUAVZp+DPEv7alKAcsJoM4qMRxpcC5OC+2
XcYelcq26Q0RO9TF26yYZxwO2fdRu6JzF00MH3ikFZWjRA1606fPjyrTsJZcWVTO
houQFVO3UbaF9qRMDHMhWqQ2taZipz7XfotAfnUgVJyqZ7zMIdEVbEN2+CsOHUpd
RZOCQABNkeGF3UIOCDhpZ+Vtw0xmihEz2fAM8514B/v1l1oTnDnzikjuybCrdoFP
aY9tT5OSVwP/bToNa9mItVSWA3WT1b6sSEVQdfqjfXrRBbpyKaqkiYEAoh0geVVD
hbr6iMHF1jSKGfKbZDRWqT10h8YxxDVEAJR3jFUEqkfUb2CJbc12f+ChdFOoT40d
Jirrp4oMF8GTTF36inEY8krPrhVIZidYADKckSDgy/Pku+Nipk/pd0pnq4ZTzWdC
MUij3N3WzUHPXEaSsiEj7Njk/LaQEz85Ng2pOlwdbkRM0wXos6ycCFktFcHPqlje
kg4JmDCO3pRU61Zsh9WKq/NR8rOVeNJ5AGvt3X3g+4rXqcDsUWgEzCtW3McAWDwa
So/M//q9wsrLOuEE0b30Vp+EbghqsYHxDoLXqdXvZBXL8zwEobM2AI9JSS33jPXu
2XHJwCJlllvgg/iayVrJc0d/4b9xUR8PuTnZhXuGcGmERQTiOlMTBe3jIwaSP63N
W/s4gzJZdBdEmgroQ8mqLlw2QdVwxC/BGsT5T3ac2h4evadccdGLjkljCCMg3HDJ
1Vzke3g3rRlZWr88fM9L7UH3Vv+jU0NWX6LqK8gbb+oe9eyKRCKCKM1QuhhcPONK
Li3sEBQhzcapeTR8Dl4bgmyxw6VcV61grWmqVpWDNVWwtHSLI0BLTHDA6ym1IY9v
Zn1SftjJCJMa/EHeYMyfFswzwyGkdvuljnw0EGLHNEaAFCY7w2f3Bqt2g/jX1Ssh
rUGiSTPG5gsJYBf2vNscXHiJpDYWh+lXcUI2XLfsuHx/Ok7YKofeB+/VXk4z09B3
0U2/i7PNlsbwqn5EKkvKz8ThHQOYZaWkDEJnryljrYHsV9jioP0dRLLB6EB1QoUt
PSHGcminzKrJ7PFjq+WKOCkA1XbF0txacrXKW828e5GTsyZ4N9h21dr7YmxeMW4i
zUj4O6Bu3isi1PBpi6bRdaL9iPnYCn+5bd1f5bqMagqZXbL+k9nXDWuDl2mFFX5y
WOjid95Ui8szonactNWgHhHx9KMlKg3ekRvV6arpJhqKZwrx6pTc7K68eVFYqVvR
yYgkiTM447eOGQhDywccdaA2pKHdrO9AJ2ipDH+0O0iLw3uqoXY1niVAEOHXDUIz
4uZ29hg+n6PmfzrCrsX5za12Uv68EWNVaqId1wB3Lg1bMON0kfiWya4tRF4gsXgB
odLgYpWhm+Yf1QkfaC80BPu7wqjaE7kN+a9axfNHs1/0c+cVf75PYhFmdSU5AQNe
JQBwml2GrU5lbyQvcYlIgYi3K6+q3aL6t6Lrki0bi8QL9d4pDalg3ycEpkhbHrFi
SAct8fTAU0zSAA7ioW8myaFq0GWTHjdiHADjqPUyaIsDgbgaqKFWpi37AtaLF2N3
wOkEOdWLW1WMRLBLKbDm4yQlYs22WxOflHPrcqWtAdn+1AEJ4cV0/Dq+9pnZ4f7J
IyNEMJ6pkyDIuQwa1SsdjW4S3XDqRbKyGr9Y9F9mH3xyCtg8gHX2lJ4hfnmolXTu
WXf+o5rXvioGoNKkq5//0xpyO5OVvLZHhjnV5ZX+jbeAUZU8Br4kwQ6snCc6OAlj
jVSqkA9wYazHvh9alkflskNmdPIWbCD5HauSIojnM2SPRrPo4U2Qw+WWU6HSd8WK
Z27H+Snu+/OHkv1vk1+c17xU5IPWOnDT0G9eNDVINF0TlwFyubLHNQmrT1ujGsHI
OxICt3+qG+7afG8cJHG84AavKbXSGox7vvhqLtykLPnHN9r1tYeq93hsHvdst4Uc
JSPxOkn9L+h/EaxSeL+RgG1JlnQ4YnhfMxwAJVWv2uY8haX+uPf9bZiz76iRuchA
kgRk8IL010yO1mHjbrHjDcd8eS8Eyh0OxnrMfGPxBvOKj+E5FL8qA6ORC53F956t
ScnQWbKp1qT6E8IlnGLTZNgJi/1Pp9FWKPY9Ff86mD2eqglxQS0e1aEA9/l9GTrs
HU9BG3ypA7YsEBsNNEBSJcInrciM8dNp3JafBxOEYS5RIv5Lr7dmy9jMrlb1CTAG
rcN+5TyU6NCeZxj/5x0u/MCzxw5l7A4eBjrvczi3SPSwZt5Di+I27UytxqKzAZVP
L+dAAKfBGj4VaXtYNMem2grymK8ftbOQBd7STIt8V621USKq/jONflEVnRRDgsO3
RbvMXGGha2wZGvb+CB7H5wbIPRL7C6rvpyFjqVF578uNpI9Z1+YJHweARABCnQN+
ryTDop8KRdUM9Ut/wXAPaM8kRvzb+OdVBBCCBwWUOVTnEhR9HMBGwQK1TFHBdx8L
tz3YguwGGLq4MPuzx55JhIJ1C7D/JttpiNLG4QPU65O9Y9j1Vy9sUsgOOF/5aZKh
lUvHEVB67LrQrxgYW+YYwnf1HuojayduPmh0c6fuoTiROfRJqu8YkPm96L5HSlkX
2M9SM+RoPkR4IugJXfFO2tmEC2QpZMBXn4wT/aVoE637Np7Lkxg2RhYXJHCj3Jp0
kpoauh7JdyKW01ifWZNmyAncd6ktgIUz2qFqqQY7pQn9G3IzB1NUsVuKMKJDUOgW
vgD+hzkL5p5PvGdpjHHR5t0hrPePEnKvKCRBe/wVk764OkQLAxBS1aJjpIOBK+K6
rCYOp2x/f/OTMGPfzzcU8CS5h60se9W1l7b/aaQWtOTnvHVpELvk1A4zf/nEmLzD
lSYNYTTb/ljvcofguJHR22cBcvG7bMNXzOtz0vpO6DYETYSo06tvAhXcmpF1U6tj
1xdHNP5Hcqkn97TiSkIpez+klbNgjITiwprZeJK9PIW2wNpm9PYM1RF6E7QCYlCl
m3ko597SSuSyVGhSsxcsDD8wiG/NxMFL8vws6aCJtdyGGgG8sFWfiN8jngxqNrun
vsO9lc5SHh8jw1WIb7MlvLhhtcLYOwAZzuzm68hKPPirgE594D6TXXDP8nQr1BRX
PBNYW8P9Y5hXKxxv6qKiC0u2wJutxWep+2geyqO7AyUrzSmeCQgWQviY79bb5+Pp
eHhjkSBjuWiMNOCPWiA/TTvepLbCzhIB3riJmB9774NCbg/5NuLkfM9f9AiNg2wt
S5GM13kFla/V3y4IfMfwjGHCyqB16EoWFKwCiKjyUKPDW3+KdwWVguhYxvKdkin4
Z9C16Dv4ZKudxWHxrHPKw0G6oDGgGh+o1nIt1PwLRbyvtYhroFY/i7VJNbLNi5S0
zduyul+d1NXV7surPOmgJ8pD7WovqbR1afEUNfYp/CZGQ7p/SpP+QM91KWWghS6F
wE496DM0lJbwmhmgJeTDI+wFEVN5jRpwtNhz4iB2j1T4h5zo2wFMuaILIrkbMqPh
3PaZDwpvoi+d+7BPnewqGDFEVauUrV++c1J9KNf6pFSAjps6xCLsmSXCf8Ay0dOF
1dAqAN0yspbcgHXJRm0IzWS2QUN3H0jeER6OIairoZgO1aJM6oWU7BHENqEpecsf
1YC+GSmbEesBwZs+WmNglef1exgDjM3/tn3RJYwxZNQnGTUvBBB5fkyPZCqI0T3d
DwqSLXlwx44FAIej6YGnEI8W+CMMNSEMylciJR8tHo1mvLP7mQMVc95uj6vPpT8w
PQe6NcTkx9Sgcqix6gi/JnggrVPC+4Irl2lY+ezNgpLK6sc/TXzOU39V/n4Gc2Av
78w40T5MnUhOvxbcrEfKck1EXOQF32xMLsc9hm7rFeBi69tN0VvgmJwr7BteJDDG
kU81XZm4urfHCFoAGZpUTclGc2z4Y7iLR4WBs2OPAQ7dLwUtwaQoc1WmCV/UlD3p
8Mu4/HIOGF2vC7GlPLgYPt+c0wVSMfoaFKdW1Nf1hiacZQfrq0GTNgjqSBCKGMrG
7HkCdZn34bAZMTp/oOf8pYT4qJokaYTJ956e4N2FEoG7t9+ERwyZM3JoDKPldkcS
eb6Z963INiukQIV1CspUYHcS5z/YUM6fVDdh+XBi3XUuNn4QAuZTk3ef8K5QsQ0o
OmxQGed+ifKryNHoOaEHhVw/uNU1Qe2I0NSMhXIJFQDY120kmU5kCMuCC+tOG2NM
dCOiPM9l+HOq6zKr7EETR+rVsxzrw27x2VYI6aLZKvIWvmVcsSGGNXljf5Bs9fqv
EC8T6oUUFBiPDp50oM4cXq7Yan8nM7axjof/p9Rlh+xoH7vUrHB7sDHkXyVaHAF0
azs20UlJ8ZBNNqViA8nZJCJip50KR0mUYS9kyMA3RVVGmtKR6hqKyfuiQ1RBNoUN
OPFB9DwjvZBs/GxmJu4IG3m5EPK0nodjUXDJ6izjtr4BkeQ1H6la19iMNMryQpTN
nYhMBLGGG0CRz5UA5a5SZ0l9+mp4Hkbr6PzgrvYV8ZLJwm8B4uCL3HYPrz3j03y+
vCYujVjS4P7bsRQMEuOIqkfyWnggvG8M0H3s9bUgafrXPe3o09W4j1D3O9Ny+iZx
LFIavrowpe+qV0KwIaEfRkLVEKokL+EQVpJgz8RbOakNI0+yDAoR+JMMLiNWQ8Ly
n7YkMxq6lrP0Igf7Ajr8q77/G+Y1kHijL3mEErgtnTcJQo9H1/VeNzf22rcD2pgD
c/R0S5a3dvw0a2QgY7sDZr/fi5jGaV7oCfdrWDdaAihhha0CVVtEG03kBAyepW9W
H5jMVUEN9GkDEZlK8dG5Ky60mdYbVtY1aa/tPDk7ngcNlJNcicVO3ApS5X6o/HSk
floG+bNV7QGxZWx506ui/ZdEyCWYKpQHYFh7XmV9SwQkdYo8KKvNEaMDz8kc70vS
dSjMciVI5L5yre4k9A/0jdes4Sqx3Ln10aMUM03/ytWaFKJMUII/29Sgshsky7Cw
zeVVZJvRZvf29kSBwZWI6MP86fHLR9AgYfXc+y0b6ECJlh1qkG//ozH85wwXjMeL
9N/8Xqj+qb9ksnBwPTl4d8CYxeLE0rZ4lmzkqFQJoNBISblqwyCbwuoTurdEK+nU
JbUGHlq8xbHh4f3+07nPkAXcLD1+kBjQNeuuf4Ep8DfjTxhfVZMB4MK1KWJz8Jb2
P1ti6YHsg6U5uFtXjQWkmFAIHCeeDuqdeLUsOcNbpjKpgvXRwYK2n6Om1W/xt8e+
oFO6iWQvlkaweH5TkdsmpZMR85Fs/ZNgZtVvgG87FbzQ2tjhKRkax5CxxRyWxQ/w
aebtqYxNhYT+8bTC4TQOkvgr+CFLLL+qD2+PNYkjCm8xgLu4yA/J+SLtAxzePEJ4
9duv4r2CM00YnR61JA8P5XOmgHm+FMEi6DHrjUPqUaDuAPVXMjiw935Un8R7pudJ
N1avNpPown+3ibG1ezGa5PnaNyumF7BoOKno8QoGBbVyTo0aDBfYmc/pcoEdk7ps
0Kj1WZc3fJTyf4gY2PlMLiQ4gvURMTGPm2g8ROTbvtZGhfQtQuJ5kls41lzR/oux
RJa7VuAO+1BJ1SNeRyG7ml57XwHVdFZU/gjf8tlL8jzVhmT3IYsOfVvJXQcTuFgD
tb2U64fX+BspoRmvo/cpQH+e842E/ht333lbsU9bCVKrpIMfaxJPdVsmjXy0Vkch
3Yve58/rGJg1AwCmScoh0sGjlwa9zOy+UzedLsXSsVJ2DPVc3mDYDnRBnDHpzxjG
LC9qrLN7hwpv19iZDI1iNDpsmMOgXuQIRzsd84wdKrmiQm5hSOSv8V/wgPI3Weui
wUoCoIvjA1LgxPayTlOziq8fzk0WS8Z8/GWyPy4N2cBMXXbkinoyMlj2vLK5bfdX
aqX457H49inw3aORjOymLzk9UgAbqFGoCkvJmETUezmcucan4fVgImHrGM1NVdHD
uXZ6u7v7EsteLIe6XOFMLbRQThdaEH/TdVQqZvVayT/ODW7X/hsfnsyG+C/T36D7
ECkWlZq6EeyX7fqlQqIEgP/HPokFigOhbJlAYcqXoY6Q4PKaSwFIKy1DNpKVHFAg
F9FjVFaciDob0dnPmAS9MApooPw2tk2/pZ7m3XkYBaPq442+OMFAd9RBRejsjWwi
h4ygdDD8D3dszJe6vcd0DmsDYJMb49uL+5MAvmKKB6k4V2GP4OEPNHqfonMtYQmV
E2SiimgKUb6SwSHBTlAhCEr/BsHUTFzP3BW+0bO0N4XMAqEFP4iKne1O/mlBVQJr
XSH101P3nlLA+P6iqYFFoRxbKUUbbJYbV+d1gPVoj+UvYEnmXHPEipTbXDQe8++K
0lOal/02jI+wjCLtkJj2yOqkdQkd9mqyKHwT6lIorPDxaes5mwZkor7Eu4hEAzQb
hg50jNxDY6YLincnBCLW6O4I9aLirBi6zSv9VE2MzNe3wYYmOE6w+JUoV2mAIen3
1ctJObWuv8sW5s/UKV2Of3Nx7Pfw1lzEfGN63DRxmsQplHaQPecws//tTzW2rSQB
rx0gjS/hRNsI2sNNhaRllGThah2CxrJcgegt+931btJAdihi/TMHZVkZwDW6OroK
7xcjrUXrGx8IQTm3sdM8SoP8k9/Yw5rkDPu8l2Uu6VXE4AdimPKKb1pMJDWmgP1d
zMjiUgrz7sCP+jOaxC7E/MHdd+QQ2UY52f5msUP/BQKeVbB5sD3T1VSy5mWjVb3V
N/SvNLFzi7iL8aNnl+xBQLWoOsku5kIAjpPX4ixBWdMiiHbQh5KGI5DQf1HRtQGw
JRcTpvjDWlTR3UQldbY2s90zoDx60focTceXqkc4OrjCcLTIpVOvVnY8ipA1g91y
TQxRo4Mlzkxy0oHCeeBDE7sgqB+xidP5toqtSafR3dcdg+i7xecVLU08myVmU2ha
rDhWJO91FrTTIRs5c3x6PSSQxlmtvrIRZXPsOPR9sGfxMJPXSdFQdSB7CxcOnXFB
FSUD602qY59cPtSDfq9XhyCrjXMIDceeyFNRRc7K3HTDeZ4a/kKxJ6Qa3emN8KN4
6HwfKWU8Y82HkrC9NjTLJEfU6V+2fUgtnTe+Xy72Auh8u18N6N2mFiaEZu3tTh3r
/HyF0IGQpg7BYVEkKAAf7D5WSSY69Q6S8FibZXvKhao4bKoeinRFtwGxsOcXnMq1
qGtxvCodNEtYaQ/Sd4jkvmxk49X8pJwfct1qbHmkBy/FhUKJG9DFyRAkh1ecxM33
2iCv4BMqqWPoX7wWbcbCJoZNQgxrn0ManIBdOBoaxOP/a0zkwKSR6cUakNr95Rre
TKKbAa/B4X7OJqOlwFFwttZP56fCWdnSoFC+2HZ8Ed8zTZYKMJIMx9Qk8rcMK8la
a3LuBfGtAPMzw7TO9p7CoJKpIKW0s7WBOpT21FIbaK/7jh8MB9aHWCDBZaDP2i4O
VimgN0GLMZb9qYC+jx1rr8KZ3J7/bkLjaRvCmUfJp5xNMfCjZT5RNmvaR2DeO871
uuLVieixB0uzjgzDE4RrJMXo588MHqBmP11zr9hZwpGGvBO3N9CIkTEnG89LJJqE
37IC3dPhU4+phDTv8UDO+zOpfPNJM6ABrpECzYiKEkAG6DIieTHdpMyWU5ruiIYv
uSguoDEpOsoU7ixALAdMjLxjj7ZWjQGPmjgTnpmKe/zWeL91mUEB0jHqgXjsk+95
0MtpYAX8BCfwJ4FTGEnUse/UVOUQZo+woOaj4DWVuIjt1A9XiRb9WK20spk8DdlL
OK4JJw+PTNPWpFTZu+OdeyVslGvVSrzm5cm0EfVEWD7CThIPyB2WTMcPCkbt37jm
TMyzmAUrwdPjrL9gvji99yPY2Wc94mImvxjwHROnV7BV7VgMhdLSGBTB073iKt9Z
x/adnDC5M/Fb7Wxbd3kCzpwt5NgKcfGh2heeYJI+pT7vGSQk+nag8+C42h/1OCmO
29D3wAYXT1znWn2+p5qeNHo6pNK5HZRyzEdcpJ78IVAFhWT3f8+4hc5zkdUutC+0
fR8QZiaT1Dw1P8w4dP7trmPRyZBmMgKmiSrn3VwQCK6ewQb1CqmBUbV6kj1VqX6D
Fj5Obz97ig/OSH94ytAO79Lbxh3FOzfm+8uQSkN8J082D+0sNJJV5Dpda2rdwi5M
lgwULKnass0kguCOsVmvigvrEDuaMdMaAMQ/JlW6URB4MFnh1/0nNx0vHXcuJA7Y
kK+9NId83OIlmIBFEy6Pth9brrnBHbEZ+OUSUUPredEvG+zoaxxzaBH8HEBLzf0n
lB2nL/Cfzn+HFIQKtuKq6gqCVXccfXbd1G0Uc3k0+om4oi9ts1h2pMgQG9b+L9EI
9H5H61jXOEyxHZb0rIrFbL5XV8ihRcdWUez4NJ14nxRZT6vWNer2rSLiSkig/Lsn
7fuOUF1FDAu6cwa6ACOt/lCGwmind/l01Y2eCS1mYmDYUiW181m/5lVAwmJIr3kC
X3DkaUK4zByVAuAK3gyMD5oo6tRnrB/yGjmAyDejSDHVoTb3m0olgYY9/Lu4H3/n
3brpyyiGpEnaIhjyLWhmTNpcH3zjLxPW10OZTqnAmUwY0YVlI6hYeRSsHeSC+h5L
bmMdvl0QZpVWRtp18w0de3l8KWmKrdG29TPj00GTYq7WIABviCzynUm9dm3tfWEP
Xd6bicclFlqhu8NYNKps6poCqTaTNncvnayMC2NUZJyQgEzwKBd/2k6nM1+Vmwnn
ftbNacbA/5grCK70JjVKpUXi6FmdkJc0KKTt01JYXTU9aEI/217jXx4x5KuBCzNv
PUNZ6xPFz3N4PMDnYOQgN5XccQ05MRSpdTPuSlMsU05ksdwtjlE4ATJt0zaCZndm
G4p2W10ZagipxZmzoq2wfJokx8TVgH622Z0TAryb08kJd5FDBZEQ/EMDpYj9+sLf
rwi7DSc8XVYlttSbdUykTK6N+lD6UreUcYYIQATPH5jiWhzdW7Z7fuf9BZpmkOyZ
44m7e8Bo1++pfp2bUsQxadqkpGCIeVaxRcMfrg45fgy9gkN+Ypsja/gFT1lW7cnr
kd0OnQkSoE8WLfor40HJHiqHH56yWhMfFKf/ahGoa3SoRNwP8ygbY0LsGHMBl38O
ISweWNgABKcEJk0FP7hhPrkY8J5Wlpb+KsCrGrhtEkUbsa9/oLSyxoUB6ERxduho
mbqREoBI97bYkuFtAaC0EWnE3947pgDeiCK2BJRJmRQQp98OriTbL4gcWwXN3aP/
w2jxARmncqnvFTwUTibKa+x/n+sTxaLNZaNU3gAVaFn2uwkWUQGC7Wqv3UpRsJiU
auM1h0bkzxJOWNgkso6JrEa4VPctKHo57lQd4sswZfjsFrhskDNGHqT7yvKWIpIy
jebfwxFcgM19k4NEKy9hNBwzM/ly5RJNywZwA03EwHpbY8I+G8JGJOuJPxT0YnBt
ZdAOu226GIsLCpNuV5sX+dy7J4kMsnvcAyJ5LKWXzKOGgF16A8ZX/cEy57RyT7j6
D/sIC0RGurY6SPl26FsOZNhn342XazmX/+GiEAdfOK7khnRM2xHLnUKaenRIP+HP
agUmGspvzfJ1Bee7f2iwjpTkoTXprow+L9BVP2FFngdmVgFaWPGc/l4aECJ9DSeg
RUFBKiHJ4jRlGc4UxOyS7NHKmNwRiW6X+j0WBSD8Rk5IyqAL/A/c6IiT6YwUZ0r+
Z+ak8VHa4zENrYvJgQXIcwnklNdp9YmX8Qcyzz7l9ip+/7rfJdMBwgSlIjDBenBt
cAvMXj2p8wqz1cYzpogRXwUOHaZGziUpRN+q1stSEALdAp4uE7Y+O+tuf2btdGRr
ydoVKR4NrzYpW/efeIbHfxLLs2GGm8WzAbfZ951+hy0vENo6cnQsh+AnFTjfsmyh
OwGv/Q5k9oUvn3vLeqUfm9k8yVjvayWFB7lKR66aERWgkITjV9zNgU72sBy2PdzR
WjZzSibKrdHDffY/O/Uz6ruDyKG+v76XRZqSv4e+d49hngmjXZ9aRIN3w9Evuc3v
cWfioZgCfQdFUnl2+H1MfXgR4E8syasOEfVImQ6KTLaD1Q9QvccBN695/O9OB+56
8CrmnXJ3Zs4/fb6FIO+Inmm+DhbN4Fm4AmLkSawAru4ToJ/WOlwOfvpW/WaqqiS0
4+dZ5FEnKkzJXt8mEeX8+YaUjyM+jayRBy49hK13WK6eXGqIZcQIvLgB9536CrxL
g24jUeKeK4CFu+G1ErnHeV3ncRzOkequk0rp8MO/g/fIsqrAzaodF77+hPAqfhML
j6o4qUzkD38P8IdPNCb2NfQ1E2JYbTeWQ8jRkrfrX0rl7DHlk8vfOp+ewZWeXt58
O1Pgtq9I677XQk5FRYCq8qO/etcu7439FjhNuAN2kqzrvWuTmc7wVLbjlCgo2LBv
p6pN+gk/kq+Y3KlF73hAgwPFVszlSbQUK+Bw7qbacthLD4qcdEDxS84uA7NV3btd
OVTHVyqXzak/eHQHN+yittMqICZY6TrgW7onOsdYClR3n0WcxfbONOfVqcULYlGW
Ep1fg1TbshTml68UGae7fXALWzX6x1BtuF0k9u3qzUqCkkkF6pra3jY8mu1OnL3M
bt3SI5wkzMcecxB1RoQ63auUsqOkWcSKBwX1n7VmxNQLONwiiwY5IAcBvAFiPM5z
NE1xk/0uTtlnXC+jCgQQlqgzFHjq58UWDEbPT41ERA7cmgQJsIIXVBrg/0id/h3M
3hEsGHsjnLGTnkOJBG7neqazV/V8yJNpTLf6vcNiD5jSfj8+R8r84sfEJFhpTY97
Q+E35XIk56NDc6h5LLxfNU/+lG9W8xcJtmxoC/ZrXcsocmNThEA03YFoPTzjp5XM
2gsujdoq+Q+DkvJinnUCi7B31FSXDpk9qfCScRlet/qbBA9zdCxmt4XphQWeo1LR
w/PKKqq2H3zy3PkSDW7CrY3+vs30pR6/RkIOKfAH9Cncl3+msZLpSCEVw8qbBM+L
dOhVJV5LpGfUW6z7umpk/9nLpdAkksMCQI3bQ7VvP6pj74hMI2Xzl4nafRZhhLxm
meY8j0D5tsPpeIh7HlnUwEUO5ubtBTQ2JNChOTm+NzovcJ5KzeNjwaQfYdMy+EaZ
k+Nk5p4XWdMvyWPlc+tWPICeiHLetIRGpJKak7IYmSu76tRJ3ANiSpMLJB+uyl+s
Sd30Cvx4hcYoe5mJvWEPqDsJt+LTFho9ah68MJGNJRrpsptHH+QZ7+3j6r0dKoJr
jfwl4h3Qio2525CnWPKuIHcEAoWVmySYAUr/fEaFcwcGMfeFuv/eQWn0c0j9ETlA
oQLNvM6WUupXFEyM5CSTs3exmsbU2srGtPuBFU7PmpTAbzKPqmhCUpJ6Z4YO4zZU
AIhNv1R6a6gbM5885hgxq7qqLX+WxgrM27BUZwTtEyupzic8A2z1jzBiQniXmhzE
BAJFYUim/4WdlKkDqvqTXvokQZhw6ejOdp85wS7FiVp8TpCiHZQB0o3pJj8HAl1g
vMdtact1B/J1bOKUfKbBftRxEH/9wuz4A1TOXSO/bHNuorXg8hU0e+65Oj3v+/7D
LPUbqbWGG5w1zdQ3twcUcbyn8KfWWPxYBxTTPqQEPkyEMw9XFOM5ocKnSmggqRC/
Ezm3ZIIJe+3lv9Yn4UkqIbXaDcYIeopN3BMlBPfkvG5f9+5g6WtnqmFcWWUG2d7V
rz/A2gID3APm1Nwmj+LohhUQZ6bz2x2R4cVbf0mvttNmeXgfXqWcb3BM6R0bTyKT
1HEw4JTAaKm1M1Xe0hyJt8fxB1jKLx/6Nsind7NYuqSUzaFS4wRxQeOaZMPFv/wJ
okWWNHbpOK+OB8Jhhg5hztNbOYkkSkvKWHTalHrAaAba+KIXHsiA8SvKVhLi2fD0
6tfirsYUYIrn3+D0mIRKQH1yyiK1tabPicVmSwVBWTFP3Yhq2oFFalowMdfqE+wM
WTW1jqaaJMU9w0d+2HssYLZ1pUKeLH53Opy0uPVWeaetB4nhRWoX+5KspZEnI2Gd
oTK07Z5Nb30p5AUFp2S3whCkA3Cdbv5FYx87qTxy421B/Drv4fIaSIeR0bhs5ReD
l88BTfWl/CdrOEKDuye4e3nP6OKP3mJ0+19eXHm8/mreSN4DSEuYhBdjjuY4s9Hn
rpAaMgoNjmxo3R/zwgSRT68gmxaDeUj6k0OMK8O6vVppZIKrzv1ziXumDCLhsl2J
TIJgbhU4XVOb9LN+RtWYfRZvo6BzG8TIe5kCulQ3qM3BNTL8C0oxxKqWC3oc0zSD
jGGIaqMfvKq0xg3vd/m3/6cmNxXwzJzN9EZP6JENMjwTrR4AQwllkW4CVCwpgf0n
P3Iq+r4NqO4BahFiMFfoW0Zrmed438qCW0XhNLsvEU8bqvAsu4VK5hM7fixVHyBH
mYmeVeMpqY8Dt56hJBzygFQErvUnScGrKEUWGL+wQDUao+WaVDvvCEqCLHzTJHYW
mAQRnJmBGulMo4YIu+sYCzWiNnXnVIHI+/xBdP/+w1AQa5eHcH/tRH10diNfWyEN
h9C0WGemqrXtrS2f1dexb2pU41qJwM5mZzsjlcO/jplblhh2NbEYP/74PAihHNYI
vX9znJjzzk3SZahjhQjuLX38kLe10mfz3TxJoG06n21A1tu+TNfGISDqmNgOBNop
L05Th7tEhx9jHwZtubaiTZtRxwUzWcAyRIzdyT3BC/8IhZu5h3fWtvhdWjsmhCMF
VKdquZIAcfq7O71yT+cfvYDcQjohc1ROsjMGpvZw/GV6toiY0FUG5ESo935PM2gQ
MNjV7zJIKLh3Alv2GLPi/eyTjO9UXllN3W8Gq2MTTB/4XZLL+CMsyaI8ZkvN6Xhu
hxpEPiUBiIdQK++7HDJhYzT6I20ILoArzJGs0elqre4qyQM1vNPPIb66t5M59zpV
zVo30Z/0Yx5aCrAUFgbyqUixNU0hZ8qr2J6SrLjlXDH1PxW82Skp5VZc2xjG5K1l
kZbCkT/Bf8DaxdrpMWxEVwGXqKDzdm0MARHbSasUDcI/6KjdwKzJbgbbAquyl4yU
5JbAdkwenoQlJ+TrS0TntRlunR1L7MFooKletjKL38ua7y+QpnFX1m8W9vZiFlQp
WnG7Q3VLH2fsI849K5NzBtODkfiRhcSao0fP7QkG+vzX3f5FpJM5ctWa0d1awIru
8WyYRfrfLVy6nZFWYKa60OK1RvmxT4zjFZNiG9JMvrZwgsbHm4wy4PBmCYQpsdqh
pn0ESrAFY0bCo9hyEQtHLsPLE74wHNslX4UuG2XWhLF+9W8jktiIxIZvJziw4i26
gbgyxI6A2FX8iN10qXHWlsYWEEVGkDVbBQgyGYMVqg6ly57D226jWa9ZWxu01F7c
eYhI64jsoPy2P3E1fImVgnsPVn3fdGfOpkC58ldOfwyPVtDbETlRJ4RuDeUMkSbm
f8kUyUB3ufGxOzxZQFDYx5YT5BOUZbwk+Y0Uwb6L+sz8kXQoNQkTXXYwVgvUZ1p8
aPaeC059qGM5B6XinOg4W7B4u0DLrMVtsY6bM6E4x8n7jVhae7ZoOKiA3pS8Pr3u
MV02s9zT4nnjjewvu35YuPD+HySqM3slKZ9nXuDgQnEWiqnBbb2NiERu0S9XQ09a
Xr0H43TzsPLy11IQsam+uOcodsVbxnR4ngKf7NJ0oW+yGfPZma5BXwHvGXqpXSVY
VRmeEBBNXHtLInUriPNLiDxNmp+5F0tmo1X+YDHOI4PU3HdaLQoz1WzpbbPwvBQQ
QiHaGFmoD/fBT5JBPDKyK/yYoLvJkhPjWrtkE2ZDs0AZzEqylcNzhCI+psrlgS37
abURWyYWATXQ1RFRE78QcM3GQjqujHq2dbX8RIVC9ljmtuVLHZQKTKHLQ+t2qQTh
qXFYvY/ZHiRN5e+In3AT8C8+a4aTtkmBFsfd3Hzdv2fbcfbIh1khsG8bzk+6RV3n
kUyFkyF6hXaaoUoh6ATOX/Z/vCFjPDKAD/yUc4/rso68gYMWq8fJeCBwhoCdGy1s
Ugt1uxDTu6omvrHlnPfOjQ9vbW45zUQNLHWVquEn564Oa4J0NoAkptP9qI2PZBsd
+uNj8WvIx8c/s24PLsZL9XRHnIv7RagQICcJk0wg0S7gKrTkrlUnVPW8Asyp4JeG
vGzz67jlJzwzzSe5nfiR6b3lzDVLkApDxUDSpWoa/C+vuf79Jzbqnpyi1JxQ8taL
PlX/cnKXDof2Xlz48CoeTr6JrZp6GD+SFau7GI3CGx2m1ZER1g7TjezHIrfUs1C5
/GQj16G9aS9PMoHYFKr5jaktFyv/xdr9iLK+Y31NedtUTZRpyYqRuIfHPgKEKydy
7mR8YwRmQEJT5DI2u7q0Q2Kjfg/pV2ITn1E3PfzW+8Lm7c6SW0b+lcl3jvCl62Wi
HRneRLo13Y7RBHWbRl0EbYezVIp05fH2DQe0YWAjs/CuOWSa/tJRfBpUAjHHvvrQ
qhU336ICkM43HMq/tdq+LagtWw4fuA7oVPIPHiNNPULElKHpwRQRx9ZinJlYIIhh
tI6luii8zkHS66siSf5NyyN0k17wUCcjT785zdC/vPPDkdAXSyyNx6U+ayhKFRRC
L9ZSL6rWLVlI8noOv0un1y2qhKCCI2/fERzNd+FLCLgUpAcK+rt+VnoiE6vbn6Av
4R4mFrAeOKLLcyvv+dV10GYdcfHHpZy/8snt93qbD2yVbHBv170MX9I7MpWccot1
0QImxXGhCBGU4IcfgPQEKz+nbj/YODklVEpGQA3NX6El1QUeb4Q/n2mHxXoFIAGl
7qMMsBW7uvtJCwAjlmJElQO9xwt1aFRPkb0A3OIHeaanziwZyXmNZ+1ND6KztPEG
a93wBDn23DLR72rWmCJTRBsjkedE3NCrvyhAYHM0W/hoDy1abspyUY5r1c1j3E7U
vQpASWDaeFj/uvlijVU1bnuqTlEI0Eo5nDwa+CvyopX71K5Ct/0viRWYyV4IwVnT
55ZD/RBPL1BtscX6gwPYObfePBtoSPOhPDx6xhRu0iaKLYNqzjoxoy7GfsxDWrWe
zPyNS22TnjI0RRejIweWiGfeibHWp8I4gcbC3V+s2BnO82TlJRD+xB9s2QrAkQ9O
z5ziOpo9zkpojzR/ea4Zd3aXsvC1neBAUoZ5V184XAt/tDt7InF0vvcOqx977R5L
wLuCGcz7MbEVgQdFbb7xM/anqpZv5aIT3APxSHrloh2hnG3ICljRRawYTqvAnSDU
8C3S8C5+7S0NJz/sXoTt6RXXwnPoqP6vIowzZ4INISAyjlVHAgjSXdPYjVB0JFr8
GQQPoOijKVxgDbI++xkuMv9022x6X11OKq05PW94AFlKMACE5hCj/JSbOGeZssJn
umTF+Tjb4TdxJXyxjXIzDYI7s33v5NgtuyuYEJKxjv19nn9TXKAgFFkt57SQo64D
JinEU5yoRv2q6Vgl8ydESFjf1TQ3yxw8rTofVwA3C/oXbHCuXfKjUaad8/WqckN0
Xjfgga7qVAEKAu4gPGqCyuCX3K/unYoHvXsZaMMnE5JZ7US5taMNP1elljM4HQ2L
Zjho1lCoLLZIb00fkxerRXIJd4ctKM8lxcPZc8E6jiPiA9tg57EjcZvYnnpWg33H
t0rBq7+ZXyp++pINMC5AlGAQdorvDq4jNGrIfBJmxkFBBuRxlXgM2Nq4tOg4vUZ4
z2VIxJHLrmwQAkKWRHmh2fhVJjD69PW2qBiRaiM7ZGNo8UZagjZbKOoITnVeAmAY
e8RFW/wI2TrhnXIgBZUgoXNpSrn0cmDwxoHYC78JvcHsFmoKNTfnOwIvaCHZ1uyt
d/sph+dDmjKIYO0yWC3EFfF2qaTVkxD5lQ3wiQbWYkagHqr1bmYqGKt1g5S6oBaY
p3NqAhFUqfxfPHrdGTmF9BIz3DGYTLFkqdMn6KyWdGEHmaQFytLN6a6jU2scjlX8
nA5iKSFdVKow5SuaKujwr8hIhTe3uEu6+QNAvBqhl+frTVGVtjeceMYy10nGeuOL
KslukdtNJzl8GdPzS7yc28RlDJyKz7RxPrvhXjbEds6sWuj5qOIk+mQlPDE8zmMz
KdPeh3nCLtbp21Gi4jS/eKYqVVBRgZGekFEw3rnJZFPFubLhgcRi0Q2P/q/mOJOf
LET7QbTqNA5K2R9djuq12kOMH12iTFuy4w1c4A9GQL5klqtBshbxY/FgAjLYRqRc
mSbMZFTV4IOKxoGPA+5C0nV+vwt1JVIUgr7os2MYEsf/tGEBgZHFeOnCxcEM1o2N
y98aESgW1zWypu6PPHs3uvv1EAuk9PuvnKmlGRSD6Hw0wKLG3IU378m2eFiNiTiG
+4emqkSwGl4xQSciklZnzcwDl4+yG1vS2S70NkNZr1wP9LPW2BT8Y8gS0x2wfmqp
1xgnJ8djYyoNJgUnpYlRd/T9sXLhCGIXQPeBhHG2iBTZBIbrUgwY79B7VOEEo6Dv
Fm2+S7p3iwI9udmlUVkkeXOmcgyLoEOsT8HctK1vvhkhFArEKYUKsB9jgqR/b2yE
GenneaG3jfWRCgM1+TtTBV5TMM0/pv9JqsfUYjwh22TrfCiUOZJslQnBvmD8tVrA
mkktUrg9gRdX+NUE/+yHG8ILIrKHShjWU10XCvACTf0j1H4gC94EH0+LWN0qDghz
q6XbMUv2XlH4cP5kZ55jIzfnNYK6DYTYVQQyftT5mO/OAV3qS9fd4FwBH3FCLse1
2z+8C8FJ2X9GlmwX8Lq4Un9VdXoIo2YLRqYZEtpBBqdFteZdMi+3fWzaRi1V61ub
HH9ynTCkjZFhWvRM85yM/av7uDPnSHYVbKV3JBHfYdtQfRDbfFHd6O62Q2YXHd9N
vo4xy9fvovxEBA0hLEjWheDP9sE2eHXQg1aeWpT9XOq04Ig2ESniwpNWBjVdZXEH
fLJJpiW1Y3YG0jRLMA74oIPQq+qQCRyvlQAGJH59GrFeEYJT/fG56HSkjEluXiyK
l78Kp+Xo8ut26vj0bZtNi/d1FShCxgOD7O83y6PhSu/4QDYQScO6aNuQgu4jciY0
ICYtaJSfwuYeTgxrmdUd57HcLMVDSN3MemjlaB7B3Ak5DBxl0ORJngDWuEMpyfLX
HVxYhQYFybpuVIdWNDl6cUrNgJZjWA8bBtPSat7ZEFyesnc64bk2vJojbfHbYvdk
ihDRQioGDjEfGSmG9GEmOagshpg0ww90tR53EaXhdMCtmYWRq8+eWdT44q4WHD0Y
ENOJC5MKYw7kbk25U5iW3zVG5KsuUhvndY5lEpOq8OfiPN7ncWJaNEecCAJN7C3K
oh1j2W6qnfumq8WR62l4vfVBfbq85BCd7THy2IKKkBI9Bm2N3HpxDYkIWtGgZabV
Cjz9rer8uIBHYKVPIyvb6ajsJ+9VvafCJYmzPgu1jL/SlAa3DJqo2R+q92JnARni
PmrDckwqVeVpMb0ocQy3hizisN7LvcKuwG/az0gtdss9Y1F6JYLEAmAmbJuAaH9G
jfwdOwdDrKePiAb0+pKFvk5p83z7AH04xcVqHsFoMFmLJeq2soITBau+XXs+8DNL
qbUrNeCuy+mhTigg16C93Tmj9hsbbAdSZ14Og6+Jlqx5dLzyFKj87yXVxRmik//c
syq7LXF0myjGLW9BuYToPiKL/KjDY4obF6Yl2HfKfCW0i7zM0CV5sx1DnWLp+kMV
YUEiXQ1fZC/S8+4V5zvXfLjgtiRO9oElSXrcpFkUlDKIy1cW2vTC+kOCisLBZVCv
GWYI8ML68QAljJ2yqPjkdKkPYlfxQDZq9M73JMzPegCemrjBhVbd/taLM2rHuqlT
nsz2OCrpTOc92AlRwo5Bsw1z1s8naNV/G4T85+tUWrLNKthI3WRvckuSYhy8t9sT
oxyPUNj9S0M7ZXkesMoAb4E7QiHlswIFx1cXilICMoHLgGzW/EftNOy2ZkuUBMN3
yp8lmI+08cZfP4WTxU/rZda39I7EZezI9Kde+teGiNz+np3DKPTfsg1fpuqdh2bO
QJfYMTQg/drG+3i8mrLndKbWQEWCZMwYFnsnmqActLNRqgYWgOoIdMcHh+Tsaony
m37KHlFLGShU82ySdCqRJ3SsSCB4wKtt10oRGJI4yDlyLZIidxFyGN5Q/cqXEmAb
uEfsVo6HkmRAxvFQ7BxnX2UXCO5UH7xO21NzVhGatTERe2ICzMfAOFfQjOwjE30C
qdLFL3eiNyGVjIZWx44TBtuZFL7ob+FMyh5cgUAZTwmt6gH75AYZAczFs7xZCjW0
f75qNgtOmc8LhozsHJAUiQp7pWX2VJceTs2MQcojHu70I5usW63eOtmT0g0SBP5L
WrkJbB0bWwF4MyMM1wUqxMR581SuKTbyMGac5ML7WjDVRfIb5W1g6KVNSGVmI5f8
w3XhfrhkPaM1G0EEp+0BDYfITNgWDkQZxtr8J22qtdwj9Mc4Fo9Ev+/yCxIWJJDK
IaSE6PPuSnDuWxRxFUfUqYrP6Jl7qQqXSKiri5iaG0ig9kknQos0F8rqvZ9OaCXY
k7jHKOQ51MQLgnYJqrKkwx9ce88IVdXntbgUIt21slBbIQ4xjZWZPQTHFrv9ULyF
PX127b1yJZscEmty1EeaefgIyFm5qUg6AiR6QDKuY4FS9spPgIOUbaN4yiR3EECh
obWRSmKUk9yogpXuDWdigC3DN1xa0Jk/bB7bz8weUdf38urkKnuSTWkhfKOR1lTK
haSeMH1B6cJMhiullTuZdlMD7lP6iA5Ej0qgWHB45fdptbuVa40NsZeM1oD/d4hY
R5MiAsPwQas/jbdLfW1KIWRQ1q18UK95hV91bQjvozgW4QmnnpwKZLenV80inrRV
xLuUYcvv+KVDMD1wbCPQuID+gccJZmHZ2CEQj76HaO+v3vRi/68TEfSBUONIQ3Cf
TdGPIk9P4NqNBawfgFb4DBFVqPvfiy32rM+f9bry6CP4nLeHWN2abtWqqE+FVqHM
4rg0/lSYFdTYR2IQheONCVCAi8DidykyhdOeS4qLB10ntRn7S2y0WPsIEQi5CEzY
MQcOhjUjujcHi8lagLL6+Q8CeyA/+kjg+U7v15WaLW6cYFWAHRq+TekA2O0sEwhl
wFq7IlOsszYVwkTDKS2ckV8dN1DJBuB+bE4n8ZlrSNuFicoFU9aSv9WhegS24fBt
5iuL2GAIbk4oo7lesQ7mqzIPIsvlORbtTpA3S72VSpLcBFFAvV1G7PDyyVGIvwqn
on8zbLwVFqk/WEKoH+IIuUHzMMiURiSDxwLA+wAp48anTNCeezh3Yp32LFWXopud
E/qA8Puqr3E6tvPGeBNqILpUzn+xlS73qQ87hMlm3NL8OOYTVXDM+imCGa/3m4oa
nv7Tuh17DvTFVLtn5dlPeCt1H/15ExgQKqLNMJgpYRQmagZJUKtC035Ts+Swh7Xk
eAL0DLjNeZ63uoUjp2seAldJvVGzQmi8PIRqQ7n0RINEqm1izHPVVgtKxaS/PgPf
86lOHwULLxdaZJAOs48malYQ55PPKfu5dOvzeBkDIHK5UH/y41yrM3jBboHG9zas
iqSAKpi8RVNw9SPaQzkmuzIhPQv2wN6Yvmg7UFGSDIFKbRpszD5mxZrEnZFxTwfD
4OLzTlpHGmnRyOWmKFZTdnZACZHhBof2EPbJ/wF7Fkjb6sAsHH9yfkgp0q6t90P1
5Z77pEPy2KUlypgY6kaXGq6haDifBFEqo8vYCxslrzCYyYzcy/NByXFGgVhhHgso
Twaq4cFgAcL1IVxxdd+yl9sokIVtoTWJ56wPgLqbDrV0qOz9W3hZ2GtsTw6dYT6g
ieIX770QushUltR09oH8UDK0pstmzjIqMCJPhLuXVPEy0FKeBZ/+vnxuquzx4rsB
VcrgBc/Le/N+h7kZlfAIHh3PXMhNQ6nqX06AqI5jkWxJUJc68GY4NPwpTahnxN1t
/s1lwPnyvN47MwdghsyBmvDJAZ+TnVCb/YaWfsr+CSVrEUF+/1g8CiI72EaY8YPr
4TZtmvyG+fgt5YaBmn4CPiItXAradw7aI5iDT7uj572fRm/rSHFiggYP1mQGHN1X
qUy3Fs1uYadiqqdHvb3tnPyqTJlx2UJMSrIkLPvXwG/E0AnMH9HCrKXVyhxAFAbi
PKqbYF009+ow8UIZ7+rUkZlbmH1/KVktnrwuwBnqKcN/eFN9O45HY/h9Q9ktxbo8
agLwH95FC/V14hR5EX6wZSvz7F5N+4Jy6eOCxTIGgijbfZ7c5oI3FQ1duHydeqkT
18hBBSvOlWCDFEX4rqe+TseLFTSnrRjcX2w3AnEkQDjVzxf7MwHqgiQnmRfinb++
ynGsnSkIrlmuywqZ0mfMdBbVvB7s8CvisqDxwu6xhD8yQfRfBnwox2omLx6gg0YT
Wn35Hldk89AWHyfy7DI+hYqJwsSq0NTqx+IHnNn95Y2XpSKgG38YCeKhnjZqOzTb
nqolokaFxLr2Dra9qYuAb8v0JH38IgS/Fhk7S/ZcAjYYYj6c+ZBpwZNKP9Ww+TGR
Q0Hn/oF97o3rmNuQL+bcqF5kmOYNEoXJlDd5rKkrdGK0dtRC1iA8PRk113gSMXhM
u0+XbUe/6FGD3xJlCACqKhhOOy80Z8TI9iFu1qewFGUvI3eIaOht5pV90N1j7CwU
pIRV77fizSLuy1w3H0V7fmGVOCcbPlAkWCFaJQrm0swajAItyJP2z7r3ly2MHIPJ
mUMNYuMgq+cZO24HKSfNkzDdvNJkdsEZ/gqNRzaZiTnbM+09XSpPbTW2mNU6ssW1
3hEKJuqlhuUIDr7qWnRMIs4hdFLPqL/DbyDgXGJ7a1xY5+k3f/eSqBHJoWqVXFsP
wANUii45CBJhjoWGMz48PC6hwmYWDxO9cFMMoZ+JXMbiGvZEfAxARqu+lGN+bcFC
Y1HK9RiUg+7c0BueACfoPbj4Im5FALZIHcyXj9CIa0oTE3E2rAqIlnVc9CI8Usmx
Bzu3O2dVeXewOho1l/aOY3rMl3EezQ7KeOhym5oO5hfFLVIpe1VMyXD+vw7tkZF7
Kmgx2QAdDBLTlI5azpPOnL7yi1LzF1iFQ5yXJL+lccI0jj6O4S0Go/4VA5C5Q6Wu
JlBBJlkGDV2kx6lfB5zoWc3LIbGUxai07stiOK/8N6sQWLIEeiLOGLpgdj0cjU+Q
osfZTIZYD0RJqKG8aXGOVmraPGgavlFauTbeL27n5j0tQVI/9v7FO+3ParKB+reY
1hwhh0ZklDGTskaDkM/8RslY0La04qrFP1o29//grtaOQKt0+DQREbXK5AlceBH9
dbK/UHk5YAIvM1Gop+YcGvXvJPera62r2OdxrYWsc7meDJY9omga7agD9FxSON/j
D+/dFmP6xuB4XIlY5/EEt08BY9oMdtlrGgQ7r2QfhTIpT4y/+Uqn2KIEWV2STXiD
kyBair2QhArgMUft5cFgeEmIq7B5+Es+nWrA6r3dAAZmRqt9QKouPP9vVS4oe7AY
ieKor2Nk2ERNHR3VoXRNkufUZK/dvfsuc0efl8Wr7A+90YJ3Lcn+Yr6ZU79vmxds
yFRdY2oL7hnvu5K7vLsF21rMuueaA8Gu4qqF3QAorBZ/JJUJsIEyWqLy9Mg/9eOg
ZzEz14Krb8sT6KL+1XIxIO2lFeXck9Be/t3Y83X/30gOlKGo4cPO8+risNCqn825
c0WCqOzZtoN3WcI/UDmM+n/mRMa9B90oAVrfLAMjWfZgixw1D5QaFkU9ZiG3mQPs
r0J1BmZXLFLlcYEpyhzL8sfoIuFJFXO/GDsz1w7TroT2m2JyAtGff3ezLYo7l0/7
jykp0Z4dyTpdBjFrPtk3c+oEV6o2o459RgPZ9sQkvDEMECjY9Yzpq695SFjMLoKj
s0ffjP7SzPeaLaDOw7tfBxucIVRWMj71XuBrvPqfH9oGekoN8aRF53J0S9wcIzV8
WQjtclNkWeARK4R4lOYpdMdJS6m+3Fc5rzMWn1ccbhsjvUkJVPHFqbX5NHVnt9WT
/yNH0xlNplYLuMkTWS/pPRzFgWATDkm9mTq37de8n300w+Rg6TR+JV8u0ZdJju9e
+BiYFfKhXIwKXgZ5CYRMcVNpjVzWWnKwncDsk1VVAGJDGaibOAch1kTABZuOGOjk
H1WIaUEXJj6vPO7ORw883BTLvJR4phIdlm3q6UqEOM7m+XwK6DGEMt5weM4zF8Zx
JbD+E9ohN7rdLmUKDP3AENEK3iOLVKMjh5QjrBZVJq90pCKF4gBfcwPhFg+QHF/t
w8l6SPkvd5byt+8xvBZbdc2LlgAsOrtnWeBSzElR5d9G2w5z1yJE/FT9+MScXtFh
Q+BVCsJ2JoXx+ERRwmRSWfT4qBuWu2S2lE3TABGaFT74E2XMkTvzjhX8yDJGyLTT
3SQx1SSe8G9qO4EHOObosKIKdUQT7zNZmHhPTy3IksURfzjX+6iHC7bJw9uyiDbP
BxtVmrE/gSxmeVC6Dt7Zi4duNMewlQi4WPY2CHp5lsW6/f6Ze/y7C0eHJE2/Ld2A
XnfanaFmINNYdKBmdYMwfG7kpx9X759LcWExkYm8h7+/RRl+7Zz9dffzv3xl8S5d
nV9ApNng59r6u2v0+3r3b2l6o/VTrc49beCS1O8KngyqaBAMqHx+U1Yw4UUiafB0
fth1EVyONA0TiZVT79xVQZDNRsurQFjQjZPzYPMNfor8E4V6hna6i1XDXbN/W48g
fV2h+g1jWTl+OwbbmwIp1PqPmCG3i4YDnSYX+FN68izLvlIoGhwhCQCaX2Z45G3w
InTytMEBQFQvljU5lWFVCeYKgaL5S+kaknvFJYRnPY6TCFcryFDXiATpmbiwOtSJ
FMoyuGrpWg49d6pq1mZrxNZEI/9Z0ClgimSut6hzAgfnFdy2sfjrcvIyrj1N3ho4
Lr2p+VDvR1mqbeyl9J6ncC0s0mKSCSbHCzvbnTSGKgxhuwwdcZ0AgZsKOM6pJGzg
JzVYhTbRXHlxgwEAupbB3ZIBu5IyIxZCWFLWdmBpJkgD8yRCigRKQ5TVHchkIxxo
oSgp8/uIp7eeUKvLRh2CPTaJKWD+QorkW4eUR069kfJ1j/ihtA4fm7OzEqBUquOk
VQLNmNQD0vxaYHKjpSe3rBcMy6tVPEQ4qcFfAjJN9yKnp5Z4dthYwRW7W0q8ugy+
JsTEiXi6UkhZMGzbc53LBqKeYafrHfr/dotgG+/l/gXyLXr8BlW1xyPajkKAOV8J
7szDvCYh7HAJ3eF7x3mQoSrTcUnLxyxj8V4OPd83xxfBsm15EzaFyLuyFcHtco2A
QFX/PuPdpStPvxKrl5G0k2bkXFya4xKR/Vf1kdMYJhFk2Wy8cj15qjVZJAT5Dfg2
Ud7gbwwGFSZrsgqa5XLp/510y1xyl/89+SFu1SAjvVuenjvl+C8EDVzh91Y2BerI
RAjE5YL/rMvs2hIPnXEz/8hi+hiTsGr+e7RgqDUqhNZbJJacKyWT66Lf04YU48hE
pr2M6t4B6XTGy9d0vIN4reiXm3mQr6nLzlb3wKYUEWkYbL5QE1U1jnY4UNGBSx4N
83AbP1rDMxEbdVkGPaNMj+8tCU3deS7DJwtgETv2hCgPxi5KCPaB3OE/t/svMdEE
SNUbo+e76QV6BetEQ0H/b8NgJzmstIYvArIgeTk3nf9BwlQF7QLpyJCTAtv0AB1y
5XgBTDi7hwu40DFqY+ThkCD9ygOJm8xcHWUiq99julp5LD3LeCtgW1diJQXrAb+x
l48tCq/RqoDm4dky5TI65pLj/DjtonoGlqAYBycljcnbR8Gp7k5Ab8vuWuRxprhb
+K0ADpbqpQHUYCx0MohFRU58x5Ldm66TxJ2y8qAQCSGVhoktkT5EVG7FFMwj7+ft
NbrzK74eXTntE8anfZR38io9qRv/bdRmnRd2Hohffu+Fo56Sf9Hmc34Tu0+IpEob
9EqTDQo+DOulO0g4pTr6nv6Hmu1ntiy6ZMfTOdeqLQYlXLqbVKv/ZF8cerepS1iN
18ELwjgeIjU959KMcNn/wBpjL9EaOQgl/I+knVFR+jVGyzFhnfXds1/CUGNhyz4e
vOTKsD9UooeGe5zWzjCWPNdTlgcOsu6jAgoPH5OEckAWqjRBS8gXUHuxUkKR9G0R
JUNEdEUxlMg1gUp4CLUJIdwJLQEJDqFgJV9Snxb7DDjsqjM5GEK7lDCUCLngsgJZ
21jO1pq4wYHI6vnsMgRAJRlocFMPORt8ZjzBsdIlTZac2I7piOvvHDxXhb/8Jnrn
J9At5ZsKNs1vtN/WsZGpgesaCS1/phQkM8H//yKc6AR9FzULytxKtUV2FL/xQqG4
pOSXp6o6GMq0JrD8EeFi9UWTjBQTrGBlm1Zj0iwaAWYyNWGe7Ms1FHvzk6+xQ3TT
+caMbUXp078ebHyQrFSVTN/y4lR7tXH0eOoKnnufGm6HB8Y19o5SsbTfIgu6E6Jv
aFTkJ3a6Uzfw83jaKQCbF0RBu/7Yra+s8EP2vD6vbb0lRaofzhCIem6Y9ZzRP4GN
WweyGO6Xj2ER4D3d68hXC8DPDorrpJpwItm9pFi8jq7pGR9d47x/neJjMXeEwN7s
XgUNQKnruZgjeOTdPrnNToHR6cCfxNYsPYA0VTnUl3Gcw2A0PAKnqZyASBPLJRts
GqGwyeO+R7wK4TEeKs6qq9EH2Tnxpa9commZttmpUpiHJWPpEpCgulal4QFOVrKj
ZJCtwRvUqF6sGyOwXDcWldQTeax0XtMsW0v6c6x+rJK5pazDJssf79Pt2YWwZy2g
QE9imABJkr/VU3wmNZSDX/uFhgeF3wIino85uQwP7C0wFV9SdLbQIR9HNu+kq7pk
7RBj/eI+Tjyn23m5n2giYy6Os1yy+1E6Vh4k/X3weJzuP5nIaHR5t7LCFtklbDYP
MzxJ6Szy1bOwUKm6lh5PlquImrKiWgXNAMXgmUHxSAOu2aUwH3x47hTD3lNkvH4f
oNC9gKJpEENHExxhC/ezFtkImDk1EuLcYd5AmI+uPm1RfIvFurT+MWYZld6g7uPC
poTgslD1M/9Q9hDblRfnHJ3mp3uVwdfVxKlg2CaASp+Pvi4XX/TF9kPpOeESm8cN
6MswXgBH8GQBKLUgj/uR4d93RblTaSZ8Th4dDg/MMiAx1EM4/mqcEiZJ5lg7z25e
ygjlfrFt8eZWgptcAd3D5EwGEfLwcwQbfT2U+gv95CHQ+FkvJr1m3AKYOn7xQ/ZN
wpuryZA30Gyx547jgUm56zXNjGIVXeG6brrfAYAmp1WcBHDmgUoqA+UQIsnd/3op
1ezAutlP9ds0qE7Ag5aTrqCFUFny+rottyupODOkRfX15YUE6R5W0RMKbRVohKpz
DFn0k2F0oBxlMESkmjs6V7sLKYdwAO28Bjmp1AJOLquj8R4vBH5DJXK7gyjt4im6
Npe/FOM3HxiWRsZ3tU8ibLQgXPIU2l1mRoHkMPnL/FERj1yKysf7va9MolATkotg
pG4rJ92T+NkovwWvWoS/LVObIeMpsQC2Ys4pHfJcWeiwKC0QMa6Njj/i7Q9Mrlvs
RnQkCfVa1T2AZyInlcmVrv5MY94rTsojMkWXrjDnON9zcMMf/f9YWjDNmOKSGNy9
yrc0JVwo6GNfdXDjMwghz+RmsiWE3a4wIqk17v2bbE4jLa0Oirmk9Tx+aeEqnP74
7Musr17ytfueNNzNDCvof8jXWxbIB+ov4BQzhDda0L/H7C43QcYVPr4wlBsSjyXF
ulD8GbSAbifq3QJPui+twM3aS+d1i0GdwiKUq/JplCOGUbmAikjQ49WGne5lrD5/
o3PAnXyUKDkKHkY49PcCVm89hyDMnxSCAwZjuCPip7DWDS62M4FSQTNMsAPuVib6
PvVQ73uT1rz90eaAaTzs9c0ByCFU5/EC6n9f8EmA5yb2G46nj+nq3i04xkQPjHEB
v1VcqyUJBmWPT4pmdZNEODvXuu0ae3d6PoVGjuxK09joGsqQFgBBVwBDxr63xe21
EDQuuKzbGCbtD3GC9LKhfR77SEckfrttW/MbY2B7CUiU3RlyCyfya7YJK78a7iFM
4mTIjw/kA8dibAT6Ne/+pKx9yO0Vj8OIhNeGoi2EnU8Pnc53D7IVH9JhBUOfrKSv
/TsLG2NuCG78VPdbwQzvjLKEpptGMcDgVMVa7BpF+KH+6z9V499sfDbM5CdG7/Rb
cNOCd1HmIyMxr12MH/JrRLgA+aZ5dLmuUxAEolAx5RJGHDpq+F3PFieXEkD7gmfq
YjSqfiNrm9iWC09NpRJbQGhELi71rYxEBvVDVE+YYeuE7xDYoQn6ZYhjeFxOsTj+
31OMV31rUqxIG2D81s/rRNrc1N1DZ7OuwUZmtpLvMZ9FsWtoGz3Z9IMhyb2U6lgT
1aEdC7sfCjwydeijuthKM4GfJjCo60UnpSiZSoe+olbGQQ4Inl7fzeert/lWFncw
dqFGN7/ovVLu6TSJm90e5/BESZQGNTG0C/5cDRWeGW2dXBPpQwKr9m/ECDxyBnlY
wa0I386IwB0ShD36GGCMrnMwgCvZWC1ZgTQ5tAXwFLxSivo9av1QFgzezY1EaHUd
dUvlA2ROLcqZTkKTW4Q/YkBNZ2GmmOdA22hMd6pSBUop8URoL8Q+mHRajY1/dRAM
Y/x6nCpXUNzyqM4N9fy6C87M4e9I0PtJz5Mr3p1oqj6NbMfValfKWLYfOxw02Kfr
krGukZJIuiuauI9Pe6Dp9ukdjdKF9LLnPVIZGIgfOhdX27xEIZ8h+qbUjsmXxhz9
Ajuye3I+ARs5zqZfgT7qVDpKq7S92d6o6iFJS0cnYOx6O1If+IOEasnyOkYC9TNx
/BxRHrhRB02vfV/oZA2PSGod81wHYwMYyUVwiGSzWjQeU8ayTuWEa/3MjVT01EJL
XYI77I3fdFLaj1f70mrl4wDjeFjPSvq+Pzz5KyjtAWLl3DQ3/FGt0J9DgmbNand7
r8/CUTlwzzz5Pa5/r+uE9GmRlhln4k/ENxJbDZW1viHRJpRFzCHwRdGYbsXMXzOT
piWyMrtomnKG/ycNmbnM+qV63EQpHPJDq/C8OYW+c2pFWYGw15/o991XpO5ereYd
+3LsbCiyJdj8oDf7QB6aQ4y14x8kcKjxBzVBTDNlGAByGcbVkmyMqfMsGV1IRz1u
JfFm94wmzIBp6FZ9CvsHywJC69sWPQzb7YLHQhPWrxruWpgLZRXRBf96Zjua3wjL
f85MccP48hhlm9aAjF7qa44hDaJifqI0s+8jO+n0cG3XRbN3jk0AhtXwkQajCzJn
dWbwRjN4Lhse9MxfEgrg25vEYqaX+33JE7RKIfMOwcakMt9bJI3hTtlf+pPSHPn8
rjzV/79obeKD0yW4RI7dOK3AW8I39Qo87ufLF2SG/PTh2E9S2geOT8l7HDRpRBh7
HxrjoTapBe6EGmqUkogqUlLBmvMpPeVx9Ovv8rrsPoo+k2V+R6wu0IqF3+PUdl61
CC0QJXw0kLyKRmk/KKZy5/0mjGP+uRPybvDSiD+4E7+3Iu7pp3nsmffAwN2PsvG9
zYk8EzxuWhOSI2GmvtojUVYEc3+n0FJYznmJK8rMPKPhYGrQRn8ZC7jQrmS5KpA8
kB9bRde9dhkUVadHOKSFjTuGdtFDMlEkipTO8xichrz2vFqCQlir/y1VUQmhSwMU
7XBzaEEdi1fmVoCb4xH4nn4NwKk0AlsYtHH+x111lCggdLV5iW7ZLk5fkDrI2INv
MBKkjsnDUre1WWEDQ0xXauBNpLUGLB6NJ4DiiLuEmQr77w50Fbxk/maouPcu1LbU
f8nB01TS2uE2ySaoEr6ze9Ij91zxAjEni/8/SPAcysNFeKGi7aCG2PPyO00KTVvM
S7eZJ7XHQhkZghLtAR3grpA+njWWtGVFgsOfZTPRm53IyAg1kyvIZYS2uaV89LbD
qRtnwx0pV+VgjfTyIJsKUxsL4alKQBQlCPJ6Wa6nUPZICcJVC0o6D7kfaevMZq42
zM7iq7z5aM8XaMQbTWjZz0bHWntLF8kG+cW5a0VOGqBzZj6gstCTaydppg6zrWJ6
qNCMITnXxq+ggbJCtKSd6m27BUOfO1LN5aSDyeEd/G6v3zWZvntiy2mcJzfgKM42
N6eGRDcnrMPs20PlQL+9TSwpiABL0619ipHHmOXPLIEzp0XP8TJf+vpImqzA/ThF
ecG3fNEDvUlmX0uPhMrdQzU0JqeaH015TvADswuv/+4VEAMx1bSGY4I/I5UzwGoe
GOuVMZpXfaISWWpDPnip2hIEHH4W/j5lyYtrL03QCpIegT/eIrNYo4MWipNaJ5A8
zVac4dbFsOOsNBXA1z6+wvcuoNAPD0QtTLjwH8F2WCG5vb6Rv5lV8+wVInTl00C+
F2WGMiWH7hNUnm1mO5ftekjR3ugvRhZ9n5MBcIAvZUrZjs6X+FHEO38kku65GbnE
ch9uRaaNAdoGi6mqWSX5NXjSCOL1hToPGkmh96sPDuUf8DupQzaQAbBfhu08W+kJ
kIqr1zZ5htao9DURwBJDpWXvkq3S4lp+niBAOL/OCd27HCWrzsd8H8if2lOD4IEq
Zm3fJjyCOmCh0Dh5YSWwjLU6ZDhOw0MnO+ZN/IbaS3qd6pzWZjP5ANTrhkhKvCD3
OHA7kE80y6B8pst8GF+27zAntRt0AvYsIYs/CgNnMsS2hyR2VWEXrUOyYGsqUlSy
WqnVHynWGOeHszGA5hdBTO8ja5Pn3MsSqmjGEqr/85X6BXeI8tXxoISZEPH8J/sO
Eq13AwfkLbjYg3jMaOjx3oxh5TAlX2SED+MmrrIdDFF5RDGEIoOT9V8P9LhuiPcv
7ubwctnEBtjYieaQWc19eAgniqJ/UZoRbU4Bj+ot5/p6UjdQcPnjEXgz8tNaGmZZ
iAzDFHROPUbr2nWikz34/toSLE5u89LUks6TXbLV2b287rqr5D7HmLb+PXzYpzPD
pEIQRTjy1YcUZYVdSZUwPVlpJBpDnq9FsSCTpjdD8XV/I9JeLBAeH2K6OgSLMPNM
vXnWOKzZreD/cNnynu44fOCkZK34BKOHWfPyghBd1JyeXUhmpetzQdwTQqn3VYzk
mNuRaVviTGkPkYGoQZuDq85r1CNfQGegCEV5hSnSvI+Y8JhESpueZiznLQAcDRbp
peJjwnVCuO+ftlzRyX+dx+ro8eYgwxtwqrbJwcvtpfUm4ZMWuxXE1VLJ+xc/m+vt
e2gKfvyMX7wml/ywsdfluGtMzafPC2nYQbmKfHLXl2aMgC+1dumZvQIYw4Q1/2wm
IrXaNR10f92Bhrj/kV9e0rZsJB/Bf7yOWX0sHsBt/oHT45jCKGHikYap1nnl5m+L
kgjhiat7PytmsiGDvoBljh5pntqZ5mTjhARR+/kjIY+bTnQguVX8HgYUS6hW1dlO
N39muuXFhzj1oWgjCwvlny1TkHr/6hI3xhrrMOrsRwMqfq95XxePpz8MyYet2bF3
fJY7Qw5K0Vymw6Ih7z69pR8O8Pn7lxPwO0KW5DSGpZplJP9fzZEnzdFiLNV3rygM
1Ff1q0K62xxSvDwgz6ScKliCWRqmCUF8gpzDFvwK6+UaWpBPPZXUF984htPuScFL
X4TugoCtpMFttAu7dfc3QO5qUA5m00hZP/Pi0gNTlR8KtHz0E0ltmjr6pBEhEGfI
F8KPhQtHRB0e9INEus3dkdfO/lxAiFTqZvBQVnDGSJAodfQgKodInrPUAnRtvqZK
hhNq8vbjSNPZ+7Z7+EzGmZnOyTxqt9WeAff1O7zaj+mo9/LvQ05LZrj8Fitrvdvo
4q8wZJ3pE1qhNnMqYj2JyY9Oyy5znBDtyTy6iENMX4QWgbKPD1dmtUgaR9fRn128
M+AP+E8eGDhuWgbwoXK9D7so4RwyOiJ5CJZMSB5TGaDmiRI+nRBqRZ+dYCASTBxQ
17+tvpXTmoVC0jFh52jRhLXFh4RCiHCATZ5lw3rPKZ55EhXPGZU/HakkijiB26YK
VXq46qonsLDZV0DCvJJgQG4uKBlZI6U/I82ZQaTrXpt3XlwpLWkKonEOG2kxqQzD
Of3QkIoiCFptXIhzpsZ+6JY4Y+nscc5BSA9/jhsXcTp+LwqgpvwkPFFy+jI69x49
Sln6OzGP8Pe0rWOWyofQ/mJ44J51a2fBlTfkUaA7VZ0gXEsPecQjCn/EEwcn5CTq
C2z6pdCVec4bK+DKw1cyl/ZydtQKy4CV4q44FmX1I9RwDH9a/mBzhmQOQDWv4gBc
J7LfZEv9f8ajZrbkim3s6EkLIdb0h8qvVFsHxtJDfEcapZ7YdqYO78Xl+hmolVtN
Im7e7ZTKwOEo6wOTv6qqp1ploaYF5Ld1KDvSeq8X051flJN+eKF8hkjxVt36EzAu
ntDCnRLSZiR+2Bep9FdSAcLOMHYRnL9NeacU65FlXDtrWe0S+YNQsysHFWh6UZGW
DJm1zIK8URcvgy+TDJYVfjab8wRrzpSEZuSFAMMues4Kdbf4hiQ46u3JsUyBK+vl
L2dsx7r/VVPFLvL3qGoSAs6zrvYrhj7FjE68neaNh41R7PipWVzrMmSMWY4dZlGf
wwpJvbWPtieNKnx8P7aHcJSnboRpC9QABbNOBnBmKMTx2iJk065A7zvueYKnh0Gm
Ggjm0SuKzHSUqMN6RfMaoKReiaYmvyiHlzOFvwa66Zf4p+dMBNs/SwkGn4nvORi0
jXugUngehdcxDfTOkdWu3n4XsdLYKG4Q6ivxMltFENUq+vNv7vPy1RaLzflu6z8l
oboZKC6ad1dAvFuXKblkHELfBCigY4kqe3aHT//LkUbEoOG11W8Ydsos9h651aGj
ciy9OC0ONwWkjFw4JZo1D03A9N1ItK8Yti3Y4P7mZlH9wf3F3e49auj5KqzErQ0i
NGJ5QywqnLFyLEEHOITjADZ4UQhYMfwlJpkFaEu7kKz+sx4HEzBu58GgKGP4uX93
Odp2ehv9xNbUsURMBZisK2KRjnakb+sK/BjGecWO9BvvZ+6479xMwTKNukaBY+5w
KBahLHZD3f5aP3QKFyiDsML+Usxq+dvNJg3jCpyec9bNfNxXnal/8QHFaQJrROMg
o4pLNWkqRMWOdg173f61Xx7dRpggWHSmCGdH7TPmV1CSdYOXPwGpbOg2nqZdh/Fy
sQjbk5nN9IBWs5PHVTXA2F/RBeXwPEYzCqVJYWFTMkyTOX+qVGZvKSgsWJgtAXQ+
3JGZJtWlmHoYm3XFIRg6j6M1F4Z7BUpXw0c/iJ2NbckDXT0E/nNNb7kGRQ8HbYPm
pQC8Ov6FgI1l9nRYiXbEpBJI/ce/Fc5sYd6PchJq/svdnFfFzYw4dstK2jMgOZgx
34+c00gtG5nyg+mnOdPpkMpHUzA/IYBFz0xcgngCuff/olV2Nlquh28RdMeYnqzf
kOevC0+k+beAjYNTTKJD/Kwlc8fNHUiYWbbFH09P+KezuY/AL/bfoHYOh6uiI+a0
YtL9jaN2KoLEyji1Uc11ZGDF0zs41Ti9aVbmg+mUysxONxkNXFg+zzpyD8rb1a89
yoK3rwv/TXtZAvBR1OKRiIEzK1mKodig2sVjgt7sIeTIMTWL9fmgObpXOhyDe1bP
+W0MfkdHgH3TdLyO/XtzoUeBmpSmdb2N0zHx/WVKurJdc05ddCsKo5wM2tjn93hJ
L94q30LJQBR+5gY/iIVGQxPzJdqZ3FdJoqWI7kdNaYdEw8QchSMvp516YgJYrBqZ
5L84s5jG6kvuutMqEIsxZbDzkBLUyDGkoHtkeIP1L5cKhOu3R/pBS5tJhk/il8Fe
/hsybkoKdftZxPGWOq3EEfc1eUo+yYH4AKuNr8qF3CPlPe9rBpo8NA8L1PZ4Ud4B
cKKpHC/bZKGZZntDtN8VBE/8Z3Hhcky4Lx1ni4n7inoawxxn0CpBa1EJeAIXJA0c
olMKupCgar8eSeCwa044dCNF5bVcPBuVw+XJr/O2Dz/izCcqWWyb04/FgUcGoZuG
fSwywCpR8DiKNCNekV5tfxIOYTtxscmNn2NqjEYTkg2sDP+Gn+mRlPe7HpVgQ1RX
zKCHEqFI9hSRIEkNHypILuudm/dZVDjn/zJF3oK2sDlMnMcXHybQ2crtVG/2ucQw
OwpIKmNmaTLqbtrbAIg0hU/jrnUbyJlAlTYzcTCn9kh8lB9OxXMhinLFXzAxCw1o
3re4tWLG+I+3yfsqxaIjVCtp7g8xpzbKudf6E1QAOCmGzfVGbPhlwnEuNk26UZ61
SY6diFVOPxWcTmx2frA666YwWayKfH2Kznl/k/H2qMk/XuJoxZXj6jKHbcCdLmjH
9lQ5do2khWaWrSbxh2fHEB0kanKaIQxy9SDtCh86X3JWG58vagYzExSMRTjWcRRv
7whobR6ZXDSleoN8xaly4LYLPHPGbi+M9ml8jgDMywbF2bYvYUOryHQ4D1uN26I7
kEMK7Ll5tUAXPHy30E9cxW1JQw7WrI+byDvcslymTqEBSessY6SrhNOSLt9QUnQT
XkoPbQF9i9XLX9YlYST2dNUH9+O4jKX4iKOHASDMWtRknp8/q0PHWIv/RpQPti5i
cyIu1rMkcNkOotC1y/MPjx83iiw1EYesgyBNtlFwe6OnBBxxwXBghDrH5MgwYWZz
rxN69LofJm+bfVc0el4hoGlgbMlijBqUtHBDaj/FNSCwhZq+ZqtLBRDx0vZX9aNJ
kh6tU4SwG9Jq+TlPdSFwteaqUdJh8jVnSCd2FzsOnVLJ77PsQHMsmjCuOCGhILqW
zup5Swv8v74OsIotO789YKHOHKjSbJqdeDo1RoVhaFvCm8QrnbpiMDFw41Opagjw
4HiEa80e9G+unExrQKmbdrpKPhGUa+5vtNUO82Mh2xFGc054fVFrMKOBlyH1vCV6
kDydxfJcmb/NEKIv7nMIoZwIWAwK1o8mIkj/zWYQGi3jg2NDweCde58F2dqMX3BX
xwgmI35DecuN1mfMayvX7fMzJ93rBQaZDbKrWdv1cG8Nm4LxWybjTJ5JckEnVOX6
u1o49v7O5eaVprjigLPhxtuGGa752kajJl7KbKseJfhO2TChR60+cdZvcE5Un4cY
G+Gdn2Ot2IfmHswCxJp9APqVbQoRHFXEhaHjWfWBHSMcMjFgySmhHru+CBRivw/w
8Yzw6oYeFJH0mMNCf+MptrnYiB87M1BwZa+svjbdPDYotx2e69hpivkXZw7sO+pO
IcYj6uoEFQUWdNb5g1XOFXF4UCZ942zfzXzrQUeFWNDXD9njfyCw8sQrepKoleyV
QyujRLhEE7x1yck7g9XdAv9X6rtF9uTHGVwpwfZSg5dUiv3UrTOElcWzp9Lrenwc
aXWwgRb91L/OYweNb2fiwOTSydP/cLA0gnhi9DbRLzsvchfw2wgfzRcEt6WZdwGM
tghZhfWKF5gWxZU0JFqBirtL5ow9Vn2+KJK0lpVLB2I/HjV+qS/WkHSEStZNx4Bz
CVdo9Wz1AZoV0pGzembR42gLh3UjHyY30IaIzHN8jJ2H0xsf9WoPa7Sb8FtUA3ES
TT+ANu3nUant1+XrPg2iZSsOxx9TDQ73XqWqlll11eSFpIOcTunpwM8b6371SHBr
vTTn0WmYJo08UARDr4luuzUi0gE5BRr122xKHNDtFY/pxowGQI2MNPY7gHiOfT5I
6YO2OoxpRs6emcP0f9SWQ/5ZyCGKmO2aTlta91nnu3SMTB6y4FduHdKfBzHAaeRB
VjMo3aElG0qSkcZJ1eEPPqg5NHsLAeDuYINZAKbBbUqJRgL4cvSL+DquGwGSlOtp
JilFvsGCjFdP7c4dsMssfOugaQT88rcz73sslkGNtk8pzV5+CZF3ri3Csdz5WHCg
g/rcduWkncNWIzKgHWWHaDiTcLHpHBjTpud1WayQezMJYmQcLXYpAg480n9UtNG2
RDloO8y9bCTn9DJUsykODU/6pKdCJwjnp7og+oSUtgqFyzwCUYf0qPE2V8QYFxs9
fx/jHV65FaVHuXbVSNAvtpjGq01qGEP5jQ4rmHWT0oip/eLmqFUegZ+5HfAy1t6R
bX9t/ES45zpuMP7IJDEiViUOItlPOK0hNwfJNLy8CInpMCbgBS1YVhHYaj0QLUkh
n7NyoAWF3WqEzTG0DVHQzWd0VBlqBgxpdpWwLF04ikMdABHnj4nVKlvZI3YrJA4z
dZDvSmPZNxeshrLynGPr/r4Ez7cILMRGSdtPAbDPvqr3ffvqzj/KoSiKWQH0rj5A
EFOrqKdggDJ5cCJ5aQadFKU4IcoxLSgw/p6ZpUi23hSpvgv4fNvz4vxK9+WhUakT
p9+3DDqGMCkZCDrkPouuxRxLVllLIGSfV+fvVix1aah2bNrfR+lndV+wsKUU4wF6
mV2JemrPfQmpVALQucN26gYbW4CpQJ4IeRB8ETFYlXsN+6n8q/bSZFoeeytZVpZr
7r4yiau7+4nJEQaI0YNAb7mJhfZmRvDhck/5BjEW5Oyihmb4M4+HNr0FXeOolVuH
LrWU+sq3kEboJt3QEFetS2F0n2pE+IVKvz1i6kgkVpUlWh3Z+qELVhSgkWbQQU72
TbHislz9kgiATqFCQ0x9B0HA5t0kYtrABZGw4Sih/HCp2kF7EQxRzdP0KwaItFQV
tCu2JzAkR1IJBOYM5ynWy8AQ3+S1cV8ayFB72eMGJu0qgvOP6z8Ax1rGnFERiZYN
dIMDq/5t2rQpu0n5K408YcsK9TlZht3YBgpyP02Ypp36O6ASK51LECWV4nAT2nIP
6HpTgRrNW6z6esGkjQvCefhvW9aQ93ZX0C6HVDFBzO/cv/6jLWYy/DAzRySGcjcz
hQM7QvIbgRo6q5XLrj9/4aQ161lBm5Kr3VXiC4E+Igf4veqgKs7qfyArQ2p3qBHI
5D9Svd1UbRO6JdmIEldyJOEzdebFt1iBYjROOGxYjslIJAppXzivlMahm9gCHrlY
fTGbq4Ncbnp5rwTPjMBAfcLUHJ0DlmbMpo3/28tQV4wdp3OEGtZbghhRdKnIqxoH
dv0BTnxEBH8v/XoM7wHoB5k/SmgguKJ/qN5+GHh7LFap/0Lzrv+y7VVsDLRaiCjb
7DJmCjVLnfyZLFJ2iZ2KY52D7+GGJrOTLNy+zgdFeRNGPpb+Kxq9FaBe02A6gfHd
Dhsj1IC90ySe6hgqMwW4aFc2/QV4fZcARtZ6SjQBu2lztIVo7oIFrPDPaJteq8mE
h4u+/FRjpVxZiTZnUHVQTIAunSB7ND+6BAPuKv5D4wXcsT3nG4Dccyc+yqBB68Wy
GXLiOoO/nwcwdXO4GAn8pscfcGgc56Q3jowKgP0TG6tf+Q1GXvto46Qkb95g6BzF
/hkzJthQen3iXIl2l4IqqfRrE5xCv7wfMWlSnlo5fxj2YjexA4fWlDIG0IxKkYp8
kdI5MJJAgjQAzbwDXX2QkCqoEZyVm5kmxem+8UtXspLuHKmuoWKfFF6B0E/g9RJu
7JiKhkBxCR+56mATrzRSy0PW0y63wGHZpzgo0U+mu1hMGGb3974zyu2K7aJoUplF
DmS+ZGP684UQfgWg+GyeiIDoaObnaej4zA2bcDwGhB81ZvoaQK7oNUAD2ux2mCKz
Ak5q3Z0FamiURnW9n7E1zP2zskXeCIEqedSUVRU9JQbmfUIJk5LPNrrOrhsPj2eD
Cr2N9zBGRyiRj9hBRV/wBV7Rd9SI5wZlBALZczri5KunTxfmXwM2nfeQAbzDl4HY
xro/wiag7YF1WyIM9cPsTBCaHqtwTfEzBAb3cRdHXBqTRa0MF6GSYOjcYZsnPZGw
+nlgKh80/6ckGnXEjuypYe3JNqcR0ypKZ00006JMOF5HCeeDRabnhlPsWHQAbP7V
4T1DEcx3dwLja/HGtpMTwlVj+xIiOB6h5wY2SjbTsa+jeXIlpQmmEA9EAzQSdN9Q
+YiFBRdsgfy+QI+l+tjiZzI+fRr5U9egsGBapC6tbjaBSsyvNEFH+iL9jbnHBV7e
ROfE/Z2yq1tWuhi9yf8auQUxQst/8C4musbVYS3AGe+DqjKAm0IFrH1WO2jeI71b
RgN+n3E4Y3rgmyNeuhqIGihPLK19O8v6QjGVXN5hn9kpXMEftiNr8HOYC5fIaRtZ
WzC8u047su9yI6S/XvIWkk8mwkOL6xudIzxEnzrNvX2bVP8OVhIlF1gZ9ZP2nQqA
KCNSE5twL9vzNftAWvAfMEQ6vh4cGQlqXfuqPT8EILsjoekQckVzdjVHEnlh3y0b
Y6EvmbwtmL/KO7StR3VQU0QpG75CPKmLpUQWfkC4zwAXnC4Kn9VA8VZ0NL9auXQy
NAjlTt0qlhraVwK2VtFv5hAMFzxZDupUJECEAAjGy4Opu0HaRiR2GjTqktwaosSv
KQ/9KqbZjOYM9Hdd6jDQQf2AOXwSZWBChhYCJk2a8DfInyp06vATTkm44NR7AMw4
UNxcMn+HB8yh8/Lbt77s+UFQ9gchfKXgbSWYL6Ws8LB1pDam+132DE821695r32t
j9VoqCsENfsHwMsTlwPGCQRaNo/+F58JP/og8EnsMmnrMJ5Od6ipAXjyByRnzxgI
TZwxs60WzNBmMXxxjeAVoJs7NB6L3y0ONsKRfw0tJpTG63aUhWQELsYz9eNURSD1
/dzlgaq1t8kTZ66yJQYCjrnIGoQbZUDT0i7sotjPcvWvvnHtSU/Jskiig6pHgv5N
dd2/NdXeTyAIaGvSiHCB7YRSqxllGtWsDc/N/B1Mf3Mel4rFhkt4nrzyqgcm40sc
Zb13PLuuIwqVC1zEc7fQd+TvC7Y+gqPs++0Pd0gosAG+gv+VCY04PdDjgekLjJn0
FTVaYV3cR7PZL8HypXf8BYKEvPx7TTdaYFEzd1kUYATUY2y4FBM9e2HAE6ziBUWj
/GKrvzpRABiFFgxim7giMjQcWW12vvgvFMEXkZS3splpWjWDCEKcGK1l5QJadQW+
HkYzSkKub7328IEs1cx2OG4WpgzUDE5j6d0spagvMiAKygj4ntmto0idFaETu9+I
zE4rYtdVpEbfxegN2aiimPW/Iwa7iq8KvDwrGoT7yHrFqz9KkE7ciI0z0Uk/Ytq5
gZka9mM0PoGlcFu8fkfQ4c8dcwfXNsDuvDZNtExN9RVoY9/J0oJpMd9IzZkmybkA
vdOnsexVltyKuZrs/zSyt7t+GOAI2MamV69ztcVVfAWd0/m6yIwZXXsk1kGygyQn
GHgLaNuHhssKaWhWQA9juzTpKcsvnwjphDxkJHn5N31DbkYXNFvvw+mIutIhexL4
xUY+hbf+Xp7BuG0emCGNA8nyxkwjXl0lyPzj4/35YRBGX2709Y6Y011rliJTGMDz
hRFVDMc8aTUxOhHIYR/H8JzzGtOg57sUTZ6PZ/tdAEH8Mktol1HTLdq23fXIiqbe
BOaQo823fzD9ZJF25CQM/Z6T/1BP9S0xYmeMwRIsHszhSQRH1XQoof6nuQP6IK5N
9JSpMAwmMHlEKrZqsjHwLCms9faEge9tCUjEzHPFpFNUvcrYMjR6Px/0TdxZIUtg
VFDh+B1K43ftILH5CKeqX6OhMoF2+A9P17as+6P9qtd3+DprdWDb2tMmjrOCXsJ3
9WqvjPEbg9bpjvV2AnMoed2Pc8aCji7AYdoaCHvKLv1mzDZ5c8RK100882mwP+4L
tzGcCdANDhvoKJRgfTt35fGR8BBOw5MNvGgxicEMkZjxcdel0aQDL57r1NTIXUtO
TXw1Na9FS4wtWPLmmI0jqq9vkDNoC1TzxZm5I/E0bMnTA7clE2yqtHIYtVMxUfyp
gsKpW55JyOqSU///RtoMkruVGsN+Xmb6gsSgEf2Pwe7sW+sQ1D0gS6CfhuiNhvFV
SYCo4j47sszH7+A31tc9W32w2jrVZdKW+BoQIrcjn8ptDmlwpJ2TNvMz6PzdJCHB
DQTEN3Z/Mvg/BTj8Vc+9OQQMkYLSMucTsBeKhrYDpGVbFqbXC0sSDKBIFiqbvEDZ
xaW0cW+jXCmMJMfYEqrzZDER+UsQ2jN7QU5m9kOaQdHGm6RoBqCFmlnQka2QqYdW
ZEMSuqbedE8O/jUgcZTapw6aqxuHHt8AxtVitcbQZHXv0nJ5S/MXwvmpKuhrQQo7
qXrsa6lZqYezIZCn7Fhd/f6RoBNTEto3pQSxzln17X2xcjfDHtzMYrNEawA9/Dmk
O/SakX/aHGsgnIkn8XWOCiR+ku2BYytbgkLfrcI/geMZIOk5ef9eFzz5jk7qWVJV
u4ClnvxsweHV0OJnV+Bc6N+gi4UBj4NIJNbSSiGiWB3llY0pC2cgKZ1M+MM/EAHN
/TrQ9nSAKDO+ineqUAVauXP5dA9TlNhtkZvZXyWyAUBw/fF9CW1XAurUbzAJSOSR
3VeeLGtKmv9BWeuwbepnL3YvAO/VZJA1dz07I9VKMnZG00/LWDNyojZ175KKUxut
ffPF3wFaFamAVIAQVwwfBOxXNqRyD25AzVPVG4Aidf/bzktszn+1ySDhFZGDGhy6
UnpvpPg1A2JPatU5zLlysyu9ll+9x41iKUPNtGj+cQYYD/CdiSjWgJkt2Z0/BlwB
4HOz10p76SV8+rqBD9W16d6ihQv1tpUhTZGtLAyd6uwsk7wq+91bXq86XIQYs446
traRGBeo2c+OYCtzERGNeksv0lF6cz5/0rVlLnVuwZgRNi9jQcxhZLG5zcJCES4A
kd7xtj4CdqeifPchUl5Bamf/AkxgojZKvN34vVP5j4teKCxKuC4S33JjDwtPgxHk
ONY1I5SmWsBsJ7i3xmJxSkj7pcHkNaiwnxEM73B98J1C3Y9GBuDvuH2vumtrW52F
AdCo9hMS3IH9FbfWFTvXreTpcyIk51JEC3/GhuWy0ObYd7TBbs8XZzSQ2FQrAEY1
kUyqM19KfeD2cEGniJuTUJ9vufP6j1xIcTESivKVuU7X59+RBai4dAQ3lpU/4Hrg
zf7zEEQZQfCKpM+wWLITkL/OUJB5X7f6key2cIA1oHQOwO3uJtbTxaudcP8HExvx
ZZmWJ6mW5QUr9sEvWFDgocjdkcfHaa9N7ndY5odDOk1ioJ2ReIIY0lqLPtRqv6xh
+0Vq3BZpjNIirjhOISb5Zt7qRjOAm1xn3TdoVvkjRRqt/Kx3oePaGrhJSTI/BhUw
IA4dchhoptnz93Xhkat9WD0iheasEdK0tzeGhPIZnQKelWsqCB35liGEYG3DJFgW
x63StEXp3I5n44h6hhFQuf2+ZY5qRiRv+pIRsXaxvwMe6kPdYzeOXAEgLK1Kt9zQ
H72PCrN5lEn/kQxR7ARakDlHCu5XNmoHJc9jgtNk+kf2GmJvCeWARJOsNRXwg/rD
9/yNmNKZpGBqBsvup+eqc0uYP2QfJTongM3M5NBlvZYCaGge3AmJPbEmRtF9DxJJ
lvITrBwAwhpPIWe8BFeUePrPo4RrUkX5x/km4NY3sp5S5awmaMcCnSK3Vty7RycZ
HUWpIkKySv7MU26kV+RRFmiqRS/U5IxD16i0DN5S+XYOOf4MWkN6V9XrQvXYh/jW
Ed04ktEpzJOS0e8ejIadWNo1P3JADjio1fQSGZKJRUYK1id4wQ3CdQeTmT97j/I9
LF5pvvF7DidG5EiSS3IatQfacOKe2ku9Dh8Q1//8Ze/JRlxV4GRvnM3GvIZOkGir
pBNx/nv58G/N+gMGUCvnUytHtHAR6eEPgzme+vrS4F3nHhCdGEK/PQT8YdPdakYa
db3ceQYw3cBaz0dsfx48qRjF0jh4/+Yg5pEHScCSMsyy2cbxgJlwLNJqD7bOPkGn
f2I3wVlcAzqUZN6lvWFXFzJM9jBNaknYsTGHXbEF8flECDIXMQBrahQWrzFTcn7E
YlL1QWq592CWvRCFfCjscfLES9n+dcKhUh4Ka+MnB/cbI0gcd17ljzaFYKvo/2aA
40OGiqzK9Cwk8Y3mZO4zuk3+d1wtKrx05YPUSoT5rjLFzVOdzLCIlGZv/gpQG8mD
mZx4AX7YRXfu3Waz+zBYdjK59oiGhBVUNNyMNoXnUduP6jNc4I1ljJPG6D9oESdv
1gyV5HnTn3DUzAA9K6pCQlNiVCuFisI1bbR/YN4OhTuiyi6FVNTXZK3EHmWNFiWe
nJW1dn6x1pdtbM7wy7igaOh+pMCwt+jqA7Wyewc4EmcT/XmwmTVDFsYBeXYuee9A
9mfDiulk31wl58wAG0QP/CVBS9NwFt9DZW1Dgtm+U+3hguCPpMMl63eIFV8iLUWd
ycN41CwMTpt0ciNsoT/G3bRk2rNbN+MhiLgi2Ba1MW9WSuHlo1Em5Rj548TK2jCO
iJKgMn2sqRj9NayoPfgkX/hCVQ2keHdnG5kDi6/NmUnM4prDzmMhEtg/yAaWPvUd
ZvziZerc3eaCwsygzlScfYm3b6AbR9/7k0X046qM3ReTjQhW+WFHswfqm0r+qRoy
8ZAGYs34hxiSbyB1o9k6bbL1e1nFP4jt25FG3dunc+TT+b2zWQDVrPESiQzcr+CS
eLzLdAVbvX+o7xs4GIAwgqjj1dHWIWBgXgml+xfYtPfWg202aL6zdMdQFhXMXbr2
kcLGJF/RIS0WqzDo+ZIr4G5wpubUTmoOfhnvSqlkUGu79AGw9nrp3nE1Spd9PCJV
LHHqPS07bQqm/HTsq1tGCzFEfalCTUczq37SISN0RrQYUZLVXzxmRuvyPjl31GzC
FG+WkTYps3poyCCDZjJ7MQwf02s/cdHer9zZXdyKnMHL0TyLZS4lZhuNQVXyDCT5
VkP362hTD42HoD0vfVr5NEa0etDcdkQjegfLiOVy32zL20EZpYZtbI5tSIo4XZge
E1kQ8R/8WISscjfO+powdXjyjADfEIQ5SEpJ1BaSCJOqgaaKge1dd/f5Bh8cTj22
bue402NUf/YsNakAdMzGCtOyZu4Iw4ph56EZG4XWLxZmxufoRL+Sh0JUQTBpZz4r
0+j9FaUaDCKEK+jizWbFOp0fH7bIWjRCrlzzqoO/8EH4p9XgUoCZRrYRvzborX7X
bCRuyptGI3d61zSN1r8Hs23eukIAHhGXYPof/P/NQJL0PC0tHFbZnF46iaVR3kPw
F1y2YDNAyxdsYTi+OM7V5Bg8CnfKuK6cmRj829SZyPz/rE4grC16J8UlgzneYW4s
l+BGehT8tQRm8tbv69OQW8Yg/kOjoDsNtKQ0jCF4P9YNSMjXWhmOUngO4qM8/EvF
Sj2Al5ubdLxvfXzZxqf76HFjHrbIWn7eYZ5oCSUoi4bpFo4uVZFvEli0AbQwafKm
M+xGYIXgVn4fBfuJ14o0bAO56gDef9T424aXXCSaaAdMEkvKtRtvBBf9yDfgZOdV
dvWeig+a4a5IMOv+Bx8u3uvO+2uoFncrY/VAuisIGSmAOh8zOueeeblHZOE8zB/N
RIC1J2nOMQBJpmklh1yy5OH6YYVqz1xPIJRotW50b4x4t2voRl5M1QkHu7F/+Vdo
nF1Cxg4qDo8h5fswkDCXhqcqrmjIoxp5IEiU7E/Vxetb+iRFmVlxO99RYV9gTK6s
Lg2XUJO+H4q9XsNDS2DFis/EjTD5/BeO02sIlY4XN92vngVHpI3Tbp01UAIGoDVb
GDRg3VI6kug28nUyvuHF1UoaIObqo1Ez9hgUMFPrmM0RrYs02fImNiuxybz0KEpQ
W6WkKANkZO4RG6IqcZrzcN4YbIZpmI8tboRFE2mvdEOWXJj1VkfqT9hV4CHhNmQH
Ga94EHwpk5kQn2mBGLaDwOj5ox1InWMhFNdLfZWGVnnAvhzQw4LbSPXYpk+FOUjA
Muig//t0U4cjplAzyk23UN80sG4Vmc4VsrCf+/yIo9yRLHzGkj7AkViygX3S0BfZ
MGVK+oerfXPJwzHOgv2zuReRD4KG35j1+98ops6XXrzT4DF4smeAF8bxfGL7TCuT
BbT0N88ghgvDryOaxNh7dtH0dQrog9XIltOHgEMUgnIRNsZrQbjoLgUGPoCa3pck
u8lz2Foouh3rEnkwGv+89dzrA0Y+zn7ErWjVsne0Kd6SrQbObLUdH5AUmcPNmW/i
EB3eUJh8YNmMQ1WWAQ/lc4vrRZGXh1wxwKr3RLwQD3D4yYvfudiDypqkCl9HAptB
yYpYvx3cvIDxp8cdOFtlr8O0mDgeY35RoP0NNMjGH0exwpUwCcelX5563trQ49wG
XFU1IOtiEq+44F1PXGdi0Lcni9BYZQ85Zc0UGE8Yw63/RM9ug8f1DLg/VXTqdi91
/Pqbi8PB9xsI+icapvaPcZA+kNOH6Ag+SzVwGQ1r+V9jVqBJcqt8fv6zhDm6N4N4
Xfeu+T2PV/c4Gkqi5t1eT0rlxvcuK8ypSvHijXTZjYllu2MnWWuAAiYYdbmn9/F5
2oeGwpGoTJ+7CQYyESIGUjnXrjZ2uzOpzHuRlnS4mN+YFC+CKGHuQRXzcmEdA4F4
+l5qCBzr3mtNs0rLrqC/UoS4bjr2D1GAv+VwXfYcZI9Z6hElgX85sE5qkPYogDGc
U7J64IXmD5XsbzegdkJcWL1uviDEqXl0mw0vBy5xfVZmhlcME2JfVZeqimondoJg
ax4GB8NXCLwrBwcoO/2iFFusDh4wh1fn0Qwd2h8dn9HuSHD/hd05E9oda9w6gjy+
SA7tngL/T/d9wUvh70L6iiuYRh347d6zJzoLE2WcwPTcukfIXxzwfZKwifEc3sbC
AUqKpm/tuVhKBr1GnyVRqO8gVeqdnyuL5dsqL70VB5sKaYdLjCffkc/441pAMIpU
4b2kvpRtkbERTbvwjQdVrqPMckiq8PKhpKrkn/Ejv7O7Z24Yolo22j16cWvT4qvi
WhqDgdsqkYeCsdWTT88zuOZMRBn0PAKtTSUIC28dQmIjnTYGQZrmE3Rj487YIUmk
g63taYmzudG3CInLwCzCSFRTe1O1bMp1Pzz5G6B7gxzdhQ2RLNTYtcejHZOsh8mG
pAQrJmcV0qAtFAzhx9gDdautNBT6LfIeCAjP674S8A+NZeRaWePFGRp0QrMi6Dae
sRgEsnaAV7Wkksscfwtkgx6oAgNm/5acTYEocezooOx6W89NthsdyqkTQ4LdDw8B
/wX49L1QQcf4J+icDBsBOeLa/L6C3P4FNygekMpt4fsY30NwGf4Q59NWQyLKREeF
I0u1CkBw6t2CbOeGq1HJ+tTJxqZOMxBVcMcHsQMh1Rs0js7MzmVTI/CV37g6zQpX
IELSulcV92+/HIzTMTI4kuE0iJU3jMF97d4Rnag+0rWFLDDr1CUhonOEKU0xvifI
Cw/Xxnk4s6yOEUkJtuQklcH/oSjBSwxeivCvgc5gykg1wvTcMXiSxGagvPhMIh+1
5QMj99RWBgcIzNAN8XNrn6F4D6aSoxiFL36MERVw9nKbNzhaeFRiIBzHjMA/ujBT
zWTY7BJPCwRHxn0GNQv8G1tkA17gYlZ2QYajZ52KcABEwQ2Ih4plzxr5dxH3uGP1
S1BarCA3fNegnGNV4Rk4CPBAY5Bl2LqQF2s8FoVz4uunJc94klMkvfZJZqNuChpL
lLRxNvYvmIP6Kgj6iiKZUnRUkaqqxwrR/9fhIay19sFNOsR3ncVz2gXY5Lx4xUxd
cNctLdvUUiChGQdEgzfiFxtAubOGKhdKM5su+uOicjxkpr6kmlrjR7VHEOXIcj6a
f1IwiOO8YP/7ThJFtiHwPJPrKkYMzTN5t+2UbDHttZJ/xyUc2u47XPkjkxo8QklO
7L/OUB68lDYoz0M8lWXiCYrUVszj3JgtRG3naCNC0nP6z84LW1NKMsGkowZz8eqN
WlE81YU3DkK685aa/W3vMakSP5FRKbGVvFFhqmp4uIiadki86Lz4dZ0l4+c1/qpM
ZEgU38TNXRTsOeNel7q2bQbBu1eR51Q/vfb/Ug9bZ2xi2W58PwXDV701YY/JEHVW
1IOrctra0fYXC+IVLM072KhjmoNWoAI0Hl02RcdxjygA40o2iiMGHccvz5tsy3u0
AzRrxZcXPxRB5b+3KmiUUJ4U5b2/0lxX02cL8SGiEFjcZ4Z/gl7kcG2Q/4m4/b1G
7G7LE7EkzU5A2F5CbauFbTnghVAc9zAfpAZd4uErQraJTFru01Vylq0lHCHmYoTA
Ic+rmn5yHtrPWBy9ZEBIFF0ToDDZuPsFBUoxwJNiUPaUWMXdPFlOJzsD9AobX1En
rDKdC6UllAwesgXPwK7OhLqwLrim8MTOAkAL2cXBVco5x4i91WAM8p/teCff4sIu
3E8Z1SHnT6KG6FNwzq8n4FM77QLelr253/3l93omiLk0V5pDXoIqy9gqdzWSg1iX
oHNol09q9smrUcvvkFFaYG8Y22B65muLqFbOzO5l5RdpzckYXs/sso70FScRnImo
YaqPTdrhz8++NIFvbhX50ltfcyrWfciJ3qtv7Pb72R65IPlZoLP1p32hqUNGJ2wk
LQpZj/X9HG/wTydtFwybTJ4ByQkUEsNjTdGAs5LzdsfnvGNu/WXItPqPIOLyyoYK
lm2EavmZB3IDoOY2xgi8i2DqwQ8NVISwAT7R9VSsAE7e3fvL9X961NQ3Cj4a6cRn
SabYHsH0bnzb+T1obkbnrtt9QeNpVhEsa0hmIF4ZC5OoSTLNn1/wwLW3MMBLe+5c
xkkKpMEOmVxxgP+ddFyJF82PpNlRmUH2EGDnvmz9cuYIQE/2MUCbxGXH7npjrjKx
HThX//divGsYXU6OVOKrdyqRMwD97Ejollb4RJMKGyudNtdhte7BaBwezAJWTbXM
cTJSV2aXz6Zuf61VZ8GeBpVV78sKECEFd7gmwC11DChM5JI573/JWpEKFApgsB0e
w/Dv1sXnBiJi309cpHkKXhBnOkKcu+KsaZHqk8ecbvwUyE9BBegFGq6gHorq7vm/
VSPECIyrK/TNsqiar8lzdplK5z+MmlYpGZdeaUjqQVCXpPZAxBkvrJBv9KJ3a2EL
L8TPl8s7sHYJJI97ydqq3V7oyRvackBS+U1RdzBJRcBB9BYOaDSSBMlEJJaHEEpk
i4hkx8/39Ijv+zLnRd6Pf74Nm733XiA4DCph67uvszf4arRomZ6bvAuCOuwjhgHT
WCIO5Dwn3iQeHpPQpotlPYkiFb912qnoErXxPK0WXwoGLzfCwn5ERczdBYJJPDZc
bS1cm9y55LBe+3XplsDA88YEIoYISUHwtxaNN0fQTdVwDwm8bbCpauk/9Cbdavl+
UmNIX0juqXFCQ226QGKAkDHsdt9rla0pONUFesrlj/UoIAHcfftwBVSdOyJ2oz4w
worqe49ESIm2e8WQD8hf2XioiC7VUeD8heX0KlaEHhk2j5UkRV7/Cyop6aW1sS+d
g9++i4yzSdvjNOkqadNgSiQ32n6a3q0VOxjuXFLGuuBeXx2k7kNhWw43lVnzgzaS
m4aDlu+TqzdUWFnjM6SqGTnl5IY3Hxr5Mnsmam6eG8dtbCQOqPjo4B5xZyqUAgQs
QV7GFKBefjpE3FVJLmCewfRJ9bdu5y0CVvEeZllGSOqb7lAgKyfXmybGLmPiy0x6
2DrtQ+D3Bpi7X0A3vzXGAxFax1wbEgXbOZ4iT49ARIKrkChdpy+E7wkrYc6ah83i
eyWbuzoM7rkC9jXFAB0ZSPSSBPfLGAqEl5PiiMsCModPsuZv62qs5kdxGzEQsDZk
+tsyvU90KNSSQbyxuvjMoRXiwwKAZI57AoVtvpP0T/wU7NPy1j/ag+Bej6FVostu
H1ixepk/5Z+agKvU6S+KtIFATMnP1X+wQ/A//pkjzqIVOhFHQjYRqitHD6/jNHux
m/lxMp8SViE4pipV7o/MUgJXDaXAasjPzKYKkEsVvktZSbJ26YV99WMfaB0u6JbV
Z4CBv1iq93LVCwqd44UPLuG5YrUuh7of9VY5xN+mSDhFJoqO+WmVHqK0+gZjq/HC
HT2mRUP1/hfvmtnsFE+9X/zXFvReVl01VwOC5gqE08bc4Fj4fD077HzVMpOgTOw9
0JpvRwvDdMzb4BeMEHlW02P7P73CtKx9H4lhSNVbU0S93wzO+bfkFs+/1vpmOPBX
aEPfwrFRAeqBMvCUUwJC4FihcnTsOncgTw798fImJHiYy2iA3x8B0FPrVSEkSFRg
olQtpVoGxT/kVnzSut4a+J08jeMyTmU5Y37FXVWAOpRO/9GqlM2cZTopbI6/TszE
+X3y5mMPQXMJLRLjKOkgoncEoBvEE9NAYAxxWJOgu+gQrCGuGZZMVZE6YiHEpewa
ma15hMVQ7U2BNKmiEmBP1QfU/nB/UGCzC2ji00dWyL1oN6toIrcDZ/VHuZaRHDJE
LLA9OJ5yVSH1tEFQSlEdc0nPZ8aroDgmz2Jk+hMkaYZbma0xczfgHvCFXknwQI04
KJZItVnGqllPNlHQ7HRylv7O2sFwDjjy+5HwkXFOkRqUgR+w68JRARQchzOs53GN
d5mNWOHslCd2+pchchtUPjpGbiNU6298WzVjEm7weh+3yBrgXcnztzk+hqN0P+4L
PD4XpdOdq7EuEqJrpDLnZbV9M7K6g2NOUBebw4H059iW1bUnDSJIyl1V7GMyHrqo
VGDQMDD8PEdF3sovX7WDPezjTVQXo8I3d/tzKTdFMAaW3ST7CExcHObwUdcIDEvX
vFcbGONhHv1HcWlbvo7iUuYfJFu5PTRGrsKuqpz7J8DGOAl/R4/ordqG00xt+uYJ
Wr17H3JcpmJBILdHgwV4pR5a+Sh0JC2tNH/O33fagwYk8lu+RmLqOKJzzDMo3L1S
nq5SWlrG7kCtSZBbPwilhT2m9sMLVlG40g/HcluWBzmyVR5KIxrfdGNey3MDbGdv
hmKa2n9vo2eGuu0BOMA6d/exFc/+0BIBmURhcmOgpivRSbSADFzmrwcMEd0XwjkW
UKHQ4HVMUvEv9iTwXrypPCqE86BeDORpHnRUG5qWt+Y7rJUIedyJgL7zPojPhQT6
rJ2kZFO4cPvC+trwjBWNYhApt7iacGcoyt90XSwMJMA0aYkSucEqcqioUSIFUCSf
Bk5Fqahye4k+A28B201rGNQT4Sa+XNSoqIOH8N19lT4ffxFSKY1SJ2W2/TKHbUnL
xH+9CHF+Rn5W4kZnkrJwdtwwroqO61dAddE6GD6n3euQka/Q7eg6iQGPZJ6nh5mc
VLi4sFcx2LpYDbqP50D7t839EXYbh2mQN5/dtR7mxQGdJi3i2vN7v+9s1nF6hEFp
/XYY20aH7cOp77qu72mWz+q/LY6T8yQOeCHJxVeR4CF6qzCyiFs60uByjwics6Wn
uIFwUBip045pzeu0jPAW8HxQvdzlDdl0zidWA1Wwh+cuk/dvJWI4DtOFWxqN8Yea
UZlKNUj1Y1nIs0Vlyh0nz7L4Z0yFasbHfAanFU6u+uIv5i7mWfgOMvnzOo97VDKx
TigtWVMizg8MffYd276HnO6CpWsoFQKIOHTbL3koL/ZzQ05Hfc/kXVpr3tTDNurC
YWr+cFENhQ/FS/Ja0ZT3x2gaB+0gH6OFAaAm8ifSVolkU2DQX0BvP3zwzs64K6D+
er08tNfBPQNi9FTh7xTZCX5D2xWlmgVCPMadwQU413scZQ4gZ2Nl6KqywBuloRpy
j/Ub7CpGHedR6faYk7YbjdDF524CJJ9LZ8OeYnBs28Qor6mSNtny1qionBSOrurQ
qoJPHSYWS34mu6jGWey/hDN+EdvDiyGTgXNMpYi+oW8Zvzb0RLU+1CFaSyfhM12o
ouS+SPD4Myfz7X3/F2wWHG1WtoHxfxLLV7vxs9jBemHHpBMuynQaPi7VhIwlAGFE
RwS1luvxr7weZejD2//Rpw65ohXcJIirIqTD5nm2IXVGLiE/eKX9y22tLOt+YK9x
IdvIdpR3GkIch9t0I+/JwZ2G3C5vMgZ+gdrwXSksx2r5MXEr/02dLqLgutzENZBP
kLr+21IZ2mrw/ZsFqcUrCtcUHFTDcafoYyWtLfzw/xvYKPW+FE+Zgthwxcce4Hb5
dS9qnca3jgI8VqUpvVD7fL289dsXQj6WUfsgeHAiD5bkzxVLaBWVl436uOwqHmcP
WwbSz1FbhEvsjNLhJ4KOpEpOkEiPvrtr56GnokXLj3oGGCR/ZGEXd9hO2+2QbgQQ
V4qIHRUxam2Zx7uz9R0tNx7bcc0TOnfCJwSuKgoB6n1yjRa4l0krs2CAouxYsK0P
u394RubU/xm8Y9lGn1cz65kfFwFq/JOHDe/2fbDcHa8nwgJGMNz9zN9d2drj7Igo
8bBzS8PHvMSSpd6ZpoqkcsCqw4zNU4VkvMIZYfSx35XQdx8I3hrytSF7bMWk5OwH
Ctm6ugvyuG3CTtHEuiFnXBDY9QjomI4bh3O7+2Jc5cmqs85vFCEBm86WgoyArslB
PNBsEM9Ef49QUcaa1QBYGttJlL1UH9YLYbET38rYOPzCQk5JypzdncH7wZ3CuQL8
nQ/y0llCiT1PcDzfeD9EKWDGUfjw/cw8oR6nkfCSRBv7UeicNakVxhp0oxBeHlBo
Sw3i8VWjqrii1rHXR6Y0UZ64PADCZnIbJDsWY4gcSZBL7vor9xbd/PqEAjXbGQr2
4FJszFA6VJI0hd/Wg6OBKkdguJcL3pJokNfSwdjWkxCZs8k5PIbSd1/HvBTB71es
6MpFnWujBqUc7O3PZBPDmQkkIqYgjR0On0QSYJdvZUCDlOu9BYASHGLSPAydP00n
kfgZzEbz9z0GkaIji8VkeE3cRnnT9WItU41Z79AFqUps9McQ5Iny4CV8siBhZlm+
mxT7plWxj5tT8K8GFGCltqviwzqUuQ/kXFaJp5hIPVN0NK784nnciKbexmcI7EAq
33A/+husm2tDnYGCZ7yKX7c+Zz8kKleIFtJp4FDkA8Hyu4sPtrkCuXN0Ik24iqop
SykpQ1w4OArAkL42A1LeNSFgC+eMjN8MtadyxM9HxOERjqV1Ob11HVnYWVQ3+ise
rBiiTxkH8IfETPIeNJwt2ybk197J3wZXqhTQIOCnth/7rrjMb7PP+jMJde6vw/x7
+A6++LBors1b2zOSinG37BNgiLep+QOEwo0BsG/4izqh7T03/Y6dHu+lZKtKKiRG
gPyarA7iho/nEfhKGIUVD38gBLrDeifly16XPu7fvxNN56gZMijui0hdClMFcx38
AUhS1ZtmEbhRryCyuSWSLBGdoDm2gTJwsNBj98gxDc88yMPGazBj08AXkktQ+/Tm
MCWIIE7/nhZUGufH5IA+VXdqTDzFNKTMnDNEIiFGDVvalslUXxoc8aNh4p4PyK//
U95SgbkDvl2F3Cfmll4dlB6PYtxEVxgNYy2KaURGStdmuwQXkOWoWsphhgyR3RQ/
n/x7nlqqaFfpApPwPcmoft27toWMq0sAnalB4cd/vTA/1Ji/mGmO7IZXQZiUP8Jd
WYlVTNxKPWi0uxz2TZIHihxPpBfKQX3zSjhPP9iZXjK8PLYS6674kKhRuQv33guq
uDwD7oqT7EXmWmd9JS1Cdpaji367TnPW+epeLYX1DNLrJURXhtwtcFKHb3wskPOM
mor5RIX/ojOVD9RRRwOo7026dK0QMhi7H5bb7mOWfYTYufbnidvbI0472tyWwd8R
T5jLazCCH/hzBcvDgdf9O3hljsk7Ycz2IRHnm6/R5YwLD6DrQOCUFXMCB8c2VOFx
raUk2gslRn+wldeSdeWUX84Xab52aiR4bzJLhe2yPVq9F9VYIQAkZLR3Yg//2gQY
OSkm1xTwKc1S8saZ8xuDpVVYZg41iw1QA1RB9DSfkQ/Fh79bY/ti50BO8LVRKJhy
xhO0JnhBIx3Vk+noeFYIIiYNLUe9SHjHgAh2SLPvePGBSsxwTIdWASJGgTcEq66G
aE0IpHr5d0msbTSKgte7UsJ9fg83Ife65Ft/mDh/P/gK2EODIDp8U4PiYeEKwQ7U
QZSsinYz5ocfIoT+QFDkLpSS2Z+k+INdhZO7AxP8mvsZK97MnVELQAT7+sz+JL8Q
+YcWkqgUI0qP3zRjkDLEalhVLmk96B/P5r9jSS+ImLJYU04ZbHuwQsKJ7qO1bv+q
pfyE4R0nFU8M453bns/DA9rSmcUc49JplT3YhC5bRL0e8DlBoXtRSsNejbKC0M1c
doJeX8HOPUcEty668eQ0ghaf6VZuSyUhsi4ggFpZpmfuXkch+qXacMz7M91jw+Sq
FVxoUcl1zntk5GCB0XG43/cSqBDs/XA7wEziH4ARWZr378V9evJA1vYTTGWbxIG5
cw1F1nx1LNBgY90UcQs7ZeaQFBCo26KQFrdOdN2PP83n686tZXFJFAEaXj8mpiOk
Cx3ScvoYq/yI6nsJvkHSCBQieHkKShGXI874yOQBFaOzYA7kL7OBFHqsDj/QQjjZ
lxt/STzdGD2aWesd7BkaaVmFcRZiHhnV6Uwurd25mY4acQa2TSlE5bOeM+8JrBRd
C9d2lzJLcXytjCMTw9E8aKyzu8oQObRn1FIE3R812eNSwr7r3uMwxtNJpHzAkaV4
Qyz6J2NWYYYSCb20Ttg4uuJoETcOE8IaYraCv8OoBKhcrilA8kjTqo+MSGhRCwb4
NWy7AWX4UvG9fpXTASb8ceKOqbBeWG3mYdnZQwDpZtC0uKNicMFzJP34FK4fKutH
2kvIek9bL/H0aYxU0ybuPOkf47woFzhPhIbm/OPEyanNF1w6Hab4EBbA2yf7db/+
KsEjemkIRx36xvvdqTXsKGNynYs9bkhhXLnKK7WMAgufDaXHodP/IXnuLS+SByl/
SiQ9weF3f9Vw0cvuImjKC2kqC54YBZaoktcIdZJgFmsY7DgBNeYvZU9lfle5j4JL
CeHK/35owKO5TbOZfNHC/N7ydtQCLd4GPZYFsDIDCaAOK4qofp2T3D7GzT2GQ2BM
UbwZJwopnkr4lOexhxJVkHw4MKVSU13xvayCuoJFRcAn+gZ3gKeaEHaJ/P3Apup4
yVSTafo47Nx2OeFaMr8Z32zLGznVRy8dPEK+v7O4Rzej7owyPMXDECEnr1zjLqSi
L9r1kros/K+2/wvrQK88NiyZug+BZs0+YWUn8ef64E6RqfQQDeOEaI6J/tc7PTGi
CSdwihC5UiG2ftnIBPahV9sWbHlHDLUZOw3FuruORJr9wrxkCsF2Yb4VoTvE430j
SQy8HDsnFsLdz0yygbP8cdT0pJI8WIkHWMoNQwYZygGtEh1WKW+K0i668ioXUovR
jH/kUjyYdH4KyY7OtFEbEO4ttVzcfT0GxZqmATcU0kyP347PAlfIvKsu46vtEpyB
ZchqCbEu1cy5kpjSdg39Bb/GsNcFQ3zbkeRZb6P5BObie91IK/d3KaAF45E/5Dnv
uNOuNyOIvG5TBqWG+rPkmDFuGXfSuFaS8wFBQ5GdVk8dPB4qn9NELGhRQ26N+Lr0
K/H3/wCkynQ0y/7c/yQPfreGgj6X1qcWF+qIMj3LFitFKOoX3MyPy1uY7PLpxEGb
OeYn7DQ2PYNSMKGGJOSTloabgu6Hf8t6mGfIGNc0gUjJY6YKL9R9g73iEWfnLLkd
LP+BlH4A6OTmtEkhSwotimVlgIihy3df/2h+Q1RPIp3izqD7cYQUh1KbCfzYX0aw
krK+Dp9bXGEDMb4IRxCunzdkYo59xAg3hHZ2N3livx6Iv834HSOlYhHwlM53tLF4
gFGZhCRlTVCfqVGnzBJdE8EoamPvQpHh0ebugFTMVT7prLAL3tn8xygwk2U0DeoB
dfLXrO804Img9ZCJDZ4b/odhRR7YfomzhWpqFGQVq+kQmFuhezNCcuLID5akeJnC
goXkW3oGBR4y5MK3PK0l1D6BH1FOSVTlCQDsYSNCvJBb2H7mshsGj1oZIcc7Qx/m
J8ZED5BSWmZ7ywgtRhk7wOiw5iLKbAYJ4Q0YxRmcPAmu699cklN1hf6Qa/gHC04D
VqOL3NcCqfDjx5uPlyMga25wlE5/2aO9iBp7vq/aXYyizPfznvErEQ6PxEyB2xJ8
iQtZ4sGGvIbdZB2ZpyDT5V0SLrAEDJyMauo73jeErumcLi9sHUIVum2AmFQIzplD
nrfYZ9VxFKKZdScheuCGMCZ3/mLEBXzKr1V2BPSUay2TTVP31Z6+IlaU3OUwsKdT
o5HVMiUUTZHFbMtfZirFuHt5cbk57YfuTaMaZqdjin5Q8y4akiaRaKMQP5KnK6ll
aBWOL/Z+Mzfwxl5fPW9/Kug+bCIpszgeBqwHi6WmjjA7481mVu+BOlMZJGJn54mx
Rt9+jSZ1c3y7WCX33WFfXY+Z38nqoe82Jf6H2js/4089x7+YbCXfWNTV3DFPPkH1
LNbE3hOjKzbASscZqZmqznZ/Sa6soMEwpRyKeUA4HdWGniCpSyBjauSWWxuVKUDr
Y0B85T7LFLsxWijf75l/XO0hJeXMQmsbBm049efAIOlULUa68Drru1JGvHEHnSX5
YH649yn9KRkuHGgBO40v/17fyWkAlcb6IsjnKma07aUyWxuzaF/GS24I0BxqUh47
lu/hlwxGlqlDMCQ0DUorZ54yG/IjznyzUiiTVgwpWe/spTVArtYVNrnYo8u5KS5i
PyY+qN/Audk3Ls7opBDKQ0kNzXvGlDXi6AZfLf/31elRoJgYaLr6VEuECpMu91mG
xn6wPyiF/tRn1Nh7iRBC1VnzYWrWw9fZ4RPTbQC3ptG3M96bm8deghkeVpNtM1Cx
8iSkyclIFf5gQDzXcIWDVxuH2msKG2+KZ7dGdoxkOqtB4nYz8W9FyHsSgGb7DeXi
C04CBSQIHCUyBw+qqH5MvbyuW288VVJLMK55b87uJ8F+fv/ejUkH9AReplcw96rC
xmBrUd6EAMGq9VbS+Ym2zVMNZ1WAEIzlMWLQGATAbTmL14IRJesEDnKBnD7GZa9M
rMu6WGlIJI8HToTmQoIWsZXjMJiDbTFGAjLuF/BF13t8zMtWLDWx4UaG+w203j+8
8nSf4vZLDjjkRhOJxM0kP/IhEAR5wlnfArBr3Dwymy9czmRy6MXNNqUfRy0YZk3a
ZMqJPnmcYiO70xxSYLpiXMtzXieL9gcJJ2g8RcZ2llCz3hN6DdoIYSzbIFah0A9l
EsPoN1INcjsDhHJpjq3zqzMvbim4alcEhcRARS4OrPC7hd1u7lTEvGkoSyruOWH7
o3dD2Aq0oP0aXdH/y/wGoVBxuum/QnX43mxA+Phl9tnJtMFOwWtqxJX5+1VqrvoC
HsBO5UjJvtbl5FPjFFtPkOwN0WSAhPy+NGG2JEXB/y+pRqY599HyySSoymhPyrcx
67M2PIHetiraE223S13xcRfKA3XBvlH+bmV3dk9pYIGf9gAfxve0WosFjwd7uWlE
gjl43h1ESO2fuuQ3+4t8TGvzvlfp8Z5UsYXjQ/ebd0fSh3h2/BVWjOPXFhKWEC7+
R1vwOBWyP/N1TbJh5SiEKmQs19h0t2HsYczywJvXqlJ0dx/RtDP8efqJhIaFVCSm
lazP3D0iKItOcJoH9hPR6gtJ+OBNVhrWjUDblQEclMPAuZVEtkbUgi7kFZy0Ax45
f5zuCk8z4LJkoVpvKy03eHl6AS2LuCM1CB0DcpG2y0r+HaYUPHNextbx90tonOn1
W8926DgzJ985qJvo4pKFu0k35lqycoG3JeVRxEf69KQGAtaNiYLHkhArbOsQPqLX
7MPSM1Dx6vvmBWkmsNoKFQmxESBdKksmUGJt06LvsQm4dCJ3ROr4HAE7w62vS8WJ
CWrB53r/ZmCoAjWh0N9Lc5ooyDLaAEqQLrIQFR93Aoi+vj5cjakho3HMf7rriMII
5lGTWsjB9YGOoxURBpEWACwUj004yeU6f9ZEIL+vjlmzRi48KNDE6Sj5qPxjyMQ/
usqG7M8H+tTxU6tcm1NEW5UZW+obJfSA1N04Uso3RKwPYiaTsw8yMWcRPKB3Oq01
BL/AH2vn3eWqdR6lssg6b78/7DzmPm2hHr9rQHmTSn8HgK2D0OOaxE7azUkDmgv1
oZfLOYns5sH3sdUoqWagi4xpPYx94KAODGZl0wHHuA+gYYWzZZkoLKwvdBJXxSfA
4ui/csPDBYzzd6A5yzhXycTkK2dGuyl29KwGkdCxIP5IMn/UENjaKgfFgWIo3pf0
TqpIVwYXbUe5U7xJOMY3oq1uL/45ErlV5HxrlwswtOLuPdYL5k2R6T162y7FMXUi
AVXQ32QF39etC2gHW2adudZVZsiIx0Nx4HKxvyzFYP/lNFExA4XZDQZUGapNpW1z
hhC7IB5m5sOzKDHxoB9Zs/Rt71ioy2wtK6hP6MZzs0a7yTxEFd2oHZPnTYXcr3Hh
mgB0IXT8yPd48rX2TZT16eBT7RT2Att7rQe5K1+AdznkzgkeNnOkI4RXBlUKjeTJ
A0HDwp+kvvhhrax4D28nIvUdPFEZGFw3R01uYXlNXrzRUfnsRCCfRzStki3pC108
gTV2BZKFuaTxSKMWIvZtkwIOSkdiPvWre43P5M0p7r1tRZnkRuNEsHOna/6aRZM8
eoi4KN7wHVl2EGVBNW2XFlZiBLNHMoytW1nCXy6LDvLIkrVBoJIYWYW46ikvPYDP
kIDxWUIGWgt93tFlFCe42VbbTCGqo+h+QgaUTMZlKDqvwLCuHg0mBbDFlYYi7clL
EOgg6HRGHjNVGyKYwRf/nC0wF/xq4g1f/tTUUehcMueV76A8H53ADSCpmZzWZlYP
XvFL7qcaMiHzH6sKSztFc8xTU6bNCgQGeIyg31YMTT9en16Mp8l0rrqrcOnBu5/N
Bl8PatBPdTHe78xGWgW5a6qOBbzVLw8MxyXd3FzjM+Dukhjt5j9Z7YpQ+w3FPJ38
98RBRYVvY4fYbAdUO1nPQS1v1mFwTOl5EwIQjsMmy62AGYbbybG1nRfsej8Yf0f+
vCLkPTOkk8BNQ9/nYBpngxNlc5JRNXgmFPH0E7avQnywGt4i9LwRPYaqVjhIUtaI
jHap47Ji5w7ttydn0fUcYSZq+upaWD4MolUgxjNIvNEcvkv00zjWrIxQdSUU32Cx
Cscdrwkd9HtTDsa0/o9YfUJNa/Uw20BmAbne67+bV/jqqxmMkHb7q+30aAburqz/
N5zT6k3PK/K1n+Vl8Y9Bj88W84/dGjBjM2ZB5Ipt3H7qRdNw1+raGulRENummOnz
IGy6oI+s6tWI9yYiggH1y7h7xCCUkpaEEzzmYEq4nUwUa3b+qQGDJ95XEQGQ+8zk
iOlOUwcWg5WjzRGQksVAvyZdz877vNyRZtqGpjXqaT3EBfaLJb+sC57SrOYqD4Av
n0jBdAh3s1JOYzTOp0CkY0TdYr6sDs0HL61kz6Ih9J4rwmSMYfUsy/xlf7sIkLP4
HcMTEv2qHg9uzv0hDtI3Baqt6SKoOCST8oq8ZcZzTI+UpJHf6rKWa+bIUGKhc+3y
7tCczaJMCMzygCvIwHqEKbARNM1ED1Q1v1ItJj9bB4feWN/t9NUkRsfsxcd7EdF2
Lp8cAhE/lm118ruaKvTm0OuVdfobjtFQDeQravALeZoE20xu7JaN2z/cQH/6ghAW
Vk2+0kJOqlqNiC87rTXmcqSw0yl3i65w67CS/7oGWQrBFXDMd68l8NX9VqK8G85e
HY7ajsTG7b/JdZMwiSd1KncIsS5Wj0XIkrVfJq6n4bVKOsvpW8dPGTBQwmmIkM6r
njo8jpUWzKNOkPGBZACFB50sig3r2exoPIGRwWwvDfCNtQbuXVXoD6KYHCEE2+lc
KTI50V8Lhep0Zciu5HwxHxKIteLw1L3RQXmYsF84k928TNg8yuxzIf8HXByDm3Iu
oMACfMtzQuvFhB5p8Z0kqNEQ+uhpn56fqFFsn/uEnAfWfyrv9C6j+pQuh0XAd58j
sSbpu32bF7McOa+BEjOGIJ76mmlPT6tg+grhYr7rClQWkPZ9tev2oPbTewNzqn3f
udcIdwIRCia81eLFyXm2dbnRw3rCxXCOGAP3DXEB9K5Q8LJPairrx9Le/aesjiBf
XkZdRdtNiJPBA2sxHIJchxwGNGM3nhzHqUht0Md0pup1ogVR7gQbzM1gYqJnJl9j
Vzc82ijPuS5Nm1kKETejuqLEqNsRW/ffYjOhEqEHd4c5eEc47nygcFE2kGYBxxls
AptNjzxaSiTx/khhlGsnai47UsoX0h9f7EapX/ZMGz/nGry2nWwL4KIdS+UBmMIR
tzFUawZs3n8NB2+Tv/OWfyIZc4gn7jnB2buJlpJT8SNKWyz7FPsuPyXosT1Zh+nF
PGt+JbBR1MtgJbA4aDBKN1VH2SMh0uOXa8/MOQ6cDVqJqfbVovXeTMEtvb8QzaJ1
LT8/sq8gFFDkXElS5DZDYUzUsIjuw9GaiY2/c8HVY0hdrh3xhlYlXOIhYcDynj30
8nCkRaMdvKoaAnjbKR77q88txUVmfi0NfXeuwf8hIAglxqeG6gtH3X4eDYW9nD4x
H7B/PqqaZ47/tmXRjJRtN+oq3b4xT5uS26XfhGxZSbJueOxFEKR+MZCiDh4QGeQ6
t5A0VezXvpPdOtLwZysGHaQCMvxJlrqtKrhTZ++wndhucPpzPv7X7CHg4a9WXfkS
BomfIWQynd3IZjQQKbOM4r5EI5jYyg+lnorUeaJ+PbnDXjlzSBcyznQEKTWS2En8
q30m7MqIoYHlMCeTzNt57xOYZTRCVsk0hxpzhL5EdttOEVbTwwdH6AmmrJom4+0B
nKlKBvEO9/gmcIYksVEMBX1Rotj/fWjcMWBycNp4W7FUu64hIH3YGUf6cvLod1fn
yRX8OhzwkCrbca5CFGdukFgO06uBc+kCtEyxFvYfoEieISSWzVxrS6M1q3SxSfaH
wlvji5gkP7q7foqODpvlajoSkGjnu9cnO2aIypRH8MmcH95Hcv0JqAnOUJiJFSY9
aBzFYSEDyfeNNOPgIVjsRAYlNu9yqo/GY1h4fVtdBqxIunYfWiBPQ64+Be8zZxq1
M7tWvMWUvQdeAcK8f8eHLE6/75S9ZyxUHknJhAWU/VQprEiBl2UWIj/xabfgTAm0
T5U9wfK1R7Sc1UXYMxPfxiCeWNx5gQgVxnIvJRpepRqUP3Xg0fceFHvlw6xptTdv
AeJYBn4XEigWy8AyDCF5IFJrREup0pmCBeIXq/yi3vtnf2K1rnDz3JKAApA1DBjM
XBjhXj20jOoentSzQ14KV+z57wdfU113RuqSuVgE9GYZUaDBCRvdsMFNfZGy7BfZ
E7RWUM/B/3iUZCuAxhMh/yzxSjye2S/O95N5mJ2EByECuLe9iqHPip1tZLkOpPb2
h33/JPf66JpMZ869HeR4TRNgCEsu5+sTf1P9YxVhY8OTGBYpbVL+LW9CJeF5uEcu
9NDyqnR9C2nOILxc93XmcL1iJGptcnV8FUgWQEUyFt/kDi/Vjx98kOKSKwBkIZpY
xg7Nz3C2X7/VqTAr2amS20zy6L76eufIRhBM1PSSnJyG1Wd0tt59wBvqetNPac/e
ZIhktEFjLnjBE9Z17J1DyQg7oeDlBIBvtGEWlVwDaJy6E0HcU5LIpYAZnGXAB9ws
mThItN7ETrR3gUgyO+K2xJmpF+p3ow7PAwFnsnQmCQvDYwFM9iysDcxVhF235PcY
70gmxVzan4EaZyQETVWN4pc3mqQHzmgjrjQZ/V2WzZfC2mTEy8cpEy3xVR5W7wpI
czP167AKm35FX2cqgYxaRlRcXBhNMk6ypPSx1UmZVOsg0UzvWBw00dH/WwjwV8M6
5cZxqXUwSKLIVXHTA0dpc/EnI0D7Hu9S56r6kYURzJzzPLszhfBn0oUcc7UwCjHA
/0dm9ZQzhR10H9yhFBhWUmq79VeH908hOcICkA/SyRs+Jg0iP5WdaxDkFST7wVd2
k0qW2S4PO9CjYS8qsFfDXyE3JxGPBYnKrRZNRwPi6jlJ+5lDv1Ae3V3gF7+b5wYU
RtRCMtbUgeoaIYmlodfGU4ndy/hryisu6qavKTyGC37zoYeE5TFL65CwnUkbaL6T
SoTK78oDW/Rl0hGR5NKyS4sDRe289uVuDh+himvYzM3kNYD3V+VqUPtq4aOrX2Wk
yCxkeaVO9YF8aeshsmEzKwbLjYUVOl8X40kRM2QIRHxSF2ub6JVQP6Mz0sn57e94
lBR2Q389k2nOEgAagGRAANaJ7glZpS4e46/tauw2QofgY7vTZ9erJSwUmE7noXEs
1sKNG+jromt28o1ojr13MmiaBj+By8RjvXQfBo1O6kzkx8JZaJx0Xqq40U8EqSHP
NwN7PMHLzIoDm6vpM5SLETozEpqSXPLMS9CJmsLX54WfLSbGMzltv4Vmm5l4pgoV
mKRI5o9LEwQIlDV/Hn+5gPgNIyD0aVPYgwFfFOwb/F9zG/X23ab9p1pg9jcTku1U
LrbOFwyJWQvb/rjXTO4if0p5NgvrwE2Q+bcEXrdoT+pQxumzKYA9L3haErm2JH3v
iHGybPOCWUZsMjTQPLWTnKPTMUDaYdzTGw05QFkXCpfJHv3eUS+nuvegQAAfQJpC
zFpsmneAGt38T+6DmZoHVq5MbMLAm5SM3ZvH1rMKZklldIAYPUct+0nJ9mnQgv5r
E/KBqcZoDLlaSbVnavwTbz64Qbqy0xqDnENtFwjdaRN2Udwa+ft7qgpuO0R2GivQ
UoOLX6lditVQJSCtz/w1LoqYTll8/cmhGs7LeLUHsUK6cGlg7I5i0QyUzwCQ8xVt
plgMc0ptUa7ptTvBwMr7NHosu4BWR2LDNaNqLEEsgJEFB0XRJ2Q00YjmWlLlE7Z4
GXbUDV/gMabVouov3x0RUzzDZKbCIdQwrV2/GfodaLNxE0Bk5q01uLeEkhw00Sq+
eRKEDLXuZSF8bvip+kaMafCEGIvGjaXFt/cf4yWmMgX1sOV1dvRG9NEXa9wj7Jmo
NELDyGe80KDJlCkktHbxncQQzq+ph6hGBUvWM3huZxBTAydyYNZtkUuDnk3aLxF5
PMAum45qZyZ6eXw1F4/ZABtvVamA9z79oYlArlBcjjMxO9ko+5Pf9gIztlkaBMWI
F5n4zMx2rBWMsa4gOHCWbFkikU6UEAWLP8d0Gu9xwFYf/5Xx8Jjt9ZhIZaudph8k
mlVLg9CWZyvapbpXbuzLIep4CvB62q8M6Q/R5ZvbfWuIc/LOwwFsgSzIsTFbvelc
5Vabn21KEr6ia27I/iTZvYm0DDodWCQTo/WLxF5nETmjo+qoBbtjn5eRPO9PiC70
x1hWBKuXynRRguLsaXsI779fFsvUvcc/FgRcmnTL8U8df5FhJM0hp6UgulVmHIot
ONwy/QCpYnZZwqH3at1Rs1mWbf3OciIoCB3Wa0A/JKPRxHjcM1tjU6fFrGKKbR8q
bywF9ODNwDEiQ7NVPee0WXgdKsDauBHOpWKAlkebVp680IB6qTF4n//CV2ETA+Yq
oisLo+EAKtQtvI2LER+8cgLh9RYXccVzfhRc5t7ReOMIZYihRXgaM6MwH69W6imj
K4ZGS3Ch4zJMKTurfRpByP2tkEVHUmK18OXd+6iqyp81A0HOSHF5pflfQ7dJwcdD
GrG53wP7Yz326VbCOoG+g5FjLLQ8JBp+t3sYljm6w8ooqIvL/yM1ZQYhdx7Wknw1
XyiGHKcaaDCczQe8ddja6zzzQq68TA2YCJcqg9wdauuOWEvZuZD26Mrbc0cjJPJG
NH7srnLve9QiLavHJT7XIq1RULWSymuWkVDUUln5v7VSOMMRnt3twPp6+/QCM1xx
3CHfLsOt5Tbirf5jtDaJo51wEOvGW1BONez1swjpiG0dvNzLsB28sv3jFhHyZ8Zm
AqHAvjVk+2PnGT3ZJ6IN7NhCVjcN9VxfLsQjeSUfOJty65VfEJJI9E+Edtr32lXv
WQTcLGTb+Zn7B5j75EnknT/9wDQBftQkThRK1Bk9yNPnNeuVFgi1xVo1rC9YJprf
2vXGyYBmFIM8qIVnidJUpfn6N/bbHbom06g9yKTZnjjYH4mgbQgrbi2sd1oMcT65
I/IZgdfRtXkdKfk4oNPxd55NVjrLPKfv3czICkt/AUHwZ1jwJd9gSd1VvMCHQX0x
cYjL+3raqVeEwlsiMsfRW02ncu4rTbv/bGAiHImsWPQGED/UzWC5NoCR+bXSNouX
SwvS5s+RUgoxyxDeOMU5Ol/qJaNz+ID0iATxAjP+q6C0HhnJSxqxxW7Lh976PEQh
yYAo+f5rmEiUWKlSlB3IaZlpopgQg30RK6IgU/rJqm1vPhYUVX21YUc4X3+VBMq8
TtPUhFu6U9ZR80RQ26yl4he8h3odYMdNNjcA5YUB96V32vqfvhPijvTc2KfTQGsd
Tscsvvfd6bYOb3B3wYnPq9ZXnEZZzzvCXvyucv7rB5EIz4h8KnvwnXxuJVZ5A/pU
zIDPItZpZF09QHE9LVSRNd01POBbyB4/g+GqVbxlyFwoLnxb9ltpwP2WHhB7uych
GeNCgbh7ZLNZ+gXku2txvvFZbkRAhBZwX0z0AahEDqcQvdh6Jz6KOE3hdKM/bx3z
ZMNtnHfH2xcyiybEEOEk6MaTtpzKBefyJzhjcOmymHPn/ZWe9Pk6y3ui5m/TWisw
BqLcrz9P/DtWb8dLLilAkqeK1ou+gzxWuesWp3lbcosidms48bvPQ4muHDLyGMLn
K0eEEfRI40YJ2YJtwrInB3JSu4NvDw4xIyHmMc/XW7yIHGOtVUAhklfgswvXuvZz
3QajKsjCeB214gviVLfww2zgMYy15QeLnIsaSPrhfePtkB82kDcpuYDRB6BBQP7u
J0aP4nR3RQI3TQJYfTNFHMjWt513nCL7yQPrpS2EJwqi23MDdPGS9jzRNLAJqWKf
XYgzF1Rrym90IVO81l2cp/lDggPExmHaG2DvnvyahztBst6cwLx2G0BaVMslUnEz
KPpaVl6sKRIzAUZy9dVBl9TABJNoVqYJdczx1dgBb+oGaAUNAinb5hK79bCa8Aij
VJlNzUAhJl2V1nfipqERObCn4/3a/1cx+THOIAaelXyKmmUgnTB0XzGyNIbdc8NK
ANyu0qgDZ9FxD7HvwYj7DKGnMiXMd9FGTabJH8ApzncnqRaYw57qzPFD+TaOYriZ
pBTKzQUZPnWjUIxNBoKm3Nu7RQkxu71aV08LFZDCUjMTl7SVD5sqS7s8SgBPGWa3
gDb4iXwZW1zNPyR8HKpvbloT2X/03rfJLAwuwEgGLl3SnT4/6bMq14AxbDgUCiVP
qgEBpM/17R4IeQgWJBXKu296abFHfAQ+Vo7SYGAjuRc3yEkbFT2COvAOsn9wTL0g
vzk3lgT493Aak7MYlrFab60U+ZmygVUoiX2+sfP+vzGnryKvZWOahckeelm7e/0h
SSCZkiuOTiQaF9fW0GY0AexLrWFtm4D4yYyuYA/5+XnNbI8h5HqWFStSawvZv7yT
iI2ihkMMouFzCzkJQuc/r9JQoeBn5xIJ2xYLe62XcpaMJ/VNU8vI5FedYXrg3NkT
vl5t/gcgE1Qq2RDFX/5XmcsDBJydU+A6uQatdMUhA9TlaN8pBIZJMeOCuVleJMBc
Th6F2bQFa0K8sMeXTDkgmh1jcV3T6OCMTfS4rf6gPsOquW0wH0at/HorkwPE4aPF
b2ANcWwYD9M86S+tZEPVx6EKxhjeeud8hu2C6H4Lnhi6tVuulRN4coJkg5n0OXSU
xEyTnbtMTuSXH4QT23f2twhSq2prUtUctdlel20jvFMCTup17lGfKswc6vl/dl3Y
7Jo0c9/qAziu06JuAB519a042i3sZTBzZLWhrMi2hhc1ydtbYJHEn4jdP6K/Fu32
LRDAV892WRP92cXGvHcH4L8cx2qUC5bqE4Xsbhw41Ji1v3uUTlswePCmbuWJhgCR
xe/sNmCcSJte4oK8mFL/FwuKrOIW5TkxapyffEHI8IBoC4MhA66sTzdq2wbZ+fKR
5L6lXJFi8T4drkG520twC+HBadyucHHmbkp/sIq1oim1Zi3Q3vUGkeV0dF0fPO27
2ybrUl9IpEkeTw98+i1zC/gKyrJyHeLmbF+Uf7SRjdj6US3FAZABNPhwk1NSbJi+
1W9FnLfGZH9/hFaewbmixKU8U0ntBxqEb+IEx1fIeud+8KD4BC2wNKqLz7mt/8l3
ekaW9u1nYWs6VJILQ5BodTT1QFDCWKRLml5J+Dhz7pSAnkJmA9cvcTGY2A/haxMi
xzVDco0eOSpevYK+zkdfqTK/br/g/LVS6blkF2FsisrOcU7YikrWRDohbdAelbkY
+UKeY+SqSBqPRgs/TvhpnJIJ3wRsRjxgu7TwfrH18+Rd1eNZWStf5A0eOFkm3JAS
MgCE2snjgRENsnc9KQKqui+mv+BT5Pjx9utcYQIyxj6imfsnXiI4xwkyiq7aBGzK
oQyUJCi5hHXNtVl0dVhLCntlCVmoKc6gD57Zom/+w035Vwzo5wqDVB6KjovoeO+X
yWEK2x3QReegV5orTkLc3/xEcD3vFuBZ22vx1H18/LxCJ/GRgsN6RxC4suR8oBd7
HGeq98PhmNYT1EHl91+UbS9iPKJiu5HK+o3/u6a3N/qwXKkcdHDAmfyFSNK3iGuH
sCymglLOyjQG011JAfeVQ0DG3TNG44Slu4b9IzKVXGe15y2tzjn3BAmIxTAZVQ5i
J0+8fvtASvf4bVCl4yOWEeKk8BZUU1rFjQBvsYpgu2KtlPKtsVwZwhsQUu8gGD9z
4HzuKuboXy6m3zQpNq1DqO+zQ1Ixa8iV9AhlLLEGD/3/2pU7cnIL65BkkwKt4ghp
FBnRjUg0AQ3hxveqDn/3FavmvKIsSjQAsczQ0ywWCJDFTVY7R3ooneUid6gK9Fd+
yQzfm+qmghaxdCwkWLKJEI9adKJXGtnpRqwKkiLYpOIJJmXAifGmhJcNO+M1aeBU
uzgP0uP3rziepxAvMGOZbA4c46aOFOhStX39ENNrdcDYtxVRT/fP0GSYYgmrLxRp
47DB673BAAVgrPQulpfezg2MBA7c/ZNDw7o6T//wOi8pVE/Lxd+9JumQkTNCU7z6
F4VtqU3iPOKFgAQg0TTkwyAGXZxj7aYwDx40WHlOQPmH1fNi9jACQNkFaDi6sRnI
8OiRcWxmwTZ/aHpddC75Awit+0yYnov1xmf97fGHjMp0NGGtktJJ1EogbOdggtX6
xqZtJjWgopKIJ7K1re35cUkXeiG/UprpQiOeFpyjFsU9jXnYTn1aH2qV4xBUg/Bd
Nx3rW0mHbXyzRoUhHgGJJhXQJ+4Rwe9v7t+cOkSWAXcRPfL3eAmUFXilxIq4CsSK
v8lqVBDe6gH5RgbI/kHmilw/Y2Z/6iEUZAdokbfBTDWbw2pivzYIDylvNUH3ZUWr
dRbsmA29sn7168uhpLw6N97b8ruUmp6rqNurmyjVW8yUpPKE7+320pa3tcVVxYtm
+wE/vEdrDnFA9H+Z6/Q2JYjJwBhW0v/tRe3urJw27rYQCFvU+H55CKqnQ/QlBE2J
YsjPcNHun5lilpGdOyr0rbO8CBKGrbT+OeqvTkXIX4jMmcZLJikkuUvpfMyWV/O7
/zOrLly5ojCOHTPnRaPoaGvUUbVa78iGcUrijHZYb6t8H+eel5QzQmV3pwPWInnX
db0oVruYWMtD9EuDeTDFhFA5d/zJMkJvlaBnXNZ/Gy00bxpR+9TXfe4Pj8nM18KQ
lIoNC2zcXXPDOQnh683i8hNNCcnXPV1lYnPmfXuTM3dKoo7+dGzFayQbQrH6LmF9
XXzSGW3GYMJZ7XfXVUpySyf+NkSaS9OJxfoNnXsfWsfUZnRHx4bZ6Z3CJbJXH9Fl
rxJHjwZd9+JtwRmJnA9xX5w1jEfEd0x5bE/CDHQLOMQSsO091pXve1kyasKIIzjQ
2Wvkf5ttCfNbPSslxScGdMY87YBQOX7MA3iUX+2aOxKxnRq4WoN0fRzN0jM+g2sO
eSLgQgPErqcgPwrDN9auevuZ8rI8LJgXuUxqC+41YUawaDaTeaLGx9KzMbHt3M37
MepFuF2OHztwgodSvBBtYCdt0+9lqU1/Um7+ge7eI0Uo5dmX9rFlyau7gpn5rrJP
B1TNiGKpp6NMn0RIBDAp5b9zUhnJ6vLZ/JyFfRmdBjXsIuszlD3kpm0CvgI1j/Qp
5dGJg9iel1JW4rM27PXHARk6WsHlWxxoYqgh95PWnUU1jcKdTS0q45IzJBECnRo8
MauGm3R49gt+/3HxHO3LmeAKPQtr028UaynK8p35G0bSkEWpcHakDV02e4Fn8zND
0r3dfEPv8+R5a7+9AQ3nPYdq3Twm29X/CIE3juS5V/6VekPKl8Hi9hsHed1fZ4Nf
6mVQqN3d1g+M+ZbCU35XOT1s4imM7qMrlrkPFqmfMws4XntPMf9JQnlm8Ryn+j9I
x6tqr66E7FsDT5HqaPU/hEvmaUhTAk5B1Xqzv8fzmAbCFgGqj25rPWRH+3A6Q78/
1MEVYVOOw9crtAqEziQeMGLAwH3f+p7Js8P9YKE93kMeCA6TMHa9anmdmUHaB8tK
bl5JSArdHKbyXosnp51Bz9SpnZtkSGrDnA+cEXQDgmmtfZRlc4vIp2JEqUIpkdlt
KWf9sMbvZ4NexxY3cDeNysSFYAo0L4ZJrhlkkgzS3iR2sRpQlM4T7syxXw/M0mk4
seVhOIZN0e4zsekqLss2jYjcC+EEoqVgOIt/hPjJqHCt7pnXVquPwIWjGnAS1mWP
OQY7Nvg9c2IWpgdyzllMven7CaANraA2xOdhAO86hqHsrQGRiLbYD7L0eCZBzL4X
E1U2vcmrrzrgqBca84OqaQhKUHp9RKq/Ork5U3zuvS6GaAEI2vgqFgDSucNo/D9+
4ClgYNmhJQPKynoRKoS8K4lXCJngWBmyPO0FbuLWA1212tpBNV3dKLaSnW5lP7GK
KrMMCbgqETuaJXJW0JaFhZGe+obnOk1H/kXUtAz4H0neY+H5YuXnqCjYH/DO/Q2k
Xrrk8GcOuXok5MMdZN6tR6K+IrDfnR6UIJwbj3n1Y+CZ8NWRqUZpVl976vceiB5N
ueU1FjLFYnLtFJRWkY4Egm8ILXsWaWWrcE0HreatMXjtuVi9sY9+mnpP0gFY7/lM
WY3MjZ1x0M+tWLFopPQIBX9IFZvKWWuk1DSKax3svQ3KUublKdJBDcZdp0Ju0MCx
A+roamT9Of+JkS8Ba5bI3XhM0jyKKMvVuQmBsBTDBSZbRithW7Y/DCcH9JsjHtGB
bBcLqwjaSZexekj/h59C/XVFN8o5f5GO6noNJcT2fWh/jOkTrp8mmvXgsXu+99S6
c669zderY8/ZB1AkZagJI6foyA9ESTROXJ8UVOEdoeI9yn6PXEYTNhPo1w1eN3ME
DgL49MxEjLRGmqnjxYl4txINEcPU7RleMzcc2ekuFa9lJR4KYmd4YqaI9EG+eZzk
90Ml0GZPZrSdGzScHmI4A+vbNJhtNmdfTd2RAHSZHx68mVaTCuJwWN+Az647uAGH
tXJN6oahj2NPobLUIruVvO9PeMKbrhJeINcmwfabmg0qoIuvtZSiHlli7T6vtcMS
gHSdrxvJX9QVr2Wt1dlzQiXUEPTPEn5mizgeUzmdwFzdjNPgdRi+sVAQ5HXXi0tB
xIjCdLHwU3kzeJUe11syt3ALODKVbptM0ypncyIOSSLNciDYmJMWUnHi2aqX20op
FzfD3Q5L6c+NZXMDRLucwpxoJqEN8s9p7IljKRBrXTncfheYBfKCI2H8/q9ww/S3
dLjn4AlNh5//1ZbzTEJ8VCzcfs5IOClhZieS3cx3wRM1jIEZiqLAXxIDBeOhxJQB
5v42ZnfU7TA/4KiGcVBaLgXmCLitV519p3vt3zcLAbogWrqoewdTgwwKvQ7wyFnO
DUjpumCpmRe52qbnBGdY+A+UhtvgXiqNgdEiOqxBMPvFszieLO3csphxwCw5//W0
GXmQHKurKwgX/jkvEfwt076i8GPTAhFuxdMhOVvppTbMCtLtU4AYrp7uAwvC6MKV
08d5aJq2WdEW8V/tFgZ+30uZjG92wVbhJ+NWAkaBuNlSpwt0tXGy8nvhu3SVKe0K
QZBeSzDI07/mk0UtAAf3wMVyGBai6ZhyZx3yL9QBj4H1F95EN3Smlt1uVbsj3eyg
Q5R20He7Ffj4SsnJDPQRUHWX9mMFcWWrPwRN5Kz0TLyWhQbTyIvd5pnb/j1ovFhj
rRFrs5VneA0d5189qb1MLEt6mUpGZ7KAK/XUC3vJpZBiSEczclbClrR81RjPLjZi
Fz5WmK8OTJ8hR2jnLKcAFUNM/2f44px/V9k2eD0Li+tQhXTMkJO/+7niRgKxkJ3+
5DT5M7jgluzxqaOThvIGUby/bKxaAz25R3UiukAHy+TOIwvPTbtE4rVfciAph4+2
6ZkCphpyq7lPdDdcLZorxDUzFW4XzzSorrU4PzVNajKWA5VUcS2wpplwdHFhfpMX
371dQA3dCd3azqNjMzst+TcPmZTNsnSXREsBN7TLtdr94yxEcHANhg7k/zGREQ+o
SgO5puKQu0/5yjSc4Sg1xJuSMedhhTw/dvevPtYZM9CfM1pMSR8t/+gZy6n9UFuY
uRu6SUAOZMKvoXEWQfgBAS00q55okDLAIyKkCYehYKNmDsN4YS+jsAcacALVyF9U
ttXcFD+8zm95+fKlBq5MHsC0URrw008wRtDBDqAbxXRWpTg5n7KsNvVpwJBI4Mfw
pwBKd0EPj3gg9JHzSSXkdxsKpJK8GvvoCYr3fBvhCc0/1ZCluKUp0qbve85GCGwL
MWOrzcvEXQXRG/NSvmu0cqhqGQYwsP4hywSisLAtbdlK+kSy3vwmXtF7w7XS/MkT
ZfgNEg/agG4xMSG1cTT5Z++6otgD1SkiY3xc4/wUIf7HFJOA9mN8uF2nviaxKi9o
oaiylHDktOkuLJoZ/QZLkHnyvimDMfy7uqKQVM8ER62oLHk9D7aN+n6h2uE6i6Rl
25TSQ49R9r+iuep4wM1bxcMOAvEvPQ1ktJ+RCVeWPIhphg1FblalHSM1C8OIzBqj
ORDYKMARLewlkm2yBVh+Dxj8wyx/UEoMEoGv2kkgywflaD/kBtXVNLI3dfqMa2o0
iYlHCI5u8hzAIV77vYftkC1HBm1rzWjLs078P6823sMAZK92n2ZPqABeo0tRnP70
m/wczQ+hKZzGLGFlDHl/n4DOT7a5ATzjLBdNvpjZ5UQuv1Atkq60dMGvo++r1DqY
Roo3nz5/SHbIQScL3W0FD5H82eJRqipTvgfJQZLXTzj3Bni9kFj64Vrx5CJf9TDQ
RZUsxvMGkzbV5JdYVUUSq+k9DZAKGANm96A9+mc5zez5bocqC5Cpm3YP9mvV1G/w
m7ToRdcTZfI8f7tdGRs+FvdXu6IZRe9A5vWbHQQhQr7U4XHhX/3qC3MY1hjCH0jK
9+LVuHA1X+IMPeFSJ20pbpMXvHNaUsNHLUO8osIfqpfPXMACioCXlEGlLbKx3+3x
A8CqOj1wCja5IuaKFGq8KK2wcRHWzG/s8d8J6i2KLDi4NsjaVO69H2Ul4NUH0w5A
vzFsXyUgggiV4TMqyXpd6AC0Grb+rnxM64M/RFs7/QqUly4gi6PWRp2pKbN9lpEc
ROBD5MwZBH+M8F3CmS3XsuUFAG1F72V/jpADD9/0EkQc57YzsMx81WUDJnsWlLBr
HTmeYDOgjpNJuHQx1ZdDLu3j+Y2qg4lMd6x8v+9ZA6V/ldDLC4nNbflztlEeyffA
EYuHrfwO2C35gyUgs9a1MXarSIkAOC6K3ebS5djh3GHFdhMgDoCeChXqzALpLQSk
vCLgknBYbjjb2j9jzgCoQ3zkNu5HtwgQWnyPk6378Zh1iXgLGj35tP6arcJyi4HT
Tt5MaoOzI5wHKtbwSFiDBwpR52go7KU/Yzhc8Kx5WNYrGA2Sc4m658EePOgDzCLi
LjZq8uairhMa1grLiaKRy3qqKRV95LLRVn8hfnLR3hTbmWLNIUnv0YG2xYDkOABh
doR1z/9AFfAMLeif+U9d7YkI+85o0XdgWK4jvsrvRbUzR3JEv4f9RCruDzOnei50
YBxUsoZR0Qtu+CIexGaJR7Q1dJigbelKwft4+eN1QzpcE4x9Ye4HVatxoMMwgapG
oRjkY4qBOHRgdqHqM0rw2kuQ9U3myPGdWqd5y3Fi8hlwdeOYF1LKIb2XosqetASu
1i4LgOwXRZgoTR2Kh2KatIKpd9/jdNkHpjjrifmTUZvG6WjVcaXDHRnQy672ftzv
0l4qK/a+QCDU1krMmle4LvCBqlpz3hDwrGmAtuSy7jfIlS4EXuTj0Iw4Q8n+jm76
XtnR5pyKYHj0/QM/BWRJqvFVusejxE2IJGgDWFvz9JhYOZcrd0uvhbfbNEyvI/ST
zgntgdw/LVQuh8RkVk+i7Uf2X9pb9X5epcdWWAFpyVJl50DYnHKDX1m5Q4f7PiAm
oVzsNvsHBpE5DUfPDVj7pMpLnu5hzDqFMBclulGgsdUKAdIdzqZVGJCMpGumwDzI
cApG28Ya0QFh6PS3sPU4mTYTxIExO0o5reLQBF6J6H1Dv+7/ze1jY3zw/joDoHtY
31KVnxmOxypVrL3zEAWBTCfYv8Se/NLaT248LyIQq/vnpyQVQe8/rTrSCxBiHCMZ
+u69/7GwjmtCpBI5cJJ1EWNIXLBgrXiXJjl8tywILW4pmBpc+zOxIBNmomnxS8LC
NO+ItaoLYpVRBPm+u5fh2bgzYCrSj30X44pM7Dt8CXPTy6CcLqRxOtkZOZEKC7vD
QJi+IpIZcTZkuhXCyx5GdQHoZDPa5xxhkce+whQMxk8Esb1SNyg9jVme3u2egWzq
z38b/EBj2urxIJ77h0+Cb+JtWD3WVeTCMXhRHDsYQaA0eAxDQHZxeuiXK4rqbRu1
ki4YJjfapu+HRM8Qt3ijd8y4qfua5AQDQeHephBw7hDSUXEw3glPP25TgTqG4xbN
KEwo72n14s7LBm2bHzCsZoEvgqEipntKjCFtAAhBO0y8LGkRovIVl68vtZo4gjmN
dMkMyaZfQ442qLLcdcmWJrWr+Ngw9ZCfIBXpUqBAQEMFxovmNKKQ8msB3DKGMbNR
3ghFl2T8vkBPzfadVvkTdVb04S+tjY8IwBQ9sxdnzn27wwb4ygi5wb2I+2SYhphG
6V7KJrZbAY4EYiGIeqPbDmLUZBUpsMjKo0jdlPAys6BxGZ3buE7XDIwR9ELs75EG
xgyem1ucpIcHIsldpvyvdsDaL3mQYVuV3spT2JDQa2Ge4Zi0ieUA36WMcRqEnmSz
esrjR34Vh5Irvzh/IthkbQvLgIGxWmaplLB7egWOHbqWOntA9QLCqVFTxWaHDppg
TziJsLVLKChIAOOg+SKCsgm+BOCTSsTKdUO1PxGUi+2gnmFVnSQvL2thSs8JYrTj
WatsL+fSPR/EnSe57P7UEtHweZRvt1XKur1hcsylNk6UU0aV8DCE2JlHTq/3tAM4
tk7+IO0U3aLlW23PkYJaZs7b0bZrw/YwnV2FbPfOaaDOMnCmCOAFvwk89IqfagHA
RZCd4WxPqARh0UsZxIXf/JvwDx7dvkz65WIXGTsGp2a4+VJitSTD2J06b0TPgWaP
mWea9cx+ooYv3+gp+kjitIAwSALUa8ce9hmITmVzV31Aisekb0lvr89FtOFdfD+5
vcjZVA8+heQdZNifkNOCcbwcK7uv93ef6OJDGUOMYBzFYSO3dGbtvn8btPIzpUad
2ZHal00cbG3Tr96uT1VgVDDwF9CV5BM9bcBfd2R04da/7ZEuDQZaPC87ISpWHtmY
FvvXaaM2T6cP/Ny75y9kIWXuYZiOPQpGS/S7VU3x2+UE3NFsrtMDhwNwvTneHHyB
HKtYbFfkwWh6KA3er7cq220u8AlumzlPXUxU13RNq9XWdXVrlhshq4MXjwbNvg4a
j1rqG8NDO5HXBh4+zVfynmyHJKV+h0MlUc4Fg29fTk4KWq9BewYm0MpPXBtFDVu7
+/yRO1c9/8i/TktJciZzeOJgegUNS1YHaxq72R/n5K5wEzvbx1imcLQ4PzoqH75U
taDX589G6m/v8sV8o53LOPvQQ4FEjHuceujGW2Y9W88aH55sF4qiKEWRq8Cjo/V8
/YMNPyDxmWJtPOzfARWuGMdgsIzMjpJ3zNHLc9WJogp61GpmNkOD2jJoYQ1dLqtT
YAnMX3Irn+yR4DpHlZVW7cRhXRjy2wYAUkoMx6l5ZGPdP0vAsdJHiYcYxq0/sh/i
7Sf0O3ybE1m3UDzxZmdg6aU2x0/qHrz/DHU8An69WQTZKmEpUGdqTGi9xsYGiKLu
+ELbVl+smfHPxLWF8yn8IjuHG+RCMLTpSEHyVG55mMt++kducaL+24kEEs4Vf8wQ
lgMNGQ2/1ZiNu1CVihTmUbL/lcWpClAS/IoYAaS5SgXYAoRYMz3vpxUXznyjRgIa
K8PFl0Mkpgf2r3tmPFTVx6qGL5bGzVRpMxcMaJNuVx1rMvGMNsOZxDLhJUIcGeP6
U07lzqND/i/EbYd0ruReXkNS9lcENW/K4fZfIWG2rgNulNpn0VO8i3rZLGjOwZTD
yPewnQdCPvgTnplqYvExRsQNeTqz6XTJ+2rci4l47CJsdpv8/CG1s+kfqvmUtuPB
eS/NVJtkY217X5fPVZhhyJ0TeY0qmRZrp2g/UIWOlxbD3zowlM4ZFnIeeaQpZWF0
3lQoEMoTMjgjF2ZjsdwcdoWU8nolcKljK9apI4i5MK0h3L0mJikTFCq0fbccPeFJ
Q1iYqWhmS5znk5TRazgGUjKYpY+FLtoJhfmqMWb9oZfzFt4tONYP71WEq16bN++i
wm9eRAVWxhIYb8xLEs81njrke001mv9fjc6LEAVMWLN+s/wGy/tXXW3VhlgmZcVI
7IeSSBkrJkEDKX96LXYkMyh2zwIjlJpKqQeJIbDA985ERiFmLaEklckHc7hp68WT
hUbk3tHWuwPmdc+S8ChCounQkUbrmVhaUNCTmb4SoWn3rs/ApNC4ZOZORg/eLetI
yRtN8veEPAPbv0Ir6XiOfXR7xXtDs9iW2QAv3e6CcUikROkLxfMETPinIM/15Z50
uHqryZRCyG7cQ9X4WqpJlHm/PUKIv+DP9SmLYyAQt9EfVC9wZnz6MxBe+WWihteV
lGij35ZpKSdsUxHBIy7A5EWxzA7MQvloZV1MUjfjtJToVm3qZX26tVl/Bc3c+rdC
ptreI8YEZ/AwlzcyqsS1SDIjxKBiNL1P6wU7r0YYisC8Dq1YgRgZdaXpELtZGrhK
Zk3W13BLzVHfi3Qd3O2EufL1w6mriwZ0Cpp3UKyy6lHfSZ8GFCS+DAaHIvwLxUW/
qJPzM9ib5HRxe7bI8RYDhSmG4MvuDpwgQxeOOZGH4SDmbqopiIcozHn0ciPrvOsn
JcWyvK+kqtd+u1Yo0gtNSGXesrfQ3uwv7beg5ikXdUXoA/+5filXRjlkzkA/4kV4
tR6o6REwpbV4u+1NTcmQxo/6vOyhS0gg6uOLcJbj3/hKq/9SinKgp3pxb/O2hb2w
xHG2i2zYoErEkiPiod2rIo6haLJ3JxbWhvt2sKhFvCNC9/O0ygHc0JDBKigVIYuK
XfEiaDnOMocZU3gXfC43bidWdQxhOWYpXByKPniTimkMk4eFdN+AOqnCvB/3YRQR
rm2xQOljXE6IrbGh5lRamGgwJspiwOX0ZGWQA+4NfO0zElkY9I6cC8s2xTe2vtKl
Wyf/PtKrHuXSjcVvvhkvc9+EhrKVgbqR9G+BPzxZu8QDxJudK58DvwWiuHuxHa+7
TlDCf5zTr6gDdabvge89ENF72WHZ7+AI4YrZk/eeBJEKB3hJU3Jv/8GtLuyEFk2v
YVLzKCeT8bNerpzqkXX2ZOPhbPTY/tz5eLZug5DRlvUy3/iDdZgwbWLU4pb1GHk0
N+6So101Z6b6S/isQkp9x5wvAwROxdy0ZofaegPtSjIv7DEDnKpSpImbwvinP1d5
wLg5Kxu6Vs+qW4TeEXGSV8xGdhb75xvoMo702srXE21zdHnTOFRleEwBH7vCi3/h
5rHVamq2umRSyhxOAds5nqZul1zvsrRkMeT0JrwvGSLF6KF1TlEqeEcwEXKEYCro
ZRmT9wM1X7cLFnm/G9oE3PGD42d9BGKd/6uewkBB/3ix0aoUT6FFSmHFceF9YfGJ
lambr8stclMV9j1dWPuVeYQoZmDoZpC88qpLiT4mDohOm5WlUgVAqAuNQdhwydWr
NnahbRvR0Xo4m0HIv8HMQp0oItg2Et2bCVtpD2D1QFXqwuFcYl78S/Oor9FxIE2n
I56nxPah8fczAEWecdYAjSoTxw4+abIzgzoNrPirlKHESpmk9l6ndGihHMorP+kZ
2b3IG9UQcRUx3q/YxfR+M6DGc8O8CaBmwhUhY3SMg0nI+9jLqSfbZ9bzd7L8a8UX
Ebovvd0A/MPwRF6AYsFsZMlMq8qidNI9cgSQ8TM9TNQygjXiBRV5TKgvXg2tsAVF
WUN+DuSlgDFevN/CcCAqbjFA28ZKbnwSRcaTacss4HNnal3tq7L42jl69iL/JN4B
HDYzNCFC6p+R4mjoHNhGM/mbSakqIE5SxbHwb1CGK25QLGaxVhu3Bu6oe6gdpLO1
bS4hHOgJL/5mqqSPmjyXc7ockg6c+RfpGNtblmTSUZIOi7sTu0jqkdRuhjI0fgZC
eMwDcD1ydGKTwkNQAKHUZUq43y7RqiEBQauSZva4FO3wxaTU7lst9OC3zL/wz+E8
HoU2cbzH3HU1GmhQPxG+l1g2tYdNbJVpij1lVoG4bccR+nlqOIItDZHCRAuVQx8q
3lQus2ODpj11SuO64y9B/DGjRCnMVZ0DJueUdDHiIhV09Kcy0wQQGtbcyifvGbcW
vBPpjyl1YLL+IURi6xOCdY1vAgMa51rkDbBKNTYgdfyZHUzioDlBcATxH9V2aXMb
A8+MVWG9JpYEPJtE7wm3jPe9jHz9v0sjlV8M0woxcg7HG7ov9tYK6qSixrIlP/cz
HioZEJ8+7UEN3iiEI8XGLYnVpufYLht08h5W+qCGDeTNf8L5ETPutvr6KO9wTsfP
Ml2EN2f6yeaS7ihpn6oo+ds4v19TmJQFqPSGBbEGtoG9mduuTWaBa0iX/pYPJhOm
4jZ6RxN9BjEwKVkz+5eu662HWZT+3PuJKkwJhoI4cAwIpuXlndXoFPMiJyrC8MpF
lX0pWvqrd9lZaZ+d6FQwbKs8sdU4Al2tuEn+mvoWFigycT8cnraGRnm944h3Fx3x
XqAXFQ+flPB+874SRP99ajQkrYmXKrlbCDT16qVjKBjwWTMVCd8r/s3M8b0hUYai
AW1fjCajejFC8KBf+qYNEKRthmZyECUPYsoRyOK1iJZbRbrxMWz+nRlykCBKAXFf
IXn0xVsT1uH5QVlzcmS81Romx4AYogcp69ZHadYSaghhJLy5TpEng1sVSCUd7Qgf
s5RQIzjlesrS8Ekf6lhGFE6Hpvitt7SORmqs3dZwpy13JVwWFAs6P14gXRgxalTh
HYIqi22wX90xAwAv0KMUZGkT9MzO6xqnK7pR2mRMjUenhvnkugnC1Xx8m1yVLHv8
79IZuG3lXqGLG/YaIjIRtAAVMIDGIiaSLk+YV0J2Vl6IbGo3Qaf+Fvwgkn4KVQAb
TGmR+Kh+5Ct2XBJ3Man3Qun0LKPEXsbGT34T2BgG6ZhMylBnhTGgMMopcp9pHhIW
y+WZaM4mmKlAmVvwWuikzxTO14Km4Zn4MXDLVoOZBD9YtJgk/O2riEaafacM3XTI
K66thzuCCUPeerYdq2R/W8RFf0iwgCpN83rXaLh0F7p88VwLQk3PEtm3fmMv2JKP
IL7vlOqCA9iZF0h7l5hRilAVful5MpZKS9b/NJk/SS7uy+N6a0Y90WA8WOxZy99P
lPKoG57QR3SEUUcL4akmGnBbSxoluD9ekUzitFTYwELv9WE9+mCWhxLLNqsmzeE4
QX46r9ioMLOzh1p3Vh7x1XCoynHrvhFeeQ79IalYGuKLYAMV4Y+RdRt1d+4wVZ1G
S6ZqvVINGubEkYUT5qqfCTy7ijGxZjDl4slc5vWSXVHl7MkTtyJw0w5S784hmF3G
Ltze4jjyjAhtrYq8U3DSqWzYa65cm6ZQsQ4Gq6jksWuINKzpu9T/Kw3OFEy0rhwf
fK/qlI1KZUwtwiW0UAfGYYO1SZZ6C+ftvOMrGnb/+ojWZ6ck0Rs0kN0VEBERBEAh
33nwXCzTEStmFWQ9QSbEBeCbZa7xe1ZLisevF14MNlkTIZ3gDX6N0DlAmogmbH5I
B2ctanKNwI1n3s+O0qiLNbKPOdyMlYa750X/jBucK+OwAg1Dlu0DA5++tSqZV6J1
2Pv1y856wR1b1xCF9GcpyI3a4Itck51O0MOZ9hk6GyMqNosqudoLCET3n+XOaFlY
3lCOxxKAHQMSFnjbK+sUMUDYlYe/R9zvhJPlZ2Mtf178MbLqjjHf2qLAGAOBL693
jh18meGz9kXPZ2Ru6edc06yMS2HOcFtAfNhxTGHS3POSCytBzH3xMoaa00jbkiZs
UVQk60wNjyoFHbTo54A1V8Zs/88CURBolHJkPeqK1TjXdubiBG4vDwwGrPR2KM/g
23isjcsL3TH4Ytclpdc/zo71MvhDvqOj4GQSsnvXCdCMHyJTpoMVqDUDyBHZUl/t
F1LEAemeLoFIqzM9FqnB+HNBAlIN4ZyskJwOyOUlakTk6JQcph7MksZ3VN4GS/d+
UGw/gD4wVSqeDMukohkRdPksFWL/L40EkqcyTzeUc5dVyVM1MWL2VnyCt6eNmCkc
3yGBdgaPFb2e5oQW2GOeJCzVbui8VbZfSJXIv43qFUEN0phXVFZmQoGxMR4vW5+z
YDKxJ+sf6f1UpEVttyoWrrHxo/67Z++WLl9r1NsQ1b/10Xq1SKblQejWA+dDW7QG
n+OtqcJIheH6rXI3AlSWH5CjulWmfzsb4zLr/VFCzwRJVATuPDUKkEl9ud0ARP7h
MrE2xHKYC2Q80QLukuNUHRKgoeau9N4SjuTWoKjjyKRWN84YORluFdW0iCfHtkpI
+EuAr1+p87cvbK26bDEjJegvzwg8mJ8/Oo1tWCfg3iQxSasu205JrnWrsQsFPcwj
J4F5RzaShky7lxa3FhGj5kNLLTLo/sII0Tp2ctTM0e43cBfA2ciJEO3HrvnANlFa
ht+a4r7uyeW10+PUJcCQFFrMrNA3p66FHNvQ0gkI5yS4Zhs1H72zqYgWDxy5fF+6
HCqmSqdladHj/9HKJFwprgWSzOGNcE3cmaw0fStKYlnIjN/ZhpG8ejOYMe5Ea6g3
Sqakncz7Rb1p6B3yNcZytXot97KXTxY7WDhsqDua99C10iVNtrUsfkoYRppkI/Xw
UH9gL3AS833+dpiVlIs8uCrkZVweveJbzdeqe0a8MpyO+wPlqqfcjljLNjtczSfb
QN5lh9rTgzpR3nGlZXr5WjqB7iFwl7HGF+uX2btjEwcf9fs430Q8FtS2urk3jLyM
Ft6i9QY9f1y5xejw0igzuRSbtgG91mzhUNaOO/eRJ/s1NBkqCnqVRhNdj5WgaksK
0/IPPAHeZ01RcWoK9wMpqst++s2bL2Xv0Tyr0TolNa1U/qpxEVPYddvVlPcEQln/
FICBMmxCRnxM/hQKkNCInPeSGdnytCigxF67n7zmRkJbdc5njhc9g1hbswsB7Y7P
IyjdNiq0znbDwE1AmrMug2qDKFZDKhlLUKdGC//ADqcICl66chrZMap8dq8vI4n1
hmOBv8+Ls/7gcHjVIsPMZNmPV6v/T+5WzbcZ+V/6fSZoEuN/z4PCDT8kXnQNvWP1
5nEf8h3OXYiJz0weKhYpd8dUlpSSBeuFBr3HZLPzI1YAs+lXvm7R2lGXTfcdcaF6
nc6Vz4z/TYjJR+eQwN5fGjykF25HKx8D2rUE9Fd+AjQtLmNWJuSc+VgcfU9hrWOE
sLmHWlsi6h7rdihhdJaD9GSqVepVLz3l1qrXKbXhl8ARG9St6IySjHZn+sCw4mW+
bv9evnLJ8D7cOJGrBVNu+oRsSbYK3vEfKtMd9rPmXMvkageRNUlscroiUn2BYfXY
U0CvaMXCsimPbc28UsAve3nezlz61tKXeGfvCO/TEngm7ijKyXqNEVr/AZRg3cM6
FXsu8uzKmuEb5qnyYGC4UB7bilmNjpAb3INJ7fzKHPRwzlMOAKsKER7qgF4fmTTD
6wm+gBLunPRl9qgv1VO3G5mnkg4tQQsxf8BGxClfQCZDzq9lyHL7uVnxrVLGFgNC
cHd20PiAKMYRKr1ncOxHTjH8RQrL3U7xUnIkbJBmUyQF+64Zvmpp7BglhQ9o179l
4AqeYIBxwrvJ++fuH0wAUD+OvCQQzwgyWJVhh9auYL6xVr7dQfvOvMB8EEV59U+b
KGPgK55MK6r+uiIUWw7ERAw4wivAZ4MqI3fUyAQCCh/gPqhXe/u4stzE4lSsqYw+
vXgrsxIJadlvLg8vaU0n0i21CYxQfG3BH+1fKcttxehmRA7ZHJ+RGqf//gQHuvbL
MPVINOIErJcPzYJdogx3O4z/Pqb9K91uwcRKGcDLuDY+QeOkFqCHDK15tWVA/0c7
7LbSSdZX4J7PNVZ9TKMDiJrk1rP2ivBpNfe9aa5CheAgZ/ffbbeV3oRGBjJPdXee
2gl5mrCxXgWWjR3yjYG4RW9M2Rck1QwhPM+nu94566X91hZfQ//oDDc/AcEOyiGn
qHJixJHiopP/2xAp0NJyHMtJdqe45ej5NZZu8n95nJOunBlp2mdOft/SOC7rX9u+
/R/k78fWhmM8uu9Rtot7dbM9tnNg17g+wD6ZbEY7RUInzlsYTYih3XGAbSM9JKv5
VOtojhw43xPL74p0Ogj5wP/qDY1mxLOc7Hm+pJMpFCvOsJqyNBMQo9rjEsWX/Lrr
BnERM9BvMquJtbKRorwlpj88467+R/jdMwJM4iyN66fxMykGCvQmBq7a6ACD8FcV
+cL81WtPgyyNbT9PrIWYoh8pnYVeP9qUWh0cGxiNZkzy00oUK5tBqON+wJBx1o6Q
F/i9huO8/VPb+zQ9kbiHBfd27i7E+WeR0I/GH0cKBoB5Xslsvy5rmH8Qd1B6BSod
LdLGZ8CCY81pF6uBLBi02r+KFI//dn6CwN2XbOmZf4h6IvTG8mPwqrszjy3D/S6/
0TM4jIxIHU6TtlMmhHsqrBo18pQmzWQd0HbLH1yKQs2w9NPbRBV2J3FNb/ov/WRY
MKmX08AGnPbaYLuWcAurLAnvd1vJUqPoSGsW6TCgpxBEVpjKwlxcXgQ8p/xCbLij
1Ay30RMDFFOaiU8l/y+V/9Gv7AZbtmxkMUDST29UHJeJeWhUzzDnwR/22atmBmuq
QK90m8hUTGYlWp533+IjM6EZ3pxA40dPutPK4iCTpeITP1BtDdGQlm+faAgqNbFT
elF9lYJd/lpZ+OTnIR1NOi4cLAhEyHcapZJLo7VQyfhTarbanSvZBnFP3dGlPj4C
yayo+095tNUVdrCehmeCVfHheffxhI4egiFcQLRsiOZfjB1pTJhbzKbJDnlRNGhm
p5m+JCJAce9rO7729SK3eDQSnDs0KU9jPQJQAIIlCmO5qooLt/9iFDwt+waPnBlC
FHEQAsDfUIOun+/NDmmU2SKhD2SkXyam5wCujhkdWkLaHx2+kW9XMF5JvWQtrLrv
9YWBUL/qNxYNC3uMtpQcdyfxFK+KQqbQ+rU2ucGwT2QGhCBxMERT3noijy8lJ5RN
tbUUdRDFWMRFUz8MA8OArXlDyDTPkP46WGfynpR3fdIS0ed0hrq8Vrr148apiAmf
5stHHqubOMZJqXnE1PBTn2rR0O0fX9Nely6Gg6iU0LtVIOegJPvehm9pAed6O9iS
vnMx5MLygYXzK1xy1RYGsqCGYeFthlW0DbSPXk/RmfOrI3f/ZbpwGHUB8NhP7Ntb
2BNLo2/Rw1EbUeH95o7T5IMJ+AzPAQZD2q1hpWQwyUcAyRHFlqLwvLu7vSNWWbGL
kh5oIhJuckLDY9PCRCKd0gENF2PzyEwItHKnbRzlUCcQ34wQVdDbqbbH3f/nrX4j
A+YlYWThpi/kCVk1ULEenwiAAE+aD6BajCHNlQZAljJ8ApPaQQjQ5NuLSj+KJ9KF
it7Q/CcT6Q19VPupFAZTNKksTfZX1uiVJHvtLjrY1xTZUiJ+7fcNCb0mHkL7qJuF
DPd2yLX0z2DesYc18vL+So1NbVV1KR/KMr95dL2e4rre82GON79aubVobMWFIPKD
w7yq9lc7IZNfcCRTq2/QkbqU7sEo+zqPOfBxcJe3h8hP0IWibOmKTBLj0HUjblxU
Jsi3hEAIprtBgXlYvJTkxILC2+zAaXRm8vyidcUod8Lovby4/9XpL7i596GNZb/C
/xO4teSUJP0WNIRokdOsWbCWehj8pXD9mzJ8Yy3876P/81l7P3DeB6fN7isYWPcn
74vSer9NLh0SxiMtfNrZhnlZICRH3K+Z1QuULOe3h+ERnwqA79ZzAv853LM8Ps1V
HVYiqJWvMBZRS7NkqHvQnlBynG9+lWA1ql/ER4VObn/ML3L/Bpf4KfVsnvM2U653
MLdrXKVS6nihjrTu0LqlPp3b2uGSFzp2oa6LYcNXbNkRZk32r9O4/RkZV6Tka3UY
zEYZSySYiJGyve0UsD1GydP1dK3fJ/kGUPmlfES4dKJolq23QUtPl1OZpCyxpxR9
u8q+d1gZJWOnu4yMLk+/T8eO84XMj5PJG+yp/z1zrN/ne8BlPI43LVzd+KhqTKDV
Paiw2vd44G2BVLUtVwwSuGvU/8hgn1U+lFd9jRMV7SVt126RW7B2LIN3zfwsCk/z
1Pi/7mkEQzsxVwzDHyWuwN5IIg5lN81Jn5o1vxNk9O4QK1fthSiA28edYPfRUpyl
wW+8cWEG7lEQrZlfDZftLsZqigEDEWMVNJWsIku6WyMVCgnizeFogE2NWsBC3nnG
sNF7C6/S9oMMBe7X8S4mwA7xFCVlD7g4wFHdhSbe/Gq9PAcEWbucN+o6E31TDQ5S
Iy4kE4fazIs3gvs3LuUPeSf/TQPDmQ2gi6lbmUx7DkY9PruN2wX3Cc/d/5n+nF6+
zmKO3oA0AMEizPsKLDvakm/ZW623HuhMCoAR4jdelEh6dLigi7DWsdqhtUhP3zt9
vTpZn+tZvZ6pJclI7ZL2C/TDcyq4cJBE/FGizPQey6ZBKXrWN45xZ/JYQZ3yNWEc
rVm7IrrXkGpzFmYbt7n6WVVk5/pdRitMkP1sBhN5neycDGaPBIXWUzFyfciCFAhi
ILK+hty+fdfYqCfyi+DBNVKlXAMLCosgY2B+0eXSaMLG9T7fuFdgKJJ3Z4Y5lTJO
jJ+jUz/rywRe2CeLBpM6LPRCVXuqWAb+Erh+tvk7QOMmAYtJVTYTUSwM3MVtA3JB
qDs/gR+p7MvHaWCO7vJv0qOCFsGa9eLotgi1dOsNme3ZvbITdWrD/LVMJ6GzDVuD
qf5c2vxP+qvfovVypZ1KO2zmeGcFLUsr4huYApapFs1Jt5YalZNjBTY3MlmiT0jQ
IcvmeII8viNIQswcMU1wYQ1JxFM504aqwrhOyquhkB0JCjYcu+C/83shU3CTfspI
heUg7nf8En3cgE83s7NrnluB3MM79q1rzCkq5sQYdPzIs/O15MtF1vQkl+CjzgVO
oLiW51xb/jpDrAWT5GpqOr3AnwUJ1AwnLGPCY/xOGLn/U9f8mDteQY7jXz91GTz3
xi+1qYb1+GzWSgkmOzb1arefFbOM6K9hsDqMMQlqoo7BFH2B9tkR6FkBPy+5Bxjz
/aILSAs4nduKUoPu4+mNKc/t5Pc+r3YuxdFKTDISIWIHBmq/FsyLUfMZ/6Y57ytX
NOePuhLjHW/6ynjiqu1tbyzuSoy6B1QNwYA6O3e2fl1DjCb83I7n73sorX8rhpu+
7ZCmOJwd4CBtC9NOY22Thh27gPJlKC4IayyYRHWf0yKymAbbR2bl17IuBQ3dzlLR
pGEmsgsGC+x0xuqgYuAK4SvJrZPJg0UQZByqY1d4/IT2BPebb2Urcccoq5W9PISy
GPHICAISVgZbKPWi++sb4pMQSFJKpsNGtxVvAtJykdLupmtoxm9ULhjhZOIJUYxs
vBenTyzPKrU7bQsV4fqdkfv23TorB75pujKZAWknnZNgQ6LhtHKmmbeIfG70Zqwl
MLqtv7VNK10PPTyhKUe180XjoJhDfmM6p/u/WvOeZ9+ZU2lPRjlSou4Nv1tA+tcV
YEUxC5qHtU1etdRFd8XPJ8PiOsqD0Q0oJ98FvfU1CFqXm/JmUIFKc0KqSGgnxEMN
KEUXLtrlXmdo+zdEePABGUqyNgwhuKeS/9MmpghHpU/okyDGXG1T3iNZzTGgUNIw
zCgGAUhnRJpZ1TpJ78In5gIja5/C4QErz/pLyV+B5xF5O2613vdmnik0UqtOdSi1
7sGddVPOf4w83HU9XaOP3FOnww3pzw2eTtcTiIfEbeIGHM52dl3OHjihze6g5GGR
BQwUBkTRo9SN9trQTWykc3o7TtYDkWptK+t2xNNQgLfT4Hs+IRodWmj6QAOghMSE
uRxLIr9SUNLa1DNqIW3dEdd6QkFQycy+CvgCGQ8CzLsXm9bsmDfYiEOf3D8+QlPY
uazTiQ37qnhUL/bESwFVsBr4i5fayKh/n1Ci7iR89iL9CUu8Xn1ZjbqOIRvIyq92
abvnfHnp9i4J1hEv36JeN7AjMZ5rNmNrV5VUrWZVYF8VA9M7BGhzad/Uw2CDd51M
xnOXatHhdJZJPq5/86RYH9DD2ut+DbjV/84nvfUxQExthw2vosbCHS3Be4c5430l
buqEdrBC/ja0jfuvwVNDSEoYMBSzhIr7051iZ0XYa4t0y3xp2H0dThFORGb89VQp
rdYjo2Ybzyi0/n5UZgQUimkpiYOpqM5umPvHGwTlP2x4MIOjyMtlesw3q2ehD5Tx
Ea9ziU6JUsF+1XYSi420zAYIwWRIbwnz0AZGAEM/kLHWfmU2tvUNunwW3Iq3jzkC
zp5MfNA/Ps9ctP/q6Rb2O/ND/5OC319cnqvOJ6UVgdxTE61J5IIofVricJcwBrd4
9qT0cDly+SQdkIV47IP1EK069bmkjHq5bzRTpEk/Tx3n4RnkDp4DoQxeGdf6fUma
ovKHifXKQ1XonJ4uYk8JNF/G+agNvYE7E+hYhuglkyeuHTirCXd9RwfTmCPxME6m
oLTuUv1R9GP+d5KWMKly2sBVsQKTVuZ73LLqzdg1N1+G7XiOCxWUApgcGGPJJ4+m
x5R10LBCHmMwchI8kzZMHrLSD+uNqcKdcGdjhtPr4ThRJ6yYM/J2jr6rS4+eUPMo
K5gZlVijPUjUvyi+zV3BFoDwOqwwDRzn0Zr38LXqj+XQbzY+JrUs46JOTq2ns8Lm
vowmsZ8KjWdEekN3DR25kybH3cizSf3Kkp8ZZLZZNDutr8h1o11i3fZhZ6FEyBTE
ffs+H9LknWj93o/DDHWEKhoX8Uuv+ZyWHRa6vxsrT5DjVMojM76pFosrWnRMrEyt
+20TrJk/+G+EvamGlgyFWx2yh76jzFq7exKxKbQFbbZE32BTcQQSMcJ8AYkXD9Hb
bik5F9gOK3OkPlumhVl7hy2JDOomTOWPKIQzq0ODUJ0k0jWnweQxvq20LPn64s/f
elEXhM6ktsehFKECN9uyMWQKDHdwzy4yzALM3KUXL3dYx4vgGWeAafyUqaWnhP8z
hrp/P0JPW0ATeNWlMmFKoaLUkAA1RzyYqKo/A6MYYY1pOjON36hwxwe5ayIZoRR3
9Oni15Ljz/O9aSpkbvC3EUYFqg2r4nCRzrW3kbcBmlVNKA/ulp3IWPoJisGZHCNQ
XnXOar+BTcZlRptgdmnTuINNrMoZfbmInLJKOkAqIM8Vh7rtrnKskJi8I3CzcOmi
jIqt+6rjR/+BO/d8vtojqeD+JnubmFKxcIGURUaT4l8TXCbVXU7jEy7qkeqP11GU
rkAsMA6DbUSkngoIErYITIPzMT6JsK7ubNwcUxQCAo0qs7hyqsDurm6CoJoYf8k9
joZNOIYlHlbxqye8i7xe+aj4zBf+bx7DRYVRZJADn3O/uOaE76a6rCjXGyIe3VsK
+stxcEeIgQt69V6U/jko9XGnVuLaNNgQ7nd2LHACekoqQCJWSvgMDqQKJMbYW+hM
9UuZX9QhIpYq4WYJsKgve+BpZm3opxa3ZGxUHNirolLZDeFb2YNwV2uzQ95VMpKl
zhLwHkCONQyj8EHK4+retAZLngnWeKuCRoUjAwASUoqyHYouLBMKHlB/VE7iLgv1
LDXGlslXFVet1n/NzQDVclo7nVuWs2ua7PmDaL9A+erdmjcgvrefzrSGWGkQ3d0P
sdmjXN+3AY04dAC/LByCr1wgb3Dwy/yZo0XxuWygslW4esg7DbjDkRU95gJTQzLs
2M2fGosvrVxdFcp9Dgju28+qdIUEcC6y/7ZNHBsjJOhwfkbpizzbY19nYHe/tZD7
Wu8/vvXQy/YJ+LGsNP/OrIbqJcIqpGo9wxHDmvAnMBW0Xr1Kr9tzYGdSCTvLs9jb
eFc8ruFbiSIWuPqVuNVUsAyXP6sBnrNXxd0lRREKxYmR+WuRKh2OygAu9qyIXX+5
ThQA1BnslKKImZ2Ld8urHG0FlH/xRLofvCAE6QW9MY15fNtYhBlFK7ZhxcebToAX
ZtdaI4hNj9oR+WKwHBLNKETWPPOEqKMXS3IOhrGsMqDmoZBQ5CnE92c/5+nM5FYE
ct9U1+szHAChKP6oj6NvZwQfMmrM5FCfXubcXMLzXVEdrrbMx4Qm4mdQb53lYs2U
nghRWPRIPWC2HKmcnHsr6Q==
`protect end_protected