`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
ddtXksX2+yylW5zu6QL2Lhnb2d1sD00763mmSITNX595NcHTEkwn0zB1Dry37fOW
FufOhVzEJp80NC5qZ/+F0Vk7Ik02dIR0elf3clrjeJRK85K4e3Hoo4xn7YbFUIms
l/8VZSb14+JVGURjfswrIyCUotIzlzVYZ6gzoZwDXIi5gQIBf/gI+KxNXPaKV+PQ
Ufys/12rjO6aI/pPlqSm0hCvftmBcnezN2hk1UeXgOIuKZnogjOsf0iJVX2aOOWE
6pD/psybjbnsNB6kH5uFTA5frkzIzkzl5d9+YDm9OyC+k84E83I/7/j+rk4L2dah
QJOvksSIzN867/4Qt8qYTQ==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="MvBXkzurAa5VTw+1JJ70nePUfoQXBvZOku/SMmg4TwQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
oRtzZL4VJ4iwysPsC8SXYCzXS8Fw2gtZTOskLcDV+1B9Nzn1zTyNtlo6lNICRmmK
ZRVu2BmCc2G+fmzynYlNTnSa7C0Cuel6FYpxCBlOuk3OF2tzAmLAuDyOH3Z1Yjzk
a0aHuoCdIRKv7BrZCdALt03JeUmXKPdOmIlkVGFl8yw=
`protect rights_digest_method = "sha256"
`protect end_toolblock="Jn9CQpRhJt4rnzZPRk+dOpzAubz7omckX1MrFd4p81o="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 4832 )
`protect data_block
gD6l00tciPUa6pDNTk/+t0OO0nC/UTtBwLB41d4inuAUA3i/ALrNyoJVcBnAmEQW
ptbcNp5fxEUJjnOxnedyZEuEBxWRieZFQnkRdF269oP0ohOcUT6cHeC5AGJhWCuj
AnvOZGcuLYBJ0avxVVThOmKNZ7gZR274AaWqPFlhxvsl33sMd8b6DGgFUKgh/jJl
uaTOy2p56DNlIxaXfAp2GDnyM5dZE/CFiwW08O0i962JT7fDPXOJEoHFHin4iFbF
WLVtS3mwKpvsjO6bk3MYSHOEw/tvfPdz5tN/ppqh1rMAxm6WF7oJIl+oKR/G697q
uXkL38QoBp/XhQ0IkK4xePV7iuwyYI+txOqg22sTQavu1JbYIWcsqzRbUjdHQdnr
AOMEsY9z9yAFi/M4e+AUog3o6VQFcDoYoNcnJu6Ef0sNv1+cDXIX6tILckYTm80K
GNyaJ4vfWq43qPe324wiQOEsSDWqE7nDorNPBem/35DQqBiw9+qD/tHEoFy+0ic0
bzU4gtsEvEEwWo4nBc2/k4YYh78JVyvjthuBRQY0Szrcu0ig+RoZS3seSSi1Cnnx
zM1jR0S6f22XfgxXKxg7tFIv4gcU5QYXuWismlmGAV9dGkpGnp7hEPxtQc5O2zo6
VdNfFNzeZxDA8sKkPfSIaem3nkGxf3wvUR1yDjiYl7+KZ/tV6/Q6C0bnAM/0OGSK
cr7qSTXDPm2rSbFAycEOOsluJRyMgn/zU50aMqpzhK0EuMdK55XQeNl/ekpNXfwE
fBmUYi7l1SoJRLIlYY9kWUcXl6t2iZHbGga+vFk6Q+SJxHOzVa//lXDmg9+MfkRj
BVlPa1sH36tfNRzNnzjhHoEhk33cU0/ZflrVGJBGTeRedjE/DbauIyadXdymSUrN
QVkXNoOKnR1y7Vb5F1YBzgllm4ImXnTb2L1q7gj2/jueXp5WoxDygAfeVfq18cC4
VVcvlWPl8RGOzPbQXpjmVTsL2BUjcHArtjoW+D7QwvL8vh1RbyG6OkjzEKIZvXRg
EdwtXPmevpb+Rq24yrl9ISbP88KpVJkiRQQnqqRyHkR+ms3JEQP38Jy8FcqitUw1
9Yutyod5jDVm5Y/uHx/WrGftFNiP5poeeJoFNmXlUMtn8OmsyhWShqTeyZrlTTlT
uI4cCkSbazMo4NtvA0v2KXpBnRu1b1ecxFYQP3eedwmk/fVWYn9xQZ2Vd+VIDRGA
o87orRIWGZTQHaI4lFKsSIOpaRsY0cD2P9/tv4LhvdmO/Vr4dz6PNLswGGtzVJzG
StVFSadf0dmo0ai+rwRHu2AJn8tOVg1iB+4kMnrfGVMVyRLnm7ArBgcydavJfB9p
VlmIgsZEqWszd9QU3UAQxSlk35oEoDEGPIyF5Cn1Sig4QkDdenn7vfaNJw+cRh56
jauFAb6chexGIrSsV9H93EviNyE7JA0+PFSZi8KLn23xzGnun6hsjW6YphepiqDn
sJ0gcqUW+7MFZWYEtz5nAoTV9ftkKxTyBHNacaSicrmeWZBn2/Cdt6RGZjfYPlog
CM+57OdoQItTjcibkaieu0F61hb/9kL2knKT/E/ukvIFnCq+oECkrXBXJPN2Z33I
jKoBeE2W5hbsvbFgb3eTfWjjj2JDvm+FHUYogfKkt51WEnUCFMulfd7XLZBqgTN1
OVtdoqwBfdGhWedpIVL0Kr14b8XRJ16gYhbZtjOy6vzELKhmMNaVe1EipXFt/AkY
+p75ZOgeFixW+7CReAYBkrKmPNvjF6z6VGF46eMP0TVxvoVDTO2lo41ceC+7CYPs
okFPaGMcnfeF/VonjU5DT7RAdptriGrrnGujc65oBDpfjuE5BuYXlqNct+85Q+5i
FQ2Fcj+DPieYNTXrlsxVXb2ygkCjFgJmws90zkQkYjhKiQc7PB2mQSUITX+vcCu1
WSaeVbwBh+3QPr3uhi30eHCCFMKgtxtdegaMe7+BVn+Jxkb56thpY5yhJaxvlQwf
TmDPXXDtY+kmD/mcPW6bticgo4HqIu1jiY3ZGU3tarahm3XIr0QMXrUhiyqwX0p8
fptk2K4qy0BGxvCQCZq8xkBvU35K9CIyKYUw027sgkoHJ8uX5/WxnDmctc0+Phfp
AAOcH8coj1yyl2ZrN6Cji2ABuTx8iQwrjvw5245cBb/X3QVxkY1GNopVpWnXuqC2
DqDOpwcRZ1lRbmZIS2PpDpOcXRdKR+sWGEiAhK6fTpieYnPJ7ag/EdAxdhH4En3a
T1wjliLnEyH1+61nzYm/1WrLNc0dAgCLDcJ7XGP5obSS6N86mO8mKcU5aDi/DJNN
0NN1+55O5+m211H0wNua4ljUVgkEMhEHjvMpynNtexBL+ShjbQ4wDTN3KgWpKPxx
XwOHmIS/MRgtouHnWq/XcHa/5B73fXETVZtC8AwN1FiwvjZsKZaesFcLBuIYIEYR
ASMcr8u/7/fuUXkAQ0qEh7u3vX/nj06/s+E0K5FHMs5HwIMXgF0ocLyW6h9B9beT
xORQsmbLhQdsdJ8YWuAzpoJnqeTEsSd/q7y8qdOpaeGf4zKFmfB2MWliFC7eiiYV
H4YnsN85USIOuX39W1vfy8O0UVqBe7wuvkMnCdlLTqBsmnu/zr2c+41dmsD1Zl1X
3Aw0x88BiZpqCSu9qB08ikUv0daGsLsHiZ/uOMCcOk8ivDlE/DnFcnlgAwpBneq6
xyiCrU3pyRwp1FvwjJ8Iv0cp2G09Zp4NCIbesTJ986gazltoTlrgoTIVa+YDCsk2
rf6Odno8Hu/XcyM+DpgUio1wx14Y1270ZfP7BL6jszNiQxITMW9iDxH2rvv5NYBx
UMxGr8wV5S3JKdp/cDEySJ/Q8PIMT3L+44SBFsAnt2o2HYR3Z204+uOxW+vHk84e
Cz5i/UJS6kuinHKYxOs4Rnd0rOmm6MqRu+IdfJSYE1Tn+gF+jwqcpsZEuFUQHz2b
EErxbHCADihJHUhip+T0ktq+qR+qWkXeZg1iEl5AIKmjKUWzmCuqjM3HlaT6llVS
tGQ8MPbikekjQK/GI6vyByp2Qmv3GwuPYOH5GgL8ZVf8afo6ZYMqgbgjHDRZ7jAw
C6+biFTXkQA69Rc7HFEBHeXlmnZcPvs9OnWYZDOAQ3vcLhacYGWaYJvYz6FPemGN
BEvHAOKZ4fFZbDlpehFju6RFO1rF149QVUMYsViexlrWF8CBmgawR80jU3uWuU9N
aLhxr7kTTJq/RVbaEGsF0zC6Be5cUf+PBgYApP+aV/xDDeEBPuYIWujMMjCBOqI+
rZq4FIgTmtM+9mQ9r61vfvJ2ogUUPnf0KGNFknH00Jw5AyMb5R3QjQxv04k4StQD
ItFlEwrXbnX+9EyXIgFDG8Dv+4VmkCoSP/0Ap+eNtbVFUn/fsJc0LdLoVmK3dO/b
mIe8+8CNK21nUGBFofXviW7wptctodLaAgUsa/xIhbHSHGnLCZMFkTGE1C38zmC5
pLPHRIVsLJ1AZNuMK1ga9zqkO2n9LnIfHEbDVGyVPKxT6Sn0IRu97c7UKrcjNk58
v1FS8PbSYAstbwrwATp1pB4X0uwCza76x+HyMgeXKsSjnzifZ6ao91b2pp5kuWFE
SJC04I2V7Smcw8uyvzKejPZD0IITBTE24mn1Y7imO7qoAFMzg/Zz9347IQkFzl1w
1KA2YaxuGb7xs8VRAwJ8H9rKVgiUSc8DF02076GxJ/VusV4gYVQwkosfmLqyny8i
Wkqk+JhO88mw9zY7DMrZoZ+YDmsdbG0Ds7z6Mp28FnahyipIpduJM2k4M1VdjjDk
FB3FnAflc613Kv/kBfsCO1TaUH7DzrrtOJR8a/JZbxtXe2cw3KnAY216BwWJ8Ydt
0pNCkQxPiDOM35tdpqOpbA2Mpyrcxr3ca3N7ANo0i1BJoWDTlwN5dncQmno5Yc4T
nCueRmj0A63+kzcgIpbaxaHnpquqAgU+zW4bgrCHBE1cndNUR38EDYbZ7YZeBNwg
l0aQ/A/YV+pceEvMEicecku83KM0/YCksTaYZ7PyDVesKHE+/cLkyH4zcquoeCcC
auRP2nK+yhL85OzC5LXZmghR7ONZYtiVbmTY4uMgvsPJ07JYq446+SEETGeCefyA
uD68f1apakFaGu3/MTjkOjOYcojN/G3oVLYUgGgCWSEERAVI7SJLhFLitJFiYoPu
RYEplu/i9HuuOqmSFmHnYLdxLJLOVOPEDKdssh827ckSzM9cd4UFnNwcxEVnPk5G
cqUstWYvr5sJKHdz9ovczFge683i+6o+EXs4bDVqwvrgpA5KRCNnnhn1PBwwDUmU
GFc70N6RB+vaG9RCl2s8rj2H12/0nPCt2FxKyhPZCvVzyQTMr6DWb17gEs7cIawB
1lcV5Q1bg2AXzIVVWhpb1jLHfHJfGQXxbftwHsTfc+BX0Ewi2MiLbpO0R5ezmAcl
f3VwSwzcjhQ2fHzrdx7j/L1G+BF5NaJcVaKxZrATadWICRF8FNMxmcw8ApFxPmzj
pHrmZ7KDBBbmaR+TBscmxC6JjDHRbGr72AoA9Fkejib6CdKkq730pCYKt+FKOh4g
SRLKBu8LUiYpAI87xm5AAgb8zD2in8gt9M4dEu98RDJFLjm00wgSf8DcFk7nEw5W
QdpKQ8q8v6upF7Ox2IMAIZ0mlGAYHU3YSLaqAHNmgnN61Bz9bsk6NRFi4ePiNl5L
HWueUAsnoB/ILqiLMxKhzDlwz/INoMjqTYq8i0hFJhF2VjIVe7oOMGObzTQj/c8F
djyH7jdAVl6x48EvfhH5sBGcGSfWlF08Qc1fW3UWUOacbU1NA+OMu8uzyutB/ANi
8DhJcREJxARyYvSZ/X2NTjD5uXOj3yr/pRveZ46F3P85lk2uUjBBPBSPUHdEZmuh
ACqitKQvKNKlqat8jS+6DQOV3GGVizPLYZotLIpqLkA+HvRwxaHoCO2+wgJVcHvv
sz6QiIPiEfwjDW4kGHEN5pua5AsT+Qi65ZUAZ+a2GJBSuCMY9G51zeQuSjwpLjWv
K/5wmgxS8hcgS2ShnjZn3s3fSsiBmOwZmsVuLOKI/C/Vc9bLtpmHgR5veDlZYTT4
O3l7qEpwh1td5s+XOORBK4Du9+YKkYUd2swQLYcOuDLkvVlt5GdPGhJdnfZJl2jR
6/25srI/Qphntn/ROwzknV3cCe+JIBpZPPheBN5rTaTfCmrzeX7fgDPNgH9NaPnr
x1zqPElVfqE27g3QPo6vAw+6Y74//+xjWzxdwpgWj2wFF+5rSuibM3zBe8d/m50M
D/TvWL8wOfuSf7EeLDa5KfZGrzKMENIEL7wlwg2BFQxydu6xbOc9d3Wayqg22RHw
OBhHmYbLR/gfgsiOLZO8/lg1+sGwLB8C0zWEqY9ARS9UtLT3/Dr51SuA9x0kYEwq
YpVeR6Xdd4iszey7EGD+2dvhvClt+4lC5KD0Gx+PvXcIh8CC+W8/3KhAQNCvi4cB
01oWFHHjVz9jNJRaL5ja5mFKyUh5QqIV43O3NzHj85jRqns1JzCkHLkEUG2arDsD
R2NRZq3sy9f9ewpywXbaXjCUCT3Io7WiBk10iW9OSXJeHxeRw9AFHush7Gsjh9ij
yeO97T5baIz2QCcAwdUzIpH6S52T6JZdE5h06PjVOysnvc6BN2IKrIasBPrdGlD0
jnVZ67KwxYbX3yVBBkQM83JqnfhHFcSIw7DZD4WKEqnXYZpyXG319U3HoJaZBIUh
fotZlSsPSejiXom0VoFVWEXc9JDNKN7j/WwGoz/VuiYgS+0J6jic/URwYwPJGxOf
AOPyXVOgm6ybGL34obnFgNiJcBbr0dGIYR4qJAmQzLtMWm6N3dzrcY4TJ85qlBBC
0P2p9erJWRYN2PlyTB9wMbaDI4/NJItFnQhwRHDipnPQJ7a8ng+tCkAQkJYNR3Qn
5Xiki6y8vOiBt5d7VQNcbetQ8GtD/9CM0tc723lkEthQZn3DUkGNGYECCqAUJ1xy
GQbWLSUJznA05LjQOJDrODp1AFDQIreo3BzgtSLrzKn6KsMGz5MYkq1/7tEPj7l1
8nvss8/duIPat1UJEb19kWe8mjmPnysVgKo8s13eM+t0hC1T4daxrMIKqXUAcgtz
/oCnRN0mFZC7MmtEhLQkXvEcHuMvOUo0S+3HRsRuNR1vHUVJk0D5WO5Z8I5dDnNu
rTpZOyjuR2g9qn/t98c2fvndEoSoHaYV2tTUwxqgk9rL8seyF30AhQbZmItMTfHE
QgsVxdzXflpMcDBlz53Cgoyq0xtYr6dEEZKnHNbJzrgkWioPMDJIj8Ae9tVKvz7W
4LZQ1VoXprAvbklAOZTaDkrrCMFNsvx7VIJ7V2206hwNCO6GPcqKwhx8rsRKUUog
V9XUOuZOMzg+Y2gbPZGeHkU4y2V7r6nLN+5u88lE9STQDOyKhAVgqVk6KvjwJd8T
h95lbwlbNLtACViu+08U/k5+pI1oyqRRZjb4GCqngmw=
`protect end_protected