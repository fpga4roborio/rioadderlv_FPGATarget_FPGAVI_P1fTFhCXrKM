`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
ddtXksX2+yylW5zu6QL2Lhnb2d1sD00763mmSITNX595NcHTEkwn0zB1Dry37fOW
FufOhVzEJp80NC5qZ/+F0Vk7Ik02dIR0elf3clrjeJRK85K4e3Hoo4xn7YbFUIms
l/8VZSb14+JVGURjfswrIyCUotIzlzVYZ6gzoZwDXIi5gQIBf/gI+KxNXPaKV+PQ
Ufys/12rjO6aI/pPlqSm0hCvftmBcnezN2hk1UeXgOIuKZnogjOsf0iJVX2aOOWE
6pD/psybjbnsNB6kH5uFTA5frkzIzkzl5d9+YDm9OyC+k84E83I/7/j+rk4L2dah
QJOvksSIzN867/4Qt8qYTQ==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="MvBXkzurAa5VTw+1JJ70nePUfoQXBvZOku/SMmg4TwQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
oRtzZL4VJ4iwysPsC8SXYCzXS8Fw2gtZTOskLcDV+1B9Nzn1zTyNtlo6lNICRmmK
ZRVu2BmCc2G+fmzynYlNTnSa7C0Cuel6FYpxCBlOuk3OF2tzAmLAuDyOH3Z1Yjzk
a0aHuoCdIRKv7BrZCdALt03JeUmXKPdOmIlkVGFl8yw=
`protect rights_digest_method = "sha256"
`protect end_toolblock="Jn9CQpRhJt4rnzZPRk+dOpzAubz7omckX1MrFd4p81o="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 14640 )
`protect data_block
gD6l00tciPUa6pDNTk/+t0OO0nC/UTtBwLB41d4inuAUA3i/ALrNyoJVcBnAmEQW
ptbcNp5fxEUJjnOxnedyZEuEBxWRieZFQnkRdF269oPyXUCy0Ae4Vbdx+bu6U0EQ
BYNKrEDx8RrFwK7LuX5qQafmdzulBPHqz58/VWrqfQsLsAwK291L/SbwV0HYKpYS
kVxMZ2iDpDp6cDi/YtJ7SyFhn/S0g448w9JhtN44sPrll0C5ivtQBkSk709Rl/aK
wgQjIfV2mvL3gS6HsG/5gRTEr1e3GbQ+f0uB25HaiyNGxXLXJ5JgmyjT09DaKk3l
7kId1cjUj5+N9cxRoAZdC6kJskYtS/ZAxY4SlO10NI3kluUpZ16Uhg1zczpZsd/D
YsCHxJ2/rigO/n/0huH/XaExrCx15caOFdRnfGF/yIjI1PVrYMLVX5YjdEoAmVY8
qoeTrRpHdKvm9cL6/fRYRl2b7eaf9aEB6ubMOUg/4Sfa1+rxeAfEXFUlp9qLpXti
xfsuSlSf2xECWwL56IbVokBrwL6z+S4GOoRIoz730I+PEYX7afzINK+QW+1r2ouE
dvSz2Pkcx0ll5vZCpbscwnMk6bjzWmXDbsfJHtWwKkEEup4WHqBr3rGko8J51/IE
vS9G/+bjbzERof82nDPOcJ5BtGqvkYgySd14KoWNPgFUFOr+EFY22YJOn9NyUgUN
bHsrGDsO2NqSqcGWI+yk3LfZieAPXuUMofyO6+Qy4DeowFxYOj3N80iUZFLKr2Ci
ffRA3ADKi60gMmlxVq9h7aduls/5jOtGoEQzF9Ao//m/gu6hx4f3iBORup/SUZ5j
vmvo101p1lJgvmjdMoJHGOxeaF/BRjk6bA7IQFsW59J8gsZTBZjrCb1ZGwX02zKU
EExgWIGW6dlp7fRl5sGHxjM+RYZbfLfMzdc8X3pqwPuKewymRo6CAgduK52qh8qM
iiAh/7S3s+Y3mYpX2RdP5upgv3uSwaD+mOHM3rdmDjX7mGy9LZtvWByXAnkufXIT
iEDTU+M/JKr3vCA8CVQnL1mmFvWSKAcLP/sa7NvMX1VU1J6tg4g/8MDY6M9PrR83
fnbqasXsc1bWuBFcLuInrT8ZL4W0bmqjuTQNnNL6VW7lp/xNkvaEIo8GX1bHU5gN
SMrMF2AzTaXD2HoatROB/IaV4z4pmU1WK5NpHwyWjEPn4yzvww7HqxtLiCPrFlyT
OROyORpj2VlxMCjmvQBX3yuCgH3OkY+SS+Or9r71DulR55Wb2Heg6JqWuTQxYFeK
eZ/5PyZ9TTtPHvs/nIAoCypnTYA3p1/8uIPKMWsyDNFrmQ58sUD8eMIKrPvQmtCp
TfrXn6Agi2mNyBbRM6cnhmmXoN+KWya4Fx178mYmFqMin2LglPBPpHSomI1PcmVp
D9Lsrg68wCGd5bFyvdkpXqYU7Utq09620rNs2LKleQCX2ZxcbdZGcUl9/cRw93Yz
lS0vluinx1UmcFUKC+gMEn1EfteRirOrlxXOnMEJMQU0FRgjHbhvOQZj+1lMe03O
ko950lkdllLsPmZyaGJZ/pIk7FvxwsKGb8AsyAdmuv6HHqFL1/hUtS16cAwve8Fy
3r6VKp/CtgyAPScNOebUpFpK4Sh3Rt1/MnjTdnk9t1zuvP7E3Q4tLMMnWXYg0kH2
EbTd9BsbdB8noKTkS/oOUz0JQh+zVO7hZkoZymgOU/+opPtyit+VPEQm3f+Oz2nm
ZlLZzYP+R7nSqBimrKPoqU+/y51clnOnBQp2OoU6FT+oPEp7XfsaIDCKk5BFrydt
H63SFOK74fMBVHMM/1LB2pQY8VndK3uO0qxPzrwdCEyY9pjsJacd7CLPC8uhSHm2
6cvdKdL41szOqa+axTZe/nvxpX3OQfCxNg7imxLkm77CMQevIyFFQFM2B3qyzuFI
QnLYxX5L1gnN6BLXGFADTA7tWVCMK0HQEHqo6P4t94CP5Tuy7i5ebR7UEUklgc46
tCQfrA6Gm8D38vDf51FyIKKI3UpabXx7UZ0QzKYMEAYWT5OO+BA7V27Y0MBon/mg
bQhAHim2QmEGSXJ95SM8R6N2eBgArgAptZt3/BmCL882hySIjO2XgEDywnPZOJBz
jFS2jGlPy05NVG1ci2SfMOhHQ+2qKwMqSot6pNqry5rEQm9sc1oE8N83Jgg12WjN
DJe2bQKjCGBpmHYKl2Viz4O8+cusMNu/mdcumlURKT8cR86I4bgUyT0m5JVm3g3u
6oZNZ3T5svCJaOHyJWKMIJWM3kIETr9RDK50vGgOQGURiHRSoxHI5f7r9lv18ADO
6X0WY/p52XuiUzhdzLbm40NBdPiZjye9kvq8E7X1XjlMi23TdstVIp8ubJigOtMa
tja1nOOioEW+f1R/rxesPA08se7C6tLUkoe0Wbo+qZYPp2PpkWrYQ+/V06XX3EQq
EwCM2aUz6bswtOjAjwxxmkq78h7dzol9yZ+rMDv6mUp3Ok6TmT4yETZXktZ5gsHd
fY+4tgZVADd2IudL8pcfm1/3BriUBD+MpkQhlrc3n9s20uoZc7NEed8BHRO6qbS+
UQP35azIsiBcEjCsb8vgZnKjhZeYuV/pRVbJ7PEB/zKp5yPmmWHMo+KyoEf5KsOg
/YGymFpuVspRrCei26C2yEz8aD8+tC0mSyPP0QvkOTEJl3ttUR+IeASzF5mJVenk
B5ym/SuJu4mRNzeCzMtcorCRx2otJMenqaHR6Qehby02pEzG66eizRiVF6dDKdIP
+rVr4D9AYrANNGYXF0+cWzlZrwuBRPlteLCstAUjYyv4bWI37tGlEzZRHTttScEc
aCzLFwCDvJAqgig4fvdXe6nrC+UUNhGFR9w1uerJoMETOXsfdNeKShsM6BIfEiKD
2/LE9fJXGu9/q4jLjGNsIs2T2mb8NfZT97Okx/BpW1ItWDUKSOVNy5dHjdhcny2B
OhhVC/Z8ZhvpcYUF1bonGYBr0uUjzrdm51PtPwP2QpH5CWaf1t1XIOYC+lJ8EWq5
M9pDYUisvZwvYKxudezJMgl0FqUheLJYbUvlJggICyATSIn/pXcRoU7TsOVThEiq
ONArd81BO6E/LeYzBnPAk6CHanC0cSb1xDEy49ozq+cU2ftGotZBpjxFU0Ykeamx
UIBH7n11JsG65eU/gWwAvCcBq9+1xBJHpYgLaDtAHI7hqcyGH0Er3svajt4UpvoN
B9ioX0A+zy3x9AXbF5C+0hhYFLIZHhEkZiZYe3srvSWVEU/iORSzMuRhREm0m8Q3
8FJPJvOSXCU72PzpEwfaVYxXDwSfOx+2ssJFgAOJGmtZIuPKX7HLO3HCxh+OOOzt
HgNu+Ir8d52zc0yUfgATQ8U4iXkUohhFWNeHwQdSpPxT6ymSBtc9ofikLV4WaNL4
IahcqMuqYoZRgEXy3pFTwdMLPEgSIXOA06se5Id+NAAXxTqqNR1ZO3bUULXFoty/
F1xxhuAM3zeFB77m2TrsWgoSamVAgBL/CkYwdHiCTdethWvgYSo1UseOHbTZCLYg
TNIgN/TnAgunR1NDCglKNJeSvwvJ2mrDQ8TbRkdw/NMW7vqhipEWL4QmNC5t0lmU
Wb3fUTUZUZN9O2hpl9+Uaq2bUDosxZ3epN9+ynFWBox9zqq0W0k99sm+h+sj7RA5
0vfSV10+l80pwrRLWIl76lGnkC7tpJKGMShSdfkWO0JZUzsKhuPvwPy0xBdi8cuP
33UbJW+8V1lU51e4i1LBPN//3slPL6e2I5nA80WFhUczoSZoak6iXn41VWIDByPt
Nyj/nVbBaVOAMyIwOgLrvPkm6he5WyjzEq2KnBfMpS9a9TthIa37rouuUsiulCfZ
9sec/+UKSKRsV8IJzj9MPBboApzfLq28PNB5cs12W52SfazxKJ7yolG993BpvRdm
/sRoCXpgdDIyyy3f0hULVhGKz0yR7Irx940/sH7TlT6cCOxsAx0ubUZoNeQ6Me9v
266mhucwWBhyxhpKxBfb70cz9OjI/aZPLZtYJtO+p5FwTjdUdEfFMSmo0uiV91Kd
Jqx3Oqa5mJZRs34SpXNaMb3nD5U7Y4gt7OFg0Yvd938+HWhj5dWgf4mm+fsx+4fD
9//lnzDzIqTGMPuvw/1uWY6acR5ctelMjF+JdULiZDeBEY93CraFj35EFt57Tdks
quLEamPMGKukkR0Oq5W9SsdmfL/Ng6rTmBiIUHCmt6NTO9XufV2Pi/zKdSk6cCQ1
C7rGM1tgGas2C5vcqeBQABQKKUG3gcrebZ3JrBTJaVrFH9pubE55nAOj9rxikSBC
quSWnSmuViXP4ktk2c1ZwIYwfbV/2j+uVYl/tpJQ5sIHByQeB9xhh4hg9RT+HWwl
V0170BMGRl6fcNBCAtWGaasAS07uniLUez2RQ6O40dEijYU4Ud6d7mh7JPqse/kn
h5s5bsAWskEccFacN4JV0xRk6ah6NezJCllt5mr6h1EWf9HoWY2sjFRxViT4HSxr
TwgAmLrkRrl5IAt+PV+5II+/n9xNdOjrPrzSnlK+OtXFIpsqDxtyWhTuk+bA4Dox
bNpcC2m1qPdCf9dXr8MEMAfVbYs1EeE/gtvmqY+sRsEOjC7aynUxuXtX1XfxV8JW
cCGpruVIYMWs3cavr9gazU8OaaKtIhNROy+wQqVujhXYOZ3Al3q0LuZGfWKJ/8W8
kUivuY6etem9NFRj8ZH+zTnpxJqIXt/fA8Y7B+6olMwmWcWJQloAHfSO4ylGt3Go
/DNwDCkr8CDi1GjJNS9wP327LKM7rdSPYcYIDcBGZ2l3BtexUf5GXpPqTMHA2kge
1urumusc0REBh9oBZA1lhAqN2suM3Q+hVxT2/lOtyiZVB8ltD6kDllJg+w3AJwbA
L4IWgT8KV/Uyj7e8M1n9vo6HDaElWAnnf47BETHNrjO0Xb6AIuXwyWPYhmD6phDa
30dmAWFeCHVluvj6IwNGIftHh/Fb1wtX8VMyY2y2RUwwLv2QzlQqqHOu87fCuX3p
tFWKhFiV4n3zQxjpjBye4VKrWxg/mRiMNc8HfOEHQQPbsEMFLA0gTNKSMrVVNKJl
HfFyojng1dSsdZCiSe165ckQ3WUdxBeVDdulsh+Xdp7vF3G/dPLGIZ3Bddl0Fcxj
p1yrsXuzfZRoP0Y2XEjxWTDGbV7ukpmtCubonUr7pCbTtkeEy+3FgK1On5AuPxxX
Ro7iAPbyEhNhZ5d6VdtQzjSzydQEOiOHzW9iQadUQmAMaiF0i57d4mnzHuAVWGmS
vcQ09aLZLX+WZBaVIBrMQCAM6zlQgFvKCVKPx/tqekSZvcnlK3Kfs4lqVC5V9b/V
RJ41OtqbzUiYTOlmyDY7KD7XDLbPpBfGU0OCTMS8IS5vSsWYPmbkMU/q/Y8SirqL
HIae8NaV//hKFucMJ43/JE6cj1naS8W9B0/F7dKTfXbCVRKqaYMuElzfYpP8wAh2
ypk1QR7mkT9kE+8YHSN5u2lCd8Ybkgrg6XUlNxkSyesm3vAYXS15KHGY5WuSVdI0
9PjDsGjc46wWXxqPD2J7Tnugj2Ex0x+6BcRK0UbIYy5rjuMPOIlAfcOOe1wO5Uii
nuqSrWahP96812uZsNEjUv+KgVIEXv+f3PAzE9aCxaIREkz43rLIT1PPzRrnGGBF
zdeYGo2ONznUPhPMEn6wKPr2Hi1sPI0p7yUGBrKx6URTIzpJMZhJnqj2F32WL1J1
9abkrXH/vsjgDpEyh7ivA8+RmLFjRYSQiGfihHEHjlIsqlblxUl+TCybydQXyrO7
biYLg2rqaoPY0KSE/jbar9aAtVc3Pu/HqKCM00wmc/OoeuXfXjcagz8SnYLlUlkX
5Shk/ytFur8rULv8GgbaTmBUwCA6oeNegXvIAG5yjXd6/yI8/vyFfGxCqAIOZxri
/QwbNQH1ZBXd/MWkNGdFSvFL3Kn2KM7nvIQF3A9wm3Z7ooeZTycFWFqVXpGkikbC
9uRtDYs6V2drfO364XdATWA1p9YaK89Lulvbf5vGPdt7DpEScaexmDoeoiVn4tvU
uSWBbYtFc2DIRv1R0HqQ77oUGRFEC0C4yTfRHycZyyzZ1xvB02+GXy+m3pdLuqaf
8K5eOm9gNGbc/TKPHmOAif/qKIH7veavCP4wqhDRbT9QHIV+tp5JuqK105zzh6La
rtE/v3YXCQoCUQ97RipUwqvFytDkgFR+3WT0ylShYBNzYytxY1+FBbZhFx6+bvZV
DYyBIMd/OWEZ5+XfmWHfRtd91B+49+aZdGkrB2iq1FmqVIW1k0VpaFyu6HW/e51j
T54CRvvRnC2FJ49mwIC8QA68Lt97bjxSApCjD9L/afA2E4wpyKaDxKai0cbBBnTT
gkgO+iolU5gZfjM1YLE0jhWv17RVmSlZ8PgpClqumkKJtIWylbkSU3wwLkVmwRS/
CnAl6JCNMs/csjI1OuAooQ7xmCObYI4TCfXz+97vn8uZoeCKJV2LO0hAnEMLmeOt
njTreKR7ZEjHX9BkFy3bEe+ZqyxjjSgS6MVwnZq4GT2xrr3ivoZ2SEf/wOMONyIG
Hk0Kavhw1cVnkBfh6ML/7HKx0EugiNjdUAOHudXD1rhfFAiadFbcuL1ml5SxsjfD
wznukkPElmUsgIXRAlgdBsCvxmevm6bJBLIheok+SOL8uLP6KO/dXtwjTKf3or7w
qyvusTRDg7Vpm8Q2ELfPm/lr/Dqwc4M4IQYq7udrm9FaO0C/R8z9Q2Lxp6L5PzFP
6U/4Z5pv8tcn07yd6pDLkclxfNUzdgMN+xpcLZLhXCjxv8pI7PjsV/Kg8QXz27lV
BqF6L+YUt9KuTwTuM+R6M79E59gIqVOfyJR+WYA89zVy+UKr6lTg8U96tZ7vOFWi
s2/pSrb2y0MG2TCk9AbL1es8/UIkIL7GP9sOY6REP9XiXQU9v3BJ3iemG9fKPRpX
0Zg0LB85GT5C7Pa9Lv1eJvfA4YnmJkf5M7zRc9JpXCtEp3CekstCqIzxbnv5tfg8
YU7nVPgWYlGRwEUWAePuFEgeZENhLK0F/euBCOfEUm+/hZvnqqyIYlR4U/Oldi6s
nkCyroz5y5li29tp5sLGijOSwYc4wB5Auju6q+Lv3UtzR5X8VyPt/CZOOU95zfKl
5I6QaDVbPj4hNcfHbnWFleBlB60OTUMZZ8WGYtS8+TzwaUN9LGI1BnmaBcc2b9H/
ergvxScnHCL628tZu7AVfEFgrojrxAYp9INrc2ennJoquusb8PNO0P9Cx8OUXNDI
qQkzzaZoUC52VZSHF0UChG7osWp4rA4cGALSBiQznDkqTjCUaW+QiVl+aprJ6i38
ca2Cp/Ema6lO1ea6oyTurs5fNd2udPs4EIb5AVg1soy/e97Pfc2Ret6bc0y/wYIp
8JJnAaHa5vIFNEqeHsQEkmfhKp9SuC5+lyX8SW5GbjG3xUZ9s+OgjAtFIu0sBhlV
XFB0JMD3Uh4bpTAeCLfWNX2yw/NwEj3pUN5/WL/Q4208aEWobxw2kHb06CBfPKKp
aC3h6M/EUgTgXTvK7lG7WNs7LDrcTfF7+pRNyAVQOKWjMan/4AtN79IUWIuGr2xL
LRk9WW1g3gPdD1O8pIXUrQMtLQyQuG2cHy8zoto6D1n5dobheYQYs9WBqbPg7MnO
aKnG4ZP9DmixZ6/F/HWcCOAc8ocr8ai64VF0iupZMp8aN3F2lSfy8GZr1AYOHYkH
rlwViBsC12FTkf0sMk5vcJSMjXCkmdXsge6MAFnu4ZaYz1/6QM87/Z+x8Z3DeUne
aXv+/L/ZD8U5t0Oo5R+GrAF7QcUbpo9xEEk1OSTQtt/fH27VKZnxpytrCWRrBxEd
nA8p3g5zO6jCX0wa33JzYwYT9uRFC2tJaVQZupxZC62U0Clux94GDS6S0b8CkRHk
tqCrwkddti43jiyNYGdiRQHgdl590AXiLVyAOyqDUJEkwcM68AkZzPyxlBUz5y8c
vGYhtmYem5IS8WtJV2HOlECdPZohM+vtO1xhJGIQX5ElfbFt9cYfswHoBZUhszan
NA2eUMGKRAN3Rwd+39NtvpqFs+ws6bNGK0Yrp5fVRoJleMTFKCFhLbALeFewmr+W
Z1vsBBPy5TrMkBGTU/fsEAj7FJYRGNmggJ8NsCQYe++Ad6PO3p77dixJ5Xj+f9ey
BD3uQ67RATaB7/b+IYpB+4M/+D7RpzZ0oJij4N6GOnq5zL54uY3vhNyPpeT7H9bU
Wpi/DktOcRDC07ifikcKbN0nEOgUjs7pwYWbdDXI+azfbS/PJLfR585G+1Lyu7Gr
2riGQvsSz4LTwolDHR1ZGl8V+PaQRWuT+XlFlWmoGCuAhEFh0fp9KdgSs0yy3T1s
TkWVNcLI0v61rioRNtpuO43+1Xz362tXyIKfg+2XKnPTA8AyETnlnAlkGbVjH0Fu
Ju3jehhExVxukRWo7xuM9f5uVc7GG2hhJrlYFTgTu5ZDpiShi963bqXa3SpjSeZ8
OHxvWY/BbZidJU5WnFuZ4StL4+kIUDxty/uaauT8z1G2N9TcwDkHbduZjZCoW/49
ypfugWlR8iTy5JRplYKu04k5vq/+O1zPMueKXyDhSN6GKZbmKFUejvN0wl5yRzjL
qOZQSvrJGyTbWPeCciU/Cvol42ZBYQpGdn0PJ7YjYl2pQ1ysF77gIKfhlzIAJPK4
kOc+eWSD40JSUmD8cV5GKu09NCPM1aioi1UZOzR9h2FJUBOrPVtawYgHF2OY7BIt
72NfTtisb+qklU6D0ISrX2X221c3kf+qn9BR3XasDwBi+5rxyV3ehCkT0cvsSR+W
FwXJJM3QAbhf20zHIajAyjri9wg23sft8gB79WkY/FBAIyDraZ1Z5VtgmOM5CCi9
8zAjfD0x3IAgwKIegkYZUO5spDWtl5C+UWE5t/vyeXUcM6A400tLtuixw7SFS9IL
OjT0NEUcs7O//x7fgYb8ehnn0/w03OGTyOCSKdbY0Ku7oUDgvIpRTVRv+WV4bqnZ
EpwGcsAj+uZy0oCtjmcYSUdjBYgpJ+y451dpZ7igR+49GAKrZdMc7rvk4CUBwoF0
U4s3/v+a/5nXzIuMV/DcwSpHMNMsjFZiRllHGXh/xphVjyoBh8vPyXzNW5CZRWzY
ncvUapn8A8J2VatGGjbYLowMunoC5YWpKLjH5Ls3wO/7APuq2p4P2o+hmTOOLGZx
EU4JrbW+naOYfgk0E57DohhjxqeTctMiwG1dq+ct6+G72/YxwiS/KzKuaVW+XyLe
U0Ggw/5dSjNkNwJM0pS6hn2g+JGlkXDvYc8EF2dmEnYp4/Wp7abzBqt9iiE1FF+3
GvQ0gbI2cPGw4qZ3E1SA+9BWgJoYeAkfGYRyHKLaVVn6L7F6rCH/pyNV70UgYsM7
YZNMVhsQg67hHoH7LayFmeZZEYlJ3iIQt+2rL6hBfMwG3XLFw38/Byn8MwcUv8ZZ
WeWlTKfabo3CTlKNB/xS/enIHo+NZj+vw74Ctqsznkuzz514HZ0Ckhc86ROvY3Ro
m4FeFo4LmJpXjr2qAqH6CiY/6jYCq35z9Dn9k2hZQI7CsuhRUhx7l85hBXJnccf6
G+OM4IfQyuX1LcN7xE4DoRFNQ7+po78fGWDRLTbVzP3k8F8FJnDjdTsRtfeqII/c
szbjauDyCgPrpiLwcmRZyDCtbt0qzaWTH9FEf/ED1b15JMMOS/n/3tZPLkmK3/eI
Plo4uRuYpwzvyqMEyjJFuu7s2OUoOmdsgaSbMR8D3U1AJTYLYHJhvpysKHbioyQk
zVxJs+7pAEBYbidbGSyEov9KRjhp0+wEV4YhsqnTVPWzKvSmiet/n//JQIhScFnY
aLeEivv8w92w4tzR2ubFMhyjzG9LIoiiwFG2tP2N4w/bhpYSTQd3lA3v1lqGlOOB
kC/U1h6EP+pqp8qZNsEyCPnDK3vIovjf/e6PGgSxzAmN9sf8EOtTXTLcNX8SYdzt
tRQYz/E1SSrYNezRGv+ydjtwI0lvQZH0DFq5HwNX+Soc07NL2tKWldv7hamkYDjk
CcRszL4o9siOPbP8GLc5GdCxfKejcUS6shOr+mDx3+futHthF4PlEUCTX9Xq7wyu
T5Wk7pwryzUoLTkidzo9r2z5g09WJZyntRDX8dpz2F85e3odW3iHQOAKFM6/+9Zu
ioZkvbhw8pdIXZCNCv2deuP0kZn6c26K3nWt1Au06Kvt5EdfVPitbJzdN+7F3VpD
kQcEW1j6hy6y53xj+u+kKYQ+ebwcHI9xpQeTyQItF2uXtEFyQ15PYIEtRnyBHnnB
SQJCC6P0xvkZ83RPhk32IltqO82LOYOcmGTwmQotv6kvYomIgRST2bkazfZtHuWv
VKBoyAjL6bXvPGieDMH0+CPSeicTFCMYQ1MHC9folmHMp5j+i5Ozih67dpLaJK1v
OLJb6vGOLu7snDZdFPk5Tr70dhKFbvR4L0um80Um2eJKhyQ9EuBokhZskDeLgO+O
abj/mj92+iw7JkZvGAY1/OyIWVpDdvdgSdZ5XCBiyIAMZb+RytVIgbxwlXVNDDa5
p4Y7BEsA8pyEARvhrzCo283Vm4bHTExvGf+7P8oGy+AJHCibZZWQc7M3JTRT0XmA
C/6Ja0uQB1WqBxgdDxBvjK3X96QpK5kdBeWQRWvFHA2kBJEz1QvurJAU3slcIs9F
LVv0ZFtTO2BURhEX+O3XwsYCH8ziUakZDWc2LvMyVXZDaf0hzO7pIRPbKEYRgEQ8
BvciQX6Z3/BInAcIYJ7y9tL06Nwqatjqb65wyNsMC+2WomRaz7wGWAXnBaGItR4E
eS9gyMOlZE0mA1GqhLLr63tzbHBaegSArnDfsH+wfVSzf6q3ftI5lpQoYseI4KsR
/+bxTQA5C2S7HOhup3BsMUwpw5WF3dTcuBh5vhEX/EsVnnfBWhIpRaCg0tJBnIdL
vTG6tVxdfK7g79PZWm8UR3YiSC32pIMPGBjTPbPwmq8RJO9FAFtiS26kNtKhNSG0
oej7cFly/nCe6NvjE5VO28+RPFY7yZNdZJxM82QmCoMlGkqfI8qzEIAi0rS9Dn3N
a2QfPQUdxHknHhqWaHSgPlHjj2BGARAmMTTOqAR1l54imh+j1NCErhogjjQfMyXq
/S23uSkGpGVU26pEjp/nX3Mmpor5E87FimUs8/4dzzVrzD2DcmJ4pWDPNKikO0TD
6v1S1a31bSR0UHAJnYt5LSZsDBTDuw5v0TMKYomw6vToJtxMgK14n0E8Y2F1RpxJ
gpkRFSTUPRtGtVtn+8aYlVaEGRWQWRLplnn/ld66y70t9Sdi3yeQgSBOeAPJElBE
ySuBq9zCvVTBBYbsoKRfa1JpcJ1FYVaDTWYzZfohWF1XhtNvNCCzBwnyJdNhc50D
V/6HG0XXQvJREJ32Q5UVo8J1DcRAEICpj8095F0ALDTznHQXO5AhjBPDQi9IjxdC
iimeeQspplv2z8VCN7DlhwD98AGWCYd7BoDuwczGYJlsnD95Rg+87BtYAu9PJrGQ
Tm/rpQlrj82A4RLMzZjSQUo0bbtXWhyKq4Jz7ZhhuEM6LIt70j9S/IlqHb8HK5uV
TOJxsMJTZ9wq/oV2Pw4Aq67WD7uZ1s8CUPsT0XKduI3v+KnuRCnm7BWbiWAY37X6
rd5+KBzE8c/1ztI4lFeDLkje0arwREgNPtkVBrAldz96mANlLLrSUmIybcw7quLu
mPVrFyyqV6tAhJ1csPQGFkaTY2AJxz/wctLrAIWcG5Ixl6S5QEhY+ei9IPPUzvXX
cpdMFEsbo7VY9VZL70sxITUJcxw+/Ldql2MRTrhuUDQXgVOzAta1ogga3/WB0Kkh
IpcZCnwnLXqaqElxliYIRX0nwN6Bp5IHxQphehpEM24FG6XYL19QpBdBYwKUShQ5
hvUrv2m7kLvGGKr66Rg45diV+9m8mVhbVUUBgsPOhRF0xSXky+ctyppFhdWATwl/
WwmhsYJ5ydbSplbskS/PQLdJNgIGoPG476/ssvNBujVGtiWb/e4Z2NgNymRkp7wG
Eo9Vm9k03XmZEuX0q34NhQFV+mElt7nO6G0TbyQk9QA7yQPcqSzQrApDCGfY/dZS
ZLuM3im0qqJcD67wjpV7Hm31rhb3XHA7OLQ14E2/WZemw8ZwhQye9jNzY7oksmJx
8i9BNEbB2d5dwLQwxUDgh8NdLUVDrA+WRYrhtf/oeX0sgTyEvFwCT0EJ94oPA+5u
uBAxEjhQN7TWpr1EzjBSoRobAuA2FPwzkAANk66/+2LvIukKivDlMasatiOsBX25
H/74GiHyZE30p+bnHv9VnRVoXo3MafH8uFnyEViVQlC1X8Gioec/00nb+Tyb87NV
JnENlTgt88SL/snOG/j/GczOl8JUNjUpewemEkpu59DBrsllLct2guILY8Brl5e1
QBXG/ckbNsjtBRxyT97lXj+oOXEyCqvVwMze8kROWwidgA3cUexYhDlvex/N/KgM
NMR9hr60pOV+sAjRM6koYf/9vuB5sUc/jDwzBjU5bqttzNbaR40olTkO+PfBtZ9s
F7Hkw+Iqd+Ia2lCI6gowu0P/pCPt3AMS9GXLTw+oe8jK8q+W+gfYH1bZb2s4FBy9
SL8VADFh/UqYOyH2bbu3p8bQNLkp0R9MJTnBVafvQULOwPk9Uj5cdunYMLAzDFfC
Tb/3hC/ozLujqE8UF8CEQg79q+/pV2q9q5padYBC79qRN4ubhFLsrqGQ9r1ia4iC
avXrusQVIwVxNU1sg1yL1Mglbf/pouT7ZKwAAQly5s8wAId4H+fdt/INtNUvjHFx
DS4Lk4jX1eo5D/pBLR2s2vqtjGgLxTNRPIk4z5uiIDBzmq7rMRS5ZG63iJoi9P8O
Hup0OFa7akpdkiqwTGFT38RlgpHDOXCD6EI8Q1AEcXdmk9yJP7/LDsxl+6h2Uoow
wiiUjXtEjq87dvLExHWyTR5lQUJjISmsRbHB0zIJoJMm0EWb5yLJo9Jime9e9pjQ
EPanWIOSqvXKvgYWLJ8DK/BnPl5rALHAZgBBI9xgXXtTabEI7EcUPw5HepSqEUyq
jcZihxpfdiOzT2T7AtRxjfsIKELUq0GjrjxKJ00GcpHGtELXco78nezwTnjaeXuA
sBcnx6eLTNOEhdwCG9sSK1uSNkp9GIBtCZ1RL+PuBHNBdcz1K+6gEMnrjxA7fzzU
3PZoWk/ZeG4j/YFmKe8bqJNt5DLKLJCYDPwPHZCF99Q8gytKeVTLU2kUBDA6aGGc
WTGgIISpT63YzGYfTujL9ZTjneGO1Hvske537Wozx4q/wiopwuQ1hC1ZhZ/Xxx9P
HGT3Xbo4YFTsLDi+ZzIlb7JjlXufagRcykpqgHj6zwI/0lCr91CW00GC5HqFXKD4
3+m+cVPC8ckQkwUZaUdGuhusEgP8iOk4IBQtRrHG/61sbG70dtElDbLn/WvTAubS
8DX4ThrBxcLYAQk410SxOVI35eXcY62Si3BRoWXshNs/C9aCPAfT2JPI+brR7wBO
NpXHBzNuLT9rrx1yaOLUmM8VX1dKFRvwu4Z7XANiwQpZKCCaTpeTq3OLYLnq/Iad
vHavhD0o5Go3udO3v5Rt67BwYOGQtTlGOqf1dwy0mARWnmUUBkqBgvPbUFTtQ79o
bOPfFUCLrnNrZ9TVCRDljug1TOn3+hlxiKTZeMIuSWwJsAx9iGBqFaZE/HDog3VC
oqv0a9gQdFdNrYmM7wrFN3RANLlU5Z633c7tweIeK918A/d5FKWorRODv9V036KB
6++mHP8Z00mTXj04K/8x10CmSW3XhxCVEAlGACmtQl5ai/b4VYzjygyM/h2FWB3v
hej9tvj8nkuuWBA2fLMYZFdIQjH1Fzg8EZWJRhJRT7LSewFziYdLlqi1In8juRJh
yMugUU8qqqST3E/vXzP0x6ln69B2UcwhymSf0btGTR6JY+aXKPzJvLPgSww1O7qM
3GIRBp5jqs+Xzhytdec4YDHPvmfRGQJVv/nGn7gRZli8Rm3bExTvy8rTuyixJbRc
au1LSU5o9DnnmYtNbF6B+Yf6Tc7t6ElKy1nAUwjBp9sGEQ43NGIoQHbau3G5imTj
agMl+oRxWJTquf5vdqxGV6x7pNveBTUXE3A59Vn4sxCJ2GkfPpvw28rs1LzkCJgq
qYMlkmfdiKJH5PqTlA99d4jp3sx3/nuvMv6NeFN7eufwwnAqo2Ji4dZQ9u8wDO9i
vzN25sH2WzwptJ+IpjFlN9CVdOEb+J44U36E3ztrfleBif9rg39iiDISP3gXpnNa
MPU3MpO3XanW6jjRfM41HxNiq8DdiAl+LUVO6t7N7hSV5UPN8M54ekFIILCrJhGs
Xl0ylMIBtd4NZFAKPUcaaYsXU4E7lOeuOQIacTcT6BczSX1HA4PmXHOILF3tXLYB
UvQbT0cRCdw+01hBzyRJS2+edzxUT8wqs4Hh77zhJJ1MxqPkAg3kUGlhnhvroN2+
4D3OUSy3j1TLjRMAKmdtPwrEpxAwW7h7h54TOnlMOoUWwgd5YDQnbY2T2byNp+QD
N6zlt426TrKTczqliaJp/rAt2FHeT8ltTfrKveVRmcEAc4LrCONkqNAdYbY2VZxG
PqPFYZbKE6qgepTvLyarkE0sV0DC/hVEJYqLgo22op5fzzFdDT7QicKrydJ3E59H
J4TkwFkp6KHnFcDMwSuKh6lUNTpFJdd/jJVXGBO+hpo4+og0g93NgDZXAvIA5X8N
qU7UPjUj2bL2Os28cWOWJK45RKWx5T79Jo9SEqNj/3eySIlgTUVGvUi1ccGC0kxe
+/Umk0KOIAc7R5iHBjt0Dwgz5BSo0lrNXca6CZ7wZoo2YIIuSaS2fyy9sqJ5UnZ8
dNw4L8HXdXG/r3DKCobkEQ/R1caCq5JW38vbxiOFRhHFcBOKPFDu24ObbcUZS/jJ
g5MlD5f7iQ2Qxhtg5K+pjRHWnXEEMuJ/A7zFhMZRJTaQ/wTmcEkFFCU+wH7pAtvX
gFX3aEi0wi2Nuz6zVYbNer7KLUkABRN0svqEqHk6PQo8ExF6T7Qm3+jn29hYHqBZ
8ZI5BiwrEVAFRtJO9ljnUkQux9tig9XJskuTF8LzKypCYftP1U/YtNbtTTftRqE5
84VxGu93Xgiirs4+hyNKIJEKT58YdMBkHzYbcBBFAzdOG0aiut3Es7bQoS+RCRnd
gSieIw9ER8z6R0dKIQ6gf8naHvvQELESZea47XUKc2m0SzL816UuaCUz7ZWxMIPg
216QKr5aMqknBN5DxA9jQ+UUy4lA4z0JO5iWAMTCdsTtGC1TbJR+p/82QQWGUTLq
3emyCL4VcxNKuOpU9xHA591AA63QD7ZKEykI13Z/yv2SPOQjkc2XVEviXmTmr60g
W2hhhdmZMD1/vbCbA+dqECUjUr76e08PkAZdeNGTTtGkBMJ+kj4t3h04tYHIao+L
hMMa284hcgJyZHEEvwOB6Lr8c65eAUxW8naTRpN7NHeEk1/zpHediZ+4iVm4y1ZD
3RagEIeqRRbpibIUDEaPMw6hX+tg/ZtEOoHcVul+rXnulD+wMjOYgh3I+agLQT6m
RG3SvozTviInaGJOTledEVWlfKklP8Bc39zc4Z2ZDgpnMWmkd7FXioq3SFgmW9yY
msQHVld3caFqBmCkq7dH4S2ZkWA5AdngSoJHENfEgjEmFcaDfaTRRRenCfcRz2nL
MaDLa1yO2CjogMmkt4J8PCAqCMKeX3Vn0bIpnCTi8BVDFESf4HKVM8YY9Je48dVs
zmq5JJsjemVAwV59zsrneC+PSegQoHWLJsUJB5NPQaF8wO6kbtZf1ouLvFgkEav0
eEY1GV/L07r2xcTBSlZXtZb2hpP2D0ufGfPwEnLHaTw7S8fSgyTMap/F5NeuNsmt
tgGngjHrAoVvQQHAAPiDvYMwyiI3hIFHEu0OIm3ghgJs41XeofHsUb5A8UTxyzH+
RE1VDsEQRMVJ/DgbL+SjIvX/TGYFpxShWBvjRxswyaRr2E6l9d+LUfDqVeNl2tDM
lvpPe0mBInUv0EQo3GrtiV/Wk4ab6XutQy9I6QG7rUEr6lYWjZ0qpUuIZAR9S/AF
jEE5EwdZK3PmrDnxPE1pZdAhQ6xvpfYyR3ozaIDRTZsVX5XWSx4coBQbHXlf83OD
XHvSa80p02rvvyGIrg2LOWz4tlSws4vuZU36LW7BURtun6aImr2+gW+raOq7f2fW
2X09vZdmOnbOePM/MV0gIvAljEj7T29EPjxCyst33A8wAHwkU9sTIYDw4CacLyzz
rhaxjoO50XYx75343do6sN3ZvWTjMpgoRClN7orfH3N76aiCQ90XQCc94jZb4jhq
ATCisZ09td8DMlGqRR5dlMzkSAWfpEzkqu/cjH2+yy2dxnfpT4WJU0/3RCkiWwdJ
YvH5BO8ZdN7hVBArNvcpo89K7Lm9mN+pLWs9PCdUZaL/xFI0w/1BTjs2QE0PLnuc
G+pb05ngL4R8g3JoQ+AGNPePuSqJ6DebO0tp9lXNRiSPVbKuymhdL3+qcuVU4tBt
00Bm+wLe2MtKG0dGBqMQydMyxg5yKlk5j9bW8DF3d6unXOkb6r9E0JnENNkiKKjx
O3jcycSmNG4U+ZLpogXbH1QOQXDl0KS0eoNvLbj1bF2EC8XDwCNDM5JL/Tb73qEr
u/rzxIkh5pHlPLSE8ySP0xfKYuZMl1mFt1OekLABAPAxuAjIKPAAWpD6kRbje9rk
A87FBXXRRjay0byO3IAjf7ZAZGGThrjelZvhXhG3Yi3ck1y+GZA5uujGN+V35s8m
Gi9YCg/Tfr9vs2qbOXFteQ5lbVORJD1iDpIlCvhXy6uuK+Of6S7xsukLlnN6Mcr1
BILCvyW2gREA9DvuhfBQmGqP0scfUUAJ8vUOIZ8pMUBftAl4+JCAHUX3ReDlA0Ny
z+9N64aRDW5TMGvnDT7WXHFHwTAUVCiTRDDBZMIclIQ43oLfdjunY6YiUo1llHVD
9Dg7W01Jc7m05OVVCIfjYdRsfwv/ylnWcNtHx5wA858PAlygGu0KWLcXo1XQlth6
N+PMcboaeIaDw8S+lQt6dW0xsUrREF07AFV/811FrDhptkwwlKfEAioPxWla4ohI
0EifVmVqLMdhQHH2eBHzRs2PPl7/DXiTLn9OIgw5ciS+oCzfOOgaObV6vz3/u8L4
mRULPi1rb1Bp6REH/30qjdcNxeBzXB3OoVSOplhwt/eOLbYCRggvvRg3uyCEeZWR
2IjFXoIsZCNroJ9+tSyYgqeTPiPV7ieW0mlxM8sZKSMbYlphG923aFnU5EC2kgyh
iZkh9338d0sgZGbnnnPzrdF7c91R/5wbyGRhEoFDKNc32n8qFeKP/c4OQFr0eFo3
QGItjW50/Bo1hF9YGQXSEcvJ0cr/xrbmY1YhXb7VsUT3I4+apy1HrsqxNm17A6sW
qllQ/DZ2MWxzHp062GUHDp5RbCRU87LQH+oB4K1Qbb6XuVo9fEKYdylp79odXe7K
PvafrLls5UASKLtiNLKCwZD1KcuywpNQwA7E2CkhE2KzH9sv7hZZ4w0ZQBrv6LJ0
gr98nYMvYCNORDxI2uNSzskzLWt0B+vyAvgUJian6ia1fIsB7/TbBzsB7CWf7+ma
E0R2GiGjP3BG+z+G57ZYp8LwkU/7hySgrAqRg/f4RN+QxfNmGQv9GaYWh7f1GulZ
f0fObHeYLpabMI5oum0G/RflR/707ch7TCbnKg8i+nZ6a8hij+hyETo2ws5ZaIxX
vJf/uJRViBIfL8pw5jNw/92UYqJ8vQxHkF3qPKV1AOrpksNOnTV/Oqd5wVSuxCNw
mvEXkuUz9gYBHGX8L1ugBmL9SD/nGidlnvWgmasbvt8b0OicpbvUFqpyRXoKhh5Q
rLLyb4msC7o2UuxQhX7eapgHUs/Qnj0wns60wHU+eqMdYPo4o8UZqZPFznjozUTo
qUUVRncQSRUXdGpf6A2wRbx6UlXcCm0+K7lSL1L/m0Gobm+4ZOqQAUAgFS/gGhv1
RhEHaLzcSzhhV1QHg5WD44YLtN0aq77mH5xZrXv6O4dMZBZFLeXfLYw18BFcydtE
v0HraWbiim6b1QM0eJ01Reef7BXTr4kaFnx6RtYMXkwIippp4T9NX/mJqIGnsmMW
jEBUuLnRib9Up4h0k+8KYqspgicrZqHgdR64o9nBiLEU+JpElL1t5BuOE4RCnSk3
p2AZWeUwdaYmfh1ASG/vL5mPkSUxtDGiz00a4gd2J8gIyf8JCnjeOnwcLlMEwfI1
sp+0oFnzFrPSM9B3bzmPt5gSOXCa0pJSPMbqqgNJubIasyXdDiSlHDvDRsq9GTVS
8SL3f86JvVwSbuHUNBBSMXHzM04ilCqknV0QW2EBEUG4Knn8a6EpQ68am7OYGRyv
7F1iwSPWnkBY2oAyvpFfXh8vNc977HrfL72/WEvwYd+BLWlcehzpDD2g2nXcVaMS
wa5HE7CThicePPoCwJj+/Cy5K6Z1MQ9oLQEj375fWmjw+AmMqQwEdU/ovNQP6Bol
N5UNMS9DW1NDwjJfJyj3x0+7TbH7ZsomQCW+6BtlgJKvHu1RfgkSveQCgukdWVY5
uuLDVGDCdzksELZj4eoikx6fWS5NTps9wvOZ4xa4BXlH1c4/0ZBoJKUmc93u2dE8
bkBtGNthxIYfI4VD/V++/9wUR3Eg9ri50PoRlHPbSY+40MlmslqXJabrvFKKC2vP
TiUm53SAlEmQJzzTTCPwNVkmiIctzQfGZzQYX/8GcUMMJGr8F9mQo547mAjwleJt
q7s03yxA8W/KpIFTGDC/srBcZWIIDvF9fJuxbDH1qLX/9+uvR/9nfQdV7R9BoBWt
CYN/JjQeUL8U0aN8SkL/FplUjLvvM4u/D5S93LCl8IfQgVHN9bsk/xGpm25Yv2Wf
IGsrXOM48RKqGm9vX+/02Mi1PSl90KV1uy5AhfmkuSszqbaa+JZnzZnvCLMZU/6O
FNcrOqecNTSnisEbXwELB2fZfyw2WDaWjioxOjl1qRRQh0A3RjmVbp6N/flXjYhU
zbwU8VqiQoqCPDKFDT9v1phnHClMVdlqLApfW3DfEsB4EIkuNi3rWzr9QlV2I9m/
3rqwtqteOywk0qfKnHKDXzXiYipsvGJywAmviaw84LzlDDvzQDTE0weMWGUVrbPJ
pVWimnOKHmr/jo9S1gF/dl1TagrKP3d8iZP/8RXUiobjtzZUmjan8fbbvU16xFUW
Xg2kLIeUXrZ14PfdIg9gcz4xTtiHJ5H4SrxgSI2p2Lm5AaxRHD293GnQ7jNx6N3v
wvqD3w+9LxmpjR1894KRkt24AssMPadOue/uXoGyhyDHzRSDhMWgktQh7gIRUJXX
+kQfvYRpZk6TfDsskRtJtN//d0AmH4we/rZgYw6/voNEj+f/Yw7fNz5PHH2eoNkE
pFSU2xomFGsptayyVJYWNn7jyWoXI4Y2BslzzEv7sNATLCZ2htP6bIJoQ8FIgW4K
y4227J3G7CqmSTd9ZnMN+BVEKB8EvnqqGewUcZDJYfmMFhOSLZLu/bZJxdylLz63
Byu6+WUHGqxISEhAUUMOBhVEBNETMCjqs3E72buxqpV+lWG+KsdbNNAMYPI9TW82
`protect end_protected