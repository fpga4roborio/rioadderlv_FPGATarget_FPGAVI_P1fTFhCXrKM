`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
ddtXksX2+yylW5zu6QL2Lhnb2d1sD00763mmSITNX595NcHTEkwn0zB1Dry37fOW
FufOhVzEJp80NC5qZ/+F0Vk7Ik02dIR0elf3clrjeJRK85K4e3Hoo4xn7YbFUIms
l/8VZSb14+JVGURjfswrIyCUotIzlzVYZ6gzoZwDXIi5gQIBf/gI+KxNXPaKV+PQ
Ufys/12rjO6aI/pPlqSm0hCvftmBcnezN2hk1UeXgOIuKZnogjOsf0iJVX2aOOWE
6pD/psybjbnsNB6kH5uFTA5frkzIzkzl5d9+YDm9OyC+k84E83I/7/j+rk4L2dah
QJOvksSIzN867/4Qt8qYTQ==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="MvBXkzurAa5VTw+1JJ70nePUfoQXBvZOku/SMmg4TwQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
oRtzZL4VJ4iwysPsC8SXYCzXS8Fw2gtZTOskLcDV+1B9Nzn1zTyNtlo6lNICRmmK
ZRVu2BmCc2G+fmzynYlNTnSa7C0Cuel6FYpxCBlOuk3OF2tzAmLAuDyOH3Z1Yjzk
a0aHuoCdIRKv7BrZCdALt03JeUmXKPdOmIlkVGFl8yw=
`protect rights_digest_method = "sha256"
`protect end_toolblock="Jn9CQpRhJt4rnzZPRk+dOpzAubz7omckX1MrFd4p81o="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 17712 )
`protect data_block
gD6l00tciPUa6pDNTk/+tzLxvdHE2s3DQL3/JqqujQBC/Ei+vcAB8wM3doqg5vTg
mdfn9XB1bLOis2CVSfu295W2DNwHfMSTc/8BhCDRnTlLIX0UCJs9Za0+LoM0rMrV
T7EjVWppbP+Em6PkVKCwlmIQ7JKaifJ+Y+kjw9HCGboYo5074hY+K/CBbfsBQY86
AttQWvwZMXuzUkzKK40gKsAIYQSdb96PZ0XFXJbQgJRMcwss5YIhekNN/F0w/BxW
cOJcEOm5DP5tjDzA20ywpFLlrxXfLqR33SxDoJV5paObHHeRR0bq57JnNa8nkBiw
IahzfhurAyy5KEPMQnpVWFkPBiKPg4E12uCmqHUQUsIvvEiixb2q3sUqIaW9Qdna
vhyXVOu10SmEZ4yEtbOKgXaf5U/GfDoCpW4Fsj27JR1lMRJfLa5dtvjemvCJ3Eox
9As21cjatGk8q0WrOCrc/TvZg4uyWKqUV1zzkCgVkA54x9syLWCwMcGy7MkbAcDB
ncAxJYW9KOVTcl5PDx/31Az5+zCzbI+yebD+oaspuCq+Lu2i4POxBcqdOLKQMDJF
4+TAQho87iMW47vrG+obuUMgeN2uOKeYPWlOPSoePHYJ3TWXnyghIkxRwjoH2NLZ
yj7xC5f11GCBmIqE5JKRu4THYKyVqWNdJ3UgYYuwMvJ+bgwjiXsXjHw7XYSAodAC
+WHADUV7qZDOMkEWnNTQFZKDTG3YUZJ216zG2zjbss/ws3jnXHuCHAn/GZZqgHQG
ortiJWsaFtdgpavAwvh1afpI0sBoaKIFBayUlZPUFBimM30Zm/7yavIeEunhC27E
rpTcmiINbayys0RPe88Fch+9tCCHH8K8EjZLAnEuMLZAAwB+17kEkwvZejl1xdXh
fj/X3GDmsZ0/9cO4YX1C6pZCw/NmfxopVjX6A8FCJFydKgdXFT49aSe9fFs7DX3v
zdbinQwBZHLyCrk0/mPKD9dXz7dHN6lwVxApmlKgwTsOzwdvLmIibekrvbo/sg7P
2790UZQig9Ny6LP6dXdurzEu+mK6/hhmRq+h8hSaoHeJBvX7AgklmLySWUj9x8dh
b4jDx55o3iXECBLD2otwAmA1n394Rkxa+67/J4zhhY4iYkCG+SMXF+1IYwg9SoU7
Na8yGrpZ1jby5RrE74yemb9M9F2Y1+ZR1QTNPzTQ0YRM9hfl0tdq+RThaoELhvBq
vC5LX+EILlje2cJQnUr9stHH2ahSdDR262gSBpZbjslDdmh+GKD6r5q28Zxxcv/P
2YGHP+qoQ5Jt/UjEkmHveeeWO3m4hdwFuGL8Qj8+6iLoa+QwyJU7N7az18t/QKsN
GMmE6hE8Nfnu8nib/I3pGr+hdFmgf3xRyDTL2ad6R+OZ83IkBNcjxLstDNoKU2ZK
k+5wQpfVaLSXbTgT4bMEu/7VQkEjyKug6EQBEzCUHwOwcgq89wbzUS2wAmhu8UXz
+G7rBIGrbsiSGp9Adt7RKRO6cxE0MF6jPs6ojQqScALq6fUE2zdn3Zj44RtOrRkN
0V6FXmvPhRBltwQAdLtWXYC8WfSL2wy/dV7e6/BfMYPnQfL9NHwX8qFeI5FarH9P
55ihCOoPcabSKn/v655/4JWvnhcycU9sHZ3hcufIcXCmfr65IKly+Y1smhJYzmrv
5ti47Ae0iaDFgqlAV7vMBHumslXNTi+Nn5dnzGzy4orCDEq95pUHRrm0VsdZnWXS
/wpPk+nW5OOM3as+rmVsCvyqQNGFq1sb+EgEahY4e1uy6ivoDPS5jGXhvU/MSmhM
i+v43xnRQ1qpgeP6pDL9TGKuqD9jP9s9Rx02wI92KD8mIdehKH4HBIOPDF2uMcu9
aarA5k6ZMuz3c8s4/l8MbYALafzhIYBK0KLXlsgO12y4zcVFJw8bZxYJJx9VJgHr
E0tXXFI63uuz4BePa6kvbieSKC09IevuMNQ2N2m00quQV7y9yX1ohp9gPyvYJjmL
RnYbg3adBwIN6MAmL1fYptpIjxT9+JFyKk5Ppx47o/RmyYFcGpSGyChqJi4h6AaW
lCdEeGcf6zJTde/Tj8w8lLCPoNGttCJBwgE9JJu/P9fxnwx7PVaRTbTLeU8VZ91u
DALywO/KVgyxw6FAbmNPCJtOeQDWvuAgwA9HBIQFdldUkmlRXFy9OZwLqjTWcVtn
PPM6V/JceX5shG5t7Di1x0IBN+Zgl9WmEKGGqyYyPyUb7vFfvJAgnnVNXAMcvffH
KFxpcwkP64SsD5hDOtRHxEdebfWuStTeWpOet6aVmUu0VRaSg9yF9yCFmODAODI+
Ygb5GKgVWEumhR30XTKnC5Y3YhJQDJ988LHGl0ZbHlGSmB/DSi1z1Dsb1VbJ8B9p
AHkVzIODyns02AHHHEgNBHdBPemGKsTJduJF0FmMJaEj8691XBZeEyoEiOIIxAMT
GKHMDMdjUDNJsmOJ2rAO3HNHfxyyC+vwLTf9jdbankxJDtMb6LfJnDPSLgWebm6B
PpF3QjFMQp91ZQZudYHAYZhHxvr5pqPwZPc9II8pjulHS0918LvEiUSSTA0CggqU
OzHunIKXwDzYjK4diTi9p5WHK5QCpxq9Pv3o8ai4W0sJzovutWV0bJPvpvBkq8n8
NN5oQvOO5xcqp0+5FnvrZVrdseHBm0TBZuQ7HTDqxRT4ZM/ZrzWH+Dk0OJxFhK3z
D+q+n+zpN3lrS5fbQuO01H6cX2HDyG7LUQAkKgXn5dTTGIGM8JXi+1eSa6SUh/7P
fNF+uRGg4jTlAkxVBx4F7BH+nxOw+2n/8ufo4CzIF79PbjULpSWeVsAgeFUoFcgv
1Dwlb3z6JnVhEFAjjH1IIdg/pwrJCuxJYHVncOELcAcFDM3barYjplhEYQPTdhEc
d0UN0XpFFG2fGFDVp1Lw0Bx//OZXXBk+wjE4ixW4Ug/7amUPgWZpaOqRtEkyqeKf
gVyFKaUuU/3lFDNXXlo3PKzOoOVZWcI0KJSjvFo2uJSV+87UJ/Aws8StsVOOMqQr
1OMLAueiyRrg5x/Walx7LEjsdStoCj0wXoUQFu61hJTKKI1+aaV0dXgDC6sJCseV
Soxi5DxpxtaEl9aOtG5ST86whvWwWzk5x11Sy8oPMgL6kjVVDQdMVSm/ZGiU7888
m4JMyfYSB+ox39+Oecm8ekhNvJw8BDUDegkomoJ+HkPLYca74J8WAJgjQHqV8mu9
zRa0nF1SI4THcUCy7+02Gefh3J8I826afoFTHzpD/4xQqXrUuyzTZ/eEZ+BsvGow
jpKcIVMyA54HmjT1du2lhYvbwMni8P68SnOdAmmxU433YPPGgEETlHiLXciHJLFG
KEcdaqdUGCEaV8kHIeKJILB4NhlEVbLYNM0wiIBGKmn3pufSId96CPXVX6HKlXnp
vU/OOaNgjVYSJA2gVHXSDCvgBeuLHVFDGVRpNu7J/tk66LOQnDrAkwopL9XSwTCs
q1pXw9J6+6kGQI1KD7KRNNYuAsqFQk+1nuuuW4IVleRvPICPlVjgpsN34UxO0h5V
XUEqcXGfo60Zp+beD0DhQGJmmy/V62Nh8wEOMxori+oH+880LI3DyqVRcF7hyeB0
dJ7mu2rJD3+NB4mw/2Z0hqdT2uw7jt+X270cMdcFYobyVDt9VsnofmzhPukH9YNB
N38SWXDkhtYySTyfiiLJyCj50RWfdpFag4UxR3gWNDjEUbiEi1FkHqmqBK1Nr4kv
KcFaRTf2rNhT1AYZLqM3z0EK+CjrZuS6U5mcv0BDO97lpvnA7YQdnYfVsS1Z9YvR
Nm885H49i4QXPIOXr7Dk8ykWlsXYSVHbVe0sEqwOi0ssRTN4P+ANfZJMZ/FzIcPO
jEqT7s/xTV+b/e2JlJI92gDnMsxFrDXsm7lYjnqSDNnRdrmHkdNxisoFv/wIyiWs
NQjY4q5QY48QiEQIN5kaBMSF9swd3lHv1mbEKj8iJyX+JaFcNrYcd15wi7pOkykR
mk9ibxZUNGtNTg38hDPdZb2K426M6QAQ3h9z4f8KEitDKi0LxVC14ic9CMIk8Dgz
riBMCuhqZpPgJ9CtNq84t1j9qnS/9/p+7trIYLgBepq81hE0A9tB+SD9AtLO6y+e
l/3bm+jtECGRaUfp615XxK9yrsZ0Li6kVQX3ChySgkKHTLLKQJ69ul56WihRWq7c
ekTyj2+5Y7iCL6U0TKc3l9anuWnz6ZUC5MZZWFGQvddSx7T94fu6xtRevyet1ux6
upQU0p25a4KY3KtekMo1EBF/dA7agHcnZ4STLrgsBAozuIFZnVMlALwEyWOWwcsM
b4Pe0Yy7dzBJ3Z5e0kKXVRNGCaBEIcEonWTAQ5c3TCeEtF4LeFbYb5Xare2s/sH/
Zp9IC20NNdkZ04irXttOwAV1+h1o2CRKqiBJKl1RqhFDuHfUgcxj0BTN2gXzcXnr
zrGYLh43UZ2YCyU08HOmaymlxP4pvrSs1MybiowTKRA1ivyXDJ7waKyWX0ZrffSQ
IfMTJhYgmNUrZylsrdK5e88ho2/3VEKlYzaZ9z0Dm1hTlA3chwSXweQ8+v8Caip6
yaJDykBdM5zEZXppvsQDTYb6koxz2En7ItMyho7X2jZcIcIhsXaKv3EimfCjPtLv
zJwtf4RmVHlerUmVaLwNechY1V/7R7I9bDJxefuOcv1Dqlrf40v2G/vKZRlApWX0
t7GF1ek62tSzb2gNxXeb624pap/Oo0vidhjn91n2u5S5J9nIBjKsA/6R+/ir2rsi
xTzUp7lZSIjtbO/88ZOSj+sJn0r0FpasTpQfhB0HSHdcyD5RzTy3V478ybB+IoUW
MJfYLFPAtys92R803gtXQkHoyiZ8j3+ArU2y+AkNlUHA0BsZWkIlZWNk2mx3vf4H
gNsiQT8EJOQHuraTi0EdzO5wSUqWoUGxZh2defca+J7+TSatPHwyUW5sNs5OckOV
A73mugaSEWwPxX5Zx6hG/07yyVJF+eEMFKK0xK+1J69fBJpJTVRcODCrmofFTyd1
b+8zUrxepH+nxIE+KVNYlOfdfVSrttPpNdT1p6uHKfsRPvnpFKH9DjhRtMRhVBov
Nhrx7AQ82yMeR++Hb7sVDiCKtLFWRc4CvoA1d98h7BTqtB3l/ZAGrYDMYFc1squ5
TlRo/2kfLz1hghA2DgSAmfsOHyX00fMOboGNVirUHZpKsqrluzjm9ilWYoKlZSyH
LaSEFnh9qhRj02ogfGAGmIzTXmym2uFYjB+Nzefq7WVZjj4zvkGM918jV7j9o1U8
ZG+WQkecC3RbFYlTApVw1o4MLu2OO/JNBEFmW8+QExuYiLiocCFJVmmWcJleEwDy
PwZZpDefYjnpByAu8B3zmWNKmU0gWfyFkC+riRyBL/Wc8c2JdEoPkw2mnTIzJXs/
mXza6sFCmDGTzyHi5X7BqawuIfvgzwMBQnwc6KAGostdSsSWlSQw+5dxdREM9Kmm
cEqcCFnM11Tt6MqVXpSjLJOxubB52xzZkIyE5eehlA/t7ihw34DeqrLKAob9QmGC
5syHrykshERA1BWXBok8u6otMLGWgR1W4hNZsti4D94dcJyLYoMQSI/E0T89Hb+t
w9+RKQ8w0z3Dv0a6rvf/nH2WM73Nd0+S4JB0AQ93KLddnvfLYD2satTb63UUb3IT
MQxEPg6guwuHo1W7L7NKwe0hOyKonq/+dunQgBk8HXbYGVzPfA6WWLRto2+w5FcL
ou6JKSGeMafyIVSwTD1AtJkBxh9cm7wD2I7p5hIX88VP3Y6jF5Kde7m89NCUu+m5
3Ix/JsAWFzVMAZhGrqB0AImy8HwWiUzMNCxOlWHZ5Nlik+mhSIpJ+vZXnJU09MJ/
HFwCMnBy3HX35a7ERS75WeOKQWjsQPSa/uxb2qWG2SS8OZKTpF/DZcO6jSarxGcJ
v8EExxj5wh2ACykEMr+QAoF3jc8OsT++1wuLYgWP95GunMw6jMDxEz3uOpu8cX5b
raUhTr013IOlBCt8suuBW29TlxkDXpAjA75CxzDzCjaQ/fYqZ2WjS8P5C7+PkANw
mwVw5I1ikn8ezFxOq0UvEEoAS8d8082MagVwqFEL6FqTqYWkQQZry8rKnyV6ha4V
qgMFHV2vXDNfTPH2UBK3O6bRmlR2KZSAplCOMkNsmF676uhcIpLtXQ129xZnI4pU
rurNsrTKTBcxpWWvn2Cs4nQTCj/ayPXE4A3jctap9ifkSZxoJN27+rLkvC47d4S6
fQm2ICF7tTjL6I5/D2Djem+mDQyk+rTX3AQ9wp7nGox0YtIJ4XRnHV7XjB+kVCIu
QBVXm3mclvBrXApU0eCLpSmAQH4j0SElxdXQ30RNQLBzYtt1mUPfcovq7wUrY8fS
kLlkYKcxhfoU7tfSMMIb+ew3mADr2kN1t8eTSszRSJi2t7PXElt7q+E/v76aardE
Cp/+cxgWreUjTTIlRexhbokk8WCxHsT0WDMmpAliiE86uK9eKTgw3TPJtMpC1o9A
3KBY4kF9ekTCg8qnD962mxBkh79FBu4Y7Jap4v+kqEtzth8K9UKRBt4f3DFxgEcz
nRFoQbnDeIhutQrUJ6+v88aw1p8leBzh53nP+jxHj4tzvsso0D97GEauAHmWy1lx
9TUk6XSKH0YhLldS6W6PQ1VPB41skPVXjZF7dLRt8fI0fR1PdO2h4Wd06hrDncyS
2BmWPiVkvI91+5O5jwj6Aa27XGYFbo4MY9DhVENDEv4ba46fkZkhFOHZdpNtyNex
tfOzN98UabqNlZ8wOSk8KhjHE8rGs+zrg1LaenXsG+LFvo+/1P3BsUaYH4iD7ID8
PWIX9O5p26Gv0SRAxpb0p4OjhLcfYyc8AxNDxhUvut7pSpaGjTTKMItjytWcf5+e
mPs9YWau5RSMhfrLbdsyjuyRrKKVbORrUhHxdq3VcZrWtaLA4LTedIwREDylVhRd
pR+5Mwjq9gnFGXiU/TAZO7q+6/mfqQ1jnsODxQKYlFJmiIiE9CUvFxnlfMsKlQVU
u+g7wTDdAowaSzPpszlHgSzEY3batQPP7zET6NN0sRoBRHx9GXWzQXEtFmfTonA8
sb6YT9eEO0+WgSD5Oo4rRt+83Y42CRnXLf/q+U8eqiNrE20RnK48Y6HBB3+LncrH
T/nO1Fa8ps3E5zag2gU30D9jrk86nlIUDJGHzPrtpBKCFN6zTJzhW8v6ZP6FLbrz
WONc+GmmYRRsRgbKe0sRUvgYLyoSU1waWeEcf6tjZR3Zk6XnVq7+Zrt70gdUMTpZ
McZP1TO9leS698MxE1rFUF35B2qHPSUnpRC+f9zSxxn0bI+KWBX8EEITp4M0s+lF
WAHaVPDQVlsqzXJIKUDEaG90Z0IzatYYt1+gc3DVHakyBY1pJ3d96WECmlzYMapY
D0icsMEVfLxr24bO8lI2RyzmQrJMbRnK7Gt2SEsK4SulwhUbmoasBauITT7P7sQr
7GSjO/K/Q90VlyOfLxh/7Y/X7tQSmE/zqLGw9VK85OjcV/WK9fOTSFy0VjBJ4ESm
H7dS3X2R5JvfreIL6EnDCw4EDUoddNp8etqlZi2j29/lfXlEgOl5hRdWTN30/3hT
kHfqj0KuqIok6Js0NMMYMiA3+1osuMLhFC7lOz6cmOz7zsnve5S/+sL0CuqI5Osa
m7fFoulNdBruvatBqRZVS/PstL5cR6pjRulP5jVe9S+9w1AtAUA9MKL7UcaOFSux
g6hl79k4e3qscTJ8ls/d7zjSgKXetzz25xqu4Qtj6QkLxPq1rTMda7KJCvpZ9Mp7
+SrUahTrervVJWGhjucxoqxJXFdGyaLUUtCRszCYaZ+dCNDy+CrGBYS8a9oflfvs
P+sP4nBIe/EwQL6EYNOlGk+y9OnnzzOc7eBXeIDz602Zk6A4tEj+pkavcYuJe0uN
kNX/GxmEYUeTEavuCwVIiAf5lWPxevosTlA1vAZy9Jmyrrcm/kRt8m20fj8P4jG3
KXn+jAv18rLYlbCJiFWhAzRCYOwiEttIoHZDb5JXozynF3BIAnf210HAWYzG6iSM
75lrYzCfpzdGPbcM45g92eMX6yhAE575bAID2hXvVrmJ4Am/LEpANF3TF6BjJ+3e
9CTgGfWzqhKQerJFYKEH7VkgjfNt965jmArmXRxXkQBhV2txcTtjaZvZ+uLvN5jM
9rFugAKuNtv8CJsu8kSU4EF+Km3Wry8yKlEeUGl4wNv/yRQIFAcqIq1NPsYRz6Y3
9hHpOGjBVpteLFOOftqFyWgL8FTjaZYdm7my/NmfWIrm/cvhlE8c8/CzxrhXevbW
6gZCf08Pa12+4+29zedga9g5n2KN0U42qLYhk3ZcfS38mrG1wdJo5OvdExDqro6U
mUVaYKnQlgWT1fmqHP1TVXwzKu0I8ILSaBgcP4J6QODgIG0DgAyvSpfU7Ar0VJLu
WAaorLxg+VfcHgQqqVqsK7z5Wiq9UjkItcqvoFV9NGYEGKgaYKiI8FjL88UsL3nq
tkyguyW/5mh3QXEK9Tl1swgtF3El0D9GiM8JL6i7eqmJdaDUAq406U3gYLIz3wfO
/m0O7Vd5hN7yBST0wQRVhjoDYKaZ3mKKq32PTLJ4Z82XBJKDHFkqWydlgcB1n2ZG
mRzK3QhGZy7CukOnPzLfp9tgIXeki9UOZWV5atMuoSsdhFEY9ZPP970ZtlvD5k0j
9dpoi0Lq/K0r8pppc0W4s3FimM2djd0FLc8vE+OVdOgsu+VEC5zWKisbL21Pa7y1
0XMAT84/rw31PTMf1VmPm8+iiC6BWvjxVJBB6O9la8AqRHjPThsyQ0YCRiZhE4ce
QhqkaG658mUx3lKmn3U3qJiFsZzaZaaiEJ4W8RY4NTsgdC57L7pokVtFWYoBYdIp
RvWm08ap/Vse94Y0D2JlBpNSivAudc1FSGaE7CITYntPWUslswUtzdPVk9OE/vHf
ZV5AzMr0gl7tRbumsMR9KUhcNomraGRZmcWT3iiarSuBP6yS0woqjjQXg0p58S4R
P4bTBY0Pn1sumsE0L7cl61k3aD0iJaI5paO1082XhozZIhBPdEi7MV4m/cwYNtKl
uECGdAmy2KM8/wxNUN548Qt7ciQod6LTSV4EulD/zYxWVXZbxdKe0nWT3mulszCH
KElPgDxFCs42rmKKiqFJE+bgVIT3/JALZv3vbD1wsjmSa58lI7/ied9k/L9kBhMI
Qhj8ko+mXU3G0uUD7JiZeIAJgnoOMh83jZgRsOla/1LZmUdpZqw2m15/e6lRt6+K
zfljI8Q5Km9Tn09T3sAtdMDGAv7k74lofFF7FHOd8pBt+DHmGptM/9n8Igxov5zG
6EmyIHoWeicPkZEXvIv/PssIcvn2paCjvJIWybGqu+USPgrJltze7yZFjncpzDKP
Xolgf29cgTtBLfVsvvE3fYitCzib1oeaWmNgzwg4gTYvRWg6gkxOl4/A3E2268sI
VZcsoshbVrkwdVLMcHFgr4U7aIhI2U/axz6ZBkQN5gCjV5A6S0vujk5sPGAqwndo
G32+P4SHMsCu3kYWDP0pFXqbuL7BMSV+YuYpFoqKtW+6PeuNursblj8oG/eMeBaJ
0qm/eM3s4zsoc3iEWY3O1RqueLcA5yxk6sXB4dTabe+8U+FDt1nFB00/y7PjL/6O
Km7QDcDF/UgJF+WFHtflr7ndo7Sg/UGy+HbCGpRi7k3U3lmnOMrnN5HyVMQR109A
/Ll5ChgWRotzmXad9eR/0XYboZ6kmGrVUMKUpRtlYZNHy/a32oDrT2DfKVslPqt5
p4UO5AHGhaGka7R6CEv+8STzk6PdpwtWWKPp9aZqebFYAvnb+6MS2WKxK/4y8BfJ
nBHyEHrSRVAgVVIWJlIJrrWWLg0ibW3OaySMMj9Ka7rkg3ESvzk5gEdeWxVAIyd6
jZuqd1/t9X8XFIbNry1zyL14sFcuVot0xnRB1vCbvJuWlZjyjltdSFS8OmzOsqfo
drMbTJTPW8QE0OMuBPHqjDrRLxd3mESaKicjnuhciYZMmmVALkfGkmm93MWekM/Z
+Tj1JopPu4oWP1YvQmX33u64CronDbSGHJhgWgz089JIrggfKaSY3OaMXKKKcXin
0AaNMyCTYpZfOIBqIlGxWAxb2+khiroSvGuEqoLbQzMfl0plkOl7zMoruLfCAv65
+7DVS7YkZc1WEUmzvGhg//XEsmyOmLQh7f/bUyrfGUpcOgjc769dZGk+IdCSg6BG
8XDkhMk//WwbducdoNwFx+iV1QQVF4UXuQgaH1L3tPfe+Cz4ytObAX08EHmjCWv2
uUKJCQSM4JRJU4I6445yicUKOutAJJWdgw707bIT3H9s4LbqIPxMYLF1fXrLaqYE
hm8XFttQqUJWQJ59I+ipRK6VjtV5YgIIoPpK0JOnQhpBewNcqTiMJ4aB5tsDxzkC
jS3mAj0JjVVprNT+2aPj4BWl46gux/tIjOWHJMAK5SfVlyldqoRA2qYLcv8APKxn
UX4juFqZ8ZnoRnASxe5Ouj6975KawurSk5bm4bKLoCuTVNFQKLJeeHll8bjzCmFZ
w/kOqwBzhhK3oX70KCkKav08xZU69dvwg0kLnl/t5y7fuHQrVbbBecAGEQ2KkWM5
R9+GwFWhmjgasOEJOvTbeK63mZZYynL3I36pUNXlwCgE7uiPdUMOj8vezNKNCzq2
PTRPd6FsYb0IFmzbi1Ap6yFTeE/OEebF2WExZoSwyzSMgV8DeIxLIThFcEpkWJwM
QjTJrQSPPtki1168UJLUZOcCUhTowJBPX57eQyKgl3LgJe//KJPZvL5R2hwf0+9Z
yed9TgaXw76mO6RTfd1FDuBfTO/njyo9LVd8IqAJTbv9RPX/YIpTBJ/Cj/iagkn9
HRZeZlxq5RgVGEkpoQ5XkhfzXD2WB1/5hKqxx84xoOgT7bUTMDpD/P48Cw/B56VD
jeVUqcl1IpnRW5HGtZJg3ecITTU8vzIohc9CwhsDM1MqwVPVchR3pOZCl9TRI24H
Ss2IOwRWwJNl5MYGxds7kqhEZPUiff+sMUQLLxjrF6ojiSk2Cbga+9TpYHJYO+9G
PymkCrZCIDMBodIboxwhb33E8wnEETWZ8jGc2lAhigzu9TvBwoilBcrFau4b5oSo
AmupLqVVs8qIbo6IbZouGRpSg0oyzexQuEcV9dBkn56YEfgIHG3gDc0JTpCLbJF8
S5lmG4Nwsc0Gdo71E3PpXoKNMycaFy1A6jYqMzzyEQkSpj0rBXKN8iqiQnelEL5B
ssiKWetRsnLYJarn3x1wEKRvP9H837WFeWY6pUi42wR/pJSE6f/sNbenLgso7RYe
IotwCU+2HlRSH0TiKmVG3UdtIOuuYin8/5eqdAsmRGVqQdGJ7/bWdP8F6TAFsFaJ
yh6aq0IxLRj0DDrTKGMCEXwwPofAUwIxsmjy2MK0m4nuTQ4oys2lOU0fWrW8o0ug
bbZ3Z/ZQsXc7x7cPUIutef0l/u0vyjW/ZTHoR/978qZeiSJITK/ECyy4KBYHbY8J
AmCbp1N9HDrBi9VJcziDK0ZCVoUzkBNbEvO23l1YjiuBaaL5vtw2Gp0uBhUOhV0O
dewWcBM42gcB6HDGrDKLfPgFniif31lFoC+AKXEoLWmS3FzZp1FR0YS55KsnONNJ
2y00aAOOYvSzTG8kN8mC5/H88hhDtUEwCEMiNpzOwrOOcjVxfpqO077T/+M8jgUp
f5tUMd3hK1DPYyQHvjFe2vtuU7InLVEUWd4oHdxFuatSeuGo2NtC2C94fpmMLguu
gN+71OYZH7yYvFI9/t92w/VxEhHipdR+5RoqB1OmoRIEitoVoXuIg14W2/d0yX4v
Y5pnK9ifcvXS08YNmtP2G5Zu6LmxjoxMmTjGiHP48h8Scu5+ldnWhVvMBQZcIkhD
JKkz1UNcoepWVIZ/gZ/EyU33iQt4c4VXKQCD9k97NcAsvtJl2Mv4Cab9ff/vBnDx
Jnrj39lOapvRX5vihZau1BuNAueA1qx0gw2Ewh7TN4CvDv/pyOEXyPVbpFMPksvT
WFTamk/ketD1PezPOc2Dyy23ZfbV1PtUTZkckWljgiQ6957kl5uqOAnk4hXUDI7o
pfggtVyXgLI81LKNMGjWWOOFbxsewNuufc3GsyxZwSn+Uuv3Eybm4lTtlV17QrY3
zTBfiKc/tyObv6aEPJs7eJPRRc/Q5O77p3Yt4KMmCy6ozNiIKS0ZqUmj8gGdspAo
pC1f/tBXliysGYPBNbJ6WjcAbW+shVEjBDpmYGiMxUuuGPSvUh/wbeEfPXL7YdiH
RZ/GE1Tz/3hmD2ORVZ87WOiVYN3z8zGIfYItuVEaspnXzgRt1EsJpJx+LWNw14Yi
C3Ra+nO2RHmV/xTg/vjiB7aE3cgbSlzIJ0DuuzL+Z1t+Mvn45v2bochQMfEZNLNH
kUrhDjTSJ7AeG9NNhr0pDHTG7xxCmeDhlWT/pm7/OgyTjV9G8tcswWrPnyjzqCJx
6xncbrmbd797oV92r86ItqWe1X3s3HtPSAa/BPGWpTaIRORr9u3ahx++xKKshn9f
FW3rCfprTH+aFnJRWA0z6Aq/Q20UXSNDPUyLNUViZCzmATgh1FjQRwvCFgi8XQTg
2g0iKEqSMVquMh8dC3LkfkhvGOBY8ft9p30ottX1f7qMOCi2J2p1EYFIZaiGNf9R
cu5pEGeiXoq6y8wjGlv8QoqLTiM0Ja3vcMLsvTIgFvpgrHm4hSwWg12llBpotC2i
SeP3ThzjFKCD+Z21cVNMi05tcdP38kDeKKCxp12CmTHK2oMMtMaqlfnuvSetLEqM
GRYeAe8/8wx3s4TW6Cr+H5i/cmk8vJWBuOagShFpAf/Qs/j71mqFtq7GgC2uMU6n
wIzK+vw1atzxZX67h41e93NuLZ1u65qvrTWQ3IQLDfgA4rhqbJwFs7XEjEpjxjfb
m0IjwcZe7PnREOvteAIR30njnJNVQtFCzqibW+cE5QUO/iUdXjTp7H36ot+FL0eS
eU18/3vVuacKP42P3oUVdJmtgpnbYrIDtoqF9p5WAbssaE10yLldwRdCWQ4ZXCHs
ZQaehsPtRLBUJFZvCvneXHC1dTM4MJoYHDsfbbaZOiBrXawYaCEaPwTIBNz/kg66
lzSGR8V6EBhqDq+Sz9zw1XH+2dobmGXVkiAEVXfHZtGr2YmX9U2QgKxKvg/bZUeS
WS1n4A5iSe3YPLrmyI0Njs86pPEe3D0vQ9PLKUif8ZeAEWJN/ZRcxgrHPmwtV6xZ
9jtCHZoTcFmP/PhznJ0vdx393X4n5J6fMvDnylU7OV+bbxQu6JvgxdyfC6rLwvv7
HzWzGuKA+mukstKUchaDysoUz/tr4h8cPdIJ3bHD36HdWOUtg5zrB6rC6J2QumTq
W9SV8UpgGzbbo7iVBgXaq8K6ZApKAuWT3CwwtxpIg2mE1RinY9ELHjwX5kKGrjWF
FgOu+QIq5ZVs6moGHPmuObfjOe/YTvDaFsKj7Bc4rJBgJ2rxkhD+0Oan2DhCXL+c
Yzz/saITqtKac2fT5Z9zm5dIathdIhUYgg4UVd2Ii8EzhwzC15kpcwtqnjUu7FOW
T/QZeF0iaSdvib7ZUfic9iNcbcUs8L+NHi8eF60mXmq3FKdbobGm9nS5kxhlsRJ2
CGeUMkgU6Ifes7/X/6Lw3aQ4f8WuRdSq3WeJkK4RXwL7heAqe+y2wZYb3PfnxaCA
WKGRfl+8uPsqfTtZbs8rREThPkJ1YDjx6RRUo2rph1WYhhwB8VyLVqK4U+ufyACe
x3lMzUZXtNDKG18rUv4tR2i5blNl5Ju0zZjg/z6IpNEo1OkEF6T62UlUSqLrcOic
/U6uQqof3ueSezI4DeIoAHTIlm7KpMp6HXFiPpzAu4FxvdHNQCXQDWEAErjFcOM3
QhXTju6ycZIcj1qw0+kFHVlS5QdjP2sfyq2SB/sYFidtkB5TkQvL1h2q0twX55sE
EDP8t4YAV87Rkbp9OZDCPNbKIiIrVbYfYwCLakrSRcj53LqW2Lltj6/NUEzxtwJ8
ekRXXOuvzErFFL4qMTYoflznfao1WbWE1EwvTZlE8VmQuP7FsTUDhqfG0wNQdYAC
RVJv0mn2Pp9UpvvUdoWSA1PfSdhvRgqE1iokRhAAvkOXa0jd4W8UJuzZW9TCAcNv
VHkIy3pPkCGitquTUFkX5/iIrtYy61svDtlCUx4teoekLJQLz1lfNx+fBHJ8vAVw
990ymB1pVbaDFu8YLAsyLd/gF7BM2yMrmEa8dUWUda2eWGU5mj3zmnrWbUT2GJMa
wo61sYk29hvjRz6SM4GCRfraqe1KeCpr1xKjwdm2tmcZtDYdbuxZdU25LNmIuBLT
lXp0A/T4BNkBlAWjAXwrRnbmYEtFycqlRZRRg/Fh2lhsoPLi/dnjU0gK4DjINMIv
y1K4Hh+HgH47fQKRCNCnjxWZuzSdKu/+i42NO+JUNPWV6dnGT3YAf/uV4KM/pe+h
spVPb0eUhlx72vfpF/4q2UCPzLi/+UzllqmRZyrUiCrQKfkRhaPB3QFztckgcuWZ
QV5lLC3pynhQXpEEJ0mmBFCvr2Pic/yDVhe4iC8Mr7YeLQIUh8ogx9Wy9ycAzM7L
eLbmDekX+QrygCgcW3599blZrOCrZyn6ciU1F09ZyMrHwKw36zqFN0TANBr+VFwf
hX+5SCt6elIQHr8S217B5Fzmz+kw7seMnJ5Xn/GXqJ2ezpRWdomoAwHfljefsehv
m5vtDed7DbxEFe7EPE41d+mFWYLZLgYF9h2ofAUPg9lVWay48/vbRduZN1IkiwQh
lwSwcNOQuYXLb+TvAYyqs4qa3UFJf2/nfjWh/isRgGHhWb/hapuAf5M2jxxm/RtX
yO9xBrQsL6k8YGPLl+tk1wEtO0i2m5g4ZpvcEHexUKJhyR13G9keVLeD8lsvFIIx
SLpDdEcNtHyrxSNzWtQi/cR1Itae7mIM4tRDJRSx88E1361ClA4/svhOOiyrxOsL
BYKlLY1zNKUuu1nEwOhr2yC1Qi+OL7fWQxszgMantt6C1ty5qGIwuXDW7OP1abnW
P2TD6zg3JliVBS+kmX6ysw21i/Q+QE0qmEsyz2Eh8+dmNYQVofSZPJiAlPXU2828
eO/TcjPS3Ofh5p659f9i/Oa9efbVfd+eRoQziC0YOz/oC6xQuwNht6jwCb2FWYso
E9/n8nX7AuMN8eZpXLREzdvKa1wiHs97tm0u3jLPC/ON3gLFXKqSwwhqpqgc+vfT
WGqiq0nyO8FH59lqNrFnwBYxssdfX/8YJ//KB+X0k8ZOo3EcKh9EPqWVGIkGoFOV
tZCxhS+O3v+DWgy0bQe2X68Yu9MLQ+ia8FzNBNQNYBBuZh6cx6GWrUghxaoD3Egr
45xRHIGMqCqpToc3WWK6+GNOZhkFVF6nA0smmTgoktmpy/I+BDuTxGwA8pcY6ztW
efh5mbKbt5KA8W+iQF7ifIxvWlfQsZGU3z1EncKNfmCXcNKP+4XwVNPpxyiTlOYW
sYvawvUphxo3Z0yNLK2ugHWKZvUpFmA3CkA3UdsracDzg1Lmi2R3epDl8yvqEq6V
D2I7K46dFKF21fxqO+HTK/VFGWZy7XzFpStpC1Q4Fhjy+0Z7Uil/OTyiRlfl8SX9
/8IlvWcaAJrN6kF8hYaJcNgUS49nfHJP0sftZ69gB8BY7/Akk1cHkemdyUWPmGFl
0sOjq3vJhOiugGAov0EjcaE1Yg9KbESZ39Y9DjoLc5H1MdwGL2fqztitVxe77/Pm
bETjyIafDxNd1XJrYwJGgpy7puywozLh0+Frt2tRvDtZzquFUJfWMFQArkGmAxm1
2Kfvzp2slerXfBvFiouNPi8tFKqFRvGtUIBSiZnj2p3wgRFPJffOq3FDxaRArjEM
KjTWZXH2cJzTnRQzHe7tAKtWVXwXcoYhAZJAjpc5Tzj6RaDuaIqlun+ahMYhQ0Eg
SVOqArI9Kw5gFSeRHVKk8UKCac8fli1y1Dax2s5h6GFuThWtIBILuA01kDwjWxIg
5fVWW/JWWJ1wjMzkxKV08pBI8Y/JUX3NjU07oqCzpeBJBf9hrjSRpJsQjR4kfIfG
Iaqrk0dU4uxBZxRtCyvIgAFMCpFTS4N7h13WBrvAmHCbcNDYjbzhSK2ZEs/8vSH7
B0hhN5gYg5SCwJ4xqXIBHXAsoQTsgZWjHhjg6H9X1Tn+pArpga0BJXj+ZE7bx6iu
GlJwE6O/DcD/qk9BZbchkeYC5WtThvJgzHGN3FHjzLZmt876J+peyPuv2M0E3A6u
XazHSK+kE0ufDDhp9Pnd34qanHsYr6F87XIHvH2+MUVXdbp0FTzZmrh+jh0uFA+R
gvJhzVyjp3Vb3UptcH1nWNUiYyq2RlzvG/USgh2HzvyqlFwAA152BWzv95l4ePSE
DxVRdgq++xBlUdce34W1YQ5MulRiiPaAl4WmRaRy1FLjFo2tRQ6AkhXHzSe34u97
vJtwgswsoPMCqXDodR6VoODs3DOQfkbI23EdH52rA6eylkVPZQ2lJEVTZrJfHOz/
QBn7GofRSRFrzl+XJcWpGkl+ztP+uo1CIaYR40Zv6CdBhinP+q+TCw+9vLVOyHQ7
AVznRdDo/zPHHy6o8OyL8zoGMrD9B86cpv/Asf+LiLAVu31tSTcC9y49dwilObzA
mjcmlAJsqAgnU/PSeaWjYn+cbW0cZE9/35K2GAaYchbwqGFAKkTV229X4nEi3B9g
a+zJlbkyqPaKhL+ydGme6/bu/W7o1AJBj9btryaMrazhQLMMMkG09c6nSu8OPfgL
brBD4M9YqZeam0odxe83OQ4rTCnXM1nTCK+gfhds5YZjBvPKfA1N80Qfoy7q8gbL
FcQ55SCMYcgHmlgALbaNv9/73vPiAfCTuIfH/r/+YqLKAP0DvJCy04/miP2MGYEH
4ih3NSfDXUroLNW24jPhfe0creAXlbDoPBrdSz6WLJZpUvOIsK/y35siGkWGx51L
JsyrGZQNn/NMBEvbQnA4Py6LsKohFQkNbjRIUlDGlJ9c6KXIbwnCkW8TkTIzKh0F
J6u2GdWIO4pYBWXzRh0fkHam4Bs1aysnjowjhfOkvCAOFOqnMZ22eDOdaqXkIXtD
MnjXK67ZErr7HtGQ6553kFKC7J7jw/M5MXDQeIPK1P+Rxl6Bjpw1Asj9rdAb8Khy
PtbN9FLx5JEbY66R7kdECf4NGwdsTjT0uaQE8jbEYUwIHsY5FTKj4ekq4tKCPneb
Axos2hwjZ2jl2OuSu7YRIdM3X9llb/V6ZnBoo76N0Yp+T3Zm2TMMOLCnrPGMT5iS
EHND+edCwPxaYjSq7UiFBX0lh/0bVqZQQARQljwr9qSG8dCIpceLbglfSCo/KOod
eOGR2VaixS0VUo+7zda0tK8nxkf4vbkKabOTn09de0CM4hrdzyk71tuw3+yu6sMq
4cFKD6dc2hYjpjhoyR1pMo2FygM++0Kryv94pyRI1gyw6pSspp6HK0Ssr+KenO5g
9X8lwQmI28su2m1VLfT2lPVnYh+Y4eNV9nSPxEHma4s+ZZ5sp0KRuGAz4UxtIwoW
D3yNBPNT420TDETCZet1qsbZbi7+LpV+szQY0rdd1kv8IHjyUMmhCVeKXg7ayJGN
QQRReCyF0H18RSEAJzzFvUMBA5p+KrFj5cyQI/kiZerLFjpN+fbED2/quNRaqEUo
/LdI0kYtGWKIK1JuUpqg8rEd/6cVff+WoNw5upd3qrk4r/R/4jxDSU0HaOTYlnMM
R7Yo2YLvPqXkvCvmERotVX+jxeARbZa0l2KCoo29sQ8VL9Ost9zE9Euqw6yDUVmq
jHkxWrMqGwVRv+3C+5z5HOzRkAvTBw29WyTL01CPwTLwB+ncJQfJBLms7SPqCPvG
obhyuL829F+3bFzX0JNQfIcWl41RXZi4Dhm1skYlEvMU0tCw2FGqh/adMBRmtP+p
HfkFx7icQC/4AAy4CjBjNfNioLThqZD7vCceF5Y9RN3b43ayIgcnm6zc6VtRkN0J
pSvu6OvLIeiL3/gLpfbOOoZwV0O1j3MnQ7JVY8ZGatbVftFb0dgd77VSork42oyE
7LRgaxonwnwQBSWnpBKZ34EK7O3/z+R4NcDsx88L+4AvECqA7vc9d/iOjFgoZPtL
45+d0LI+UzUo2QxXs7CjLJNF+YIOOojhTP216rMDbQW+ILesOWU4KwpPXtrESJR/
Qbm1Sr2OYKE1/lO6L+mBe2MrM0UjV5jshlwMXtSIUddapxe9aE7UFNk7pZAXe6Jc
L07EP0r6YElLUTVk+Jh3uO26vYRDkFtMl1JSdTt1W8wjJNuqRUdTts76Vp1vI4gC
zr/AOHihs85tW509tDvFWhqc2pZ/zLnHhi7R+StVD6/Zt5WiUdSrMQuVE2rurX0w
TpFVp5kb3rSJ+ZOJfiT9ebMzC3lthhua1cFqwtPgKN7ovPGfDgYhbBFF/7sKC//1
QTHCrvSaLu690cj7VLfa3SPlqIMq1y/Jm+WiI4NEXNpkMAU7y1OvGIFFShvQ+sAZ
Ard5GL112WWZu2VHg/c7pBhdEqsal9GNdRNsXC3wcWeI56AJcacP3Ur1tmrCj8TI
phg/iu4wCTsSm8WGPERK7ByVOp+w+me2tt8G0+iZd9bt3pJ9ZqZlt2oXPK7kbX7L
yDnn5CN2GFwDfB+UC/EPqLt164T3aIKiFV9ihyOcdxw+UFz6mvImi9bt9piK19Gw
pgHGebGqEx+GoVy7lkWnMhiT/JziLHc6spiBxW/2JKeyXunHTTBN2zWmkoNXMbCZ
oBvQTXP+3Y7lDMq5tcSiXLSGXDcJBmxhyknjujJKkk8Swwar3a9LAM+riLeM6NW+
Xhe0MiVu4l2P0xh5OHVccNo4dBIX/lfdkJgqy5MWhAZN4Xo7CAfrLOfZEgzVOmOX
1bmtXAkgGA7ikBRyIvjHLyTX9hN/FAKmyW30MNhHTKNitFq6UgYI7/eT338KJt07
eBr41+Ljv450gbHq9cqxHeYmK4oJhOTy1G6pXCOi4QBcJkzzVGhEQAJA7n4/lEHh
ZXu2V0huWv6PlYNA2btN4MRe16WT8EK8OLaNdlg9jOjxlyrfeD+uMpK3C5YPjZMo
JaaTz+oZv3H3zvyXQBs4+QhvrOM7zhWnY6PudVPpNjraNCJ6pfwGwTXROZ0CBOQP
ZVsO4s4XfjlDhtlXZoiETe763tG4AlrMC5YGismKwhPnoa2SEcUOwwyghL4ThgX1
GX3UWtzw5kqGJSklTSQR5Cve9ZltJZeTq186sRyq+bjHZ9mAPqwgUXxHBY6qN4FJ
OEh20Y04j6pqdzkgAaJuWA9x6fDzyWsH8BWm2i7i13UY+IpWbwnwlHrvlT6ehHCS
iZWA9Zx0xhEbQZ7vF2FZjpOu+TmKAJf/aHxK/J43bLc6nJbWLcKR6XMQNdQdiVr+
FTqCM4ruLBgn3j/ZOMu5lCEnGBR4LVpBmK+HBoupZ5IdQ9CCsqTWkxkytJGuUE6m
RVHmxuYvl8mlnG29vWMS2bz5jxbgK8bR5acKohJQI/JOfisKUjpF3bNnqCSGLX+0
eXKCfljXrKo8t32a0V8b/v6C9Yc1iv6Wd+giHU6IopG9ModjeoH8+rjeveIoIAXw
vVqLveoQbgMAAhiEsMyhB9+l/j5FF+OZR8ktX4FpaR4t3fy2/b6yXOAb/SdNiYEn
/F0Yyr0TflVZ5H/jKXiWVvpM4aDNzdENuUyWVVYtfSlxgcdx//pB62+WZ1F9wqa4
zt+KbcYLYn6ksCZ3zmrQq9UdRyCXSPZdSjsyhfU1Ed8kTPzLKHeOZ/eTq+VuoeR7
u9iJ93ZArfLy9hjwNakjY0rQ2x9hPTqM+dGeeF6I8IJvG/FXsdYIr/CPkhvsMIzi
mNUy4V1rB+yHuEd/SIf1F+SxVFMdJ+Coy86/xBeA3aIcJ5NRLZe32DNgFRIFplT+
MyAhEIu7PE7FqVLR7sYzZvhErncQYyXk4o32GIF+0JKZI5WiRxivn1KeliYKdVgS
cD1KfxKLsPkzXPo+Dmje1SjRqRX2r9RlWXJaCN2ZA9CzbQRo9+0BShsUqAehAITK
e3Tw+5yraQFT22mSg8R6TL6qKDWOTARHBD0G5EBO2ewAiwr7nSfSY0GzKGISxpI4
vdnHENyj1FLsPMVoCCMWrJwsLrFbSV4PS+Vfq0mfJAoKEB/gDllf2LwSBt3rDx22
ALLVNp3q5TL6ZEu7hyMhWBNi+UlbIUMMZOYvVUFfH/4OPd+Cpxu3cx8FgHChEgIw
q6jFb8Reh6QCF4v5uImwz8oHmnHxpn6RGUP9+u4TkjuRB8fBxaF0DUdrkQD/hqfS
XQgLAuobdkbOO3UkvN/7YKl2pJp9ccdL1sC6IdpJ54KQ71SA5eQIac5ppHElc40A
9CL/al42nqVzUftddW8LLeF4yF5BjUtWAbgFz3ACrwqCfp0gdMOTcewhis5IOdkP
1C74wScT0oINXtHhUYi+5O6OmAMvGHKNdTEMLbmEO41klEWHKgpoAZcXu3J0d1xL
Bdyj/UTf5X0tgAzqBm/Eoubk0qrHmiNGv/82aKCs0+e4eqz0zP53dfpg193ClPWP
HiVZ13Sc+6s4vFxELtuOGDYvFqu7XQG4J7dMo5ZV71XThMtqxdqd5cC0Hn3U7W3H
4GGPIj9LCFG1t0Xlm1lpZlSoS7TYy+v9gdvGnlq8GDQ/KYnDfKcB1KHChqv5t/DV
r45ZJ4znieXuHT1+axb7V/HVH6hTUayPWZpYg420vWlh2jjD/RHVdGW4gYnYCwCm
oUdQrPVFU4mxXI8gDFjmS9/pqahjPPtsmkvvokMMMLYx+kJdbqyJrogegLIh2y71
m5a4CDXd39HhQ7mrM6Ra3SHh8yJO/Y5/veL9QUEZYO1zJRxoviBHMqdIKMZk0vJR
jEejI4KuslQoKT/HO9vk8nnnvYLFXXCv/D3SRKHdh38cE9iRBr06z4oM3s4B2Qqo
tf8gGQBskpGnZIy9xJaXfb6plSkQPnbo0aDutdJXV86Kt053PxA9M382r2Fsxu26
h4NOPpS+4HHNVMdK59Wa2YMG9aX/sIaiOFzFRLo1v+etoZ0RKAHpAaQO2pMGmQp1
TG7GPZSX3Fjxo/e8FSgHGoJehnL3VUr6WCChVjaOGL1/v+Wqwb6fNOm0XnOdpYGT
IzW08M0NGgf9/UmVLjgoMegcVdVr1sEbnamq4XTf0QEypTa1lbq8SH2zy84UsONW
IkGiHwVKAtNydjObLzPaJS3CoTnrloSfaw/x2XrtjXHDN7/GS3CFA5azHbiKTOAV
C6KAS1CIIYXPV947OUkrOmOYNYh1ZVUGssolKomww4vGdXP39lSc5zbB7LUtQMR1
mt6jOOaF6yA+YbswmCJ9rVvIu1MJMAwvzYh1Gc4SUYKxxeR+bMGbnJO9eV/mFSeb
KFhOjIMF1ime0+fjdvXaIyG9P5+y77t2OQPBgENd5RQG4DAnZvjvvJ1C3fMPfvVH
LmYpc05grK9PXoyHpKrBbBHkD/XOcor3gNe/QsDejK64suxMuf4OcksSALVEPNap
xiwvccD66LgcpSY3oDfG/wDWe2wVkYMq34vr9GOpG/c3z4BN/R2a6mC07z28cGE3
dcQI3uzYEDfie5JtEt/bfKaP7ESZslEj8A2+mCVndjdSxFs+UXNO0nyUXzix730x
3PjTIdTSyl1VVtR/5q2GXha4vbbuAFnldD18xzkFLlsC+vKJsaWwaAZiYVajFb+f
0scYU7a+RXYXqCaP/nAkwtF+fDZRJlKJXfcxC9LDdDMS9hoqI1SCIGRwKG/b3ucE
/adzPgzXEGm/qWuBvU1FYCoB9u70Kjn8Ee/GxfTCx3yXzaYAWXzH/SKjgFDIrQBN
POG4b3jTrtwUL7NEKzpaYjyYFeZfWAlOijK1C866DKdHb5rdixjsNfBQ7C3OmDFR
sxbmV+xVvPk0rDZBpR0/PyQXIX51rfMEsfhGt7+vUqEjWnzQNi0ka3LcKxvpXUBJ
pl6dnkXbet9D9xc3xTVLA81VPomQzUB8JxzzqYg3tY/VrOkWj8g8lT4thiX5fW6e
b9Ekm6LP3OvfUQT6w7JuhXEnhoi5CAtcKIGpShNZLodZxzTQaXB9o2Wwwx3gjjhA
4AO5izcUnVQvjCZf0zSe3cdxuSuxoDhAB1QRRVn/X7POEVcVLsoJ60cZBXsovzYi
XIvrzGJnJnhZ7E91RqmjdR0cclZ2sG8Er5l32LYJGTuMuYGQ0WvS1iBEUhge0sG3
85d+ikiv5cZDGO14K3A1bRr9RAPFAmLT+wVdqCRt9Sad1wkmOzZqhIjjHK+61UC5
u+oPZFUI0nejoK5IYYSM1DN4FpWs/2xqsoQj2A2OdppM56VBQ2P7ACDaJhgZtAFN
RT2GwwiulQ2+7AHrC486ff0SWAiexpnaHmn2h9xenImy9bH3X3eRW5hiyBPcJO6p
RRX/JSx+FLWYV1uh2/6ySAL/wSpwyiAubJfSG1Q7gmMDVusU9XZ7vBIbosBMoSv8
ismlPPA1iIB3lqcuaqOGsSALfI7h1/NctpOd6emSZlOvHe+d39EoSJowLdzFLpHA
wggo55YDfDhylwMROmDqkaRpQDelDn7gW5B5Muq7PAxs47FmbtY2ZSS6rU1Tl5Kj
5R4R36DdrVTXDq/vDSl+ymF9e5EHoZZtOniyvf6IVJT10NMZnb7CHHHttgS/+rmp
QlugFrE+kMXXlDvdmx32rJ3R3VWViR3iblyWasdqvRn598MRcQe/hVQEDqy8cTlM
cMt8lMaYoMEmda15W8JmZhduCof8FcuzQ2LKkcJopuyMwzAqzQw3R6d8bEGPjF4o
B9SmHJA/8uBIawTOSdOYgPUAMoL6Fd823IJU1veChhfpyy1G4c3127nBxF5558AM
+N8OZx+JH91yOQcsdUSpQv55YXJZv/TyDioAUOi6nKWeJ8Be8+9I2nu/s8m60ZTb
ZNURiK/KaIte7A+wfZxKm0yml7DoNHND3jmyBGMJXKMOCsvb1bthsnngCrVoTSWO
w58JX6wCbABvrWBBNA/x1lP6IbslByADLuhHpmxxWhsuLW9lZE0pDkOLXo0MTIuF
TjhU95SziDk/8/ERY//CcYdNRBJwi0BKkZ8JGAo1GcaPh8QDujVIaZcd5rrwkM3+
nAERDnVww77C+UwKYfSvBxEkr+eDA1PBqyDMTMLkqBJ+xZc6Dh4exL41H1u5INNI
UJ8Q/bawMWyWUN//ah4/hXDFZ5phx/9vm+TFA7ErLpmwVEls6HIU3CDtLbk+5pmJ
7YaSV+Zr60/rRqOnuDaevXSS1+6dR5ygLxPNdGH72gtybfrKs9B1cB67YXhhAnZY
5nB4ShYMYXF/IPchHjHKTAAm5x+XQysQvOA2dKXW3lGiHO1iGS2wP6mZQ7/ViEdG
RBPnbQfRwIl/mLEAGfQ+n4g1Eg0SgEO1iGb3WCQKcSxA+UMEHB8iGBwTsC/jHrXd
ZQ3Kx4KZL0aifZNvRpIuhoAoUXj8HIyBYOwYXsd5hKLabBoDFvo8xZgiXXEJ5Oli
rOntvi3YDJJ+64l0gcX32Hwp6iLgxqxnLrhUQGNYqE8Emh5M0qe2LznpFnD0DHuM
qNCStz2dA/ShsVDbUkaWsKku83OMDOuxiWCWo+gMoASPiwYLJcFksSMNZDr+H2aI
E8ZON1IEHdkqdZnaqb/ElCZ5xU6iG8ApZJGzOBeS00aEzmm5nlpSS8cWn2VWwAkZ
`protect end_protected