`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
ddtXksX2+yylW5zu6QL2Lhnb2d1sD00763mmSITNX595NcHTEkwn0zB1Dry37fOW
FufOhVzEJp80NC5qZ/+F0Vk7Ik02dIR0elf3clrjeJRK85K4e3Hoo4xn7YbFUIms
l/8VZSb14+JVGURjfswrIyCUotIzlzVYZ6gzoZwDXIi5gQIBf/gI+KxNXPaKV+PQ
Ufys/12rjO6aI/pPlqSm0hCvftmBcnezN2hk1UeXgOIuKZnogjOsf0iJVX2aOOWE
6pD/psybjbnsNB6kH5uFTA5frkzIzkzl5d9+YDm9OyC+k84E83I/7/j+rk4L2dah
QJOvksSIzN867/4Qt8qYTQ==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="MvBXkzurAa5VTw+1JJ70nePUfoQXBvZOku/SMmg4TwQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
oRtzZL4VJ4iwysPsC8SXYCzXS8Fw2gtZTOskLcDV+1B9Nzn1zTyNtlo6lNICRmmK
ZRVu2BmCc2G+fmzynYlNTnSa7C0Cuel6FYpxCBlOuk3OF2tzAmLAuDyOH3Z1Yjzk
a0aHuoCdIRKv7BrZCdALt03JeUmXKPdOmIlkVGFl8yw=
`protect rights_digest_method = "sha256"
`protect end_toolblock="Jn9CQpRhJt4rnzZPRk+dOpzAubz7omckX1MrFd4p81o="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 19424 )
`protect data_block
gD6l00tciPUa6pDNTk/+t0OO0nC/UTtBwLB41d4inuAUA3i/ALrNyoJVcBnAmEQW
ptbcNp5fxEUJjnOxnedyZEuEBxWRieZFQnkRdF269oNL9/WPHcjtoK6frc7P/CUm
1RBDKJ2acuXLw70H/JPR+WQ7DEGwMl7vQvWwo6rRcfl2fAVJ/CLw8lOgsQSA8g/o
GCXe1ktGrcO31wC9M2dYoT5FLx1x4S2UZT0GLTovleXqQbiYq6oyd1ShKiBNEe4X
XAys0mKOjWMptaZnQA0BIKsEKQgdA8tkYqqiMWynRrPKwhDvukdw9BomccQGdBjK
RvI+EYWbH3vDncxU40zf7HG62Q8CohERQvIwFcw0vO6VB9PS78fWt2lHjlVR4TmJ
HOlxLyhxaaPmA1RT0BDcpcnRli6cGli6Ua6mzDERsR14gI5TUaSnZQxsTkpmiHr9
8vVo5PWlJxM73QyDAyA75rJxVwCQSxSPZ45mXZQ92VlKQZ9VfdBcqyhveVn8OrQY
QCvya8uHiMmdQneby3jwDJTyTzJSAgblsFxrY5AfeTDVqQlK3Mv+bD24mP11KTCX
0jJ0dxScf/iP0h2278Q4lumst7Taq9KJB51wbGRQUKmpCs+S+ZDhvdLIMnZhpNAh
emSuSY3gsNRSDqjFN3ahzWlTNJCjhlO0XsWuMKzD08/4ojtK5hW5pgpfph4gD/ib
L5h0pkXc4Q3CD96hi49Nu/qKIO/EVJoHOOU6bdVBHrPZoI0Crle4eTmHyZVey7t7
wTaP2vdCFkEzLzJQ3P+BWO5TVMTJzYhy9I8wrD4Gp9P3G7YhKduk9cJZW5FlK/sQ
DE3fztO80plWul+Y/zw7wGnOLSodFCWCkaC9lmZ2mRLeJNoMYlpqqAP1CrqolLZW
fVvxWMeTnUJrPxksdUSM8+n0EFhIbgCJlIQW8iy2A18io2WsWRlZBZbplak+tKix
yir2trJs0ksvlqR6BbfaeEnq2FXaaiVLbXxiNDuEygdU4uKBwD3ikcy4jrLNPrAL
7gCJ+fbkcfmVA4DwT3zkx0if4nB86z8gmzY+qeTYjCEwkZCohvGSI/aEYKQggNf5
VNnronULCw/IQhH8BZV7hinxwC9IXJkpNS8SLoTuNRCBIwBX0JBph3q6MVfWdfWC
rxPCqpN/b5X7AXHyN5vYilJfXW/HbNKMzOs4hbLS83WCuSieIkk+N5K0EaNHf6X5
+c48FLWgjUI8LgwFRv/0Ah6kM3gUICR2A8Jln71kvDS4fE4LFbspht0TjTlLkzDp
ah3X53x4+VUtHL4wI41uIZoEEOt5t8YK8uRPICLqvDDcpX9ZAcCssl/uvy2tD0/B
qeAp0hNrD1AW1o8IXLrLcJQNOjbPlrQoalaIHHi+nrsLrLnuf4w16J1cmc05YPPo
mU1fRI6+IkHxoK0ni6WF+KXLUlKl/RJDD3D8J05BAiXdWWRXmjGbxLAkisXQiSFD
bBfvOg4Lf/TJjrKQ6bp7xdhTIhrrCVwzC6xsSOUhW7Ud1sddujeBglgRz/nlRbX3
gF570h/JaO7SU/S2JqaJsrN8+Si15YwhiyCbkrITXfebLUqn3OYYHiticS812P9F
rkwygR5B/VMrnnQ113PFEKauEvLigwi/5AAWOvacGall0zc6X0Hw4ga5iu3D4rSq
Kv70Hhgk+e8N3tjneRwGv73VRaKzFxWScHjSfwzackA3EdfyoEb6nwQWPBt6XZbf
jaGF8AAWo+W6vKsGlzs+fYRoFzi0R5pPVVHfFQ38zqVO2zq+1Plng81VD83ip/65
Zldb+Kb3Gsi1bZ1ApYtw6NtHxDQYKfTpRUrFKrx5gjjpfNgyczy9HTR8Sgj52bqH
0rdgTLiP1yd8Uvx8NN78Tw8sUCGBvR3j8omWA0sv1cp5f2Z1xXs8DZmY9ybcgB6/
4y7jBOH20muv9mwmxthBcsdpLcR5nHJ5xVqN2p55OypDzNk+ArZr/m6EhTvk4OY3
qPr/QveC8Tcq+PKTpCzYJA2VDfqbAJAiiiVPcipT4l2dqtn+8aG07YSkvyW0AlT1
eLeUf1+hqEhnmOSObwZhveUOD/hHqUlZ9QA8dVq9QxQmgKtWaEunvPi3qvUZRynY
1lz1rASrzYRpuh9HBjay1C+mTzHII6caYo0q7HSNYFb/W/O15y8ooL3sWosxcbIC
EaBxSRPAuM2bYI4Li3Q/rjrkFd3vesUBSXXqSKnUBaYCbee2fIvEk+uUIdQc5yiq
t1fq0USd7ZoaI/RibmlA16/EVLn5G4KNMMOlSF3ugVWjPaK12dWX4I2w6c99+c1d
0MWZm4I4H0fo/WyRNmUQyMimjJxh7bmcxKotOp0X1gbqH1haXw8LxsgPUKV257yc
BbrJouZa16wLhi2nZnJRugIJp2juYn9LHzzLZFaoleu59ZqLmDG/hKCNzMsa4ETH
0G7aL3fGSeJR8CFLDSvJZdtVwYNZhZLX5OUvD74714bOubAJdwRf2qjirG4/P6sZ
rR3Yk1Lt23bMORjDyW42DqNOocevfgoUcbYPuct2yeFV2QYLAuVkSqA4II5lRHB6
lELv/I+HRsGvCQZQ3TfUDq+N+5bzGi7wIzwCoISRDq9zRIxRcxDzmz8qm2arCDUP
KgWijvCIAB4XEIgY7ujeQhEbiC4r/cvfa7nFyt45fZkQgps1sf/XHVcEWzrYzsm5
qScD0H1LV292Zow5OAn1fqeo2fElnueKmvOYz0H2LO+gJe8l9Ui8PemJaSiEaiHI
ajkV5Wo5WnCvN+1kNxEufgmSkE4lfjpBxA0V5td7WgeFUl0awPcjD88GfA0qraLB
bEK5HUmhkyBgQIVAaJMbua221giPYkaSMrLi1+V2Pd4BEqUEpv6YcLyvk3/FZXZA
jaN14U9o00LySmkn0kVa8H8LSRYqOPEgL0GR85uvHLp1E3i7bXulcn9YwgD8RTCH
qpiIbgArZAoeYOM3R+IimsWVJ5cUKYmjRvrRBOyMN6+azQdNX6C9SHuM+xpv7iod
wP4PJ+jwrw0uyZjfVM2sPOANrMV0uj8OaN33pzKHgea0yl952QCwcn0pUjMNbH4C
QT6DIkFLuRCVU5BfUSFfLYrk3LpnzqFUJHSyVRd2TbcFewYvHbpOZq7HEbWhe1z8
g02rXEwKuoibfnS9joO6XF5+CmcmtwV80D+wamjROYtZh2Q2lozZQ6mdalWQh11n
TA9uPaWlD4bmVyQGK1oQhn2gEoxhk2ESTXEdBFJv9kYcvD30Z9CSOl1eyb8F7zWq
T2eNQALO04qSH2R+82GRgRwaWFZcowHHzXNAAI683/q9LU5feuWzj/nOkWIh48j9
gT8bp9/rYEju30YWFtF87wis4aTsyLHhyCLvce6At7tjNo6gSJVFpOPVyStw56PF
vu4e96N4bd3VbTy7hQoXjs+zuwxFm/su1MB/SsWJZ80YbyeBAa0NdycOCm6JnyI3
7dmZRlAvNh+yC/+Lc4XMfLBoGKlEWlUxouAHDhSO5abfIy3mb+AXXL92CixEWIm6
pyGRQ2S7dPqH+mlgngm4HvTudCeMFZt9f82M5TSQldLlB7QAvh21FsRez6DdOyUl
Psqn4InLtKZKqQgbNX48zZu/BPCqauRBbu8kKNuSdmFdGk3sz0SL8ceRh41dX5te
pWs0ztQ53iM5gEQ03t34QJ3X0ixgu04PVCvn7G8vtVyukXfm3GQjAiR2lJ5EMGon
ep4tBgjTMGyq/6WrfPuzYZRf21jYl29Fw4j5vAuGGEFroOyEBIydtXgyUHvo3SyD
NDiVdyp2XxlUQrENtcbLAwcO4CetXx8GUKQiyAEU67jnlKs47e1XY3iBJeS2yUN4
Xacq3G508Sz8xhIhuMDs1a3ZdlnQPVhb9eC/WjGA3VyrGTB1SoNqzGZGMMsuR/CN
FDGu+dFxt/HshSZ3AA84K8QWRPrzsM17HiXsOzPKB6N3tfSVNuvY7TV8e7ThJTmk
Z0pdrdN0SVlSrjpUDgpT4RqPTP9wrxUHk2NT7CXC/iJlgq1kR2jfMBPJIjfK1WXW
JssvN9rgrYowpJEuKmZoQWYMn2DF+YnlVVNQRwGM/CxmGUYq9zEhP55uVaTyvqEh
ctg71iUGI4ArClhoo3XBnYhoNtJ6wBABHciqlcshr18wNAvjePYK+RfVjUJZGt/3
4nFRs4Oaw8dHj5+CumZ+mdBMg8WpfL7iN0k6KtpkzZJnlm7vXhBEAWOrd11rnh8I
cQvmeAY5WS+vsrSKCqcPo9z8A7caY0CN4jGkvLtgJikYIdZtvPgGg07BL0g2CQWZ
j4xixaMvJLpaGRSPRQpyyzbnfsg8CLOG6xBz65+wFxGnHAzyE4ijb0wPjiAT9Cz4
zdOD4G1GFj8lCqbhYvsAaOsMQK9MJbciF/8vw+j4DxedWTuiKzyxljLiPb+yKpIz
aAjoy3oVFWgtPSsfmPwWdS9uUXHg1Sx+d4eNaKiY90ye36MRGEJ5vI9WWEZzZVdD
wXeMJkfm1B5ReaXM1J48dnKCxjoPasHz2Nz6jgduH6fPuj+pYwKkWpl6dwIz9lzA
06N85dbk6Q3qTqslk3hsshcNp+kSPHZ7wt9PoycB+At5blwS+r9JtlxVysvK9Dvn
N2ppJkOpZTiBU+LbWbU3bSn+4LiJHF197kV92gkMK85QcnnK0/NjFDpwYa5SJRAi
weRpHYMJoebitw6FPKcggyR4cN9zcSdKwCuWNowpbwbLAtPx5KhB2GydBR9Vz7Jr
x7r6xt6S1onsEuZWuVB7Nvf7Mvztld4YnxsNZJ3ot6ZMo0a8KDTeBbR40sFznC0T
YIrU4/SkWxxajpSPYrlcJK9wWlkG6nPZLXleldDCaeVaRyCPFCfVUMM8XAzuHITI
jmXqOhLDUYOpD6BQ2RNtEAduxOiDYqUav87pL4Lz6fe6l7oqCkFv7XF0/zQUEokr
oa0XVha3DY18X6i08Ak3W44SwR0uOpLMspcCnPeHwzrFrTE9q8CLZdbi0hf5ZJuN
DUEsiL8NpmF/jVQqBiWVaM/n9de2ThOAjtHOPMdcK0jyL/SB/T2w4UX/ysXLBFKy
Z8zDg6QUgYCAMca3CJKpQa/uyyyvXGcoJx7mVeZ8n7N7Ctybu6BSQRTylsUp4RLl
p4yxYdmlox4lr1bPaNfS0Ocl1r/G7JMUi3FFenIEWWbLKSyQZoMCFmaeu1K9lGYf
rNxHH4zxDOofAlfvlpr6Q2EPWuEGbmIQlBBL5F190CVUClYwIV12nnpBa2Itfsau
Dk01o6SFr+EuMrGgDXn+tzDAoUyDPekthLiTRIg7/HXWDRmToezweCRUmAvBpnYk
2jduUhBWbp3i51sK81HlN6Gnn56UHor2x4IrUu6TxizVHmT3683tDadpP9zX86ZG
zx+j1SagEb3JzrzzJZAhS3/OONh87rFDOLjMvKW77jNW5kEDUSq1kGdTEULtQDDp
B+me5sC1aQrtb2bbkaH545aE70r1IVRua11UWsHqVVY2qKPsk0x68ln8xgZe1aOY
zsBZp8ZXGhWHytXY02EuCqzcEONdp045zC1r3Ars9bu6A2HSooGte+m4OhK8axT4
jJSjPqhbjxDHci/iaHuyWAGScQyH8tv5VBMPqJZFeXz4T+o9BdLOz3Fj9zcOJJNd
xxLFh3KQr6Qr+21fZ03GGGtfAkzIbGJDePq8eEDUfEVrQb4yC+TQUInmUqz7ODPr
vOlZIKoc6QZ5F4RcLXeXkK9ocmRhJhnyABLoTNN4mGQWlOMXMpzwE8P2jZ1Ox73f
j2lsRqeRPE19wzkX7Cj63h6ySUdxEeGE2L8p/VGqd0Q4Y/+tZHs8hsn9yCDZ0xTQ
gqn5VQPatK8Waya5jFuYONN/RroiPUmNkODGBx37/ofFi4xxIgXQdna+c5OvbHBy
UGF55RQlytvSCj5JO6IeB9BBVtsfuew9sSM1Lv4DEmMdnnqxV+3O/DSDY2cEpOcx
XZobC30AWBwXI8MUHPzBszN7Q35SNI/s0RFnwcc/8/fHvkyC5jIPPsGdK3AkyjsM
vYOr4kQ4C7VSAWrD6Z9OkTSP4EvFBTbi+drA3QnyRVf/0G+vOyUjRdQQftJjGT/A
4sGIZVFR5Nh+xkUZv/50OLe9fxTGB7UYSZcS727cteGs9hgTESF29efbfQFRETji
MTWWiLSSHe2LGczyPvkR9d1Pk0/Seme6fgrl6rXvIcWAjirBS+hXIbOjh5RkmNge
ccXrvHyP84V/fKQ2o0GyfG6jXCBvilYK3reb+7DuinymlTVbUUtP2J1FSxCDlacW
5QcWQXouRyKvr+SRVEZQpKtOPKN5vQg0NbzAKi8sXjbTrtlw9gxtHjTZuth1B41w
swEq5YSnf6tsX7tt0xWEY0Xw/VQ2EKjyRKO4rnKPZa2V8hRxMjHemHl27rf6Kq+G
2hPv33YepLKYsQMvEGqYQbchw6IXe004NQ9E5LzPNE7AnjfHb9R1BmWjZEP2rFFv
zC7FtdDDNZETYRBUxqPMxBnWaYd13VmmSu6Okj2dNokOQPnMVZfxSuQURBSY1mbu
8osOJsm04I5LRkI33IOhzWb6IXWj/O50AUrzB78HTk7VEGgLFaheP2KhHNZUEb0s
+o72KDDXXMgkyKbIHuBnEkljFSYFJPmQPsnopTtG2SMaa67QRoKNufwK8+3Lek0I
hGG3VF/MsybyZ3cOa5q3RhS8jxfNhNnEi37W0kDk/6+mrfnLSD6ys96fAv+VvxfG
4PIJqBLWJp588RRhKDAuOFkDlJYuYvaQAsbGEkYCYB35msdBtRCrUL316sslvRtG
tByQ/i29naIRo5oxB0dzxvwVuoqRJtk/wpWutxqd6RcIfHJASL4i59LckbBNamB3
EwGSP3OHotc9XEBd9Ypq91HXz12yJFqQmTwOmyq6Bfdfj72GRMdmMBCXDhsOXPzm
bcoy4xduWhr11GuUDb8/fy+95+uEB0TaAYdD4y15S6vJsw0oEKUlEMKBjh5PUzNV
YTwXu5z+6l6D6kMfd8+zGKIuP70qgrqP8iGXzOaWuglpYe4jYaZlz4iRhs9IScXy
cDceF64XshUcQehlkeLrexohx+e5kSlhdRD+mejdByhv0FSCl6Jd9Qi7jsJirH3p
7C4sJTNUSiZdFL9yi4qhZg+vzEfiSRHYl6+hERDp4MTYIseIov61Fmseo3B5o9TT
dKv38grFk8/c8E8D/L0vqdERV0i56lq7jpuGhVQ9WzlD21COtNFyPYNZ8OHIKr1D
Rse9gnLWNLDgPop8NYrOVGZ27hDktY13A+tWiYVhQXiiLMpL3quhISDOtvI//olE
frrbUwnP0ALpLN59HmGK2cbbJi9zdWPRkRduPwf2SOSz9RKcVh7ASYYUjks9Lmvw
RlDh73RFo2oubdUp8hwwyKRiuzj37achcVIyGKwWoaxWC0IS2Bp9wQZhgoqBMCTk
0WSxy9l+CF1z+RHMla4h4PyNr5taZxbSoF5PgIikbVfxOsGFY618S8xGpd+Bum9t
IgVdhDzmXVERNz6IA7aJKGaiAaonwCXu5bVHtmivLoUPuuesG9oDXiRHg2kpDqON
xYz6S/L007Evw7q/bccccD37bn6UXoxtz732Xhf1k3+yKjM8gSGA+VhIetx6E/2N
kzICCK3hD7tWeg8C3Zvx9DIx0Rp4yLzk44C4cnrS5NcR0N4RzywaDE8PvUHqKmP6
ZBGAr23Y+kROyHwUMHmVXGMSABTcGWRVzKRrT2DZd874I30CKwEhCV45lRXFvjL5
6LhNnCR/ngdQGtXAMoPOuPAtN6MnVrw13EuM1CLuAlwukp3pHuFFlHkaR6Snq8w1
/p/swo32oWjQi919o0hk/oiRFm8JrAdsmMUqugnYc52uLAlEJ97GOndK9CBd/gzv
ueOSZ5E+VtYn9Pyj7Fuhngw34WnPFoHtzk7rSHIfEVZSnT5yXWAIhTg4+dHL5A9J
yNozt958S7Ymfba8OpavBkfWt+19tk0bIBfyYmh0EtC3hsx4HTAIihu+4HyZdY6T
yOhyMsKmZ7lUvXh0/sBsEMdX7MOR4ZcwaJ0cFfpF6Dl9n/gZtHZ7uCavswrrxwdA
qAvvpDw7zj27YxxOqg58oUBNhJm//nyH777crPAvIHds3XwW98otRhUwneBCVAgS
jcdU7r2GBPZORqJSGSm+WClme9duDn5koCub1f+9TQe062u70TD4j1IoSunIB1BP
uRq/1y8XIi8Kf0w8vuPYuEHPRnYQImW1rvxTIV/xMRZwKMTdWST+hY//R8ctaUmV
uqO3pl7FQvcCuV1ZM0ejjaiUsM0Mb+MptXA5hHFwNx4yLHMqMZ/4xN1ugriITqCC
MCrN/e5f9L16UzDVJDqthcetKwSha8Hu6bUNca38aSAhTBSj5o5KJjaZczjH9iWs
6mRkdqMms0vstwWVe07dCKK8YMj27fh9lNukmliWsKAMep8CJEiCpR5JSRdxiZd3
hWcWVd+kD8JAQA5Z7RpOvzHtkYWuKaHN8biovY/qiwfovXpmDUxb0U1y5OOZMfSQ
211bT3jUeFbzedLs1fbZnj2wBSwFb/Y9cVyTPgFtbhaDcGrB3OStLhCunXLc0qrZ
VqEhIs2b8TDzTWapKHT92K3VxT2dCpec2u38Pq4YN/h6P9pTDml9sh0VoNgzkdvA
v9ChznWQ7xSEqSlz9gNWkaurqniNsspr6W3Rd/zXp6Z9i/ywdJ3Jct/iQXGZtMdw
wF2POI/yw9ucYYPP1hp+HYdIeJ7T2EZDwWfc0eTH0TRfJqgemr28Izp2kS1SBCLp
Yh1gu30//JvRBfl+YvVkIsp1OVNwgg6maKLcpow1WrcNzSh1qr1Hx1B9hmCG9M+C
6HIPTAFtfKHq+SbvSC9G0TRpmNufQ3Sp6hKO4yhjcn6t1/IE9OYNi2Pft+N5ixVG
7vQwu3Y3xTxqAcRHjXbTVxD+kqEYEpvO9BD/+26upnZ9nHvKXyqen1FDrmIENpzI
bfl9zG8jqIo4McPPxuD7QNH56buv7Lm+PF73auN6SPghRzuMIxAP+1WoEXBDU7yV
ixQXrk8BTrRxO7qInbV91OuQIxsqGcbEAkpHzWrt6krvmX1PLgNNGdrdUSiK1Eus
ck/CSnm/iMuCx2Cpun82487duok3aUDgrvC9qBpAL1sj9ZQ/6kgoHph/8cUai/fL
g7AwwAaBeVSwbnhg9TalpXx2FYyuJSJ3xcr8eA1+gDZ5L0zIbR6cSEaxIhTdvS6x
tb2yz9smxU3nqA3jXXAKW9BErcl2DsNaz6XS4nqFRX3ZhgeaJRINmGsN1vHU0UOt
OarfQ01t4y82VA7Cz/IORhj4c44JWQA9Bo0qdY3aHgayzukCLhSmLVv9NB6gIJAv
aoCvVGJNqO7nZS8xm6tXN4KPaJphnDjGEvTL9nKc0e4GUlsvTpshCNrCuhmINjMJ
Oq0/JCrTuZkfZxu+Kv3KiSPt4yMUuIV0VevMe4ZDcBmcmv9qVNaNce8dSVKLFD6u
YdH3DTS2LO7SGDjvTtd0ch72FJUgu4ucu/gB/I1P2PaoL4bBAk+u9VSKSIltAS0X
PX3S+j5TyAuiXJUlqldsxPZAe6fd5a6As/8j9UiEnoMdtHKiv+24+iusiIpoTOZQ
WH3nEJhmc+bNPe0Cyvuux5W9x0Jg91pet5bm1GneNg0D2Wk55CzMJzzGKg2BoORw
xwTb7rJ2k8SzHum+VHj/pDQBOibXiOxBA2OTeFtcI93QeIQfz4cbn7PXb4wvq2iO
R6xftgrbiuNO6GePpQbp+zAj3OGnnsdjWDfIVzx9b70JlorhnUggyBduUAjdCxYf
aQqTRcly7FWhLjq/4CA9L4XeEWAsB/vy3DmqJBU3qP6jgvtYjZv+p8pRhqp+mGPL
INR6+DanM4enRMtSb72HZYVDf3eYYmlJP1PV2EGwedz3mWbjTuKARducomo2W5Zc
y72euMQPfd99wXxMU05khIz4hGxvtjUUaqWtN7fUt7pIVkAtnpAQf+WKvA1DC0KP
3vdyw8H8HAooH9pJgKABJelRdsCFM/tCW67LGLJxkw+F+Mdsc7LXaG3uhnyxEwbL
XbGBUJRcVa7H9ScqzLXA7lEP5zs/YL0zv5KipYH4rH5kgvUIg97KthAvalepj3UC
IAiNav3SNe8sA8FUw/MwtISgSkUuKQMMSkiGX4nR/bGvBFdeYA7lp2lwPGRKSsoW
MtXqwvXPHWzo04bEIPMLVKNHKbO0jX2SyvEthQHW5yIa7T3P2WfxFG5BEf5yidvT
DJ/3FAdQZyPvGs1Q5hGGUEtAPlq9P2rUbx1M9UZkWH8wA78pOhGkkhvViiLFHE9n
Orz3eT9xmW64sYsx9RVmsJ2Swpo8NUk08Ez4UopdipzzIC6TqRqVwOKU21BRov69
lcJ6Tg+IP2/Pj6mmCFIgl4RY6ePhUiabZ+eZk9y7ulC76D/ze/cINZ1dAaqoiCx1
7rT/dKod5C1oyuLklxlHXACHISXVjIMF6THmQbGxlUknK3PvWHjUhNNRso/XpQn3
+doA082NtFno3hwmavZxHUuTYa6gsRpe0nDt9jLuQl+XQGEY9u3vgQAqXlTQ14hy
QZ4bb9bxvPPOUaRYLFFu3cHqwbg/BAWV76gSR81C/0WmHDwdNPqPgPdjGn8PTEk5
SZoPvPyJBuq0HTrEvHwoNYkFGXWIoW/o3jVy5o4xmNfPmSvZ3VvA1gCRhO1rfHYC
uJk8fUQln8q/YCg5wDIFwtNnaZSBMolFLNWustZnPGsu26qiZyK1Ix64KDTAerrg
1DfhymprM+FfDs92ck5+WvM5T1dgnUWoW0rjs4cZhJSdtLhnQksejFhxuu8XSo7E
2B6rm89j2Go1oOz9CI2gh/8uVdEtrinfeMs9G9qNefKi+ayjtvI3F3RUhkxgfEBP
zAfW95SAM285YYZMjSAl74Hc2pMKrlu/EoRHONsfa6mp7+eu0ltCNdIM1YUG5b/i
xinX31OC8pKK5Tj4n24+9jO3i14UmiDFNyGCsZ1cCLA4b56d4ThfDvVEragU3Bb6
JsIZEI8FFyqSADtcubYghci0PTSr+WnOx4XcRr5RNpxDLSdDfD1K8f4bL69g1nRJ
YSPxn7df+jmOxwALK0GbNnNIMHhesgJudEVqsYW41oOFSzDyQCLLB+b6Rd2TuABx
CbdGxLFHWAVOa76HSntVeA8WoRTNj4IduXww6ztmuYyRb8cjCxt2HpKgEZBuvO1e
H2N0AFdvjk9x5SXy0jeDAoDAKTcKYNOnAe22EuDXnw5LLnomNwFAepbQD5zjcHzU
gktamhaZLu5IpYNFIKvMqGRmZTx8m2UAzL9mU/SprsiG/Y6gNjW+rxm7oaIoxpHB
doqc2Csm4mKuttzXpHz+PumSkGXAjExX04i9H3fBm3P8egYT+bIztk45nAL/u0b8
JHeZl4gs6EU/U6dPULNQhT7tL0OoXYfl4OTGCqQRdlR6J7RZN7fCKEaXCSuntFwd
j8FxoUcC2JETxO9c0ufxYcXCjVNeOoH4IGKHbFr+8YPYwogenRok9tuztLxaZt4a
mlSntF19/AXNg8+WXFoOccj0yhOvkqYeffCK33fUcd3XxL2NHvcZmztyKQs7Mvup
OOBoVqyWIY8TCLD171Av3rNcKvLdZuYWqZp2KZw2AuE3of94Q0Uqs0gGyQ8urI7H
Dntu8t9IEnbu61LidMigqI1VPxgEyr6i6PCjM/+XZgwv2YvsvMfEcRlOwURYYSHk
pyoQmvt2DQvZhvZx6b+wNc7ah+0Gxed3zkV2UppfTRC/RTdr36uWW8H46gY6nnV6
wSze2LBwbB6J+nu02vDL8zIbRYWBWu4KFwh28WtutsV5N36DMPXRzrIEVnHQrx/r
MoXBDiLUwruTsoBNPqhC0/adYFsG4flFLuHhnHWkApxedKC7AyIEzIQcbxnS2/cp
+lCFLoXahvV6VAUYXNClh+vrywLDcdxpIKNq1Tn+ye3Nd6EASsWutxXtYDlqzWxQ
2FBvRsp1cbsYXOpUfNGsCXWaquzCuBESRD2kNqDTKpyRHm8j9LEWa2PDO5uHwxg7
/vNiJjK/5++BT2XqNMvGiDgZVqYT7QZNNdPK6JcdPf+KHORkYq4t4xRQXAWT6eIJ
yGyV4A09FSJC0wVOU7nu5kiNyhJfzvKf1d1VBtdpV4P1Q9w0ITEyDPTxgjAYCez3
PTRUYvobBTfyn2uMoO8PhOzrD09KjKjzjkSDMqWh9pSIG64PlLos0BzEYxGPFoKE
/ykFxTZtDoWp2eyhYrx8AmTtFoE6sVfA0+6ZJg21RMUMqi4R6JTYG4yMw8ZcVzaI
6DCJKTqHP2aPbHcTf6lZAq+KBD8ok1WkvXw+fw8DufTunFD9JqKhHHfMmjZ4JMjv
O6B+w0aZyQSWJO4Qsc5YpExvANwEUyOZh3QQkDlTQWT+w4K0AlEGt5nV/Rs0aHsc
nez0LI70FwmoT0ilRU8ejbWOGQglfTxCh//8pLjJbZni4arMjrqqJAtEC7bbgWeH
Ps4cLD3X6aTx3IjEx7BdePrUq2ONc71qbrWGOvHI9qNLsgrIEaOug+AB2eM6cmz7
eoxEVL/S4CNCJtD/RnGN+2AjUABtgVfP035HJh15N4HSgiZBKEfd8fSu7M1L3vKr
S1GzGKuYsWpqa9YCMG/+V5sThgfjay8tdHKJ1yBIB+K/sikkikAjezI/Z8e2AM1e
rfI2j0S9E6n9b8+5fRwfT5OLlNT3rMoi8fzEIEvZobB67HzdMRCF7CZDs5RVx/O4
Eo+JmGvY7+vTuO7/DKeZLZhBmtLI6brFiYStOKWG+KGrltqsMXXsRBVyg4ihYzG4
RvtRBb2el7DXuUPh2EE0EtSbKhpb8nzgwzv7BG9PjuySITvX+yRj0kCJJByJQMVn
jEZV6ugUN7a+o5fNZ4SsTlrP+7X2vN2DbjPelRonQ8O88PQ9SO6w7s3YEQoqXEtv
kHjizgyL+eYXwY/ToUEjCRtMnjN+DbAiwyMj5JwFt4R8LMRYgIVCcuIrGLrCib4s
hN+U39mSKPfJKkXLRPCgnPUC9AOI7P1UKFYVL85YhqK4A3TkEuDhNCLv59gm+yAH
Ymd8hFfYBs0jI6Dw/38i7aU3Rexrmr6uIyhAGwqjPA26q3xS7VQJaWbI2/YZSVm4
R/XX64y7SoByQ75D+fuJw6JBNnXW/hN3C6/2GvHSnw7NtKVLPruk9U9QV8pw359C
aJTA6WtJCzgvFSA2vk+wjRaTREEnqGzPrw39RTlAlaZHJURxtbFT0xpAfGE7X86F
hA4tgIG7vfs0YUyD8cFpSe8IM73MBYZqCtwHR2pTegLX1Gh1isLygL/47lHU0pLH
uVlugLjM1z3clbThYIYqqNUOPNjajizvzcZacNHOhPiD2tOAG3OXJUTCCpmHbJpI
bF/8rRZS8jew6mBAEeQjgGw2zyfmPy7uRTHP0KRRNF35k4lVwbLmXRII8R6QPypy
gYP3xxdDo889aL5rvOfyFNhemGyAPbdMpG9xoV6IZvq5dsbdHd+0cpePutgzBoJh
qTxM4/PE96mA9tz07UrUAxUiLQVlmmeRnpJUC9GaA0b6t1LiOtqHS8KJiKAzZEiS
vwNFRbZ6jvqs52jFXLCW1vnbp3kVeqbO0vAQgdrL6NoBfLoyfbwZYz+PAm57xTSU
Bc/ZYTm4jyEyXd4xLY4LxOPbltOkQMCvn8pF3eiARtnhFH0vzGYO2za1s7TlWIjZ
ii5vAi/j36tOCJkt+LMkPJ+FZ+vQUh97Xi5lYGPlTLFCBmFFWK2zJDPVn+7Gw2cj
9Hx5Udneu3PJVOL2NnNxsHsn4On7hDq67/gSCMDcCWPu9KPfuOIgWKuZgfu33nIr
stwh1X9C+f1gBQ9B6To8oXUu13xkX6fzForkuvVOcZwpuphgPCAOkQz6McHc+k/K
FPbkvwlIbf4DolfnElAdqL45SUDycmXfwl2BuuZrsO3IImF1+UxclkHe2PzMYTXQ
uM9+XlHxiL22X5ZxntGB8lZKhX/ZKZny5b2orYT9bpE0Grzgl9MginA9HXb7znS4
rVkRfAFtBbgvB3nJwZ7fuIDnZf2iJ/QKc9WcgHI7WOReNpXsfEeB8riljvWiSD7k
hQG5vbyBsXeNfljuGdiywxAE00oVIZIXZjbdk0yRQUj4WWIiuI8hU9ehOjSe82W2
kpb0QrEjLIw4uHbKvRTLD/ij6CShLq+BPrcy3bYUNOu1gijG/scw7HrHYOlgm2/L
SI0WD5W4huwad8yZBmPmEgoeZqQlNNNWDCxLmd9n6JkVTpPFdY+ixwEApFF9mo8x
ZzvBI4TWA+HoQ6VBr/PKr3B7XysZZNgSE+E6HyriFhkQNcuugcKwuc5b8O5AX9x9
ak/h9ywS7r6zp31P2jM/TWjUyqX/gmIE4PKFRO9A+EZFw9MnFFWvcHV4YndT6wqb
lkVwwzpr738DUa3IHAO9kUagoneh+AhyFk45HlakG5tSy0Dc4lJHakHBnQKHGKsM
pAgth7Bd3jr7u8aT4KC/qWsD/rZV+zPRcLBYi3nmr+S9QxpiHju2pbRSlZnvZ3sN
HfsFRoFy3uKev27at2RLGmB0IgAO6u3mV7WX7N1kirQPIZB+A2CsjF7O0uNyEV0u
ajU2KD1A100ksBtGjafOm7AD1ZfCvztkfEeUijtVatGRDtALTzv6MkbHqgOQpHmW
qyg4DxKpjJ3bRBKH0dt6gLFNV+c7iTUOXka9/fYznsNMFLB62y20lKRrtLGNz2md
1SbsumMdkG6ZiQMkOFFRue839fo+167truwpxqd1hC2mC3B7oWvQsauJGYC3jf7D
gpY7I14Zf6ljmxFYtmdT63jNNfDCZ+RKvCVahQ7Bm47HQfy1lQLumiCBiXgbthdX
V+O6swrP3ppNEmJh2xI8IXEfxVPz5911GjwPOUBOa3IemRfgin6DjTelXKTrSy3H
KBp+Nb92YqPDOmk2uTcjE3b8MLtVPXH2aJU1e5U5J3dUUQg42A2mArqwEdB0LSgZ
8rfnrcp/z8BhzyBeqtglEwyisSyGaUI0itm+i4bucFi9R5BV4E5gX7HerXtJNc10
pPknSoyRP93qYtn4T6L99n/pBJCcpZQPpe11WHP9glOWF0mQlYDri4w5NXZpCneR
GjpwPH9kdXIc2h67niPiNe5+gKVkkX/JkGIc48fgKHZfAbGJToZAz28cAqY+n0FO
dydlN5G2DEknwD82W7BG/74DhzeVF5OEmyM0KORpJ6XJI6pmMruawl9z0+SvBAIa
6kHcDfRWiNpt1ilGLCgHnTKPm4mKWtZ3IuP+ZWQ+681ZEJ8zkFmbIFeFTAb7oifX
TXwU7xg5N4l1/nqhkbeb71JqsKelyaymRe2KH7CHASfz4kV9ejcl7B10G/NEFDPl
Tn3LAwPlRKWnfTThGk+WGSzXAg+8frrOR/yQUOfCssiknIBcE9oPjQfzHMTJe5E7
sS/yIju0PlinlAl5GClFeGeo55s1ZlviGatdCwDptnP25ZBj2QMwedSh7nYHxCrz
gACqGHv8AemB2xqwKsGTa+4qvzjmSkLjashuir7UziuhAAg5p/NyEhNLhICdKzn2
Kn/4VlT6Rs1I30lcHNcmZAVonmDSx/A1ney9gjqu2V2AipOCSp1p1HEjHIDOF/qF
D2tS+SssvFO4FCrd6kySrN8OqOmIVX8oW6yU8OS7kGFSxSd2FGadoR8jTagpvfJJ
YDmlAneF/ewTkWMo0sTf2znkH8zJMb2CbmKz3tQQdpVTsSZMRSu53rrpV7s0ebzZ
SgrvdHcuX+RkqWUBRV8NG2jyS+aBvsJT5sU9vq4asarptMZIKFu73c3tIRFQW7KU
l0i/rTDtrgbILdMQoM1P1h1FbsRiCPgGGJ8Yuyq0vXSYJJ8dnVwGZWxX2SoBXk0v
JyjySmNiZT991r1eywtgtAZOhCkCyPKleFEThZRVyeu80ZwVSpsOvvR1+7y9EtSO
WfaRUDFgGF+/nth/4y0RAAt6VZ9OKP+OfDPWUXualL0Ydp5q9ifPMAbHWYRzmAk1
YM6HACs4/EZsVYWTDYkzQKrR6wZKYTvj0MJs3Kcwa4U9WqNRktJwSt/rF9yBs+Ll
twYcIQ0FZYq2cJR/CeAeWU+ZOa0nFw/AWrAOAfmLODeC/I7fF378fgrZUFsAaX0S
AVZduz8Xl5mjEd2TZ05yAjNSRt12aphV8w/BW/mJ1wqYK96T83BtGyQlPPK+j/Ec
CpOZ0I7QXqCGefNdwIMtjTxHUGH1r0fKMoj8Xx4kP6uKaKukjA+hXWeDR3ckBXmG
hYur4pDw3TJYeuUlKkwb9D3hRx3JdXrKf3dq9rxuGZqPUw527f2AR6Eeqqkx5Pv6
zHZUPeCzc9T7amg2UWyTdBOjag1lCX9vlPMPVDhIdgVpNwZUojdQ8AB7zNJJxmsv
5qIlis6Hk49O2tuL4dh9rnvRhT/G3SxD/2WKZ7pIhKFzaHc4GhBNBiWGTL235hBy
GadpPjSaTT2Z4EUQ4ZSKVLab4W/v8NFuvbZausPKi1Zs7ccJe6BCfytaAHPTYJOo
7HKIKd7bInFHJk5rYrehDVVc+cpyLpIOcNg044gg8Yn7Qpj9ehUp+xQO5PbjLksu
HP+zdwZa2/Nli3limvvHgDPG5zjQXNTOTZt3vWSbBwAO/c6wqpxhWd4GL4tPqUPm
86GEMMpHFrZEyN2n8FGtg/7iboOIzsY7izT0giHUXovhDAoRpUYu7hQAPblNj13w
+03CklS+aWRsxNO5vLohmGSsLMZ+Bxnvs35QIrR91CjWbfnt59RWL/4C+Bc5CUy7
H+c77GUO3/LT2jeO2nGp80Ayl+6WJ8jeI761fJmv/oaHRHQZ3EOwzcFKJON9vJyI
s4jjCSybgFR6JV3jqFltRsYMmZHu/s99/hXZpVjhJGPA8Uhmq/emud/rAGv/510o
cGTQMaD2rawr4azB6Hu/mnKDfpetJVwslvCIWYJsXtV77EaYFQhN0kSUplvTVIIF
e+TdyVNDHpXfyY6eG9fJ1Bcz746NeJTUZ3bAH8K3T9ReHD42xBT7dBQrbyis5pHI
Z7DlupLtIjd3J7ZLXKjuR19u4/6QnJcLd1xZwtfajVOxq4TrtvKltob4kfjK9bjD
yMWxsGZGVa4OPZTxtgpcKXgerOeBa8p/KSR96JowfhhlDRd1httpOwdH0pxTimku
hA36XGG0czCS5drLod164CLZAvRA6cETVn+otByl4f50eM0cr72roEkaUlXtuaqo
DVc5n+FN4eWbeQLDbuX7Ip4VFZcjy70NX6ZqWTdmnhBhnvaN9bNl7RcXREApzlUJ
3PISoJFNk2zZghjZDr6SKudlI9P0NLerdrCq+lcCs6eIj49sZ34JLs1X8tAhwNq9
NXHvRRa2pz73Cc3iQuSniJ/+gAlfMMxwrpu53fujBO8IoQCn7yTRqmc7wmnyU4yr
Sp87lZVBCE5eEyx4W7ZCfsSo0uOW5op7nlm1h0TVkkD0gWexNQJbRF571VHS7wNp
jhFvaSSIwFntNxmrXI/CtJEniBEDM3f2vnRaaKG184LInnkevbVq/NI01IV29p2f
7c/rV+6wTnUv7z3oELo+/skK+gU0/0Tzz1Ew1XlZ93OCe7NYtlOGhFXJMwnqvWCd
K1ModtyuldPaGbcEFgE4FOmVIfq0mG0w59+LBTo9DRr08EEHld+C6yTFoGrHXElN
6fOucLtDsZ7Iekd5XpfKheZNIoteCseIZCNLoIxpYnm/2nv8MLdAE78FY9QTlQN4
3HRYR7q7PpieK82NWDxuYm2uR7Xn2BzI264AtYSvGKsfjpbdo8YS+tK+kVqbzG+K
G/gHhsjiod/kIJ7uQiwXhwdIzda2hYL2ECoKASck7FYss9CX6+pppQRsv/HcIQBx
ALYUXX6YTTlkKz/a9Mk38Wkgz3ebKcGc02TF6EULmlAg/MoRITksBNWAgK+Jb2zM
2h2WQgCB6z9mFkSuS7BYP0I0uAt4+NP4o9f7IIdqc2l4OtxY0L8SqcO1Tzhhqdnh
K2EE2t0RSbmvR9IAjs3YWOn5uBeECWAstHvtCbKis4sozFhS64j0kR9if+Y6t2h5
3dJ4dn8WZCbBiZdggpoIeWMrNgNNedze7mWyaJ52mC+aulbYAmkp3ORUIiMqhvYJ
F/3FaJOFx7VIgjMrFzOVfRckk1+X90HKjAgocAYZgrFr1TvFU4MlWytItcgoKFeP
fIPvKEuKAnn+DFbgEBgmPdKHqFO5ssJu2HHUrUqkBz6y89AwzB8VtMSq1Nvi6NBd
HqocjiOxWSHbSyBhvLlMrnywyq0+klnOTaI77+XYXSuoAs53YrgQBHEpB07LQ7R3
tIapaGhRg70CI0tX/QI3MBa/Zln6Rz87i280PlJFgc8MvTgOzRLf/Bs2nO6fiUHa
xmRr71IbJplFP2WahP/Yj0GeHsI84JLebSxC237JbU4P7AVeq/QnIjM/5srU5fQa
0ClocQSnBzqicz+OULhY9oBwx0dxtI+dTUvViT0G/NtDogfyGVZuW33OFHoP2Kus
GlahQz0WFbFc7l1SakBSNewVIO1KKddrE9Ro3U7KTlVBb+T+xHwBRM0gpSTZEOTU
Y8GqBXlo8er8kdVF8kyvoimWra+iVkyOiu+1XSKBtII1jyMguj+sxLs5u3iobo0W
oV4yp4qqc3/hc4s392P1zIDUmeKsI+OEs3pMY4+//oWb0EUwK94flT0fwYULeZxR
3UhdumZg1tlcaAxs1htzNOccoEcvM2aYmIxjSaOM4nRX4VJm+4NKMB8mENR2uZOL
ySv5/hyXZPLaTOZcCZZwicBZhkEP6fqckbzdHnJEocYFduk5xc9g2rG8d0xDtZ4D
TVSac1/mrxQ5Tz0tZvtHoDHrki9K17UCtelHEudcsFp+pVYGcCHTemjYU+uqhuj5
3REfB6fOg6Ige0r4nvEHthylcbM8rJYAliV/e5tHZBbzQI08eG2cKg+FBy58hUwp
xWWz5h4kx/vbTjXigLae1hRPVMER50KHHJIaAt7o+wYd7IBQeu0j5P5vbxgIfywQ
gWcXr8Y1Bq8vFCexA7xynt5ZlGc3hsFRQF3Vocy9a8idYsKIGZCFP4NMR7h5il3H
E91J40PMny2l+TZ39lrnkH78JAJV74fjabnpvCaeIvbTDedH1gO2TwZRFcOIAn1/
Gwv4GgH7FeSp1b3SPqN3VmHVH9v7BCPaUTTP63QpojMTsFP6js1+TAMfv6XkGYr2
LIBjkQPtyzAKvDOzcXc4JCwp1EMEtrIRmhrwFko5ToQlDstRtEHaYX4Cqp1LRQ90
GdPL5r/3Irr5S7fItSQgVvahfjfkKlR2Cyx0o5/WbzlpJAgzlFvG38ekeJAI9Kl6
cBwMhB6HeNhZNrQsgl0GokRBnVbYDTzLHFnIOCA+6nI6qOPS+qvOzH+Bo8/VTP25
iy+fV1sRXHgzMIWmFgaftQcK9/0dFKhSk+CaHs0hkZObeR22t+5QTEmBCyncunNx
pB4G710yFJzLVY5AxK52B9kruzXvqfPvtZGq8G2X3bH4l6GvDxW/96/JaRnYfe2r
vDpFU7b83ohW4Bq1sxC3F9szhyVF5xgYlFKds023rrQlPjF6aj27eOELfJa7dQpG
n5m913XLH13m8diCrdzpyC7EocUkZ9iNIdWm9pyUe81OZhPPj06ynNETJ7VG4Afg
Ui4v3SQq8pDMJQ0/pV5NnJFXW42M2vm+oKqgi8VV008VkglanKslBHNHAh3GBi6q
/ABSOlzXRPa8TtCR0Brqe110IR1lN7NwBUjJh/NCLsvYSywEFTNvoJqbQmOC+FAw
3rVjct+Vpchq+srcbaH9XTY40KxMfa2pc745FKpklbuTpsjX4qVHjcOlCGSE5YNL
i19mkrzT2d/IN5nLG19oz9JpNRvtpgpvwsNOWNU1umVr9ZmOiBQlO5YoeDCFB3YI
iPXvheMuFV2tV8Bbyj4M5BuKH4PaI0xQi+FI0lCuyiuSAmtzn4bEImQlRExG6nIt
r3Pst0eXm8EpAJ9FZlO6JBdb+s/0s9KriRH2wUDotz7ty/RDligfaDHdF5AN1aR4
BvGe2g4PBMoPfmciS9pwRwDThIlLXfxgp8Gh2UNtsxLXAFyKwskRIs6CAAZrLpo7
CPiCAp+qeTN1BmYmGDRBqNv5qePk2Zyi8c2V76Rag+xwqw9QFDq+BF8+wC6USmxv
VXvrXjGONcBJeTM9sV/VZA84Tm2FzAuhrq0hoT+vfjzzYNkQHH3cG4YZ8Q+GFp/Z
Lg5lq/XjtjRkEf6O2ViL1ynHleYSFAypDAHWZsBZ1eACG4sqakfOyQQ3gz60Rspn
0j9FLWNVr09sCMqnbk1hQdZM3bFhJ6gWnzZlQxEMdnK0T1zgZsruc5tsYSw9hgi0
PXD6QeCdXHgn64eoyqZTVahPSf3VhvWqnUOaxrLz1tVtNCPW7QLRW+DICrsN0EZj
RZjXJ1ikMLzA3mlgsInwNjG7AkGQWKySpx5MIG/H+rzoAcG+u2zBwV9Q9oKB+DW9
UL6F7gXaJAzps6gxtwzVq5Pu7I4/fhgGAOWAT8CA4L+n1sANF3mgSFL5hqBHexr4
Faj9kYhC0Kz5M5orE2lmABttAfJIy2G2hT2fc6zp5PJdq4oMKApO05hiHMUJWe+8
HNntqx5nimRcllZpTAPwHoYEZlvmPIPYP9rzojnKBX6ZOJDL0VXQQVqs5sa7ibKk
HlCUbZNJxox5s7FhGL1Mf04/JotBlF2mptRStHk7FQmMg/S3SZjOWIZtBC8V1HSN
UOClAL/Rzue4BanCpNWYqGeOIQfHfJ/qfLnZynC5hs8ILzX2j8kMJ0f8QcsHLaYq
xq5fRQRkB6z9jpflbb6zWALgEl5rqdcKxZQVs0dCNCOqOzNT44GINboAFv3/FzWn
aUmpYh9DYhBF/X00Sa3/XnGxm8VFaTp8f9wnwZrZxjraNmH7QjxSxjwfzbutoVAr
iCYrZNz5788P0R831z4ek8U3Szwb7lADpUub9cHIkrdfTNtwM8t/hdcHZfgX2pXH
GjJ7uDnjd9HAOFmlY+ebsru4EASZZo/wgLn9sY+lz8e/YWKCo1altZ8h2xDd6Y6F
3vgHgTOZOoebgaXyU824q7Gnn5CzPluW22XgMFdTjTb7JOkRWh3YVeo23zm/M2Tg
Lxd4N35tU37FSWCNpDJq22D9JELWzrZyKHTz6vCX/ChGXND7Q4w9/9bbz71PN+xT
xidE4QYxl8HwN2loOGoLg0s+wppmWI/D+PzSByD5iGnMBQXi8eUDXHO8tZuXaZTL
eL7m3hkgDZmtepmPjbnD4+rM8bqtba4fd1efKNBp0BLtgyj8EgIIIrTT+mSNlSNK
6+wwH4YcFxARITLwBWbHpBIMEdknFmSgvHAX0SUt0OAvjzz/Mv3zT4Qc6tz8ETeJ
K9hZQHrKae5yHhdhSG3XvIQkNUq6swuiuMH6NmaOYtrOkfCOsNQclBM8cQoicPzN
4Xsw2DCeW3wOx1FFJ/8YcWoc25ouXji4CyZUjPHgWd1OlVUsnlb1gVZ6i1sgJ2ae
6g//VB+HyeNhhzEWAgHcgSBq2mCa4nA2NKgG81L1h82pV/CkrBrlUfx8WoKBMvfG
LbRy09UQEz3z4um6iu/F9XEkpRR7eg1q7f6wkOlL/qqPUfv8dKkougssO6z/wN4f
jJnZgxy07pJp+BwNZ7xnaAGzA0JVRZrVKKDe6FTkp9zJaBZytVlnj6sVT5DreH6P
PtZTpAdaUFNzQtuSrqPIJcSK6jZqRmUFy0DpdlMldrJYlbuOsKlDsyStTrR7Ktoi
fNZa4EvDmLNkK6VEmPNCFoheem2VROu6pjyNf5pQGrsg1xKomFa7ta3v40suQxoX
FJVvcBuB0P4Udm4lvLgQ6GZ+Qah2gwb6YzmHRv8577nnU6h6w0670+TdBwhc9EkY
0PbmLzawKZMMUf3TD/N0fLod5fA9SM1jViLNAXjufhOGMsc0K2Ce2OTkSk+kVbgy
Du83w8Rz0lt8h6WFnvwmhJhq1CCNThS2V8XlGUGrlir+s+t1gy2n2g5JPAJ1TER1
AKZIJtSfEIIxiCUi259lSQke6zdWazwyC0NNz1Z54SbC+h92iGiAdr26FRwSqw4I
Ck64GTr+aLKOaTpAnIypp48mA0JdAPO0Ve9j8+Ad24oSyzf+DceqOEbPhcM0dwF0
HL5C+OGrsV91QA7O9thha5QfqnqiMwve4Mf8ctXfuQHhiWtZnm85SuZl/zj1FKj2
255GO1mFKd73lBwq7ZYQB1IJBusDBYWmww2+zsbeLmwK24i/4liAJnJ+gvbnf5V0
lCUr0uwASzywAdW5wbanwRz7B/7SJ80Z2sLpPYhRciD9by8kvCZl5e43k+Z18wL8
bUzbGScORLp+5SBZz/2MhDKA+pyHVEW+PnLh2PpxBOPZOu4xpvwm6J5jxtFlb6tX
lx4iOFwDF8+PyxnI1Ij54BI0zLVbhulcrAx29FKOk4pK39Rc+5wWuF41ClXgg1iz
fbzIPSRKHoahUylF0HbJGILyCdBU4CmfodMTZTyX4pSCRcg44MBee6j2HXOPR9+L
fY5dJuLZIrBQLdU9hjPe6UqIdgxPMEmPCxB4g7NaofLcvxS/VUpJ3ND8sA2KLP+z
4uSAWjr/8UI221cEfrf7L0OUHfS9q+oAGqqyYI+Vvv8aj/6pJvJCb9UudSqKflJW
klJm06XH7i33MZOMWTPg1CjtKWwRHT56EIRx+AtYWLzw1bZAjUhZ6waxytTtyQvb
YnlwO1JvNqYGcbOUyx2OCk6O2NCmJo70V9ftdjbZBBtXS/P255SxIqOcjSjO4UTh
+WFmL+YNEU0ejn1zFh8zoDZhIBw5Uex0rkIIwgT4vcKtoOY3tvZgp9VTVsxF5v1e
q5bY5Y008mNLL+hsVLIQQHJt9tn3CFQj8bXURaur6TxSKfEjfQRSN6bpkbWPJ9Nd
tf8E9IRISgtRtgYGgl4vZurMnWGZRhUz13ymUo4Ix/GdGi4TuYt7k1vya/zUtiXi
OkMTvF4uEAGHnKUkxOIxeTq+5uTaQOipLaqPyVvCMEATcIiAgEn0C/dTy/RGk+eT
RCXTXbZbIBhrcFvjIeiIS460BCTmLA8j7bhxTBOLNozPo5kTDAUlxXxaYbSeKJq+
qJP/C0HDhjcMeSqOgYeYRp5c515qh1QXVuoxtbTQH2KeOPsFeV2GUkEbqBIG/kfG
jI4wrP4B6rCtY0d6gZqlEJPzBFVxDlGD3p7LW9aySRzQVbl1VCfha9hudh/i/iE/
DBVGlXGHEuf+yZiAb/kdbr/mo96RZlE10jTAYuLCKhnZXP8g4YtlzrDfgfDjHP9j
VsPhDC45J9v+mhn9eBGRqld5voZHATX6SuzIldFBfVSJhC5eDDFjbCI6QbmsHCmd
bEp0IKOMbydGejqiQIoNgUYmc2IZT+WavkHYELjw+FjB0JPa/rtWLm472BdR6ztY
b++TtcTf7i8ZquKXi7UuTNWsZSD92SKL6SBsOnPHVtR0Rqd9iL2OlP45JQZqwX4Y
neea6j6nNIO/Tuil2h2kIBVK9MX2pBq1CfXO+WeC/VUcZWAW0rHNdtxUV/qfEJn3
fFAPXeM+T73s83Iy05qa95Qo+K90Kg/piNnHkzHCvNzyZ1UQk7rv0sp1Pd738t8u
H7apvVKSWpbJFLFgWoAFIbpZbkS375zi60urQbYkLonLPzKu039XjLH7NzONoV1y
Z8RuyXQ/zF4K4Q03rqgIaok1T7LA0XEXKfNgOVey1mK30fyPaYERw+kTyAr16edE
Op0zuDIEOai5T1K6+xHZmvfweODEBQa65NSDXmbSnqe/k6r5MJRMoRsOjJfGOr5u
IuZjz2qWAlzsMPbJoLJF4k/ctbMvqAcqwIKbubUCl1fPTlZUqG4v+FCIIzJwRZNa
xmA7TVYtQmyWIz0ZwMK2/B8WIo6kcGgV0Fnue2LBhPwZMCYADUHS9ABx/jejyeJp
aDITXxJJmyfaf6wc6dML7oU7mJNgK98lGFdB4AARyNazoQvY2/t3aP/o3WPNOmoJ
gxoWlfIPEBNcuwYXnuWBHS8vI5EjZK/Y+4a8nQ+HcvnX3/KyNQou+zWDNFYYKLa9
dDnfq83fxXluxQbQqun3cvZNTucBE3u11VltCGd/LbFgkPQu7FpGyQHu704ImOok
1MgCgsWJ4UXSSBDyJnKcy5Tx+gB69ncH/bC6kTy9iZ2zN6OgLvf20WhF9DiYO8Mk
o39onLwxm+vkeroZHmnS20f/JkHJyCqE6Ld2vOv/Z6Elm/E1ftlEN24eppQzQBUh
QdvMtHCD39xzsNQ2Jz8pB8nXIPQxX7U+ewYTfGeqbYd+8+tVsJI3dYk9HhoRBdIx
U+q8JG+GZMv0a3V8oBm9I+MI58lYEiQLCSV8RFmhKAG5fJ2EvuaC0/I+/4fOiSCj
I/8so85zAnIQNEs3iJzpCUAZPoKLvyov0AtXQX7dbnpAM0kji1aTGTOg6dU4e+YC
tOr7UPBPWEOHJ7gKdVfGWjlq5gd+6KfOZJNz5gC/rbYX47xSs2EVjaRAzzlV6z06
1g9U7parwhFLeSdzgD3cnYBpURcD/DYSt6OKBwltR2R+wB2qytVpCKnx0UtPYFSi
ilsI1yEqf8HRWal+Vjza+Ta04p45tUKPQANGjLLZrbHjQUVB5OHHyE0kDvabCoYf
IE0vRWxVfeXSXfW4Hh68/TNOvmGwT9XFJdvsXOV+6UTkiQyhY/OSwgEdmRHk+RsC
FfXV91Vc7HtFPnfcm1dmrnZVRU922wD8goDtdmB41mY/7N/Noqa2lKx6P0O8Df20
W5XClmgTAjQMwOhNWO4UamWypclPJxbsM9JD0dOozyqRm9OJw6xHIWLTonJHcO6U
Pr1ypn+Po4qI+07r8HGC5+dkw8j9FK9PlEQ7+w46bQr4BKG7fNwud/5tEQO482ZH
xvP1OeXOOe+1dabX8/fAHWh44c4gVvO7/XfRDNyEiy+eban08YPo6tO7MW4OZiKB
G1x+P435rFxQkxHITJ3BqNHBR4KsUIs/BSzmuhBKRNPUuKjC08MYgienfYNPWxTC
rqAcDYrqos4ritt8Afsk3cC2ED1foq8lz2uy1hcV41ne746JRiSaVrfy5tz/RGqQ
gOe+yrzoASDi7o7A41qPKv5cr8A70we6pANBG4XayoaJrTjkjg8umc7OGQZ7gy1q
BCBBaBisuCzuD/qR2fWXmbjOGYFS+CzZZ8yPTVcXW7EvOXVnZvb9ymnS0Hb3Dxef
HGqHIYEzm+5/ovnaOePwQEk3kyKH7LdlVVM1vGaNIloFVxmsmyyUw4mhpGrxsAga
N5oD7enTnahyGMlJUgbbDAiTw0i1VCSn8nmKdi5mNqGhwcXEJVwICRNFYjO/bT2w
7pUKbztrvOae66QDGWEgdsTri5Nyxa8aS79Wpw/FWizOpzh/ow1AjtL63od/n9CK
jcMSd2byn4IeTkSg4hSrdDDtU2inXVUtiS4MJFZBeHQRBAKWfmNo5xP1kSpuknVh
cHZQPUV9I8/8JFEvYdoHxnuB/RiIv+dh/aHEyxyQ0X+WUlYgCY34otzbU7iyZpmn
LyyWaaEP1Kau2t+y5fVoZ3ilcaDVQk0F5iZ0/NZ4pD98BJUfGe9naOEcNsLOMcWu
xoGy6QHg/4RozOOfCEurV6Q8JQ6ozgn5U2dPdINWNAJknPTU+s0SOqOj7TB50zZT
mwWCxiJfpUIVV1d3XnUnazJpVfdb+AK6hwh/Acn0oFR1g8As8qOQgCVtF9epEcui
m0qee9nbrYHH4X5fSmMW4B4nn7letvL+cmmYZPsMqleu3sV5pYulYzPJJRYuegJI
D1QKrKhWVeQyoWHCz75Tc1iD5zaOBSZ4yFdRnYrnO6hobSeKE2ubm1OFyeGZwMov
KQSAx/OrCUPj3f+7HpMmtdMKxwQ8j1DtlD23bYoLY+Y=
`protect end_protected