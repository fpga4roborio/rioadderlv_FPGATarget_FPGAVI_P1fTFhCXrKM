`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
ddtXksX2+yylW5zu6QL2Lhnb2d1sD00763mmSITNX595NcHTEkwn0zB1Dry37fOW
FufOhVzEJp80NC5qZ/+F0Vk7Ik02dIR0elf3clrjeJRK85K4e3Hoo4xn7YbFUIms
l/8VZSb14+JVGURjfswrIyCUotIzlzVYZ6gzoZwDXIi5gQIBf/gI+KxNXPaKV+PQ
Ufys/12rjO6aI/pPlqSm0hCvftmBcnezN2hk1UeXgOIuKZnogjOsf0iJVX2aOOWE
6pD/psybjbnsNB6kH5uFTA5frkzIzkzl5d9+YDm9OyC+k84E83I/7/j+rk4L2dah
QJOvksSIzN867/4Qt8qYTQ==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="MvBXkzurAa5VTw+1JJ70nePUfoQXBvZOku/SMmg4TwQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
oRtzZL4VJ4iwysPsC8SXYCzXS8Fw2gtZTOskLcDV+1B9Nzn1zTyNtlo6lNICRmmK
ZRVu2BmCc2G+fmzynYlNTnSa7C0Cuel6FYpxCBlOuk3OF2tzAmLAuDyOH3Z1Yjzk
a0aHuoCdIRKv7BrZCdALt03JeUmXKPdOmIlkVGFl8yw=
`protect rights_digest_method = "sha256"
`protect end_toolblock="Jn9CQpRhJt4rnzZPRk+dOpzAubz7omckX1MrFd4p81o="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 16288 )
`protect data_block
gD6l00tciPUa6pDNTk/+t0OO0nC/UTtBwLB41d4inuAUA3i/ALrNyoJVcBnAmEQW
ptbcNp5fxEUJjnOxnedyZEuEBxWRieZFQnkRdF269oNb1hWYZamhEdTD+jSR4C4B
rz+t9d7TPze2/TsziIZ146gMSGnwdZEMGDjgqLuiTjTyajR+a6SJiZg6CrMJvrtR
z2x7iLisKdhPRUilsTJUK5yBwpnbRpC4yTCxXJYhNARzsb2kqp4dvc92PDSEY7uM
7LsQRcWmFDkgkpzMcW7CgWKmld8VlQg3pBBSQDhLWBoYk140QbNH8LXdMaR/2N9e
1wQ5n10Xquk8k14ZASI6lWCIMqWurggBIDdxIoZbGn9twkBlGokw+0NDpFUWCrAf
qtyYm3YqcqXfPsGp15zk6M27LiPAuoGn1HzfKvMaBWkb+TsIzG7wsC4Y8fKKFfp1
3+Ga+kGReuzv5+3ZtqWtSEKnTp3Aaa+WVcjN9sd8lNn2dHgKOSVI3WrG/ZVFfjgm
FRxe9YGY49TrbSM9hh3D0OvtrosUGcH0VHD8d/GVXtd+t0YLNV/DJKDsZ+9lXyKp
jTEvFPe1X6TlS/7nHWCKbmYkhtXU++gpxtuNoQk4uGnAj48aWlLAbNSPUbjN6jFh
J6Xr14WtkGl3fxrORoqgk8CbJz8etLIRhf+YiQiQHlZWWezGnZnfn3+/gP5LUib0
HD6ZOfdq3nFzSH1eivTpqJnzPGUs0afsrnKYwl3gQ8ghnXVUTtPwkhhi6kFUXORZ
z/u7PCRAR2JW2gMkwPOgwgnahmrwysNAXnY4u1SgAmBZeTNmmySX42KIFC+2kjPP
xfousj6RJRwRWI7gSy1bhlf/Xi1pvhp6pV4/5ldFJRZEJWi1vOHiTd20rllm1lrO
MbE7xTAUrzS5Z8BmtU3RmlJrGMLsHXIphQah2b1aWdjv+GqP+qpy1DyjkYrRLPeC
nl8liZf5WBisvyBTvaTr7sMWltA9rCLyhg7N35ASAio8nko20X4n4DLv+wHop8+X
wCfrIJKQOe0kGgIRwwubg9pNJsC6hPHyDogBpE0aquj4WzLmsKCcPehsELG+wdBA
vJiUddE+3xDL0LMLBvQoRf+62NBmJE1QOHylxmKTc9UYcO7hPQYK1aru70AQ2oZb
mVlvSK6v6WiV0ydGti+X9Hq/2TqbtkQKab7z8RyoSr1EmvvUwhfga1dFTw2r2/dp
FZiM+dUA/vmkVArtWEnZtu0c0/A5WyzeMi+cRssbMeYxgQVHCWN+nOpYKi2C9I6g
v7l/nuA/OWBn4tCl1IETQxxgtdq8smHXqpO8WFI/AfD0FZnW+jC6gz0xrw3MeKEK
aTy7SpaMCQ1CAoew2z1kKl+TTPwOQQvYOUd8M1hOG0fdbncFYg3QbEm6y5A5yTkZ
LOotOrojNlDGK+sW+p/2xykc7Bw7muzEj2M/8fBLRyHqz6iiFSgc28IaIv0nO4mt
Z31b0ZlCOwXJ/ECF74kMVTUl3eU1cpSzDYndyprnap6JfAvKcED8/pBLdWi1JOmb
o0gdcztyAEL/qBQI51ewssimgGGqaoaSwhwC3EcU6nzkFExHpKHwlVW4V9gBAaCz
OKh18R2qOWqN3W28IJmLzfKkfpcSM4RA5pQNpSMM37Q595ZPC7msQe0tqqAqhkYJ
s3sO1fJJBaNrtZC6Q7rPvEmUI0oWcByOGJ1vJgF8UgAqVfcJOevOhrpzj6WOUQi0
RyL4o3UCHZODNBqS7vvFUP6Nrfc9NZHz6sfgBfPKW254EQlS1q6UHzsQAFGpYMhi
wrWZIHTZl+OO6Ut2k0cZCO4pfUDAWp+8u1ExNeiBC85qubmoTlcyejfQmhUW7+iQ
oPeekgdiTk5Y5hNgU595aM2U/uOBALmyX04pwJFXw8FplaBPoJIip985HGQpNjQZ
c9ia6y0uOicfqnBvaYUL/X+ZYYoSKuG905c8YkhJNrbeFtsxtoSFDhD7AgQDw8W1
PkFsDaikmQgsk6oKv02LgiOre+D7/wAlPAATrXTh2kqWeQNqFRyhdEuHNTZZXRx0
n2I79JtxiA+003cSf7Y66QzfKJTCS3hgchrrm/pW45uvkOKLrlhRN51n5cWUQZtX
XOvWJkAP/iC06JG4FHr9UwxX6cFuN5WAZrBurmvCGuKSQKBLWsix8tb8jJXsqw+z
8QqFJm5cKlimOdOBAOAmzgzsFXEBjEbYxCLVD4Zkvg3rvOFKsYhx6uJ+1ba7uZKW
KDIUf9Q0Nd/XVwfs4/ljNs4hsm3Og8UMzgpQBub6kubUkSiwnaWIlxKVW57fuPsk
bYYjU5IOtnK/NauzIId2CKbVKt4L9dkt2OsHkFpxoMMDlGp6cP4wNb6VRZCc9l18
1g6P0O2TguEGB/nDNoLfSYZ377g67ofcuG5s8rCaeuSfIetBFVPArcb1B9xQWrua
PfQpTaiGHy7MsR1i1J9ItshibQrtBYQMHFDivM+XzrZn3mbVun6B6GsuimOJQG4N
e+vWZzBNUnIiozDwk+NsHtefd85fFNywESFF7ABV6MSWMFT5jCObJC/EAw/kKtlS
LlWKXUG2QhDMPzo1+e7ivbOzHnuIYyZcqXLYymbob36BLM5Zo44N6OppIo6n3Z8x
ga/0X1zGB/gg+dctzpdKJkkJby5Y6LeOpS646xnAZJHgtNsZXOKvrljetQxl/U/u
Aew+QHkqBvvoDv2C/4xgN54NTiGZ/wHpJeSkKeZm/gTz+Kfm7G30aVVziVT3Ilpb
1fRgR0eeNtXvHZzSypilb1NAE9+3HjLfNFFrcKh30+F5lZ2v9gyTgzKpjpqM0JxW
s5SgcIN7StCdSfoEIg2NJA55NBPsXR3881cIHgrOBQhAwRHmPnfS6oWYj7UhVadV
BPYS5F55cotpLvSu5WueBDtlUkc8NYknGZErvon9esSjWjbPy4Q5U6Zq89DpLWNs
X+B7Wlj7+eCJE/R9PMvjn4nkLKB5jUlgRTydKNSHSXd2XVhpKEvqu8hpYLInIEyl
hfgIMU9vVtzaFpgKx6c+A4BLiEEItFE48atd401JmFof0hQTxn7BdWVcP6TUDuNa
Tq6fDAzPbX0mKO9N9HLa183U//Qo8LnVGYfu3iS1I5mUp45t5yNk1xyIkaRZlsD6
W/2nio6YK1y1qaniwnIDXvFA/wtzw5BnAIeh6pkCi6vmW38FtHCB+h/AAYeUuFIs
vzGecoW4XI+OActYVTW0YqqscY8guN3jmZfCUqD6+5bZa3r/rOhM0haOGppuIwin
MKqffNY/uEPihAUFuqmTSUM5HZWawqD5KOE9W+i0DGLQVz39zy+Ki4JmxkvFf2Zp
4njdnkjcZSZfhTJ8WIYdzrO+IXR/qZHqmkMz+jmz9wKUMaOgH5gI4LU/yQovXAiL
JCrKWPGlO1zZZr6f2FneJ0UNTN8pxgwRNG8d/tGtM5UUgAYSU51WTf3kpICPI8Vu
sK1vzPjR3pNzmzZjCikl8mL7f13lA/JUBcRWMoTDjt7HB89msjOF9uB9Zk7OCtFo
zRSGJo6bcGElyYkQPQHGpG5vpJRK5hr/s8Y8eM3KMqlrgiiPAeTro+AI+1dpH8vP
gkkQLvelygWeCZVIsTekOquhoWfWqcwqvXwtzEgsh5r8/QMxYx8YkFz7AuLQHmKB
k6WCF8yON4AM3jSpgS+IdJ8M9qV49L5KdVmeCIxEW6h5jaqq2R3PdGCJvh1P73sq
xo/hv4rKoTIqqZ4dRuZZnaFwY+3+RAkpxw41q4VCdK/pMHHQ52f/S6yTM85k1bZY
sM1u7b8nc7jjKQN34WSG2IZxeWXLt4teiGplxGEQm/HA1iCTSFbhC5J6jiZf7m8y
HHOQucoS1dxuInMYbOVepK7r1ZjK/tVGZXe3lJKVuKIdetH5fgPrTsWg7iIRuM3d
UVGQW6/Gc7dTX5pFnTDQZOhcVXh3IfugNfodBEqzCshAAOTSjyySVDToGeMZYkFM
9+aNtO43YX0xhAsMr7Mi3SZhV1pFhi6EeQF4dqslJwYjiFOogqjpJ0FkJH7XrP1J
Ba7uVQ7LiOUpMsan8lXCwtK1Fs1/BT29Cf0rsMjx+I1nQ/dQYH3ox0Xg2txPwWbz
ffVN4JYMUn4eGH14PJX4fgIvvqPA9VBQR2GVeyvCp2XR7GCnjZKEGegvuBfZQFZz
cyo5IkEgd8Ug0lVRRf2tr3NpCZvHm+RgIoIy15rkwpaTmZUYBsYwZoPYujiFVZqP
kw0xuP94TbUpwpH0XFhcQ7lYBT+8BwvDeQaH8XJegYKHGa5tKPfpTJDQEsbs5Ixj
Rqd+nD2QjyZPGuZrj4+v0JrNzbMlzE+da/tcC6sVMmFUfUuzlAPh25+rDl4lEssW
pUF6Z/Y++WA805cm69s25MXpp9x/kCzcn0ZK22vnlg3VGlYKI8Ic2hSYKIcmtwle
H1bjbag3cIKr3ifEkCNRMFYlCixneYC7y/MLKPnu8fa7006vj+JtYKY23dS29gKf
HOiX61Gg5IraceCvxRyGFQdEr2u5zzbjbdNCni9Brn4KlX8h3bIW/yA7a6Oy008c
Cw41uMJ3HupXpvhNf4fAR9B/CK7i4GV98ZNeGOOArSOcrie+zST+ASQXlM2v35qz
zu1vPMqHcK7iKyFFu0rUMTgBYaciaz6NZdyqoOvdHKQGHGiO4/vqaQ+LTKnnD642
fKjxM0GnV0M49BUN2zHfHhKHd1XeblT8xxhM8DvP8YT814vDjFbXfmtlW+KjoKJF
DI7kDifUg9X86f++dCp86Kddx6+Xyvke6So8UtCDmwHlKpafv4KBOLefP0ybHvUB
2qKHNlk4Yj2OCtAz/bOvPk6EKyqutUV5NbfyX/U2vPvXCKN7+QEO62CITKmFNeL/
EFE3fZPHsuQRNdkTRy9FmAsfPM2whuGxmJ2TSYcKsXu//gBRab6YXF8X9bilbKIr
Htq+Slu+IG3VH244lQh4UKK9mlUl86x7im+VliK1vPsp963wtvgyLqLZ+qj7rBxS
I7n3uYcPSPX9gVUsaEcpBApRlkm8penZdxjr9pXQQldbKiDGzDOQsj3Lhl1lweLs
BGk7eId/2SYW0oBc4ZeE1jQ84aQGWwQEfMTZYcA+ocFexMO2gpeCKvRggJQ13OC1
GtZ9qvTO1R79No6YRO3ds6lBmX5w1aIzV3RSrGcBiwK8qaElfI6NlAcwU9dbYfg7
+9E9JS8qNQQHAccDVXGiMi4XYzeKAhI4MIf2Nvu5d5rm1EAtpFShX1nkHmQYARym
BV01DuL8hg1SF372UQG+9FoHEp8wZdwRUSO5WHPfn5Azp3tphoyhqxwxt3telehl
YxUsQSsVgjXH6XcWFms++3JYP/6PBANOkf/2/zDGggoHxQHotwRhvlQGdrC7XKBF
CBCHpqzEVlsK2TptfP6Pm10PFPBt/oPYpBd0+HSG+zRJkSBWmguz1Y/GTQY3ttdo
Kzz5wq0FJMfHz34pliNSlSeFC9aywNr2YLXOtncOVN1+/fak9HTPVR8Pkr1y3Qkb
CHt4H0fZIvV7uieaveyl9ZkikKHGUFTxI+4Hnubb1T8vv98uENjdVRvP9FbIet/t
lIc7bocYmzY3S5YBteJC88NVYyvCapszG0CU7FJYAbPdWcZX6pDBl9ilpdRDSTGH
uxCys6D8Zk/nZ1fSq1UVaDSQ97+Ar5fYBHpCGoTScFx2hMI/6o0CjnfHx3BpmkEc
1rPjrJ8R1HXdV5TqMg92Vzl4uf557u/p7ylt+rkeh4udpeWH4GMqYuhi72V7I2+/
D4U9SvxjhirtWdv5DU0z5WTIG0Akzx5S/c+CmPfwQlFNUzYmRhGwUhN4vMOnRNeb
a5p7rUa1cKv04EiCi0yIDhn94ITbzW6rh3Nogp+phKqWgLMCGEPXBnt9amdvCb56
MO8BtgXvEIrFAeKYPUY7zxSP+btPB+5ooUq7KS0R9iNr57NPPfpCbsZvEgE/eSap
/ARLcIILqt52FkfYCeV+qGjrp9zLHxCgMOFURyJWFxZxSJRW9QFcNpuTAkjPUs2W
oqvQRj22Xwd7ncXFBReRzdsLn7QXdRDTis/zLuYiVCRkLeNLu2vy+UC9ZF2ySxA6
/QzNeRKpEBT9W0R6AqrjlHJ8vJdeIQvrjT2PjEIgEhQk4jz4IITNUk5BvUHsKCa4
MRLG3PhK2yyKpVN+Q/VgkOXdsGm1R936XBrzED5U+OReSmnDg2H5LXxRKHCu/dN4
VoFQX86EI2w+F8GOTiV3oYmVa5gg+9fdf8hW1m9iRjes91PxvqN4rJ1zVy93E2BT
sl51eS+73u0saGCDiQRQNCo58hcnyz/wUiSOwBHq7g3ezPFACdVWgbh8PD8P1j5u
IPpFoM20M6yw0efBD7Mi7HOyhRLvAmBPDjqvqRNRZZuQr/jNA2wmjgzlK9HIfiGX
9gmgry8fZqw4O+kZip9k/lFIqBAc6JmUQB3ULn/8B2kfe+T+zGQ1OrZPk4EGbR6e
8/+MJUq+1P4rmAVraeHsqNpkrWjIAkB0KBKeI6MK4QHdhXMY5VIj9OEH7Z8EiXDf
D2uWLd/rv7JWDi97y1aBQczgnkGy7lnsP01JM4AzI1YBhReJzza34xRiEoyPh70J
D1uA+CMwSH4ibmI8dcjUNir2L2NTsXPvTXFR0GHaDaQfkA0f9OcAKnwKL7K5Dqm2
jRIFTUO5/pSBLPfAOksv/GH+LtfeYPqsZaF3Ga+Xw+Vpc6dHSQXWEM1VjLKmTamQ
LC+mH2gc1QHB6Gn1RZg6wB3P3nSdDA6OPlpy/4UJiv7dIaN5qRA1l8W3oJ6gU1U9
Y4x1I1bM+3heOpAtyXvnu12oxk6k5WZ5z7MNsxVK74BQVJQf+fW1d/42h+bhSX1N
edj7zraZDyoH3gFIFWoKSn1vPj+zzzy18R4LXPlKh2IZ3T3quUe+9sdjTurzQPog
/BEZ70lljbI7cnJ62jNq/5mLWH8zvJmuU5bAQEWzlPa1XfEq+xtFc3QoNbSriveH
vwyhUCeNtyNj49ez1SxcQRFlAsdehTVsHThL13EfGsvIJoh3K81ltMB/VhTR9Tuj
HXk29q3BMkECLB2/I2Dkbt1sZr2iXxSzcf2gIlgBYovCxIXLyVkeRg7AeljtPyeO
UKekl0Xmuc7IBtWZt11gPXy0L52zjzASx2MeKbajLv01yM04JX7tqEaXGaIdDGrg
kk+rdRFLFH0Eh2m5xK3GBvFG55MzWauwNg00VipzvGTk6QQyh+fxJxEV9Fy3VNom
dbMryPDloS87h+9BWVVKrTspNGPvz1TIKUK29ykgvBq91afTdDk03zzM5DbRKQXf
KVINVUIKBflsEauZnFRZQUy9uW4lRq3UHt2OqONX6dqiMKWTtQDrlgt5KAw/y+qz
Lu8kLaHsE44HGvLtAMCoUXjjvxXGUhYE5y1bWZXwvjY2dvrB3E1DecVwoxwsuvGr
NeUYdHNDY0nCtJTFBagVpsy9D7CtI49OKr4wDPi2KX2zO7SL/DYhXXEiKcTVDLCN
rb3QUaCWd1VJVFb3LqQ2g5y15yU1bXKUtjq5SM+E0QOrzCFd5SlsxMOyeIVFiYQI
5PZIf6siSGnsyXje7FZrPvXJ50AyspdzQ/qvr2Ht1tS0hEE/3Q1twoS15hyvUMb8
jFrBVIPp3Jnab3VVTE9VlPi8prkXE014fhXDx+Cx1sFnMgTLzZTwAtNrzxgTTC58
X/9NCC2yzgsn9DxhUxmEQ6P1BqGirQfk23kO4K5Uw4WL8raZDz8lEVbVK1KDuGxS
Yl/pTQe+fkTOFK3S/PdKYnqHxP9/QHRpWssKHwl6ysJ+nfcB+SSFDPJ2w8V64T6o
goO31ZQvjoBHsTkpl91cKOILcwxmSNl9FmdDLxjgF5AK+fSdU0MBoKDutQ//Qk0a
lzZ2EwxeXyDH0WKQM7caQnWDX8ErO9pDst3VXjZb1xJmQ8cTOWV+32u0jBnlzhrl
kwtoz2GOpxzZhFAG0Quc8BfCUOkBvRM/GLh9xclmnKS1vyyB3qp4jk1tJ1ceyES7
WB/qQHQ49Gkpw/FREvhlTjBOQpXdmD9mplPdgNLyoatqGQhO6xbpgsnSgI1oOvoH
kc7Oavw0MPAO4r1AjiJKynI1revRPFjhI+XKG3zhdz3gTVbB7iqcEaQBFIyYA1jN
+L2hmJSP8jsGFt7VYwNCLsF6CRCO5NZKORM5MIhdmmiwtFr3LAEnRfuQLXgm39Qt
5N6F9k2Nclj1Q+1BgQAp6dxRspixce1p/FOIpocdcuyjYS/NwJob/pLVA0u3gLjs
AvxLiOMygrAEo2klXvvnZJo3UYXO4y21CUTCNmt+3as8nbTmvdCvx6iACtJHM3M+
rjne8m6JNBfDIxROSrzcRw91vPfstgtX/vgPjfB7GSVrmlbfjJE2XDDVnhR9Wg8W
2GnqD9Mv/kKV1jiPcYsgSj5FypUVDo6kLRJ6Jb/UhPHEdwA659CyGPvauh02ZKWb
eBLXbTeR2Dfbg2CTyms6UaII6AT6ZbrttMAbZdcVFZcmJiHs0XDbZkdc+mHeVZGN
YXCovvFukI0nITMq3n3A026TjIOPqlvxvTPa5XRg1UyBiK/g0RK38AWfiUxfXgKs
46YgI4LAjJ+Qt5PVQWuzcJfo9jQtt61z1vlxK+CLfMcKryd90IcMt0/DrXaZxz72
O1BEbvmOJnBSHEIkZSHyVH+obyTvWBRC875rpqhhUPRHdJpRXDjjCNOFsK2pGutI
lDCPUAJHrEjlRrmvnaPtITHAMIUkEdgzu2jJ2nEZgtla+d7Qyg3hyMfvbJMRDD/E
FPUbABNXLpIQru0n/dHCqnudRkqqlSfeS+Q27gWPSNjNXn+p6nk2iXjPw7FGQOAP
kse05w1oN/KFxGYTR96qAAUZx0RGHVb0vkbymYO4FBurXivb4NYNu/Y6qntvZkma
K23LVsT+PQfyA0WKOdGB55bR99YW6D5/wEu5DiLdMDo/JUyRA6GXfF7tLKk8DNJ5
HKmCDiu0Xpi2LqnHDsHg5d2iQFkGdC0WYhu7pF7ZrunrkNCJfn4W12SZCiRQwORY
BN2yh/Y7su0FY4rTMQy7IsiJGz2KMUH1aDLOZGPWiMmOuP3agqhGWeDjRwYuyV9d
Oh1DRrc8joYtDxAdSmZYCN5nT+dle5kCg22QZP4S/Ot1OtyLV6KNVH3Azkx77jtC
fPqNDlc+SSmWXecO1Olmz4PFRl2Nwe1kMNWXCYAeenWjhT1kWc7B68/QgAekFpwR
t6NIl/rEp9pf131rYsGWqznWY5AGYSowbZF5o0p6Dm36zjzj7VVx6VGUkRIjl9Y/
vjnxLnY8WqmUtuSLXD1/B381TEBzzne9P0t66cEkw02TFg6UvZkVm7XVePh3XdHq
iyxczGhNsPQx1JrozoOlpSjOJAnX0ookxR4CVniOewpMAbf/K51xedeDO6rgDL7k
tlRF3ufFlHbgsSXS851RhkEo4lMSYwtnuvUiicxB53ncXmemUMsnN5PrNdavwnSm
86q0Srxsy2tz0OHIA/z4GwKjHKmPEGc/wueWaICF28EAg/WE8ISj+pRgJ5nOcmpu
UkcrLz01lUJ97GVuEEXhStfp2oTB4bn4yhUpBxaVRHzJS6CELUSd3ltQBkty6NRP
xBFwLQ2zHyftNy9T3m2Rspqy39c38R48yGceExXWx5IM4kAX7zOBBFc8OvtCxuEC
1xL+6N8BPb9Yl0U8I5iYUQoc8JPiJzLvas2djBqRfCE3I19vYXNEMjCZIvTDpRsr
muN++qHrF8JC2b7Qs+tUIEl5Z41gQ5ajwkeUI5j1rp92ZvgPeeMmT0OOp3vZvSJh
d9EE1DdBbVkCylQNmuC774Gea+50eef+bpxm3LGxC09Iguax5IX82QL5+0ffQadu
E8BoMxwnB/h/KILoVNKK2i/emfbJ0FFZb4pa/JiTtjSeRrQuGJX82EnDMKxqUkZu
pzlafQ9w5zO+zSX5Gul97ifwAiSd7dS/WbrwDtsF7iK5KIegcsVEGVlWyuPkNIzq
CV3pGAqOytXRWF52CZAiRMo8nnWch+hLc29BiGstpO0uXw1arCGWT3ig7hr3bwqL
lq9Pmg4GxMxRjBnMqNqRHYWb9Pt13EKGw+IkPFlUCZ5WzmFbfvDQ4Fkm+8CsP95+
Drvo7bif46LEFo1VxLhx+hpsENoc54WNQlem35PFe/pk8JvFE3THwNXjd2xoz4mk
OSW6Qa/u4tIrXvrMuH6KZufaX3Yf36HthVCEzvMV7mPRjyqyTw2O8pgZRHzo1k2o
VY3ycXTmtYx5tR7U6vct4fzrSA3CHzfZZ+Ab1cR3/X7Kas4iFOejj/49/Jk+zb1A
6zl90K9e+IrDK/Ax8o/9BiEY5ksJ8yq1YCY8p/aRzaXNd3acu61ebc3Vqx9rbtmx
4yiqNL+ufz1njaysBeQaTaSlu22ry9rxiIwDFPt3jdCJ6Xu/qkUR8/kp5h8ElQ1M
UcLV5Qf2syZNklMMNM9OBEdj2gzL1Bxhnf/WKxNialpVS65dDQKtae9+rtfZv7oO
Jz7FMfn8GYhg0IQn38L8W/DKfkEWiCLrawOLZ+3+XJuIRY4Tj+ISkLMuR/+uPXEn
/zTvl/XWQeKRSlHJ5rw9tqMavihPkaZme6KXISXAfpwCxfRM+sfx727y7nvSkDWL
NL19Y6yp7XA16flvEKCAuKVL+HmQzdILzM3m6/hWJdkboz3jcfQnk5tmFqeMJvWI
z4ald9WqW8q+087FIVMReSVr+CMfk3KkbON3TceA3TTL86gHWBKpJXj1mvWznGj0
keGf38fE0IJGdlKAjCu0QleN33C3Lu66v9LqdEMXIAus8d0MAVOaNkK4EARTzvGu
TKFLQSpzKkar8CN+tJaxPS64LPpn6F3MkDXaZtfbeKwy7zn8FLz/pSSQgTqcF6Q5
vvyx0ryQtr3O6rZGq5LHx/dmJLtfj8kQ9bl3W7SCjuiLPOnz2vjJuc8rwGJRBT6M
Rv4S3lku4RrB1UtF8KA0tjn7Y4Do0TRLZX8gjlDPDYa2V8+yoMot6YpviWZW0y0d
iz5OACwLPKNYab1Ee0Bm02GZCIoVmanrEj6Zvsn6QXGYZXZAaFxA+yt85bZkRNGH
qaa1XfTxruLR+Tnf2TGdPxZcHkKTu41zTTqDKMae+pFrfKTa7fPvUglGub05PXfD
m8SF22hvc7LmkxRDYmpPMcrYpcQoAXUApbeyF2gPK41iHO86TM3nggppyPTCYqkt
UJcKqCq94F04hYjS+W4Qu46gNLCV+ZfqcYU6nLn09I1taLq2uYVx/Jj/coRmsm/X
P9Dv6HWccCj2YV5m/P4YrVc6jLZse0xK8UzYJoAxid+5qX7Xq/0dlNZQPWpiKiHe
yWfwbNYGJAFSJmat33oEV//UaZFyl7AF5YowHV1AP6NNboVTQLSeCBtgW0JGcPHK
dEwCmeXjFqDJlYLqyht5DA8GuMoQN9AV5IllM7i+hPvBJ8yIdJhXl/lB8vpMT5+s
qirSJCLM2aeelo4cuh7sPi8P3WJ9Sn5Z5b9B9ylNKccUsWiehx/Cha2pchfMAalY
YrdOStCwWqd5sZUAYzaWcEfhL+JzplBI+a14mAlTX0NjxEr8JffjU/Cy5eRCloV8
Zt+xklfZJu97XNAK/Uso6qzJw/KgTTuViGpRwT7KaSTHnuGLs8YJ9VCwvfsMLfkl
cCdVxYWYMnAX18rCk/c1HJwLe1Ge4w6uv1EMrXwfgquupvXdzOKJ07jOPaAn/i+s
E/wS+eH+qZ1Ks+jaYeYnSG5RE9cLimw0DP+3JhUYLeF2ZSEs7xgLPsPLyf2fcS4g
O/AZofvRWfL98lXrjLH0anAobyDrnYKBYvkriGrMBnOo+1nzoKr3+hpvMbLhWw4w
xQ628eP0LB/LihDjEY7CyRrP/9eh9laddvYb8rKGH4KglVtUQFNrIxxrjtVpA9vF
9mykdAypuM67qFtJuI2BUxPzyOt0/2yK7mjBPwWXcR6eQ11/1lN9LiF164o53fSA
YPJLkE9QkcViwM8ljV59l3g43ssmW31nGrJ0sUYc1kiV2bnqFGFk3Sfvii0/uLES
YeISp83yqJW9pFq1x4a6PELclKtHrOYv2jvOKjbUTWeCUJ82Uc2Wkw1Htjk4i9Mm
IqFOFtgVZ+7RJ4q/+lWArF2lNS3l3AEQKdSItz8gJednRriuBD8GO9fcOENpnbOR
lKbnDtbUn0s9T91ck6oNmatQ1S0+iJFBFCaLCCFER9DTfLxhALo4Pxav9TD1W8d0
mqSAAEQKy+VtFyRbanC0GmAd/Opje+iL7cYcLWE6WN2F7DylVZjkO1VrCQ3ein6Z
KRWupefgtvP7GtOOBCZZk5Id1+dTlNVWXPMfBrIIPp7/w0dmTjLDiR95tg7YtFTQ
HwaQ5Fl7vxpUh3V2HMNyrt31macGI8rd+fVjSCLzYAIuRH4/aJQFlnXMYXlFtJ1h
OetouXb+km+v9pOx5oQZnjLwgidPCrH7qmIx91g0kuZXe3OHpRaSkC9Dpqxq1Ihz
08qYCZc1tR8ic10fZEJ7dU7wrMhbqmgBAnPl0CZt7JCfn1TKmrgR2xFlT+o98A/0
WMOvJTfpVnPdFinJGLrNx0M8xazUEVwWXI1/usoZb2LgIGDXRigLmhxvx5EDvaoK
MYLG6sFcBtxil+Os5H07BAQmyi1mWjJDR1i9dDeXdrjjOiQ1aU9AZnZxRrF+5dFo
D587TJ55nb0/LxTY1ukMhiv8OLicWk8sk+C7YQKZKw/gA94/IVeuC4LVesTGLBTC
AoTzPCjyxwHQlSMAXOPFX75RicHtWP2nR6tiSxtD3usJXQVPvEZC+yj3+FpwOlKT
b7hZS9IdSzmh2zM6zbtNoMa+Diy6/CrVi6zzrz8eeloY+2qWfIqASIoGIYtko5OH
Jto0ZLj88Z3KMn6zNH7yLkDMHPJAYkvmZUP1U8oDOom2uNzriiB5WBF/KWCVIsvS
cTu2LZrAoSPIw4kqNvS+KTk/qmlGlHZwpclJPizeFV566O9QLffAUZ7Fh99j9Hz0
7pF8w+tA/xfjqGj4la8/ZLePZEGiqhaB3JG3+kXHq3B1qCpNE8ZB3kF+M14nuV3/
gJOFY9JMaqmPhKjT5kPedMS9V2YAx++ANkR/QB61pFpwkYbJ4eyPhNH+ZNJVPHzH
9Vitw3gsVSBrFH6Pk9czhxoDVtz7kVmjCdx8QCZppc/dqVOabpLo8MKad5W8vmn3
4Xew+mb1cCYCBuLgK9FUDJUe9q944K9FFVpbp9tLrG6478JlGNMBl7KiGCvKB6oa
SSVk287PpyVT5SnHmCQtOfLHc1xPem7U6hpuTrUFRZZMqIL8l8udr9IQ3Tcj49f9
67oWt1x7qCImCopaft1OxL3LAVXSL/PMXpMfk4XS3idWYbx9SBOVlj3NzLCEGDI8
SxIu/8PREpLFBR3tefuIAI/gN97W7+x9iB6O1MigmwiETUPEuAWVXi+JXjc6DYo6
rluKvDiyD1iSCbLM+j0k9+BUQoYtJmQH7WILRZDWd5sH5eWcAqIeIqxiXhuyb59X
LFei2OaCKThksXbUqhog84aQQE8O1yMATsMOd+lC3crHugoMkK51N+nrQYRWYf/A
YD9DYLxTaRikuBWtWEUCXAIQl5diip48wv3uWVG40n+Zg34vDSeC2qnFkr9pzHZP
/Vmd3UwwAV2IHQ8Qn6jKG0nGVyZzv+cSWT3xe7Bu3IjremCXtdDXr0GBoPsAZC/Q
Ppyi7u83pzWLcRSirWwLro0hpVnJqQcZOos1nS7cVbiaGnoUS9ADr23YjMxGb4NP
nGUDu68qMG1syFEZU4VEfLfc6VTIq1hWJGFQsKVsgkHqnzZuAhZqq46tZBZQIiaH
xnf+WdTh5cVJ181kEm/qijUA/9Wo8SmDy/uL9GbqT4h8/mmP0NmXLPzd2bVwD9FM
7VmePdNKzvxUmYcbJNVWny15R+jCIffgdiKLrfkdxOyfMHeRGS7R14bqnsnicRvX
CMoDdTdOIzFfQVVae4KBr3EmU7HK1K399+FrHs0bAnnB7p0UBmur629gP/YMXeqa
UGBz9HqTRRvw2jPO8QaIpN66pWTEam4H4Iq+4NVWPkfTzaVgmZJgcvYQom9YJMml
+4GF11z7j7/vTeT77uso5Z4qEHJ4T/gweM5ayVhk+IiF9QaHSDE+jVvBJG8EnCTs
/q23Q1G04iT7j+W3lA0Pjgm6XS1Zkw3FEft5U/qqXV/2Y0ee2DrW7lExwO8z0bqf
8E4EhRNuuBSHT0OuEyOCZgNUpe97NJvDavdiYqlTFD9gZ7Vpn/Y/hF+DmUXsIJKp
fjpMVlsGmpoS7fUtJtILWvQnS0a7iSRfbQY/zVh7Fld8yJTsDo4IR85g83zTPh1F
kiYZJhXMtJpQeT/ikK210B8ZSM4x4DjTfx5qjo7CR876ch4OsQCnEpFLYBTKm3io
sUyu9Btdu+vzSlqTIHT5Nd92VFDTSErds/OiNJDXJHov2dyheJ+XgzDL5BiBXOvI
gLCiypy88blTGlVCmP3DH5PH/6Dah8FXZSwx8IBlL3tpjZfo4YgJPJRXNGYOfCx3
yJ9yUb3hJbaiLw2TeddYcwceizoVHG+Ytw2bgDXBNrcCB1zmP1mHqyCwJFtm3bST
qBbriHig+CkQVoTy92DeTUmWf1XZxpQunRDVtrpsa73l3xb3axqC2I5h0vwDgt0H
/DRRZvwXpHk4KnkhQtCpksEnKZJuhFQomdrNMikj8yyLdBD6hia0PyoZ029FvecL
FA2cfE8NAERNh8PuRYaEB+E6QbMind4RDwrl26dg7M6d86WMfcIGsFxa5xwMB4CV
mOo9AuNIvKzpFZPKbr3qMOO2Z1esLBbKraak+FE3XG/uVw9vxjxRuxQhykDHYksc
pdOV9Wrn04vzZAmVpDBiT3SKZGCVVwbajrpqLpdcgDe09DzvR/qpSH17iED6FK8c
Azak09ASOz9+fpTloyMxdVMyzypE5HTHW2aI/JTP3gu+JONnvPe8ckswZ/MuOWa9
qNureWMsmCuzWfdEkeYv5RDnci+QohydnJghZdDvwEXFcWrsN1DBEPCG6CPYUrOT
zhHDfKKF2odMAAHHtw+gMk1Bstxw5H0Q60YcNY1N7mdmsQHxsyh3YiozWi3z5j0Q
0fONbRosasvHtent5K7q8hCgdW4Kd5tg3qIZGVaMzHz1EeqYVwL9VAznSHeyg2ST
1mlLKMZX33vlmyii05hOqLQfu76FId/iLVrSjdRkk4dhxJUPYjtLjgQOEEmSS983
x/X+xNeUFsi+PevFD92l7cTfkiK8kzpeQrbumFzWmAY/xkwdRuW/HXmvUvpERwMG
gEfGgDCyzjKKza7496x6tdlxwnPBa9RQi24FYAkbhyN8m3lQto7ciKih7DjTMOe0
I+2DUOfWR2JgsLRt5SU9t5sLzqsyfnLM6aCFKa0ILi2gtBX1sBBy/dtus8GrQcFn
kyDpHQ9rGHj3jO7ERyi0YAWX4o8BoPChHRongvo80XqBnr/FkGwXpB97csWIJ+dS
KdjF4ntfFG0Guhh434pKuLiu12ODVmZ0eXH5BOgmfOZ9GlRVwqRDRHX+XBT3Hp9U
YEFPAGAbfi+t/w54eVbbmbz33+J3EClNoT8UwAjgwHtswMfhsPb15lHH46snLoDW
Vm3zdCQdhCizpixW3SE4RjY2ZgvuUt4HX814cMR/CywhZjWW/w4KEZmxvvPOkch4
rQi3pAVRr6GGCnBayf8C87z2B0e7Vy6kJn8eK1iDd7CZuVjlbt0Vj9e9mjoiRW1w
/M2leqXTZOq7ElcAh8U3L+BjxG47lYWSudIyFuLAO1o7wwaodkYnFJES0TdDGJep
kexrZZScTYiXQnGWAQX255YVvXuU9IknsugulljlEocOb1RNMtXt9CqAI/J6MhMt
5pbCgJGGX+4r8wvnITZ0CzUb+Y1em/VqMeUCDqtPZrJWp/b5KToWEGiTCMLST8RK
5NQbX43dAz7Y5z7/exR0vnAO3cxOJFXSjrUdhUC1xEU1O17y5iCgi9OT7niLoDsR
ySnUZxHU8IZlOZ+y3n0wfntMaKww8qYO2OnpdIELxqr/IYCohChN5MR61bxs+GSn
gsBFTzJ0mDvTDhR5U36/965sbUjRilt+ZhE7DVBckscRLm+XI8gRfRipwcTqcpl1
tYYn7mD4aqDrCPSxHwKwppMIJASuEne82ZnzqV3LuqCZzg/WOTRJjo4K3bb77mig
JIcj1vksHlbM535a57oAx+yulPO7bgIMYNFCwVbND6VFn2Jcs8yUx1e+GRPKhaj9
EAhrjKGJWL16nLXYrGwd4ff2k8cVsYxZ5SATT8TKT1hIIErs6NoqAoNn/JLmV/w2
ugdJKRAcET4rGtYzboEG8nuFiCDgb4azwYQSyY9caIzr0aqI5FZ29gK57wLsn4NV
/Mqs1ISDWMwpOrwG0QFhja8ALAATP9m3YLfphOVkfIdILzKarvpee3d4/+S0AcMt
UwALz8z1oWSuugfYXxy3ItJyysYuvwCaW72L1QsWo3lW0OkbD3bHTwUwWg8+see1
uZj7VtpUJcNBArgPlnzNEavHo2IfnhkkHhj+cqwEu33VaGQuW0z5Jrch5mu9sHsI
vJW5xsD7feCkunoCdCfLMA/k1BA3sV8tOmq/GHfTp1VzACr4YDnQS+Ps23biO8Ty
riK261mE4PLZ9tydYtrQYbOOaf+1cpw56Kz3P6FKFJ5QrRAdgXZt0rCO4Mt9/WaI
TnC7xAF6GmfSp8CEY51Yz+Pd3ojutEnkBSMl+7yulMSR537/+L+eBV3i797Kd6P7
53vOLdsAkzEg6B6HJpcunHD28EnHzbDiET+/Z1+SkSA9Yxs6isfoNG0QbHAUGyze
r2NvzauD+E1xjyFx46FaPSwaJkj2Oxf0xYi0cinzkO5ukitqxwPeUOm1h8HjmjhP
HVUQbNiFz4FLOi27yXtOyuXjuVFEUE8VDtpdpulyPoTJdYuSvktn/JeIazjQ0a41
hhgp1DoUHYFT7pqDVsVrLDa1V8pvEEkAGAi9ndBLlkL8kNHtIpr8Zdljvjw+wW8b
jGmrKiwiaAwm7xrFDeiOiqN0Q9O/HQ87uzmRKv4rhlV74N4QSWQASYscwGSevrai
rPpKzZ8hsdC41A4R+MuCrkEx7V1j63FnERX3UIMb+Hu52HJH/VtYPAkTc6bceQHc
u8Xqr3soQfGGIdRFb/3hreq8/JOo5JAxW8fN7uy0+xPZvbBN03qNUxX+wW7CRTin
/GSZCCn8O/yHfPs3WabJPmq0XzVUqqVyOhmlJBPoi8eklVEp4597fgUujB5aO10p
6cJZYEk6YrOaOy4JoseQNZm5vgLqexflwO+fhkbpXEU3MyILYDvGHyF+YYHgiEd7
weMzXXSYpfsosuKF+tGRPBLQr3/Wiv7bUHaMR5HwFhN9vrXdXd4G9qIRlt34bPb0
4fKySz24W11UnvC4gYQhmULrZtm2BUWBh1U09hidtq5RLf146BV1xvAaiBAOYZEQ
VOIWawMxCNl94YIGknjK8UaA6u+5L6LSLjsENUZnlzDRhILOt+TtgPi7P7gEGq1l
FKhokcQDvQiP57drjRPjJVpaXsPsfSpyxT3TSmP2MmrLfdEveXw/NJ8AqQufJuIy
4U5/I7wdwH7K0JsIS0h9eKasQp3q6HYGoRYo2tvfia66kIjIaGABr+QOQma29ssl
e6hmR5U4FifY6ZHHjeIted4aaHV38TqjrifZGA5IIhnHHz8nfKprIVB+PURcJ04k
Jp2lFHKnTavhUBoJKbWEEQZhpJ7B16cH9MrEVmXXXWeVTn1Q2LP7vLxx62Jc45Zw
ikxXlPvj5IX/074VtWStNKmh9Bxxx3KNr0jJE3nySWHku8CTv3WAxhqsdRMW830c
mj9N49i6Hh6H0QxnNfU4/j2lnLSpLpRpJ6Z/5D94bwEzHAuEnJjnA69GGcWYZNI3
+747qI054ayYTLv9ccO4/aMAaLuVQbPfUYHq9LwktuCgzEhfdc5aVJiVHharkEpK
YsjgXeq0QAYURBxstBjTLhk3UnwBT92D1V/2Wix05Qrbu+8cN5mEi2361eohBaja
eJeSpl+mlpcVqZt6tYHO3XMqgUoX6PHk0NghscxiSR+5FDlyx7yn0QNO9ancGEuR
nKD8fjeYapBD/MX79+LSklKj/Aw+TbiLj3w3/p73vh+8ZMiH5XXUgeqAD+Y4Tskv
oUPu3ulHRfhhyP0aTq8CoM5NQK0xHr5fbwwP+AGcdBQQboPGxTuWKepczaO9Sjad
qu32wXp9ZOltjikhK62IkS2KXo9/gBnrjnSSK7FAIa1O0QA4bd+stPWWHSPL1F9n
XHavR/GIixmAlGTm32agX+T2WvN91WIAgnB8CBVrfJT8MQnbmBtJEo9OtUva+Nxs
9MnoN6BPBgtfKoJN510jjAfMSDvTakBd1QR5Lvt2YouFpdNG7Hbk8cOwJ+fwChZ1
De62NDffW2+8mnMHvJIrWMEWzRT5eKcQ3XBAZf/eKpOlAT/NUZgtZheezKanSdaA
Hw3ZA0b5YEvRLWzwdkgymW55faPEjGR9Q6ZFAfRX8AZ6XGkCMNAAiGywGeW8rI+5
gBPk48dGWmZA4L8pHmFGYTh/ZPHnHvCTbAsGOVURmPFEL42GQm19fVUDevJywCp2
Gr7z/OLrvMs73GsM1gPmPdVElsQlJVOCPO6DLZmh+Q/IArJ8OMfCcIvKJHPNmGUu
YKtfL2AfF1JyTCs8XgMOSY+CGlBcvt1jnPs8cAPoiS/m+/FXk5kyEOKVLvuDtuOP
5aQM5M9P4VjgL3BE4Lvn0o8DHo0vViqJDjBjMqRrX6wc5v/lh/3pitGBUe3ebojJ
ffJKHtkpqrdLCZwA7isw5yxvrEs6RAW+EOQ+17J+6vzzp8lVwaoVwwHRB+pVOp7M
nKt+yApD8q0SdnwNbfQgglffs8QfK4Vp3iH6JGzeHK4/98qfVegQTpKCu7xkh+vB
QRRVbGcVVWC3nSw/jLD/V4mWxhrywxoakR9rsfOlIxUe+Hg9XnkcBj17BulePciR
fxT1l9CVyUBNk4mPOKlkJkeNaYtZniFYU5zqd55FN7/AuFCunqafTxstemOe+n7M
nqf8d0Yqk+C59EOMEu5POeLlXxfunt0c2JlGJtCBRHvbhRNB6MB/1RQO5qFqM5I5
PtzaCctp26WbN+qVlRK+Ah7nOlTedLvYcy/zxl13SOZhzZirJTPi9IAIWd2C5cYF
wohwtgC6ZMpVHyo1z0+mBOP4OlloBcNNJMKf8VYwdkxAAhnrchNdCMQZs9tLZHtX
msN4X7NDqJutF4zfwC/KWONezN7rK+/cB2f2v4TrV+R8mGC1t4o6TRFQwJKz0oxY
pdsFzsiI9uOs7wEK9tierJFImJPwQej4Rg4c31qmFoIs4arpOWX189sV+0IattXA
vc4doirFS07T+dBAGrwUBBqPTAsjpu/pGm1ufLk0jqZNUwqUWnFL5bwDdQHN2AhQ
9qXFelxSjVbJOmKCqjfM5Aw1bmHbyJwrTjEv3iZPibTNEdPMmWnuPOCVGXWSisHO
gTKqHa7DW4DsFXJkWEw6HqeprF+GfovM/EFgYXAHBg/s40WGY2esZ5fUrB1kVuHk
dXw6rBCxVV/EsDJxfe1UZyD477HrJ+U9jJ4OSew0b4okYC7xlA5YRlte/jeBOEWm
6ayfewaiRFcO8ZMiQzUVlUU5U9N/Eawlv2TJl3oO9mpvMaGPV/P+/gEFz2sOijxW
dBpet5jROKHxIZPRP1wGMFP/XLGcvspLKhio3P7moRNtkOfHzZlXV2PlbPd1ORy6
THQovmdpofZZB5EUkdLN8gMSP7h2tZvKGdZmuN6z0aNSrzc89IpuzFTy8NCFki6t
Dq4bg5KLJc2VDTEfqNgZ4YHvcKPWMbfD3PprNbUGlITBovGkEYMDTGz0hOp3/gBV
F1IBLwOh5h0pXhcnmyU6Oy6ayei2jTePgb1Fj5jt9XLr/7hzmyhesQ/aZYIP6KQH
ay8N1SlcDg+dVCYwgCq7Iy9YUUbV5juK6q71gN9mI5edQ0TaZ777znNvg+rm8NZ0
M5IUaZFr6GmVgYpfbitxOka6M+Jc8L/vthghnLtjmilTBfmvyj5qpfA+ZvKrSYus
/mld86NS5Rg1kk2mqUPBDOs9+Ai80or2OqXNOC+Lj+mwIRUV2qfTgNtrQyw8uenl
Zh5zVRWpwMEWu2JKv/ON/DiZDF0GDWr9UGa8ygy707dy8zQWMMTfekETaMf/gTEc
tC/zz+80N/du/oKYNgMBqkAg74tgAx6f4vsDPZ6CTejxHXDuhjh++nxLMbmT6J1a
6sWRxXNju/IYZIULVREn9WqdxK6JPkMSUEQOgb00QZJmoQcFfp8gi12ivfhSvVXL
i/NL9gPJs5F/tnkbHrHxiRllkbZszcpksCnmoTklmrOMOki7JqI1WAk2LlGqBEud
UQ5vH2vJEZTnxy+9bckB78zhlcbeCO/6riELBcywLEqHudEtyCmkdGMd9wXVx9Wg
DodFnXdE7orBx4dNkbRDL2+NYvBz0GTSGhTmiX0dyAQ5T6Lcca4o6s8hYDqfJ9Hf
DH3bV1mSVhgYywIRhiVEIHpmaLf6zqqkpMDKk9+FEaZPnmGMHFQbH5vK4gkX1XXn
bXPs5wVu1WEBx6n2hChlRNonm7mA2QMDGVM8o48nNxHjruiN2sC3ergz+koAcJx4
93Xgc1LhoYC8nKGPeE2vN48+sZ6Lx7uZlIlSLFU/AnjB1edlrhWMEQf1doPEL4Gc
/r8ycUfk0L0WHqcynr/b099fGb9P2nvd8iYyd+uvkqVj5YhdENUNFG6aiRlzwPm2
eNITOS+NbnwYAnJgBJkkqFNCwcU2jazFcgGHRhBdR5W/XhAI1fXoIVUztgL41bCK
dMJdXEsdlJ3HF+tZK8ECE9Xh5uEuRVJY/bLqzb5ie0EC/b1Wu3lBFDSXOvmkdgMW
QpOV4UU28PS5PtkFIsHyyner9k/QZLhXmANpBwDFAHZ3Mw9cV2Pu3Y4XO3pG5NCC
28BKxLTva8mUDP6iSSREjK/L4Nzh7Sek61Q1ccq8ub3ztH4rRn04tcobsfwDyL83
o9LAADGzniCXcFF9CWDoa3ABzziaAXx6yaavKqTmEcgUUoMJ2PBYpNRXGZHj79ma
txrLRMSLJotyJy/X9bIpAxko8iFgohLH5+pSwKMCDJfvZVoTglamRlkbkHAKY7To
xwoIkFXACi0CRuzxUoNxjkXbnvDuiHViUBBv6Z5UJC3SWE3z8xvsU06qEX5yncLi
gOq00vUyiRqPVk0+mrtaMbZ5r0OaILgW/3xSHp2qJHB8AQikx1yZtOpx17vZ17V3
IelL6GX2xMFXlWv3cO0dO2Aga3fW3a/OWKRfMX1u7p4E74RxMXGFyPF1nwdOJUvj
6xwfTzigldxBXE6oAUKFlFiHRGaju2zM3N7zxtp9SbxzTYyslnnFWRDr/JRzca3Y
G0HBR04y/D78fohSfdX0auaDdNnGO6yn09RYkKLvX0FX+hwe1zAYjzJ4xNSyjSiB
aBfBZkWIyjkLT5nLH9vLKxq97qCxmkXQqcf0k7PP+QjDfeeY/UvNRUuuqIm6DJgb
K0gsNPAx++njmgIDayRtF7yAi92oG5p/IlaaZjmjhlvDkNJgXKOoCjhOjfMmDL3d
snpc16rAN1djCRlGrvffaSDcLJOLkmcNUCPs/1d5FJxHyXk4n2THmZwDyx+J/bm3
RQPNAfP09/IPhsofhvIGDg==
`protect end_protected