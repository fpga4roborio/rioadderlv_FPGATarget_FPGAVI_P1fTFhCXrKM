`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
ddtXksX2+yylW5zu6QL2Lhnb2d1sD00763mmSITNX595NcHTEkwn0zB1Dry37fOW
FufOhVzEJp80NC5qZ/+F0Vk7Ik02dIR0elf3clrjeJRK85K4e3Hoo4xn7YbFUIms
l/8VZSb14+JVGURjfswrIyCUotIzlzVYZ6gzoZwDXIi5gQIBf/gI+KxNXPaKV+PQ
Ufys/12rjO6aI/pPlqSm0hCvftmBcnezN2hk1UeXgOIuKZnogjOsf0iJVX2aOOWE
6pD/psybjbnsNB6kH5uFTA5frkzIzkzl5d9+YDm9OyC+k84E83I/7/j+rk4L2dah
QJOvksSIzN867/4Qt8qYTQ==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="MvBXkzurAa5VTw+1JJ70nePUfoQXBvZOku/SMmg4TwQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
oRtzZL4VJ4iwysPsC8SXYCzXS8Fw2gtZTOskLcDV+1B9Nzn1zTyNtlo6lNICRmmK
ZRVu2BmCc2G+fmzynYlNTnSa7C0Cuel6FYpxCBlOuk3OF2tzAmLAuDyOH3Z1Yjzk
a0aHuoCdIRKv7BrZCdALt03JeUmXKPdOmIlkVGFl8yw=
`protect rights_digest_method = "sha256"
`protect end_toolblock="Jn9CQpRhJt4rnzZPRk+dOpzAubz7omckX1MrFd4p81o="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 10784 )
`protect data_block
gD6l00tciPUa6pDNTk/+t1gcgy1iCdpjTkA/bOvU9JA+cpFEv5u/7dp25hHk7lLT
6tYtR8HgwcLXTcx68BnPlzdPHkVIv0lwXo6yhFVkYlDWBcqD9ubowgKij0UjlXmV
p4anbpVt/gKvAYRDYe8Q5F2CQ8AIsxOuOcJ2vhCPchS4QF3n7+oG0MKU5ZyzxTu6
Mm1vk3NqQ1BbbE+MljJLKYlambVUuT+iDYnAcLnUqpk1Vxwk0ySHow/aJRBCcOdo
rYPaXUO5j4CPOkqcSVbLDG36ezgz5QV8jahNPSj1PxAAnaeW2+4GFOj5G4itCpqn
bv22BKY2fPz7qPdi+N0MxdAU1GWgfeN4txcjxeSm4gG7rNZKRgQmAz4jaHBLcfwt
Vesz82MUAWG4p1heRbRU3+aYk+rrPkH0zu7lwrCWPyX/Qy2laCz/W7Vcn2Ik8A1E
97eo455LuoeQzAq8nWLAgRn1TOuSyjEmsGDGiZp24eccicsA3Y1aE7TQ9xOMpr5h
BduB6IEBpRV0mGlKIRbzDP93yeLQx8t4dNqJXFsrERhhQQkWTZMT3gGhflTDnRom
Q3CKdOW9ZT5CClQT7hORSUq5zz0GDpPdozY6CwAO8UE8oo2GZxa9RhgHZHPN/Bzb
33+54WNBBPtVGCvc0MN7KpVw6CBGrhmS0CYUHQevtVR0wWHQ0Vi1d9ey0FlEV9o0
i8qdEUtAqb9V2Qg1StmdPIr3m1Sc2k69NpWFr65Phrti1NPII6VWg0yk/qItACUa
DC6n0+HYgBuB798U6MdXS6O0lh41cEKnruBSrR7SAPkEpYL5PRo9ui2WzO0Jkgle
3Abc8rgSJQOkNy/s38xXbZ9JmtRW4mO7+ZN5r6vlgOL6I3/eYbM8MZeL/SkngHFz
AcVtAI/x2SDs2Jl5u0G3zcoQhw3ID63PZRHYN690e6qMrRHB1nP1c0E++F5mPWPc
J093tyoT0eyNM/LKFzsrd9MAf3pLA8HkXgZQ23vNgNV36qRmHmwO3e1Cvpv+aMhD
26+s4e3Q6oI2TK4e6J57giwBuUdveC6PmN03Eqon4I/Gt86OOElXJu6MSqYiP4nG
oXDc5qEU9wbtqPl7S6gQn6gxTShMG5QU/AW74uyn+fk2ZmUn9AK0MuORcGQH2x4r
2zTRVYQPkXrbJ+buFkkxdZZ2KlJ6SWIW4fGgX/F7TqUGWF3PtJ815KeBnsE6xrAV
llkp/ycOIDOA6irwDjj5ITzhQWNphf7cwzJLECK/cqnmZ/ckhFJ8Unk+TCAYW2QJ
+3jFaiUhRJ1tWwmXKtwgCpdSiJi3IDu74oDKUAMC4/Xp2WI1GNr1Yt/HSkXJEQij
qlpcU/YgnLzh5koIIXWQlULIBLQJbVwp90uhTGe0nzseuar5WDP3pWIVdQQ/1dYc
ZGK8AGNrn9v0Qi+K8enHXECuG2NI2Q5WcLHHQBOuYLsp0BntUPHcACYwtPfG5bTr
AzBRzHiUWO00MMR+PSLTrqVNWxjwD8ZKD3LdgVT+U5OUhhACrW0uufXykEl6a78G
vMtbJNZ7nPuVL9777Ef8vgtcaGt4RTaa7GYCAlZysYnepQN5tM4eqm1+sPSPNYKB
VBRZsaqNetSQ5FnXViJz5TSsxGfnTeL0EiVJLgZyeLTBuLZOQsdZrR2E/8UYjGR6
nZnYh0VlYNZ7qka3S0zwgSVDbxY9Bx6LxnUg77NhcwXwWGBUYef3WFb5y7oVsqE6
+uMZYvRe4OagCFQiiltQ2XiuM850OQAQ57yvJs8ggnpw58SZgwbICJdry4XEcm6A
Z5JtrXQirXVkqbTilImROeWOfajwZw/AEmENmv7VqX/J0OQNCN7V5TWeqkV6Cz/8
iAwZheS7jZ6SeHzClntYIxkKZ6XDbfQzMc4hTbxQDK1ewG+Ov8J6XeHFTfw+ybss
YyiI8QqMMUFaRE6wiLnP6wHmirTcx/FLdzAhgtqyU1twNhfMziBcTqwI2m1iIGhy
+xfVnxDUpbQV7C4uYzYOJyBTORfTFMd24YYtg03fNkyRsxLmmOxlRPecajWxFWON
lHjv7RQDQbZC2ttQ3UBcKK5qQaKV0L4fz1kct3aZ/t/1z4vcYkTFwvP3Zz6yWMpp
EFw3al13Y8CrYQrAqo0nJIWE6khCuU/SkjBxiugZYDmCds01I88Qv38T2q1HkPw9
GxKHJyBkC6/VZ19iE2owIf9BCCUcm0ic1W1tT4Pl8myXeNBqtB8WAkT43Evzk9ly
GODvBfgm0jf8v/TdySgOCRLRqPBhj/X3vlzXHSlQaASAARaU/vMQMrGr2jMFwUOL
N/vYLRuv4/283+YwGqHXufxWI3X5Hebg/lfcCxe2nwIuEjiE5QveN3Ax/UjfouMA
jTiHnPZGxz408DQB/bY8Sutst0xVjSPu3epr0FIc+hh29d1tfvuz70yrVEhNUgLQ
EcjocGBdPOB8A8PClhSdspXraGivzfs7RBM1LyZrnW30jeUcFM1+KvAYJFxxjnGi
0ebJD3pc20/gp9TbluwzwKbnfO/9q7l887ssDa4/xYDJF5Fy3RCFZDO0wJcsA0+g
790Sh3GSZmM3crRrQ9ZdVimMfQ4T6YHp/2cZuaUOonOkgy+OCqUsmaTSdWdzeXaC
arS8ImP8dtPkiqMZqyZtfcO3T+ukBUXtdE6KHvz3tIKUR/RZGdnJd2V0Enk+LZxO
twqhgdqRKhAgQkXsD94UHSWd6VPDtejZsWjRsvZEfzv5nkCiqjNok6+OLoTSzecI
vycf7JFHEc/HiqNNccg7ipWXOwjUfj3jC2gM05Qmew9GH2LsDE+fDVpLET6zK+p0
pdfp3/6fackvBYZij7dW/Zhej3JOZIn73EaxLcX9khetIm9wIsGKV7OJIGXiSV0E
NLh/2QhEN55N0WXc+wnOJN4DWDbaX8xJMcHjIgps9ZdnFgJ+bNIJ8O66j3/OALZg
rE2EcaceAtWB7joj5TrWRGIBzErB7Zxv9JB40EMEE+zEbenRCongW5pw7X29JnR6
dRfCl5VjmMidAi4D1pW9eRC6yDO32GdeofzLwLtORGG1A5Q9en86I6RuSXNZvqRw
QmvgP0WhEeEOnJU6JzVtpeL/u0Ducq/IIEaSYs2ygTpu9cvQttwDlLA5WoHLZvM3
rnjjyf2uuUmeNE2TnY7LCfVZ7RThQDtx4y4X5MRDvsZl6u0AiYtxT8nSr5fllRqL
zzAqTAqZ9Yl6h1oLu0sTfj5nGQNXciFrFcZ9smfXiy5N2y0qlLr3QJeZYObumxU4
lAcPFRXyQSzHhN5BzM1NiFuAH0wgyp13nzC6CeEcFqHwsaOlGIidKRS1EC5Ntjbo
uBnj23wZCkgfha6CpU0VM1AMGG0PfXIi+sWbYWOT/TPzEn8opVaS8sKPeV6/2VpF
UYP46kHhsBC/05fCbOFX1HeikLV0N0btLlzsn1Wo7coUhOy4mzyFRTTm4hIKtVsb
v/CR0AeIeGULeMQTiAtNLCx3i9EHSx9d2jb7ycfFn+gqXWIQnpU2PVQhQLF6XvEf
3sAaPMy87BDNFOl57Vl1r2XB+Jjk2dQ42YWIdmT0W6gCwZbkjdIPatHQai1lqd2g
AShyNSuJjnv0M4QFXMlWIf5xdDmTOZcSBLTDrZ9on6hUQv01FsnAmG3UDy7oBcQl
/GCIiwNUBJUMfTy6uTisdTVQH10oSJvkmUHExheZy1sHXmtjHU72fddvSXsNEXGp
KWCbG6HUQUYgc+nFmg82Phd2go89p/lx9j75IeEKQb2XRTFjj4qTBWlj30JOdpAH
12Nnbo8qf6wxJkn3d2gvIEivoYBNM/Ep5xNTfsHQS46khtY00zps03V7un6QACMX
Rgx6/pOVbYTDLjajN8kmGPbp7T8It6+uQtFgwTBros9lP5j4T77fvX3ELbHAGTVI
nTX7Zk5GF/lGSM1LsS1YE0a+7GjKIaLHZFZQpQ9vUgx7KOimERAd3fgGZ5oTeI7F
qebiPRy9vBQA11M4BD8lce7hkmFj2Wj6G5hUdEnxn92ocV7J8+P4hugXJbZycvbc
syJxqKWJW4e8WqXvxkLauRW93EvKbxlb61nfJtxRBywzR5X6KhPgh0mMt11Cyqdc
CYfpyFxQ6g0lVFbmKmEgBwgNMJuUzYTdXAvayLuewmJsCvP1pNwsEa4Gj812Hhkn
uvuenFgZOLluWs70fMTWJ+Sa12sB7la0TrCgfnudugVpWsgnzwWE3P/Yo8YDVh7h
0cwhh0n/woCG1soFLSGlaREuP7nnshCJT9/e0R99Id5PT3pRL4w8hba0g22DeymH
pmMsQBguI0/qPv0SfMRNRLACsgJemPyd/q05eulUKYGaQAtARPNmDMevQ9zBE4Jr
oEDR9bOfPNmBzdzT+cU1N0vk/nMNW/XkkpU1LLDP1sY5WmabS+0MHMi/Wr5Us2Sl
Cbh7yqhQlwIbjS9XSgpRuYWoB/jnNiki4S1Lxd74vqPwTl24MLDKSNeNmSVCpGdO
a64+9wedtH42gevTiI1EH7Tgu1CUvV3ZDICBKijFN06GI4UKDoazxoqIIZys1Du/
iCWPQSnB7S4/5Gs2u9t50xXnE06hMBpGcneihUrVDunO4C4xgg+7zWAavAubIAvf
S+UYREBuNZL2ivhDU4yRrwjeaDWDJSqE+m08psKRDGbZL3aoBG4EZKg4/S7T6vUQ
ojuxyOzw/qgfyoVOPD5DcJxfTJbaGB+nvU5i2asyA1hbW3QZey6asF2oWGzgyDv2
78OExV43MrosQLlkXF8YnWOnrOeA+s3DuNQ+ZNqrwMz1g31m85QbjNjJ8bFCOXka
bsXG+N2+bMXEtNv1WwCktQR/PFx5gE2rRSxQ3F4i5md0Gx/XfF/mDQ2VXnO6ypdO
hnv14XosoznBhIxiKaAOFDvYOE4o8p5NCnV8mcMfZ0iBBRzNxl/dNWa/IUzzLQWi
CB6/JvFHhwJrYFJpzITgElzSN7mPi0oxZOq+U6nKqcVHtTFoQ5EJXY9hsHgLx+c3
kFzReLQWWHj8PqVxDJn7rWlEndNwyPGQjkGokgpczXRG5lzxCddYTMHF+8ESrdw5
W6DFPka4tdghpIAFu7pzhQ5tonwiOO45DBZ52jY3Vj2/zG/zoLsUqr7JHAeT3oud
6r0tyYMTxzp27HAtWA8C2UdO5onsCfRX+i1K9kBvdk4LBK3XAcxEoqQBTbW+fi6i
022G6aDnH/sx+KiODwXF/sVgeu3YEWe2UVelXU1t9N+maVOjl60Gyf/2YC3Tmlh4
xhu6zHVFxxTOOwrkxsZr+5sqiB+an7qExcs7nAHmzyXjfWN0oS1qPinH1sy53wnj
AnQytvhptAeYVGqNE3Fqm8ISYqxwiZWeIOBzwTPqmRk9odBvSKAjZOlGtPsYpTT8
DSf2uoUVnq3ULx0+rOkd1bRoGsZV21pl2jfJjZVQnj0cNiR+Puv1QxZ9vkm0tQmZ
fBSA3HP851haOUwjVm2AIZrGPP3ZgANb6cwiu8icyRomQdkYXCF1hcY9j8kCwjYr
KyNArPs1+WcNMCWUi27BpFffKmeoO5s0t+ErJSsLK3tDdYSdEgOp9M1JMhtdoEiY
CN6+50ZG/GVbl/klAUfZaAPk5IG/cvYEB17OT3pz715/KfwL7AWDNcWmFyA4nfG7
hN6PUNXywdXuzkAuSo1dlhcrgdDeKBOKfhNMYqVUaENDtC71OesZs6LafxMg8GX/
o+hVHgws83kv2/cy/gT2GnCEFmpBVHRJd+AahHHTUZ+8em5h3PpWR7y9rnMz/5eT
SXcrn3qHgtTUo3yzYy5CRAxj7QcJ41ZDa53dqF3RG1a9aBDBlKS5xTEMwjHY++6I
df3wmPjjbfDIV8zoSeCAs+eFFXlsBS6zgF37dLcjWiY0ULMf5InZf4HPqiwfxjxy
xZWIHqHnHHFBUsx1qnCwp7gzl8TE59GAgEZuhChIAaEsIdtB+KMOFLU2Iw7Hy5gU
Xjd7Y8bUxpAk7IxL+zxzUE3F2iEQqHZ91tw7KXXRmvfv/2/r7q0/b0GUHtt+nCcX
yRROayA4GTJpKL4EDVFTvFRrHj1dSZDigpNdU4JKoOvPOmI3w+DVSLZhsL///lL4
pHUGsc+k5/rzAz6c5giVEUgJlY8m+H9CmRXTOduMap4jkZ2LfyaG5N70D9xdyId/
T/4Zow3G+hx18/UALz3IbGfkgmw8QHnTfCBovkGRe/WzTuoLJJzLapGx14jqIbTq
/NUq39gkxINkvtq6JNNLJVjcUS6F0rJh00QJ5xzaXdH0DNN9zUc+hirLasQt6woq
OxhYHJrm/OSQ87IE2uOLojEyVwSSRGrxkrMlz2th3Jqfv1y0Y3Q8DqUzl6f4OSrC
9KSOm5T2VlB+Ivh9wRQ4g9SEVPxp4tKPJW9Bb84jBWIJ3lcMfAazkuJtS/5NwTJi
wR1oIwMD5uvduO7gASZUGZy8ygaWc/rgrAcBQS2i2CBLaLYV4cRSCUI4/dQxfa2H
gQq0Zr95IJn61xRtTssPsn5s0o+/CunCNMj56QswWTQBX0EE7IkjxXSJDsmm+Dep
M5TLNNGkJP0WLPUdlMTIt14+3wM/K/hVU03okJEgJyy7FV4qTAOx3E9cC2F3s5UH
oErx6OO7YGFF2GrDSOOG9oOuTpFIrc3bi6kiLnwxQq1NmzkX1F8Exs1qxzYfMoSj
ZX9qexPctlCeWZ4JI9KB+ZtgHCWZBna+5i22JSCVaS9lLsN1vXjhPwbq7oe58lDJ
/erh48k19upe8xbbc4lUvc1jFjhfAGcMMl9gSa0Lkt0USCk+PAwc05Hcp7Os0o5f
SZ2g33lYZge8r2r9b51YGC0C8NQFBBrfXh4dQTHDiAe2dRlxh8BmFrZbt3qf1eRC
tjazbAIFyY/sgcurwFrA30yu2LKmY+vRYcpFEx9IRw8/Tgucw42uzWESx5f8faLq
wbbHUSPpE7q89PWqyXW1kKfbHLSgwY7yV9AxekBAy2j5GvHzSqp0PX795Si3RhBq
qh9tR2Og8Tyyi6t4yoFMuIFSWVuSmrV8iRt0tOnc9bB+xOZlUYjrDaR9rt3iH3G6
StKY7/bfzXdEwx428lOZql7DTWeC6tbckptkBV2GRWqVTXuiFcvYhAxxdYMJl+3d
njdZFBy5m3OJQEfEZvLI3Ozrf8QB10nCJhBwEMRfqyA1kVz7uj8YitcRXyitUqhe
SVZvsNftAldHByszi0bN6BsecB7Q7RsyyOLSL9AAw/hwWHaAa3TGZA0kz2MhLQXD
ZtXIhqtuE+CkDH8TypqzQRRHob+W8ahD5RApdEgraYu3G7knnOQBfPECCF6da5P6
CCkrhMCV1A/AEwQSswRhhKhrA1yhV+YZM7aQXbqb82Zyoev4S8aDjpl6BLeeAxNt
z2XmcKUQmaERvgPHbyZFJvf3eFrf/UeZv4uPxikzXn+zZm/+AnSPJ1x3qSWD4nbg
I02j8xd4iaBUIKHHy1Od0ZEnO/S/UZPxxRBhBYaFjjNGs/dvH9ufjjUSznn7uSlR
ZnublEHs2e1kRI+pFBMbWI2C/9kjgcxlVxAOcLkMc8VhjAazuqy44Bxw/FNXDjsx
1qetigNgwZdUFFzOfCzj5ZzSIdYaWuaN0uuo0AtXHXKdMYBd7VeU6NZvx1UbCQYo
KPesP3czr7QewSL9Ck1foJ14m6rfqgUQ9jCiQMBsRpOD8E9Bck7HUuTk8KeHacfu
Etxb+gSbWgNTlHf51s1ewe5xnjhgxDgzNnpqdV8wdgehraVQlLoyEIHUGPgKcyMt
yTVQ2BgriA/qaVLYsj2M9BwuA+P+rcIg98dXxaSHL+cqdhSTpbnx9mi1u+v81ClA
n4SBjj0ryXxtGdZzZw6IDv08QkMvP5r4NAKpeUbrtPlwC5TUEKw11yjhUA0No8LO
O+RC8zCfr2h2k1l7dors1s5JIMfzc1m/XLfwAjYnNYsBkR0tIAPjs3IgAMsA7j1U
96rOiX8+Uc+qilZPLuLpSZSe5UqlMse+B8pc4cupKeImH+luJVQFd2AetbBnpakt
/iruhXMoVfukP01uFXB0wbrfurjG1jfwsr25GrP36Uhgu+bTlZouwruQc6qsKi88
dEjrreNsId8klS0RRivoh6A3r9aLhZ9FhCbG13PeuNwXBKCIGTYDK7PZNqkXD5XM
v8/qZmV4Y/XussDfosLes7HLkBh/U72J1nLCH0PlF2GUAWeT6oVIrzqXXjgHNk2c
D4KfJJwoJzvdJ7aSUtMNrtjct+xtfZlqcdy4OFhMqcJ5JOIc4IxjviQXm2BOJPb+
es2u4/l04y//VOlulMEb4htsZxoqSPRGYRbMwylqKnY0jfS0QCTP+oqN4ZxQesov
Zy0cTfFAqZyaKah2BWp5xtKWE4yck7XhrWXNxeYbVq1LSM4iCDjjs0i59x7egCHS
Zw+4x9FKFOF0AQq0RzE5n/DMQS15YXQ4V2JJqesSWCGkdQWb7yPePs9cRnrCq2OD
ZGvMh61Mnpcc/EWPpXk5Mx3vZ3UE/reVOVUiNmwEtvVm+t09Zh+IbkM3RMc7V9/K
MoSlnPnb3/Z5eScEhr9m9sRwbmvRA00LHrCNREGplubmTtl+5kAAXoZqWTgYwHMf
uCGpaBoO2kJy7WDihJsxn5xuzfGMNJoZWKN84p61XX2qWPUg+YUDkdi3J2x9NF6l
a/F+mBpzB8b/3VBYHIzEATdUiJFbY98VdAMREc2A3D83qTdRQVWzb4E0NI0CWOWs
Xnnyr/JJYZRCghDG11uOWu42MoXi8fz9NUAlvvdYlP/VnQWcHIhYFHIpNDWaGeMm
THqr97s3jcVbur0eaAJVg8RVaNuPSqcJ09301LrOtlAjVAr1tN4iespRAst5AYer
0/sNj5JiL5Qlhxmg7HzQu7EoYmwBOjf4/pGziwl4RHu8sFzUxLJ47f0gZ19oN+xC
mUk0WxA35jC2oF5lGTfZ35Be0E3WbH4SkOFZccBSjeBPyYfdz7oqYA6u1um5CuHV
dFFKbJWVKS7ZsitcPhxekR3ZUL2Q+IwAWrM+oykuCMbdjpOiS60oJMuFEzHDmwDG
g4pXLib6u/YiguK/59O37Jw50/jl3IsZLwRSVbHfMgKJ1qDmFwvnXJUgsRdKzeJd
nU6DgG2lSk3wR23KqHn7wv/LVSVVdDCOwmkGsp/jSzh09YZ6rjjL/+za9U/Y57/x
jyhADm4mJrRfKlUlxvb1BAUob7jdT568fdG21EI+DJVE9iC7oe5C72gT2oRNHqDe
J3rVLwvFZE9Om2qHKw/d9qEFPz0Rl1gqJNScpFuJE8BMJiVpWQCo3o1VkRtCsHTX
OCwisiGardmtFxykVSV3IHQXHoAr4Iyt2Myk0fWxeqaVz3EgEtfFhVTF76GcrbQ7
hSjKyTON27Vp7HJ5yqQ4x6hU5onkFHxNiLPLtOJHiFo1mwLeormP72c3HWY8cM51
n6PrKFgyzDP89dD8pXJHDgRUqKWuc5uemsYUT0ZLF63CqgtOEHdAt5UEd70gUt6z
o9GkZVkdOXvloypZV6bcE75Gioj6cDVFH/ktvDrOZCNPzS3qa2ZVPaS0AEKqsCSR
GTm4syc/ezRSw6zqZhw28WNrjm2ecIc8J/9TCrsE4yjoifWpoBeDsZ+ylcQixbCd
w15aT7B+63oAjeGAFec60+Vxehy2CkJlE74o+u9gf7xmSYTjsDSqDeE3tt2wwvR/
64caXm8k4Y/TAHAM+1gUnA2M95H5PW+GU8juLqg0j54dkbLkSup1VsHYFKV6Qcom
WHZWbb2+bD/4jC/saTBxMR6tOCEOWUAq7m/eMrYdUMb9ldaG5TvY/1oYTTWPy3c9
vg8MdCVM8M6GHDLi8D4yGJY/5o7xJoHogoaQAM5J1bPPo95ZVU5LV9ZpzWNPTCPn
ygKXRxq/FlmB69rF8FVo7erb2BzRB8rG1Nj3De/aAOulU9vB8isORGHqplL6AnFO
BM3TPpUGz1u7R+E51EEL47uOEPtNIwp/vgYiajh6cYbZTptOP9h1W0g6ZjMIK3dE
XF+v1qw79XJVuK/RSZdRlHtHuFwatLgEAN92kz3jGx+Y2FFX9RlVDqfyvNwB4H6x
R4heMraRd7ah+Y0kIwpFZ4kcuu13HamFi5nb/3Z7OPMnIoZIYshIoyZYIOOcchaX
oR4uMTT6SyEDM60ZT5BSVcSXZika78KGbJW38+ncleEtYz36x4VGKTSnoFrw67W4
YMuiDMmE54czzBQvCaxlRKtRSEgw4VapEfD6VtE/KeJx8HgTmzNS7HMJGvSI6kp4
tGaProryTFbzkEtWbjAz3+zrqZJ0C4CUNuudL2WhCaZfuJGj1vnJx/ZoqxIbnqYH
uTBa03pjh3WpIr/C7nezGVTsoMK7XPRnX1KdEOwytp3PnwcSsji3dNyIjL4wUM6Q
9D5Zc3yAlEacjXm+NQ5eUT4e19NJil7qnOtvQF5kgyLB55ojyFecLvRSrdxnjuqn
Hlen4VNWKgN7dPwOk57ZzOq70aekiPzT8C9wMBalCgMcwLQHGzRWfC+krkCf0Wxx
W2cV2mxHzjOnrO8LSDNjUad/4Pwgf+GZKEwpyKLb9LJeH42HYkZA8rqjatmzt4rx
JHIQkQsMx4kB6op7T8n8B8uG/j0EdIDxLULR9BO9GfBQ9T3RVmA3Yk/iXsepYiX2
1cs7nZ2G+JSR++5kmZCVTzAJsT9qQnYZM2OWa989ullURnP7GcjmcUUe6qBe9Qqw
KYKoKXOBAUl4P+F2aQD14DXb2Ud28bw2aE/4OTWUEUxX0XdWKrv6e/NCHtfItSQV
RMUoZN0j2ofb1m/P4V68HI2hZmLQy73oSrp9coWAhANZrp7+hkh+CYWO/f6PBrN0
zxB/sfRsakmXKa+hkEhbDelCv8tLi5wkuHzwkiosj+PHhuTVIW6qXJwdgxdxt3HT
DdIIPRo30aAy0YFYVO1414M6yRz83cLivm98wMl9QTDkkzfSEqWm80ZPsanpw4ok
66Mj657HgfmY5iRERpbIjYxQPN0RYr09jENVKEY8Wylm/qnmHk2xMZ4+1sa1GWsb
X0gXMlj7QkBHGBZwEhV7klHfqLkG5KZGXCMfra6zQFzkJ4EMgTNfNkrKXOTnynWn
dvbVlbFijxx9tH1xargTG9MRBEHN/okruwf259I7gtnhAGRpH8qhekgemhojU0VN
+HILP7ZamzNU3WL4sjnK5DXwAT/Axggb6GgROpj+zFaj4QP5yGFglGH0CRhBwHwo
G32Z3etW/3jp0uAsI4wMalcISF/v1UHt7cNHvjm9TN635R4gLa0Pez6YQIAL1s5w
Iehrwd4En562boxIQ1Jgush/EZ9HUjiLO9atg/3ndHPzBlSJHBzNb7bp32PrREkp
SBQabskdjorys5KPJZl6ZLOuGvo7tvmNJRF763BHr1X6O4FArAjhSmNVm9g/yqg1
VHSfiPen17rJMhUAhNqfRNKfQHZPa0h+nsUo0DoLVm4SIbYVjAamhScBo5jxcZdS
230NCw6yXbxo5/vT7/Nfdif1foHCkpfVo7JEJ+4lxHypZMvIxeKRLGr5dNkzIZ2t
Q2Kv74SnYqfhBbaVHeEgY9CsAGPplKSNEZ+mAItWE1qWTRfOWKB2zt1d4Fa2NMUu
g4QJ4Vgae5v6xq4rU3+zl/ogNT7hOLi3gSPnPOptwLApToU5hu6/WY5Nct68Kd3f
l0CQa9bNvlC4CeYBcN62hcZf3trv8q4LBvwWqxmxwCcre4Lrg1u5YG8ROaLMZyDi
wdKtfDfWI4j3t+bEZxA4k+P+DFAr9ddwyGKT0CLFr0AtVEZe1yqEYImxUWjI/cPW
UlWKHD9B0wfKkT5E4oS/j3AAMdtAo5IsXVHP7jPE5tjCd6zhor/qJJMBYVPVRUh6
13SETLk87HEs6LzbyaQOPZOq+pNDjESqXlczEgbmKXTztA6unwnnrsETrelpr/DA
A9KjyAsLexM8/ovM0fOGVvYosAZYBdjQTZ4qkI3Gb/WDo9FElK5ibNLWVO7Agizw
UCOUkX/t8e8QxCq2R9nCqE6bN9hJXXuEnR3zQXOEFusQyg1b4E8X3pNCxCcuFbmO
flOLcjc4M3FN8+e5mBHcNGvrpgqCfEH8A9VY9KTicnus2Ne67hPKW0StMNfgodgH
oFtZnTlL68IIUNHbcTx1ygFilCwm1WFlzZM78hg0oEBe0pyeHjMAmElW3GbB4Ekj
wEh2uhadf585mCWVI6lLyM/BL1IZi7SV9Oo2SrAQIArLXvhjAjvPRnjzJudsA8f3
NWVcuCvbkS8N7DLnGj3urMAee71rUeAWpuHhilFd3QNC0UljYZwCmMkGBsA899wl
wubblXbxusG027XrEnpaK7GZFSwyCIvM66E+1X8JwlpP1niOxYcA3k/p1p4/E6Z5
p6pURkbHNKHbw+XHdON69K0GBh1DlmqYt+6OfgcEBd3BNx4KaMPu1B8lHsC0mTg/
ptaljnXggUxozJ4bQA9NKO9TnMO9ytXzdwnPbfdFKxeK+nlfuKrxFg8NHQdF/27g
n6P6xnwXbsEc/x+OEIXhJvOsz/+j80lYNHt+S03hH8sR8Tcgml38fKogNtVSbbqy
pqIjDasRuIr8WMM3w9/RqOSIH1Ckfc5z5gWw+PSHOrRAX/+PWOVduiUlqcJ1/pfk
rm6NQRvVqlKIZzVM/efRChW8RPY9DMwXdw0j0X3wvzFR15EUGqop37yqruvXkyTs
PI2PK4lHsAULONn2/TxJCb0sAL9a0ieuXXQ5GiJAACiwaFrL/HRHE5ABYlhLju2O
7IvO/UTOgYsu+wQ/WLvN+jKTZn7k/Et1VBqsyPOfizT2dJntnoIDTIXSXd0MbhMM
+88Md/oxl9xiF04DnYE3scH+pfXdKu/djyhw5fvlvSBPf/zlE9nBDOokgygodaLr
7lxlB48WkFw+YGWhAnQvQfo9J6v2l8Wmnsx/b0WF/Yag0N0sblx7kZ+gA92Nd7dA
VeaU8sWTLY/Y/QJG00nFORjQLW3gmZVuTa9WTa3oUdVI0JCL6ziiqiBLgXzds4Dt
W3EhyzBxuWSY0OJg7svBan6wEMh0VQ5+swEW617bGLGWZ3YZMR+5ZqLTCIUG5Y4x
lVnVClPZCgINNEvtb7+1VegH87ThglI/lcgvlHQeYeBGCD9k/4B2P2woqKVlMhdN
Dk/WJrmsYW8L3EA+r24zwytdsXSM7mYWZXAg4CGOV1XiiwlzN8s8KvU+4Qnx8WVK
e976fXhjJR9L07S2l+ugTDgWmMdgj4QBJhK9xmVD++v9ILZkIGWOuE0qlRKspuZi
V0Afq27ZfwieHW/Gg6GMrOgXCbApP2/d2WmW1WXtamsgIntIB0Y699GETmZhLQSA
clCADUalc7FghonxiT4zcoPtOLE+2qm6qvEU7QX53NkX6/rSzAayw7BcY0vYzkbo
5ep0/0YvvNE5EOyzrRD9JjHlGpFK+CO1OtnamXoEutp5a06jNYSKBkAGDuDJ8w2w
1ynIuX1oZWa2diqkjaaz4+/NOQVXX6/hGdkI1gi97/gCrH+adJ8jVSKlOZKAZTMt
9ltE18B2+doxbJS3GGg18hJQD7ZiHT7IyzWw0Te+5AqwOSI6TlUJkhHgu4Am+O6t
fhYVYrscHYgxR1Ce1rCtl/mBU1ZaaRPV8V+rYxMw3N2xuY25LTUfGKJEKYaSlvf7
FmqqdJS73bgk4F4S3LiBZepmcw0hBHHaSb91g2KpiSGEbg+inRV7d+jvtdkjRUjF
I15/r7bK90hpmOGIiTdzJtymc9/Wk5KIles+RjIKQWrcFhaOVN7EYpFSpQ1UOkdu
6K+6nQsI1O4J/uEktHFXabFv7Kq3SMYkO7seL6V+cO/pg993v4Dfql8QVIgjgVm8
HR95UQ7Hb0OXXJumT+leb9sTLtIMZdq8IrKOQvoMA8ouvPFuOMwspWW1Hr+bRxvX
FNQfeFqjOcr8rNcnpvBGSSbZdOdKLn3Yo7IXZN0lIzIhpU+N8KhkXlS7BO3fjjfH
9XWvnPSLsw9Cg8qVq1OfDusAWth8+t+iUNHr68bJpa+FPcGnL3WcjmqHloNVpg5e
X2eEpxmhq7GdZFZt0C+I/+VkI3tbwGyFP8xdZTgGT8P3SQbirCjurzlVxKKEtlJe
de2EQbgLzsg4AIyKwQLfUnTanKlU+UuQL4ljo7DE7k+ImDm/a+/3uGbZZ9416Ufe
pEvwQ3EF4PCwoblLXnAx5KrE4pUWGT4uuGuM2mU+l44VwITYX5iSnH6gaowRy/sD
VnI/AdMygvFWmwZbZXSKoqp1oFgnTCGc8t3QrDov3x2s+94mfT4tqP85BM0aUGC8
PaDznPlix3ch4XpJ4dElKh8/iwr8znt98w7vfbG9g8MQ8UOd2FVlPeuUACaRcUCe
hAX6A+xuAFnJbvRML7JwNjN8/KHqyQU1pZv/ddetMjU=
`protect end_protected