`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
ddtXksX2+yylW5zu6QL2Lhnb2d1sD00763mmSITNX595NcHTEkwn0zB1Dry37fOW
FufOhVzEJp80NC5qZ/+F0Vk7Ik02dIR0elf3clrjeJRK85K4e3Hoo4xn7YbFUIms
l/8VZSb14+JVGURjfswrIyCUotIzlzVYZ6gzoZwDXIi5gQIBf/gI+KxNXPaKV+PQ
Ufys/12rjO6aI/pPlqSm0hCvftmBcnezN2hk1UeXgOIuKZnogjOsf0iJVX2aOOWE
6pD/psybjbnsNB6kH5uFTA5frkzIzkzl5d9+YDm9OyC+k84E83I/7/j+rk4L2dah
QJOvksSIzN867/4Qt8qYTQ==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="MvBXkzurAa5VTw+1JJ70nePUfoQXBvZOku/SMmg4TwQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
oRtzZL4VJ4iwysPsC8SXYCzXS8Fw2gtZTOskLcDV+1B9Nzn1zTyNtlo6lNICRmmK
ZRVu2BmCc2G+fmzynYlNTnSa7C0Cuel6FYpxCBlOuk3OF2tzAmLAuDyOH3Z1Yjzk
a0aHuoCdIRKv7BrZCdALt03JeUmXKPdOmIlkVGFl8yw=
`protect rights_digest_method = "sha256"
`protect end_toolblock="Jn9CQpRhJt4rnzZPRk+dOpzAubz7omckX1MrFd4p81o="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 3488 )
`protect data_block
gD6l00tciPUa6pDNTk/+t0OO0nC/UTtBwLB41d4inuAUA3i/ALrNyoJVcBnAmEQW
ptbcNp5fxEUJjnOxnedyZEuEBxWRieZFQnkRdF269oN5xiXrpIDRnyU0+w6TASgQ
iwP1p+FC17ctzJk1lfF32EKzdhYMbgdSTVSykvg4WPQ/0oaGwytOER8ekz1o4ydm
sMAEaEs8yZ/KJnbaeIgZxuVP8wUsedgi5hi9ykh0wPM6FzQ6OykxZ/CY9v7wy2jw
Yh5oSj7gL6i1+0gDYXQSGlx5RKAWoWFnB0z6769mTKeLDSZ79m88E6GLlJMiyTDV
gp/UEZ+zplRzdQjgVmQ8oupdDNYlJwrb1vuIzepTT0T3wxenu02u2Ex31KV/2Agw
1CtQ7gXDLGJOjmON/F2kz0PEoqgUYf20tUkHiQzWm1LwoqGtrHnC6SUi/SRpOGac
4ik/NPYe4s1GswL6plFw+rigmOZ095k7UZNuG2ZLjCsbzfns4aLKAEH+hubPcJaQ
W7Hue+7JTDyX2CUxUh9RgTHFDQfaIURleA8J2PpkHHsI2xWy0E0eFysb6HzOP0xy
0tATdFj8OWstOwKxghXcBEh599RFy6PSj4UUm5beH/SepuzrnJJcNo1wTMCrcM7d
3YlN+9P/weHDBd5sUTAHBUmNP5ORwZdGoCaYNg2d5itVRvnW2YOWV9aOgrVZKc9E
71Il7Jep4uaGLG4tMx7Bwzxse3DMqDquffTiKcZRLMOC8DzkVeU3GZnFH1qH7/sK
btTL9GySU+enQbsMco2JpzORhqf2zZprCQQsXN9y3Wf/4M5mEWsVIE9QV0Gk9uWF
YSMgyCRX5U0vBYAKPVEvr9CaAmGWhF5m4Cics4/+lGFIoO1PV1mx1MT6yEdIJi93
DcyGqx7lSzujsxTzgeZWZrJGGdC+b/bTqKjCrARg4baTeKwHbJ/Rc16Ktdyv0GQ1
2FRGT3HrUM5hFWDOan6fVmWhIfJskmGTJwdm+dZZuyRR4hkx6VY/HGu124XKCZPu
tCUvyOSxUy7mUBse2fHIz6r4fjD6dp9Wby/8rJgupffD5M3Fn5vPF/vPXrftWMID
OphrzGVZysQXAEfpgv9PgqXb8sOEDbUtXs9WVOR6wp/kKY7/5neq19nk5qaZBeys
A3MKesEzlW7wWZcMMXBuwgW9TcfE7PKn1XBWtLOZb99m7bBzdr6tlCiFFhsLayDK
9SNhVfO+yf1sAwNfOHU1BFNz3YIQ8HNy+lprWZRtPASM5l4/W9fS7o2ZPsALwvjF
WIVxB3eaQ80gkZNXTSSlqT5iFbKUpourdIlrA7tFUHzRj9vGHdixK9r5a6GgEo3f
W2FGXdq5KhWV4xwdctBGHZ1FJnLqGVlzPIwdMORNk/lRsnXKTpgDnDUrtdIOFZgC
e0/fENYzbznqHAg8lzWN/RolADykgh45afV/9T6QnHJF8tzEjmidrBJ8adUPnxpj
HXTXvig+Vc6e1X9BBBjwhbCfLQGuaRlq0fZqaYQ4I/AGa+IarxF6dbj16wEgs9Bm
9Vhg/FOAdzjxYkEjK9EKRC1WrlXqcqUmRiy21+XepLog0dggjll7qAf7ipv0az1i
IO1B4nG+z7kZOkm38gLtRTEaZaakcJ6ocPZ9hnQqrMOIBkJo6JvuBz91pqvyiwUG
xDCTRpi7uVSoiyva2D/skrDSPY36G8NPkaBlpTgeRnv0c8rxZofGir56tvlxurW/
UG+Xol+32BQKxpJ574PYEKtOJznUk3QtaZ4jEmiWYnMpe2UGR+fjdstNX4Yuf+ya
ZuT/gJGXK8cdRGOyKqoOhJZ8XAh3KEy2ncr7iCujBI9By51GedSnaDoyzAmd/p8a
GQRH9Xc5g0s0Ob8hqq/L1CiBTlfNRkASAJ1gtJ5cCmmZ/Napt4x3Es/cbxdI0UsL
ciF5iKeIBTJEKqAPICxu2uyFsLAsc62g/Vo9b7QsEWjpkPEr6NVOEix5qn+Gmk57
e1/JCSxBib8t+MNDjOXcmLmT6T4vVUg2IYqZgzqMLqFOBW8ne5+mpKhLgp0WlMyn
CWp16Pm67VKZpIqsvRRdCo/iIwkm8oH0HvrneVC81oQE1HaE/YU6Xnx10x/OFMkr
oKlHUe2p9Ga7EP2jgrB0GPEkZzBTWuMPSgXswr5kLCdKd1G1Tl6n0Uv8rGgIlsiO
Gjy915kmHUluVwqSLrvA2IU7Mqxmg0ckUk7xaZVeEZPb5zWxPQIukpYi1P+DEAWD
DopkWfBPerQSeL5KyYlhP/qtQc7wdxSeAmqIfO4YC79PvdaLY/LBYcuxlaHjLhoY
iZBO4bexEGKmn8gn+g3S+0PQchBbaomvyux/tcOu0OiH05uCH5T+I5Z7sn7rpjXq
8wZVRjZQlsg7jjPY4BaGnT3sGAns/ufmfDnndH14wcpVM+Rr2mStnLkuVgpRAT9w
obKWaxqZFig5EnQ+koD6xxp0atbtpi8gqKL/Lxib7ua/sj08LQ8V2uJujMOc5/GG
F3E+hCmbppWP312BnydLq0p0NPEgYqEFV32G+tmxgPGBEHwgsAjJddPzZy0pV4+S
wZ3tjtjMBLcwkRN0iOTgYP/1yQPhSTX/3btNB1CdBWEWgL3aNDzN88pxOXb/mQvF
okv9sNtNBvBdy9hHinkC6UQNapT7iZiV5At3/xVMHI9/mzQJRof/RR8Il4kE+eY9
dr8gIRr43f2Ci3rC1NEgYp9JoPgdbuG8D4+D2XQoMK1SpEuuTiWRuK6Op5t1zBdn
p1RJzea79A2hpy2BbXgNMn79vCiuP8nlbOv7C15/c5bOVn0wlgKytHqD0kTFeVK1
6ipZ4NEBcWJzWvGesdmM/q3AuJ1lekvyb696d9qk0j2I7JaQoWYy33KxcxPQO2Rs
yKIQciNDLz2nj+GLLf4nlyfXBTgWg/bNCxCuCfKWQ8TuREvINXO36T/EaQdUh4mH
Rc6xvh0hJEN5yDQTf1ddzt4nZtq0vMgaUXSPr6G+nQuKxfNE3ZQo3qkHEOMmfLog
X/GFySM6MXrxsFOx/KKOGMnjQbzIxc88zw5c64U5Zgze927m75g+RnSsiw9Qm3BG
X4nq0n6PKe75yAtUIrVZJVVUqxKESbl4GlZ6SgETiC6CbJY/9ZkhpQMfE21XSt4g
WfR9D6ifJNYMO+KCpEjTahu6VTHYIrSbVoT6HSNyTG035bH3i7Wpe87g9x9XFxCr
awRnI52VfPM2RaJDT+WOGap0tGYw7bT7/iwUAiAWqG6A8KMmCrRdZnSwFPleW1+k
mgDwTe74RoxmlKtdzp6vDyP2iIvMk9TEMY+ujq+6SKKQp3IeFAFmNtOcuMx2F2wS
eRFOW0X/Fngqcnq6d+w0b3WvUriJbzsdIkmjRNcKXNG//tpUMilI7k9Z8kRwnVLJ
l7HYE4/qOON4I6XMV1Nkr5lWFKKtYxqeS7qWYE5ekBmH+7W0hKPnG3eJoYUfZTWn
YPsSGlV7bvf/l3FnyRUdxeaLWVJTW0d5+CNRaHxopiWPJIzxshHA0GG2t2VRUl59
ea69oIGx3m75Bo7KSht2PNsDGWAhEdbhYKnEbV9WDAP+yV1XUEK10ywOaDprz5MI
poCyYtl2XRiFdLgEfnV4kJst0DPVFLPRlq2TJCWRZY9buV1QeMNh/NVU9XRZdc19
l6ccDvL3aXNSf3wzCA6EiD4iZsMEiayjkCivfFHc9h6yEo7c3ssTmIwJGb12VPo+
Q4m9JQfbv/De8PtAxpXoCgfWftbmnYAdUIsyhc50Lkv8FvnEAQ91qdl9F53noWN1
MBuPxCoFYgUG+ejmasHcprwrg891qISLZOPjymFZL/3WTQNkh5R6zYfTkFJAncgr
7yMZgUUAlBkw/7cDlXkUmKdpfX75TTllvzW/1gnvC3KiFJ7GhdRG4M1UwJGUr6As
V58C8eGrFwF2izORHhLIQiovVupakCw1IgX75o4KdkaABX9kGLLdKArbX1kpLMBL
Y2AobFLJuU+y0nlqF26SERBPoTTgOuFbZa3IYNzaQ3zen7bbW9ynL00oCdnnbWYo
po030b324SqFSlwX3smD4CBHOxq8vItSY1ysD1LQcruMGHw+xhNWwWgWFqteZ8pW
4hwHtiUKHXM94sKkDsR+9B2rnGvo508cwLhhm3YWpMjUPGGl6vvNYjhf0r+I+knF
pcs06iR4Pf5UB7q77bjVeWt3nWS0XJ9GBPeiuLF58Mo7xSRg42smXLkBXm8Q5kVN
3Swwe/g/cA3dC7harJ8P36avogtCyjbsji7+d5nC0VvLkljFqc9n2pxP6vv6Si9S
xKSx4R9aUttPsvQHoS/qr3HtPK+jS7eP3SU52ndk45eC6F3Y4FxrXZMF56xXYzDQ
75mAklSBlXvoLnkmeF7kduV99O8OGyBdT5bUJSwxBu1vjrud+iXkCLqMnT9kjnho
swl6HP8O14odGSXHwejSlHyV4NtkZdm5CvhLoOky3K1dkvo3uW+8oLDEd/3uEEzv
TLVonLuu7L0BiGjT92WYvBB1YGH9G7Io9jyOGMwd7CZkYhHCxjBAvkBRfSFyOLR2
WghBFcoJ2eTIpx4YEV9dw9Yd913nv6Bp7XV1ACxsXs52CL9VA+otkRDdDKPuEmeG
mskzPWwpCcDUIKh525xkI91jb4b+oGCz+aDWRjkyJYE=
`protect end_protected