`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
ddtXksX2+yylW5zu6QL2Lhnb2d1sD00763mmSITNX595NcHTEkwn0zB1Dry37fOW
FufOhVzEJp80NC5qZ/+F0Vk7Ik02dIR0elf3clrjeJRK85K4e3Hoo4xn7YbFUIms
l/8VZSb14+JVGURjfswrIyCUotIzlzVYZ6gzoZwDXIi5gQIBf/gI+KxNXPaKV+PQ
Ufys/12rjO6aI/pPlqSm0hCvftmBcnezN2hk1UeXgOIuKZnogjOsf0iJVX2aOOWE
6pD/psybjbnsNB6kH5uFTA5frkzIzkzl5d9+YDm9OyC+k84E83I/7/j+rk4L2dah
QJOvksSIzN867/4Qt8qYTQ==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="MvBXkzurAa5VTw+1JJ70nePUfoQXBvZOku/SMmg4TwQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
oRtzZL4VJ4iwysPsC8SXYCzXS8Fw2gtZTOskLcDV+1B9Nzn1zTyNtlo6lNICRmmK
ZRVu2BmCc2G+fmzynYlNTnSa7C0Cuel6FYpxCBlOuk3OF2tzAmLAuDyOH3Z1Yjzk
a0aHuoCdIRKv7BrZCdALt03JeUmXKPdOmIlkVGFl8yw=
`protect rights_digest_method = "sha256"
`protect end_toolblock="Jn9CQpRhJt4rnzZPRk+dOpzAubz7omckX1MrFd4p81o="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 7376 )
`protect data_block
gD6l00tciPUa6pDNTk/+t0OO0nC/UTtBwLB41d4inuAUA3i/ALrNyoJVcBnAmEQW
ptbcNp5fxEUJjnOxnedyZEuEBxWRieZFQnkRdF269oMQtofABEIP+R2iCRCvQtZF
3vmAgX24jBiHxWMWYX7OmBwNWCotC2w+Ay5viA59CDUtCi3yO8aP9Apno3bOPPsC
xQM9+tlIvvgaq7wezhcNu8UHvW2fhSXJyMAKqMymeLdKJa0CtiSb791xWm+N44WT
FaT5LDcOdPVRdxtAwHZufg7pXPMllnn8ruZuDMYP2EPzhHkWdK2/cljgIv5g0Gvy
NtljO/I1ffzDOkFKtb94ubioBrOg4FjTlztifV1U5C8dVaNwRaRD1D70KJavd81l
QwQPVWXZJ4u2YAMeqxfJuYHiIjoxWe3pWjYcSBuFH3JzVfqnielTyMhjGe3eK55+
9uhxZDeQfAKMCzbTUlrmDAUKe5gejZBugoaZtusqqKqG6jocmsROoKARWnR+akCb
0tp+C9pn5fBNZbYQOUnQ0kYeeOStqWU1m0u501xA/gH7EZstYPZtKf+TxvUHAwix
BPKVj4RARRTLgM3GqW6Ps5kkm6iT1xLE7QbGtjF2xMQn8fpDYF5jV2kXGB7tVMHD
jGVBNnl6Xmn0lpZqRUqhSjhTMjifhv9EdRfPbrC8ccm/vl+GfAWfmWe6k2fEDLvQ
+F3W5zmxa+Ty4wN8ITeySvMSmWQtTu0t4jYz8FKpkkoKT9/WzIANiQnCI1QoK6JK
YD8G8YG1RtVJtHA4RsoZeZxSuvCNK1yGm6zofuZy+tBYBk2hTiULKJd12SfzBp24
Es4ZCL95y8Qh0dkhKa4vQixAdMuOQlsoR9BtEZmDHFGiKf31ke18SQNzApC6B5UC
xjLo24mQriR5ol8MHluZRYRkP4kAp9iNL9Sm2uDvoK2ehlCWZFe5fx6CVlmiuARw
j5Nmtw/HELRpdP/RXtcDMqpBMVRBBNgvQ2eyKo5nN4joVaRdOrzKIVjbG8sDtGFc
wAWa5MSsMpnLfFaOUfxFGsoGWuOWCcu4cP4S7r77bArt9Z3dvqYXeqKxE/5nmosw
xUZy6tLUZSG9tlwfj4mkNesEpP3byUOloztJHR+WgSmE2gKn1A1bmDcwzOwPol2j
H6+xIKGhe/ocpKMivg/9WxqG6WSl+NYY2nhozGml+83/eyzdmT9TxT5rdlSqzzeM
xbdgsWhT9xWzwCgzaaJNkr4dZy6+EEdPziDA31uhsziIVd7vnGFWmShl1RP8hr0w
rouK7us+YevnSK6PlS+QdN8p2tuIIYeaXKTSjwmpZS1omoRGYDSDRcv66HGadZzS
btH+ys97AQTRJLm80gRMl5Mf32ucMEV937OBHt8sS6WjvclL0b0HbgBf9E5LxIKX
0Es9RPDcYKcNch6mAGiK0G5+2/b3YQGSEsqO8A/2Mp20GI4tLQzmE5uX5P6cARKc
IEIWWxLP4sn4Xz0xeiRE7gkQorOvgYAdbZSkddxE7LivRFWiJY0lDJw70+1YkW3e
MD2nHtEhliNo3nZ8FZP4JkL5FyK7JP8FXvxI9N685mZlLxfCtsg8f14R/7lpkGHE
+1D1Dg1ulNE4IjZS9K3gryJysQ00rjN+NtnHaPEheii/8ta842xdTxq+Fj9irUEk
LcQCXaM5qV1MQP67mVaqOEsMvfj/5Nq/WzxhPwT3qbhQHQ3zsMP8E2IzpDdY6ORn
j7jmWwBevV5gg+QIMIqwMgtr+M1pGm+nZzvQzZmbkaRpj4HKQOVDoGBW1VbM3OU+
EpVy/ipOPHaBJoY/K4flsLv6IJsZF3Oyz1zeMKxRChLb5Lh7CVdw2pBUUbdyUcrS
twkpD83h9weCFrwhXiJSSfmwjKTOsiHljB+8ZGFnpNFi49PFM80S0FpKvZZwPVym
L5dTC3LQIHQXWi880kAQXCrwBYxgMbLlEBdBjdM5Or4H7V5hbvZ+gM5LpuKYM8CE
Wim6t7YSDENUiKBf1XvsyeEhsmykZGtgWW8tyOOXhUgxexjdmx/av+G2jp+FofMw
l4/nwDecnAeNcKAnzhCbG2U2JKbiJG8ORdDJymROwiMWIHAqI9LUWPtSvvnvvzFE
fe8fFdGutWeOHlfVXEZmaJ5Q2AhZes21NR+sMWnxD1xJOULru4IXmo075AulBIUz
XYx+xnF6o9mK2KLI6GW4tvuz9R/q5xVG9wHGeNV/hqeuAEeJyNN+VHuF/GYYtapA
QpE5QyfIj8MM4PhjV91ldbXjOMFxn430zdOX8GMDkXqRbeTg6qIWHSivw6FazDF2
EPiofioUFvEljDy50goz/QqrVn0WfBNHRoU6QlLk/LGOeBDH5paWtX5vyySFDa4x
JJZN9gQPaT+3X3bQKYxGzfPtgtp3wWDu3g0EgPeemeaQufpwrpN8nvncxvtvTzYC
hBLx1weamdpTcdLgPDmTq9fvND+4DDVS1EIe+L/1pGvKs4ggHSfc5r6Y4CL3K+pg
6y5zdF9B49d5xiRZEq/JqstDvFcK486EIKMF636YNqXjIg6IziVxjzH18czcDy2B
SE1MuFDYNj21yXDbXhjhHRJ595glrvr7Mi6F1wW07H+XMkWOCMNQAXK3FfutknRc
ORF3OYEKJ1/itoVd0a6ZnpuVo2lHmMgt4JVJg0yG01C0f/hhJ5fWFd+wXUyPiSl6
OANWYOzcz5GKFoGqMX0+Q8LZMjshJq8FY4PTxh/BKJrE+44J8CDHZSnxm5yBzVVt
h2i/f37WWvwZncHrRGKbDcu9kK7lmqKnbAgLaCSN/bq7O0tKMsv0YEUhTVfARYok
1cRaiJ2wabs/W8cFbJnDpU/Q9/CN6uCtZ5Zlac0A7BZxaErVnWbZf7RGiLNi6KZd
46DUEA5UVy7EaZnNylCKmapr1+E+7R//GPhQ+vyrEMySyLZjC+RB2yC0pFs8IbQE
UlxqlGc+Xy46JBtT12kjKkIlBQjVM4w4/g94oOoZhBvkyzDA8OBxX0fjhDVJCETG
mR5TXq26Q+DYudDDPYwBl9ToRlFiWIfcs+6MLLF+sDVHfgkEhneMaQ63JrFANumW
u8NU6p2b5APSgyv2l+TKaWWzCsJqYBRBdl3lP8riAtip45zK1n88zOltyEE9nQBR
6pc/XKqS5Eqdjv/tjzbfykTn+bgKjTk8mB7EQFqE9MyteFdJVH63t74HHqQhOiUM
GIeJdpgx1y27HbmcUmmhZ2GztQ2VltPsS2bHAudmmMqSK6r/wUwJzgr7zegKaGBA
kPitZjvTjJN+INlDm/K6OJeag7NYeYKZZijs/yzHpMXc1fOr1JsL0Lcs4pBDpnn9
t2N4d/yLgmon2Lq8v8QQp5YnATMuWYLD/5h+/PEXKN0D7cenpL2U1E0C71gBQp8n
gbpuT7G3CYHh5FC99L+Pcj/dL/h/D/wNGMqRAWk7z4t9M6cZ/6FD0AH9npxDUVee
Sk7DbiJT42xcv6xNjsDC0dxm4L5uQd9oOoL+bpY330LYpAwfr2vasonhKKdr33yn
KaOk19Kc5QixhCSAzM6K7jPyfkG2tpoB9rgKW3m60z7AK6uiOpstc9BLGvNKJaCf
Q1SzzL/qw1A81AiBVhPf3+5cXJcWUCc39wii1We4wIysGFaSQB/K5DFixdWBcVIH
gSjveKGXgtNbXptgyW/EyGskDWh68hdHHJfGFuaCa1CdHYZMvejo9l/s7rLJkclQ
Yius8m6l6pnrVae4clfmdkJMV4Lf14RvG+X1u8kmYpdca2mloV9FmPzzNS5uzFGu
OODC4QO5bnSQaZZ0YlENj7sAsTTkTxmgOp9SzXLOPihsv/Uc0UN+efJpqvcz2AwF
DZ2XYTldSdx6tXAOK7X8RkS87nQ88cPeQukxKI4lWusMQax35OetDxpYBiczXsgO
l978xqvyK1cmDPMYxhxcr8wE9zVPtl+B2B/u4qsZECZqnrqXIH4n7b9WP8BKhMAT
/omglHWhrYnOnnaDBlGlctA5BDF6J69GKpEgEk24SCEiiM9rB1ny/mmyAfeWX0NX
fAP6nvqUO2pCqU9wtM4WIEiCXGsaoGXAPI4WMSkuOC1lZIML91VOOLfU6SBiOxCp
nvoChqhovyWW0Gi1WjcNmyQm7DBhmZwGCm+0vIVp3uETioVKHlRodSHZzZ0Zr1qW
3+Pd8QslIhRFYMfn6aoBNRqpXFKvIapzReQDRyLkyyYiv7w9KGYrC7veC91H7ijP
guAqAGCEYI1h5LiZsfv2AHGbfTWi9UufTQRhqv7LKAvPh5loWkoUOZYiFYF+FE4C
6tvwGGv80x72PE46vc2+cXtTh4yg4dViqCwZg46ai3WBP2KcdtDB6hHWBthyefvf
mVcMN1YOf1FQ/CVZXTFTEdmtLVOAGe8z8O/qrbOskklGTtDrUg+OpMBf1qfgZ0r9
NORCbttyeFvaA5yEX0c7+qD4NQBI/HSTkeZExMaTK1RPvo6gljY2G+n6sm7zj+z6
t8AmTv8c92gsGND5Vo6C8ciNgP5u2pSsATk5MKhO7tR4+kQ7X5fnPMEQiEgKci+N
GfpHzfhl/ZZ60Kh0WxfE/u9Hvjz8pk1wGVmaWixOL/E/ZSFWs/rHqtUyUQc0t3uN
j2hDB47V0q0+aCsg6n0u0i/x65L7XVAcNCxFniMiuSYqLpoqxEovn9B8qVHvVU4u
Ayy7qPzFjLmeMd5pWVVnJxZ+qPxqsZZ0vIEVustpeGx1kImMOhAAxyqolczJuXbh
BWsLlRPTvQE6uRxbqWSarJipagVRPIUnz4m1dFXqtCwfCvOqtbxi2JVZXkm8JRZW
5gP58a3NP9AlkriclVndup4uqDdyQzNh7HfHYkD5JapulsP1r4M6WqTKxeeXf0ml
by5j4mLJ7te+bNy4pO3ws9gxB0biQKfH3HPUuzNcehSxnRZRrAF/nIRfvNBgTPrz
6LYwc1va5qUWm0+N9s1MgS1c20baBbbq6fBC/hLNSwPd/sWMY9LTu114/Hex5XAX
mT+U3iUUPjqVUB5ph/WGdnwoG1JVdOpB7fGy9W1TJPRhw0r3Yy3UHFpCaPgJQTqF
UkNDZY0BGXMQ7gK1V9LluCIY5/n+q9DXceC6aYFgeUSSCQwlIaaRCWJwZr0tDjYV
db6a8hU5Rf3zq9Z1ziG9uYpto7NVXxiMqnSJ/FL+YC2lQpUAcqsplrPfQy4UUVhf
CSLxxR4trodyBbX2EVScWCJcpItzyrt8R7l6mFdig5OluhflKOxya7GFhsfpe+aN
OXjbuiClfke3T4WqQOIKF8RdmM7K23jPFmGVO4BLFgzd46d6yvoSl55PCG3p6ulM
3uPdI7hXKTlgy5j+wltR9ZKNqgpA/KNVu0z3jIVxMPsO7htigjaRbIotsmwlfiGn
j7MjFwOslSTbnlRM/3YzT2uSQn0+MUhLr3xQgK2tBY6SmBulRrYbw8kRnPbUxg52
6oXTBUHZohRwj1AlJrU6kRDCPm35dHWPzIH1kP3wUoaW3OUu1iTXhj6LwiRK6JRP
ttoVFt9qwVsIpdADtdT/CIi+5bc5HgReNDF7YzzAiVmLTBmFbpLIkcxCxWZPlfET
vE1D0APbk6rGPvuf3287CXgMyLk6BoSOraMelKMRTe5DobtfoTbpZ5MezM/BIXFG
xXlX+EKsw+zAMYeynYnwToTzcjl7R416M6pmcZ+r8rkXS0KHwRSfTZq/Zm0o9wM0
iYhCVVDL/3nXPggmIgMFiJbq/tkWO32zRm4PDDwD0xqv80vVLRJhAI9Q8m61dcEK
3BD5bp6EuqJVfZInVOaTdiAUyEjO6Yskwyok31aTBS0CP8O/vY1zimf9kEJEvj5Y
pyVkUp4Z9GzjzmhlwdTqIHar36WPfAGHTTudqYZ7H772MNKyiPZH5NctDEx04DS2
mnq3Dtacl5t6B1yHYfuNony13VLP7XBLpXfaG1yf+Tsg+PoZMC+6+e95EplmSh/P
upu2AMBkdjBUpxpgKt8wayYt24O5pdPp9bWVwzdIj3p2t2eQPDfLg8fa4FXj8dDa
so8tEY6gXQLNmJXbekIdSwoLnFWUuCPHmUkUjzoPvDfjtAA5jZhyhOx+Bt0II/7i
QsmRqL0r7jK8rCE9DLehHdn3hrE8+nvTKbxZuYhZJqQRsF5Wv3ikZgpael13fgmm
wIgEkQVMT4vcPqwQoTDjqUgt+pEAuJZg/TGoHMlomSZSfrnfPUAVPzJysw1GORRp
Nc3Hxvg1CAIgDlKHB/KJF64c/2Wk7keLjINdVRdRJuhPCf6Az1IdP/iz8SkUkmdZ
1BtuMwvLjkjWzrbpdwuHPLzgrZMzSrgDyU4jSa3A9dWUXctMtmRXGTYwAEAo2FoD
iEsmeZRRHICgXmGfEENSQYj6Vql10RzN8+pxSB+8ipgUq5X1zpA2e7MhvOegl+P9
Rheh8bI39yEHCrDSUmzqOgsPStRvrNVVAWlgNBNxnQLyu1WqgKX4JM86M/fR3B3j
ZidRNWNzOsWPND6g55uZct8BMPIwCG1yHAqQjgpqfev24mqJ9eKTMAuqTdLHW8P7
Cpj+2OTL7RR5/YAT0Y+tFu31x92IFhQYw1xA/qU3jFRWO/I7cQXXmf9M1ln2B4Ke
GdRgqcgSp8lm9ffvCFdm0/p6HZhGFhj6eWNgKSTupi9Ykqs+zUdOlFn4xk7p3e//
Sy5RGgi033X9XdtzXaXTv6ncc25yYspTQvYylDnaUGDNtbDbj5QW6UFGKhLeDQm2
sWhIv+CI8Ct1pTYI2qtCAUNR3+GY3SIeLNl77kA32JvFmuVPSVbcoX/fJUOvA/Tj
iWHW+Y3z+9cAGCWj3Cbgu4p3bjyn0slvV8vP+7W9m1DIHTDWJnsjlMVgzr56fYV+
+ilZ6/PImCj1YYLsQoeZ92uBfvoIsNt/EhOSMlXoIcG3b6RrB40OBSn1E8rKEHPL
Sk1vco5sUcyW5uxykA9qu+WIJnA4jSzS531wOVRMIyTBlof16yvKl1UxH680Su7C
eegdPNrYunYO7qkxMp2dlEp2RkjSUx/U0uA46kQqmmyKMbdZPJQxPq7sRo88tThl
ZRf5eWmbdhRMeTyKiUCRQZpQdyk/t504i3KIuA6OPqUxhI/XFPinAr04RAYuG8eB
4It90JIplnh7KRJUtAYwiAok1e9UD9YokH2ESFX70olhMqja1jC5ajHVd7JnLImJ
pqQKaA5d+4spHl1qo6vhf1NqL7S1/rYn0asQ9UyLea1naho8TWpObv+Q/xshHy81
h2p8iPepxVx/q5Y91e0easCDNZ1FJXtEboKXbbDhah6dPz+lHAhXD2yfjYfozhCx
+2r/eZ/DPvfPNC/UrKzJ+CtzQ2P5YbvWew52py57JhWTWlp3PM5Nez/HDS/wjl+t
75aYa26VUlh5SR5WkzZLlcqZTPCLKiVa7evDIghfoNBdbNwQ1bS0Ge6Af15EzvAI
XcCp7USePGvbgW8Yvwp8LJA5Pqu+GRON2I5JIV3Uv0cE8Cs7GUkbekz4H/dubIZz
CMxcMX8nytbxuLZUdJgscdzmP4tYjMSaYpyKCwXXfaVCH9Tc4PggW0E0RZsfDHHc
lUfke2PL3W8kHhg0TG2a1hopgCbAJVOwk5a6Y9oTXXKtUzFNspEJacHoSPoLpBTQ
RZz7wtwvKjW2gUa9gRj/+YnYUH2lOlAPSmIk+L0o5RdCbwDGqQtXMPd1eE3NmFm5
vVn1Sg97xGGD25LFSqblA7J8CVI5x8zmsvcfI7cvFCCh2Ckwx/JFUkGVhyg02sRn
/EFzlGACh1unEwbIIHJ/jY8t7MPFrXozBfd3Uv9BHOYor5nCg4+3a15ofKhgw59x
C4SpeuWxMqs/pBRKOeQz122EGHbcJnuemJpfs8KmqfNAG76RTi9RRpB99CNhigvS
KSVYEB2u44TCxf+TY13HbF7pyOguIpD03VqspeIn3m292mbozbwYu9k+obmtMHlr
Cimz9B1PwfpBzaE+ZDcTPdeSwv1Tv9hbO/FMIzJZyKar6muBAnlwDOWKP49HbGFx
EoHHi34Xldl5iLWU7smrQaeW5Pehd9I6fDeSUe3z3Q4a0vBn9PE0jEK4ki5JeoX2
HWChqMdD22RVEPiin/mhiSbL3fBYcEYAuandV7SuV0lUjyuuaPcN20GAecv63IIc
fkFf6JPyy24Mkp1BB5gNOq6K78zldLaV9FqqZ4c3WgtrEFuyQc57wX2bu7i1hQyU
kPXeLjpiLec18jdSLEQUxKNNXvvn4YtohED9l7Mtm4cLqx0OGu8uiUmLqaP9QDPg
SzsHMMCV6PMghHx7arLcgdZ5sc/ACqh6cY8iFw/j79e6RgW/n5Sl4MUyuQi5SoZj
bDvdh3BeC9M0HwpSIH36IUe1M3Gheb4btKfhXdySqJDRilzrVh5Ry7jfdhBD+G7Y
lo+O0S/enp9dPEIn0BcmQGixmSgWbbdnB+yB5ykwsYQ8zHZmNnC2PmRDGxUL+8jz
oI2a4tnZkS2nqqxLzv0UJ7zLkqtj3mnPqM32GGTboV57vwbPQTQ4L9A5es0f6KUq
aTtBQs7vzRn5hOS1nKLawgK3A91LXcuXh/2FImeg28q9jSsCaPCLzY3LTJCttrit
nGJS9k2O2fGMBI83dJaiL0nhNcQWdYdpJA67NxYZc23LEymTRH6cTxz/ReoIVRy9
JN0L5VgiSnJCiIs0bhfioBaBbs8zxwZ/WlREVDRHtsEI0N+FttKjuDFcEFC7Zy4c
enTaj61dYW1pzdchy/Xhe5btXHpdWAxreBeaxJDc4RD15LaILtEwhtYbWp76zzCD
2139BUF6BcK8VC6MkFk1Hzo/31HFeMMcYwce6/tB8Ynk/9XSRClXahdbs7uz6MJW
QFyICBESzAip3tmuEwElTid1tbvV/2RLkPzwE1azdzqlgITgje5Quz08N8ANOu+S
8UitzMpM94WShHQO6JneuAtTUWZpW6wY9z5Du2NJ7ll56A+oigh7sxtQ98AJ1Vsg
f3xP7DuOMj4LdWs0qlWtCYTZ0YYCLzLoSs3/eoUOUA1qJrjXPVjCAqCUByKT3HSm
f5oFYof+0Em1GcjPs0APtvfiOULaICv9yCxyzfc6g2AyalxtgwLUL7vVVyyqnSyo
5Aew198ss99W6gLarqcTPF96vcy0nzEjm1N1couWPxZPoIK8m0qA/N4jvpLH+53p
eGom5EUObRrYVqZKbC0dl/ZN79ZyNa8STjrCewF09rAiHSCRhxRW7CpAnVUh7BxU
czeFgCjP3bz90SUEvJS/Q1Oq1IcsY/tZssoJtQyGZ3zRuRlUZb1zYewz+I30LO75
8eEYs3hgRV5AlmpFJQHlmz/cF+csP59ltGQDwH5ukrAllc3g+EnSEM1DlYqrdtLM
AUzy8NSzDfeeDqcbsaGuvwj+rT0cqffh7q+xTz0JJ87N5XhfdkonOdUZMAZyLa+Q
47P+XLPK4j/Z6DeZW73Fy3O2pPRpjO6+s46UNYadB+Gdbxg7TUWWI2TuLLSGvQ3E
22sly7ftpW77bdu1zO9sxxeWbYwRhjTSeTNjkPngKK/mKUoXYkx9f+n4Z2eWe6cd
nfsYrAygkPnTK8r2c537rjUAl5BbXW8ubPTMhDnfBhbEDzPvvShusxVsb6XoNFR0
1E4qT4g8VB6b5nA6+/d1qi1bq8SF4HbeIMFQBUXgn5RUOyFO+DROYZk9XfwUMvWT
8g8eKmqH7lWYE8Sj3r4nxzp0QFNoCEqIvCez5/wUZqnTDu4jALwglEqlGSHtC1DY
MXd5F1r5ZXFF7LQFMkh71eCh0fqwuiN92jZkP/FoC/uLtqDy687kkr5F7DrsvhUk
NqS5I8BarGV5YPcZjOZ7FhsDiPsfqg9HmI++erkvCcw=
`protect end_protected