`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
ddtXksX2+yylW5zu6QL2Lhnb2d1sD00763mmSITNX595NcHTEkwn0zB1Dry37fOW
FufOhVzEJp80NC5qZ/+F0Vk7Ik02dIR0elf3clrjeJRK85K4e3Hoo4xn7YbFUIms
l/8VZSb14+JVGURjfswrIyCUotIzlzVYZ6gzoZwDXIi5gQIBf/gI+KxNXPaKV+PQ
Ufys/12rjO6aI/pPlqSm0hCvftmBcnezN2hk1UeXgOIuKZnogjOsf0iJVX2aOOWE
6pD/psybjbnsNB6kH5uFTA5frkzIzkzl5d9+YDm9OyC+k84E83I/7/j+rk4L2dah
QJOvksSIzN867/4Qt8qYTQ==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="MvBXkzurAa5VTw+1JJ70nePUfoQXBvZOku/SMmg4TwQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
oRtzZL4VJ4iwysPsC8SXYCzXS8Fw2gtZTOskLcDV+1B9Nzn1zTyNtlo6lNICRmmK
ZRVu2BmCc2G+fmzynYlNTnSa7C0Cuel6FYpxCBlOuk3OF2tzAmLAuDyOH3Z1Yjzk
a0aHuoCdIRKv7BrZCdALt03JeUmXKPdOmIlkVGFl8yw=
`protect rights_digest_method = "sha256"
`protect end_toolblock="Jn9CQpRhJt4rnzZPRk+dOpzAubz7omckX1MrFd4p81o="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 11856 )
`protect data_block
gD6l00tciPUa6pDNTk/+tzLxvdHE2s3DQL3/JqqujQBC/Ei+vcAB8wM3doqg5vTg
mdfn9XB1bLOis2CVSfu295W2DNwHfMSTc/8BhCDRnTlLIX0UCJs9Za0+LoM0rMrV
T7EjVWppbP+Em6PkVKCwlmIQ7JKaifJ+Y+kjw9HCGboYo5074hY+K/CBbfsBQY86
vD5OGgtuxrSV52NK85qhYx8VcipbXrwysZ1z0/BU/1dXH+7nlcfr1mNnYw9pfuYr
RU+xKR1j0CI2UPjUxwQYxVkHNoAWYltwEcVIEILKa7jNCmmEodxLa0y3COT50vuu
0n7MVdmdycjXNj04Gw7t4K3Kop2i+utRFfj8v088q9u309TAzsWeVRTwt40rleum
+/OZ0ifqEW++bC5zqXvROTI4zhvtvd+H5B7cMYFOSQqMujsUK4/GXq2VBznoGFm+
nPrmutXlHtkUWkDy/t3b2XWguq4o9JvvyBZIfqOyqGZB+5wE/6zODq3j/UgBrz7X
vdW8Jmd7pxLcLsoPQVkL+i2Oz8p1MA1XFuVV+hXfq1sqvhXlzUYP79+mJ2wizUxI
cH/zYo31vi1BNc8951n6y5IrtKf/g7Tnz3Oa67Dph1HeaaMqTdXsrtqxzuAe7SPl
wFw8iYSLcCdA6c5ekR+gXQXCoLv6MB9m/DSCZ+VvMlPs97DmfHsyLWJzXtfR90hM
MDX7fsvM00xvzIwYEfEnabvS5AwcrMbBizjYxe4G4hVr8mlfDHJ3LcpWfYn48euN
3SBgKlrRrUsOEmsd1cbGtngPBgmBEl2D/Q3s7habLTyYEkFR28xJGtiFBM2z9MRQ
S+5kj2/oKQpU50rUYG9HWe112qDVdkU86Axy3vmGWVYRgL0e3gXyUolCkvdK7TGM
KexhFiJ5oD7KcrHjthOYCrQHhCIVJe0i8QhRTt9R9PkHiNB5W+/4xAO6Cyp++wXy
8gdD/ZN2BHUO3KLHuv4pJeroGT25mV5AKvgylW6DQmQVObxgWRPqR7Sm0yYjpCad
DB3Q8DuVKCeUVuu/PktST+vASEb3VS5ky5s6CTBY2m/LWi5duLVGzQIAv0ZYaRNy
hiI+fMO6QPy2Y7kbuH4S46UE408ea3LxBWxmZHqt23p8xBTaq0K8o71vFoNj4cIJ
zbFTJ0H6ojTcWvcsZ6QkTO0bcjnzQxvGo0SlPW+O2KdQgGbgmlHH9HGXFt1OtSl+
m6LptBZ2mc02JznTc0oOKWmMdAEcrQxaQaxj8Qe/9X7XTmCLZBqW/bThAJaN9cye
nr1XcI9bj6EpNYe29ltvfu5BwWnobOG1K9YNc/F+7TrXeaYtCKbqNHQFQppgZBD+
AuA9XG5dgs+nQ4AoQpAhH9AI3aMG/ylCTlIz1/QcrfwUj5mur8T14HD2y2T9hhft
h9nLPxDCIQGMPZ0fZAw8NWMb6rbPuHdAv9f9tl81dOIWWJQHFmZIJbu850cIM0Mo
H2SSxHLW267oHRSySzYizUIQ6Yi6Dg3ovWInQDYbGddvLqHG1zpKLfy9R8HK2mYj
siBLveQbuSz9IDDqiHATxQ8ik8e2SYUixU2PB+XA1ao693ZQ9kPwSZdk7WK7d9s7
/A3Fzvxy1j0kQwlATFQuTRMt9HZRBGxY0erKdFw3Zh5gzihjrVbhXAq+DhC/tMbr
f2oBQO/v+2tjyVFA6OkUOF+FbCjJSft0WjIEce6qw5iL8KBWZjuMBEmJUD2M9ZJH
v77AC8qEzWJTF/7ws/0Ak56F/CFTWcWN3G4Rxj8W1OEhxCzHhW0SJ20v5i0yRsIx
GQ5ZOCYOfWMc4htjMtEtVwd+KoZzTiQhVgIShc5SvNScZPDpSxPFiFmqXPSp2yJb
IrhCrTGKwTM9MUdbLjXjlgYrrMx949J4cgjW4/LO1HRD6802xCPvkhetAnMgosYQ
fUe59tv9EvOepXXAqVw7i2xhFpiuE8F02RVRY3HOO+BymRtwO0jXBl8q3awrJIHj
d4RXP/xLSpUXFmYXHFKG18XhQDTP6+ly9uE8tS5G3flA5eyDqmNvtWxkCrhZXeDi
81oD1mXa93Dn825r9Y3TMsQK7VmoU28Hl96LiaOuA7CYK++vktfTv/6ht6GZk9Sv
nvqMUYfqWhzu4kT9sd+rWGfa9awb3qO+u816hfFVqXeFoUUWrcT/hH+PFf/1PFiH
n07tBvHjnKb+n33LjQWEapRadpTDECBHCC/FQouUQKb01AMkVPNWsfU1a1T2Fl/A
No7R7F96k5yXv2R9l4irRdfRZnIbyvGvwPUca0GeedjuKSvflCQE4JKib8xUqe0w
79vwmprKbrrMBIeSE9L9gJBWO64U/h1CgLuShf9cV/afweJio9JMSld5z9yG/x08
BPCa57zZWQk9NODnL4B+uMspcMkOlsPa3IXTUpaIRdV0kkkE9DSJpfjrNc2se1iQ
z4Oirpw++Bgr64PiuOnC+d/ZLaylZ69cEG08Uv7ssHvD0Kgx2/PsBFDj1svZHXIa
wfldquiIxOYyomaJpJTbn0RvLOuq40MvXgFaYKCvZYZUUWeU2lLsTqd1kDDIH+44
lM+VDyuaLo47VOgo8QZ8xcvKk+4Ep6k2wnVhxUw4+P31k7366/LOKGGz8YW4t6Vx
4+ktsPf8LENVL/4/xXFt3BaC4saLXWpd4zyvYn24sbcK8c0FXb3V3v/d3lGL7r+N
wIQOcS7559mrl/CcW7X4qS3v492S7hGK9tDduHCfJuDhsuJohneOhkYN/DOUj9Wa
3sSWXu9Ed4NrD3oq4UQZyLHLCQXChz1Mjxom/DKC/ebQuFgcKI2RHRhUsgjrzZMN
8tvEnBHtZVwGVm4cwySqSmTvMPfejCzKEGR/cq68cLCkKJ92t+eIkQXvg9+oC5/P
q3F3SAbedXF4d1YBlT19Tg/6zkUFH3wNDsu+5DkQl5hbHptFgNU9S0ndKCA+x+oM
2TBfdR3nsKkV4fBuncvzUhoqJLslz/r8fXXobSU5u38H4rNG5yDNwJdR88xIrvUC
ZMtGbwKjnNIW8NQgDzT6qQDvjTV/uz4f7mJeAPfjkglQc5E92YRlTdXYgS5QanWH
o+2N20932clA7lQn3CGdPKj7uzMCHi9YwChr/AI4Arb850DEsQppqYsKER2GP/EK
I2/DI3aZElk30ufN6govEUyaF+nkMBkHxOupJBnSmvM+TSO3JLGb44Nhp1ip/pHV
u1HXOn6SE1wHJBP4PHqEiO4i9sDTeoVBqHT+Tc3ZIqE3TiHQnTodejTvWJ+MB8po
m2SVXzU6memrWlOUmQcwwRF9thB4pqhoBFdO9Vr0IdZWukj0t2YZu5VG6CpuQqsi
J/0xlNgcY7j+f0oC3Sfpz6rneVCJ5drrsp68XM0TpQHWM6qKl2oo+HyHzoC3jqxh
eJyJ40bRx0XeJ75QHI0f98jw3hKAPw29+gPXp8ifSNNl6LV34fRx7+/GTVNl97Kl
GtxE3rX78//ctyxzQTC85S+USKx80m+EgTy+TanX3Zc6+oit1rzEzBrnyHVK/YSK
7UDkmkRVTpyM5Fubv6ACjyVqe7UzCG2/8uwXMsSPgm16h2hKIDwXa55c5W9aBfQ9
NGxcZl62+KKoeApML62LPvHKPEoSh0+4tb1e+Vcjj2oFyrSw5dhEl2hHpoJLFGWZ
I0vF/EJZjDxDWL2BW3xjF++kgzEDfg8K/KZ4sNptluLuGpSir1e8zeP4tA5YVeWn
22qWeFezL6PIoytm9uXnFhvwjXWiJWbplUxcDQY50UxyNoCFDNW5yvExmUFWOseu
Js1fvfGH+FGL3q49o+ibp9uU1k4+EvYTe3V6sz6TDcXwIrxWyVW0yNpiG05chv+C
IZ4EA3eDrCRHQi50FVw8Tu+DAS4yA2gYA7IhqCF38A1kT6bPJm37MHQNPXWYoe6a
cnEZ6flsShqj0+qY5j0zLwjy4PU5h37aYLfkt5XWY/9pTKu8QEQPPyaK1fM+zAcg
szo49GpupkSEIlhyDPxQsS/Gh5rwF5pTygALW1s7xNOWjrERQToqEC9znAjGE9qo
LwVKKEcwTmQQfuV5KMTTRuEVjN30syRPw4q+1J0c1AC7LScebQFHLjAb+D2QbAFA
edhkS2pwVQNnVF8xbW0MwaZSqnVp+Pmssodi43yM+1HdrjfEtm15XM+q7vKR7p7u
K3nR6RPlZvc36AEjBz2ixb3x3qufXTEir3iVFhF3cTsrfUfKAvVrk13ochfIm18a
hLkhzkkh7dcH/RsTchJE42p3VD2bklEwYlLkozI8zp7mKW9g3KxKByl2Ev5YKXhm
9IDCFLUx1rkgODtj1uzKgn2RaM1gw/AmZ6gKjKnai37cPUFmOo1PS8R0GvOK+GHX
6K4XUKpaGVs3xVoAVIFBBrF49ZU6nKrgK31QBNlD67UL+itB8/tZBDVH6qvHYC/P
raSL7guznKH4yi/FhJorrEbNxe1txz2NVhR8CGYRPN54tco/P9/Z2EVXutDGYQBm
uhdPs6qHu7IzvQwubn9OqZqW/zR4stUZZXGHBrZHgy+Ds3usb3F/e/lAHP3ysPSW
tu0EdzsE70WTxluXgG/OVYiS7ZEkkPTxHFUlh895a3fchniOUUqKMd5Bhd0cEyA5
xZCh0npRg/EtufslSkNpK8s+odNlAhAf+Zi/nRAenJ2vAeJTC6WfS1alRRP+4Ixq
fPM3XElGiEtvSB1bH+FvqDkXgUcefwLdqoOaRqDqjSA7l+6bnur1elbMMBG2/DhG
A4r6z22oin8fn4+v5WqnKnKWAY5mnQMSsKZ2lVuKclXD89+oZqlECqacLJYKKwe5
6VR4BUuTLiyCNKnk5/R7aJ5gl0QzPcbPov4FHuY4tM5yrrYcAwuNzbRKOu11p2Di
XHnZBExQvOJzDXqpaVNnnZspjhGEDXzQt9oYpOKn00Mlf06xexEaxuLf3sSN/AMb
Cf9H14mXNfdsUF4A7HJDpTjB8Hc2hYtyybT49WHgAMOi1ydguANFOEvNM+a42uBk
699OfOhU1B586USoRI4p8zi7d9VMbs8hNM51sNZz9AP8gUf305ajcEH9pw4lbJRT
arq2Y3QGUJnpuPKOqFZmGLTLEwa9uFGr3rO6+3i18lZFEpUPS80RaNI8k4E9yEBN
fzCPuo1keyfZHXDe1UECiqBB0tRU9R6SYZ7kmnozqj709yhO3MzMVVdPg4n8YOCk
BF0l5yP1HbQKAaywZIsF0agBxIdMoMz/22UGnxy1dRqQ+c0yJad+NfosCifcL/9m
VeK6ACv8cjQk+9tr/vUvfSS75Qsy2SSb679w1hKPTXBq7YAUQy+MZvL5+XNN6lhS
XkKmodh5m828jt9GGiQgHPlvLJK5HMRVmzbjk4EF1H/rljNd4Kmzqpbwh78yIB4R
Cta6CInFAX9BijdpSqWfB1slcuj6Kggj9VaMS1e3yBDyTUe03d4Vg0o+8EfVGLv+
5DkUlmfx3cnzXzGSm5l7+YF+67hb4BwUweMEKl0QGRQ7yUZyyhIGxLifhLvaWalr
K1F5ljqdE1j8TzJn3U3C8xZmgNTFQ9QiXpka9zkfrhjYUG1D9R5dwNPOaKGz1va7
0DXwFh5/nz/mXRagBmpr/swf9+Igd0ieMHYPeBc+bSbaRhKB/Yqqw74pet6PjNPm
scj8etEhG44YKZdck8WlOSd+YYSCDd3iJfJaCPVmDD91Q2hLKuby47gXathzCUJj
4y/azH+VhlKhW5rAeCGA5eU6eKEp+Hvbvy8bYRBOU18S7kfJoV98a19CkIpOiHQh
cVS1wRMFWkpynaueaKQLNuOypZVJ19asssqTKqfs3KE7f9Ebvm6k5b7elLlhmOQx
pWSBQA22mWfEPcKemVZOWO+qarOpjiBUdX+AcE7bHODTAN1drcwqFH9GYGiepHTd
CHOz+k+eElUWKZl2P137I8TOGQjVf5T5vuGDfKchao2E+ZPupzjzpOdkfDmb6jtV
AawFSQig8tMx+vGHJg3OgIyWriSJQGRrZ5BfD5dXSyu7Qnzp8o9dzfgS3xbMmv0+
ItK/R3ju+Emt4Al+HnmOMFZleUEgzpgn+Soz4WTyrcg40h2FnEjnPtLWglTBmiwY
lPSFVs/opyUbvwodjTOes6BE/UeW7ULwhKOVKQiFk3lLfeb5bDbYOwCz94abOp4j
zBUpta68Asi2zSTW74R/GiLSxwOJMildCbc4zHr88dIQMnBS7DW6xOLOeTW8PNDh
PYXGLr5g2CCDyDw/vd/OBAjrLVaTccD5SbnN6sbGkCMoZpYYgCjR7Z8XtSV9RLhJ
+X8HnAn7z6cBz5F51ESqplkVGXVWoiOzZABCerhyugl+jvfYSW3sI88CtLcI8Zpu
YtXDol2DA0mgNrTskpQDnPom+EovLcBKbvoU6G0m86rVOfn8jEqa9rj3X+AZRT0g
wqrr9X2TJ0syjP8xy8ANaMS+sDfRedOGZ02hISVbCTwDP5sYoaveiHac6gXdvkbR
bSe4Gu4X5Vh8mm+f8x//4cqb5ZfRN6sXncLyym/wTvuxLSbAdnLz10OHC3omjK0Z
MGiySR5gi4U/4EA41z6fUEMcWDeM0NgwmT4mehlRxjczdYFIoFT1NUcY04TM291c
88g7JhGdyZOHFgSdydUa+OwWqoLuTRZQzZXb5DKQG2POvN3gL5PmVb0oQiT6eqGm
7/sK8/I8Vw8KKyG0WXFvdN6MMoxYKQBk1A+0uO2yrM49C+bdVc6WrXySTey5cssE
vdA97V+37o+epssRu1ya7uO2z27XPO7/CwUKBeg5zQj/YCDoxBqwA5Rs/b6Juqvv
6SR6QfzE5C1wgBygwJTKa7TLPpylqQKNRjQ+srWZGpcrXm+ugtesq49Im8s/3TPZ
P4lTXKzffgKOQnJ7mhsmP7zvFncrsKhzKPudbQO+1mzNfuiHQtQwjHMN6zeAA2Es
CCtL0DtZX1auMZ/EqBuuStsY3K5ogB40aufYkIszoTowZ4anp4xkrbbgobbPkAWB
zoF7PwGezxBDti0erHgLa0KlrpPxWbuGlCEEsnLYUcJ2aOrxCeEF4tztR53ikVqK
ZUPwZGIzgxpgyggJkG+8FOpCJiLEPx24fB6DFHRDZf7OhlWQsta+/FlFDSQEFJsY
0Ry1deSnOwcX95ps4ZQL669TyvGFQuny+Ou66RlepnGM24J/tO1ybZFegaQC9tJq
ZPE94+H7+yaVEV7LF1TZsnlTx/5uw1N8A5dGqA5elG3uq6USkNaxRnsMrAPVTnFO
6qvVcVt+yiEoedJTNjkBqFYvJZSjUASaE+wT86Lw/vOzmB6iTxolXYheZKmhd/B+
mho+2wO2SgDYf2Af44aRPLnedEcfuCwNMUcOk6od7sTmXEsXgfFTchkl/XOMWs+4
jKLASEp2SecbfRG8/ZlAPPAOt3BiwhAZL86N9XmssY/TgVd9bXDNMpamqCinSJcK
cAdPQEEuSkeOFY/LxGpVSe1pPS27XO4+I6Q0NJQNuqjk1ryFw7wRFAh29ibzOP9g
AWqqaWhd56m1ewGHu1hTcwN/A3r2bKTs3BfWE8XrfXKTp2YNv6cg9tNmBrGrlL5J
D832Oepi0GUAAclT2fy8cm5QbvU0Ti03V3Zd75lI9ik1hWkmcwfg8NM+n86sojq0
2E0NwZSVzPbVEMkaRteF7zLckbs0wmH+JlAKhjQUVjvZMARxZePGOHInwrPdqqRp
oCVak+XK8RqgvbQX/twFaGRN9QjbTlbgm0kUBsNZIKG/6r9VFpHaa6+mEg1epnJD
LTJUktkecXG7nhTDRZj3j47VzFKM30BRU4ccJjEMYfVx7Gu5tK9k/H3N0H6bZ3Z0
TklDqZ+XoklRt15OGnF+lRc8spV75zQWa8Zt7KMY1U2U+iMTUy//y7dpHU0PYPmb
aqG3hYmHhSLAhjR3L+OjebozDnDkjTPafg47yhAF3uzdUgvt7ciEktfCcGQQzBPK
fpRY8U4lmf6x4WdPmOg2PlWDn9OlvYYDIc1gGZPhjoYug8YDlvAWSej2MJLGW6R8
+JxHhfYIQZfXUY29ETyNzxuybcQpB9nqPa47kKDkVK6HKzOP4SayzitpZzkk8CS2
ps5h0yM3zjXwuIw6UbBUTJxJ26POiQ23lJISO++Bx0wGfaeRjhZQ4v8GXwBzFMAk
tP5dNf2cZ5pbUYJpLHdmRbxcjMKEEZldUhUNm8ZgLvmFGapq6VPTIh3NGeO+yWVL
x8byDZ62/i11/Nm42yuCILs/r1sEoiNfZn1JagjgfgCLRS74Mbl9V4aZDMP0A1TR
Fgf17uHYK4RaaNqUxGC5T6bJMg8BZrK4rzi7j3wgGGhqbg8D7T7wzx1/B8Hr6ZGc
AyOqpWKXyyHihPD3I2QBRIvt7MPHYTvgtyxe8KdGG17JeDKvoG39RYkt6q2norwZ
hcSf+UhhWwJbTLlIO+K4F0jXwIFIaB2zqs53+31QYfIHRjSpy5taWChhNQOvVj2J
K6CFtZ5mGO2JaqN2LpboW8P5ZJz20Q/bXSVYN2MneHrbZpVuHfnQP4j2UQuPPLdH
6hYeBnED/siEYT1U4QuOJMCqwo4/icHeIF3SN0tl93vnca5PqXVh4qAAgZUwwyLu
j7yccgcBWpPTFsy3k/CgQm5qP42GdWA71ZZ/zzI4Cf3PaSGo4xjpU58WLUD39H5l
DePY9feUtF6syF5U3Y7mQyWCaGPWjZM0Kgrlf722Xz0c6GRw0vOz3jrrAEpxrORr
I9NAN+8JJ1lqm+zXk/lPhH1wg46CRTJVMzoW6VjAhDjdxwwXv5qR2mSjD9oGc3e4
LlKHnhyuu6Qv/h6YtYaGmxXcS0sqa95Eacsg8HP6a/zY0FhylBPVbafQlQou3Y7w
0k0VqZZK/v2qZvfte92N+9uD2vyTRcM9+mSWs5CnHT/ZYCusL2fbld+cV92dRDae
JOb7EYFKjxR7/wbxc5nob5eEvwhP08ZM7dpoXrFERG473sqxPruzDd8/O8cLoVU/
0o8RD67n/TmZR9QE+u+jXQ8y7vQvezO/OKjEleBLNSADGjoIVOeNk9sTCXnQqTBj
Loel5nZ2LXYfGNUWoCAGitONNDorW8aEEriyCjERWYPrXFG2pPB88ByIKuEj49RD
uBf9dVUiFS3bSdfbXe4+BaC4PvuCtB3u/0pr8bio9dl+wmnfdzAB2ZSzk+zJDFns
+C378hivdqXDQp9pNEbtHht4tTuZc2BqIkFm9xyIKU1UALhf7zkt/tnqd30xMERn
ZaqJCY5+rR64VAHg2V30RlrB2nUExmErQ3gkT8nppTme448iStcSyvfwBicWwCs+
R5ztucksvcUwx/AlqcqKpM1fMERJkpmIxRlxAOcCun8Bi//X+js0IMc3Uv5Hv/8c
rSEs53tA3i1Q0LSlu/Ul4raOKXYVi7ovsG/cRTdJ5pxcaN50TtEiG7GRysuID/Pm
qn2iDvX8oyd6/bHIBlXc6MjWpqssdRt7XtkCu3fE5XHf/bbQeM7PChIHyS9MRf6i
daX56JGpbFt6Eny6e9FfkVedALV5ds3fKHXltjGrMlORa17gwwdnD2lv0vgR+upc
akeq5Xa/dQ+ZW1kuJsk+iOOFGqrHCExNsFTk0IYfhhYcRwiYrnGdkUlCGf7prQbd
5Np0CRB4DEcL1/fQKsojRB7C0FcqsIJNoFFMEon2RkVGRls5J2Rk1INSsd3Y809r
mr5agIYN8pTDuKamaaELrW1vZfunr708l8u5nqepBlHJ13ZzAwtgdn3L4TobZx3Z
2LjuG6YiumMkFozUIMzIMemYTSn+FLCPNT7+75tieLYC97rY/uR847xxtcUVu0XZ
XNDSXsl3MaDuo+K5h1493a9UZ7DejG5FvQ1zvrI64g/6gJOL8xzrwi+9XdtUwNKh
rdmL/6KCZfPTyrIcz1cgHfuWnxgoOQP0tSsUoDTzf5vUprSpLKRjDMmkleGBAEgZ
lwfnFRyprtOlYBRIhl3hgcrxPdgjztJ4BzWjwnCeo2d0s3lkm9QVByrP/tEOm4Ge
hhSrg6qXzaHN/gMEoOvoJwsNdcr1pzQOOiLoIFg2DSCGz0qlex65vpCbCd2MOIjS
QFUE71W+XVaYVfbzXeh1AzcQLhl7dRRm0ao6V+Q+dQzF1B9k9xyGDm969H+7rVEB
B2tvZzt1MDriE8UV/0UzTGnMSE64UfPUBMQ9twlaTeG7xzwc08rki5arYl2rMsNS
DRww1LSWKdmK1GYJZkYd5Oo+i9EKtyYMsy33gl6gdktxV52+MpIL4qsUJUStcxTd
CFxSv9pn5H26JiWkw9bERXeh6jJLIGu07Y5AEoxtyXFiuwIKkZb8mMQr3praE237
19s92fkqKtu7dQZ1pbbSSTnSah58nEpL8/tPsbTZtJ89w/EEJ7KKxXLkyyo8jut4
yk5yOdU4BmLpUSAJTi9mnpsaqlcKfWbhxEB5JeRbWkCIlh5qsLrxyojtK3sroJcS
L6y7bI7YTKUTqtSvsRCCzwIMv4Gxl1pak8aYzM9hbxMEqj00KNz3iKK5HLbQbpM2
bGN95RuqoHsyN+jsSHiSI7gPdFO66y+2FWBJlbRfnPTfzUstSZoFPMPPUI0URv7O
Xl43HqmkBbgLaQfCmA9Ye4d5EVt3lsnWSLuqAZmaatf8Kyc+35DS5RjUXQraRhyx
qWMGwRSF32/Ow1oEiY8a+ero0TfJMtphIA+suD7FVy8lIffPVj6zzci3YmKGR/fY
3QBkPd3nWy+6NHufKdjOQ+rPMMhdB4f1i69BMaAS7MITncjh4Oz+WdpBWnay0NjR
LaeFlwldtuuWZT0imnDvAqdhE/rddTVDapDpnpub6TiYzku7xUhAPob48q2JWAr3
pjAnz2FE7bxLpekMdrdatDjKpY37L+egbKLxaSTE9fYdiopQT6U7HwYTg7tu1TIE
WIFKU6hFN/MFHIn5SbivAaJHuVNhwcDb99ONyyuwLtzRxrVUETax2L9WkTg1P7/+
3xFZ8FjxjHTqKvXAzV8+BefssqKCw5Hzs2Wl6osyDftdlTW2VaTSJpBwKpoT3pdo
AfVQ8CJEZ9vzTFvIU3zEYSwbCNbWJnzaJxh13sFqpfsKwJR6BdK/qg7AMffpeDqc
LgcKtn2e4irHe36+QHO3NvJ9rswd3jEzTHOSXYu4PL+7aC0aG0A0rTP5q3o/si8/
kDsfgshdq+1l5Qv9LSdl1vqy6CAiYS/ZByJovkkGJu7Hce9cP9xdlAKfRv67FtE6
74SHI5zVwxck7b1sZsHbB+n3r3R/W8C/+AphEAEEOJR86bTm38PlVEwDkrDOdKV9
vohdTr/j99R1YcGDKsN3XXmgLpuViS4kTd2XjMsDBZoBLxMzsPpuAd2MRNrvDYeS
h8EaJDNzbmigGmpufpuwQJORk6S/8dxLh1UM89By6wL7vwpSsmjD+pKCKbfH2wZs
iJH30DlV30cpfTH0sCX9hRjJBFJUOd/W4GJ5YStRjGAM7F+qqQ+iNNKm4TUjkB9X
dVlOe3aiJ3w3qCrDHfIN5QcfWGNUEFCLuKgQkWIAyN6L1bzxdjenMBgHy1zr4g3t
3xzH+Ak6ik+8AoPoQnHneJgv1arYi1WnJfKCraauJ5DNpLmKCwgPdpXqwq/c1Hmu
RMeJkVgUiKQTzJwRkpe6qF+Gy/V7Ok6bBjVP2XXK/QWeM7DyfWFTN43xU12QkQvX
sadsacJO8jrC7LgNFXyLsPhaDik4up3qAzur59NmUh1aVjHEsUeC+kMVUWU4W4ep
wN0yZbANcFnhcqIvW62bE+LOCJEUr46h8tHJnpuOGR/fGH2h9Jjo4kSuTI/8WcG4
Bxi9a0cYUrxL3kSkUK1geMMOONFtcO9l/Xm/n235d7Fw0GN+sPNd7EEd+/CCCKBG
5fYr8z79yawfDAq3bA0OiXAvVy5ZHxnoigqD3I/4N9JjlOVGBtuZMe+FLp3s1AAU
e+HEpS3PJSpYRD4CERGNxpri/7SwSs/iNi52d+EEyzznBF/xxeTIEerPxs0yENeE
MqLyrRkjggy4CNyhQkSKOb9iVQj7rOfuQmsxu+U62blvYGNcl8QToFsYS1oBMjpT
hNS2VD8YDiUveWJv/JjbUGFZX1RNWDNE70qEfbaMZVIKzZ9s5hbxVp1ELkgsg5K6
DBgDtv2f55TbgLYq5/88L4F3lgl1bHqSqfv3ZsoIRhn8gFjY4Hw5Z/SYbWGjtc9t
jQ0X01JkGKhGXFnUSuCw8stllVmNxU+QzIMTLADVkJyUuWudDi+1ZlaitMxbO5Y7
/ZwJdDE2VQxZxJb6sciAQymeLzCIlViQksHW4hpL+rURgw8f6Lh3c4v+5kLnyFnF
zM/HisrokiE8UEyk3JUQWSYlCDW3UzX8Ehpbu3F6zg/NHyC/dNeu0Xo5UZojmkH1
z0SjHlUsi00PNzGH5KihYtqyxOy5Dn68IaqdnvohfWeW4SZgrkbUySquRv7IyyoP
0n2w5WL5CEOH1PH1gIx1D/0vy116DRC43RqW5o6cZzS/JBnUlzt0uk2vzZZqvNew
UruF46kTeRfpBaQ8NIUPTNqgzPuYGqXARrvaWQGjKbujxcDqJtXLhNoVs2QRT8o+
eBTMIKR2fqn/DqV2nIZTOoQ1a3VtmNgdfG5NzzpRNOL3/htG1o4aU4p5wUwqDkCp
xMVdnTwE9vnxweOdj3uR7lukRTYqMF/ANxyu3SH1r0IDDWikKUbltArImucyrKS9
9ZSex+IR0cj8Ihuq5y8b4xMXkTLw4HKzugsdYpPgee69V8GMVvefSWvaODbLmPfS
yCz77FDAubYH4ai9eyUIKpQkN52eTklkD0XHr5d5WzzUvfJTuqyg1LC+hlxNbKnM
HXD2AwhjGQylpb2A2uVcyZ7gnoRN3LwuZYLAFFEw15kGjTKlpmn9Ck0IoPL4PRjG
4jEbesaPy+m46Em1o4+X5wj4rx0b8bc4hB/IR2KZIAYOB7QrNFlHF6iPtpztzLZ1
zprgHCGfEj9jE2Qaz+33qL5hjS7uaW7UdvOf3fnqs6yHWhwPp+Jr9IwCu3KgiVqP
hlWDNxmf26/Jl8aC70HyiwoVPBE+epmARO6u1SAu1OCYcxrDleW0jI1C2wVgX7v5
mc5+PZLGjUMh3MIPiyUSj389ttF4GFIfcytzg7H2zhnjeU8eq4nQVA9grJqFBMqh
YCFv0WE0JepCA1yj6hGtfwX25LVVUvw4cgI5heKeJBslM0bTGPLRIjTxzoO/DIDu
bQ7aQWNud6qWn1jFGgvmX5bigCjIziBqrfLlnLwt+z/1PB9+OlQpDE9PaKVKUzZg
BX6cH0LjAT2i0BYIwB++8laG0Im5lmHAQUg01gx7QSOO6oCD8eZuTLZ/Zxxyi2B3
0JVRXyYQBn2PtdA4bXxrHBA34dpa8aI32Ml9IWGUGqCDq+XAV29wz4djnMy0vL8S
MYPyYr42O7pnjd/8p2HxMF4cdO00PRLiuY/2R9/WZmW4cp1dXZTBtxqwIqZMeBfa
YJycweZJZOKeQQuXHDOZX5McXIyesulv+wmkL6DmFEIoy1d/gcCRsIh8CSEnPkz3
oNBArop1zpBjsWyjzytlKYePGyzh/V7DAVqpuIeCccAvruyr8eWsPlaX3q26dsja
nu/UogJSNfWn+B1A/GpaP6m+NZM282AljN0Av6W/R03sRCXFLjy21VbkpnJUnz7/
CaBkFLXpx4k1+WNuctK6YoQWV/kQ+QRRH1ZtSxQebxp/lbuuvDAWDOHOd5C+RY3T
x9IRZDBGHE5yWaEmhhaUJG+2BLPkhrSkD1u8QltaD2V9jdZcQ4MXwYFuCRmSSm0F
WKfGIxzeRBZmGJLOXEXqLAbKMycIIHgIPtvMt0gE6/IAARvpjTyo4qiNSFv8ahm3
pFVdElyLou/h32oKoLm5q3BUxmXLkRVnCxlzUatzXL4jR6BUx1K7guz9m/0gTria
aLjL3mdb01WXyQUqgdJKjTUib8/xs3tDzPUQ6VMwJk4/0L638L9y5ZDHwoxHa/r6
cqZTb5uSj8HuT6g9oVVCQdu9Ngy8i/3HFjoLQJ8DgGavsdWTXk6DDSKI0Hi0QmUv
+a4zpLgrnP4bKwJvdyN6M6W/WZlSfk3XTRiR8Y+j8yjD5LxhHogbmi8CYY27Yfz2
5OQ8rXT/MUYA+a9Cn4MDC//pMkOgdzGQU4ZMCBzeIDgGL6TP61VwAIPbUmqrlKWl
EM1dLzLPder9tb0u9pAp/+JL2gWk42wR1Nj9bzHQz3v1UGzKso8zhVcVy+YRYABG
+J9vjhPTGAL0mQNtw6n8ndnt+TIqQg9mx27UIVJhAeUfz/bce0BE/FpekDHNPoUI
GKhs1PZBD9GvbhDzntEJPRuPkPQj5nXEtmHoP5DAQn/GSei9IvrJPgor+6xOOG95
LT5X7KU+ldApToLR0K3U3CQtVYt9AC+XWHEt2VFW3Nc7C+UhZ8NQKfDIXlarYYWb
l9vtZeX0bC71mMRE2in14FbsrU6n0G2LnPNe3dMqr8NuJ5mMVlUn7jivHmuVoBQp
Zvg7ZH5txV/G6jD2UdDJ9YEbH3YOrjp16q/vGH/3hCMoNoX0q+tmGEnPQbC8a47I
FAJtzCGvkNjArit0t/eQb+EPznCLKIs+4Adp1R4v7DUvP3nQUiBTRSpNwKAYMjVY
MHuJ3cHz+nRmZaMNsI7X+r5MToG30AR1Amkqhoe/91UnujuAJ4SJFJ0fUQNJx+p2
3hic50JV+KhmgEoX8rfQIIQ8hh5do4Z3MtsSNZK2n0ejxJsZeIiTvJk9jc2GVLeW
Vozyo4tnZ+MNWs5MxBdRElhriZDJ/X7YiX4Nyr/sSjIpVec6gXQNsCo/HWSJ1ELo
YadZcaOFn3q9wQzuaiI7PeyjPSWe0PufbwSL4IlU03ZOaNhmfsXv3k7Khm9MPlhK
GWxe8/AIFUzJBDdCLGoQxgKAZPbARvKXA/KFZ1MUPLhgRtaZuTwuTuwYBhr7N0rE
XFZ/86v1jL/JdplgIo5++rUnHGAHQSlvRt5tlZryhDlTACu3ZmOuMMUw+Rojgrc2
OlK795RT2M8kG6xca8uSe1sIMUbPYcuISS86bv60+CXVQhMU0SkSOm1X0+7KJ0Q2
mmBcXgRQ2Sqmm7CeEtkPbwPM6I07/5XKVlAq+ScifNqJFBMzlb71t6mDmFsfh0gC
Dn+Gu153g+buiDBCMxNq7J8xqiAvmSs1oP3IudDlmQ/ZTofI4dz6kSlUZp6L2lrT
fED+Ad+lOvedA4mo5EzY9y/z+7OuAYMVmuy32ji/MslbmsiWLmiSyzInXG00mAn1
AurDtBIoN06mjsnNqwJpQM3eJ6ExNLstnr+R43D8ELmb8H9gQJ2eBhUd5zf017w6
Mk34ZiM3vzAKUwuN24HsK4/pm5UUARGG/EUkDUt6+Bm/vPP11BlSrQwQfg+oQ6YZ
NZjJLSK5uW+xc5QTa7pFlEz6WdVmW9b14dDMz625ZJzZ80hTbQG0gnQXqLY6Wgf8
mJO6kDviDCowkg5R/3sN00MB1XV4v1P3dhVeNfcN15CuOUz1GSkS5IptOY48G5Gb
rTWo4bF6SMGxgQFIlydKgSyutDOC0LHafhPXP6VxAqtLtQEw+BO6evFQjxyEQ9A4
6O7hW5f6mvmRnQ/oU86apH3sKKmPGyyYkwq1UOP34Cfdrq1mdmnyna1S/va6U2/q
nledP+N6W2SMXgzqB1AxgKPT4rylHMC3U1MJ3GJEhDqX4CgWUS57NuzSJtjYpzT1
t5CjzYlr5StBqr/5TMac6oKf1K/yHHifoHUqGY69wJOuKXnA4jjM7/YXUzexrxE1
RF0ouCrC/HtXrd8ZfiKLrF8cpYZY7V4eei5I4b2jv1WatvZzZFup9P1U9TkUqL0v
`protect end_protected