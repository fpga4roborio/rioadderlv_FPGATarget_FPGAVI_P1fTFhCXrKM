`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
ddtXksX2+yylW5zu6QL2Lhnb2d1sD00763mmSITNX595NcHTEkwn0zB1Dry37fOW
FufOhVzEJp80NC5qZ/+F0Vk7Ik02dIR0elf3clrjeJRK85K4e3Hoo4xn7YbFUIms
l/8VZSb14+JVGURjfswrIyCUotIzlzVYZ6gzoZwDXIi5gQIBf/gI+KxNXPaKV+PQ
Ufys/12rjO6aI/pPlqSm0hCvftmBcnezN2hk1UeXgOIuKZnogjOsf0iJVX2aOOWE
6pD/psybjbnsNB6kH5uFTA5frkzIzkzl5d9+YDm9OyC+k84E83I/7/j+rk4L2dah
QJOvksSIzN867/4Qt8qYTQ==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="MvBXkzurAa5VTw+1JJ70nePUfoQXBvZOku/SMmg4TwQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
oRtzZL4VJ4iwysPsC8SXYCzXS8Fw2gtZTOskLcDV+1B9Nzn1zTyNtlo6lNICRmmK
ZRVu2BmCc2G+fmzynYlNTnSa7C0Cuel6FYpxCBlOuk3OF2tzAmLAuDyOH3Z1Yjzk
a0aHuoCdIRKv7BrZCdALt03JeUmXKPdOmIlkVGFl8yw=
`protect rights_digest_method = "sha256"
`protect end_toolblock="Jn9CQpRhJt4rnzZPRk+dOpzAubz7omckX1MrFd4p81o="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 15344 )
`protect data_block
gD6l00tciPUa6pDNTk/+t0OO0nC/UTtBwLB41d4inuAUA3i/ALrNyoJVcBnAmEQW
ptbcNp5fxEUJjnOxnedyZEuEBxWRieZFQnkRdF269oP4ITahSzD0QNuvEbePo8to
oJu1o2MsPigYKhdgr9wbeZkSq7wQm1wqHKN+5x9SE99YwXcQ2G0MIRroW409T7EF
GjGJpR9hMtdTd/N8eOFj+IepE349yMwECyZcpT3a6sqAa0a3cbNr1OqvvRVfSvZc
l8wBJm6EmloWMmYfIYHf26BnkY8sdncAMwZX9dMDqX+IG0F0Pxfr12wdRynneWRe
8Gn/IvYuBeXygeU0bIj+4Qa7r73m+pAKfZbaHYBRGJzRoPHdqPgNTYT8fKseU7xa
KqQ9lzVaER/T9537WhE/kNuKN/Dht7ujT7AHfCjppF/xW6X/sISfTI4FJnHeLHvn
y1Eq4SFS3LeGM4Q2G0NtR1QbQKJjOI1eB/bqhNOfNqV2SwC01QKSDwWAI2jiQdVn
2c+4mY3ImMGiXWhkPM1IcMED4dP61HWQlEkIWkezR02DxLqClQhqA4tUw33jzCMG
U/xe4urgCf9Pw47pxR946sEJuO5ZCUHYQhlYXbY8wE3Ba04+eyX6JyJ2cwThh8Vb
YhcQyj+8yNcHpP1ESL5RhYk7piUXxfBAgn2sKRhNtlb7ci5wesc4PHU+flA3oSIJ
jBZOf7jkRnjp7tUu3KP7VbxThZZ4Nx5XKDant2aeQ6sXOJPuIEk2vGIEsDhRBFeS
OesOxYg1ETnd4qlr9clA877P8g6/rbUTMVYaV0glAPheRPZpunFazA/NZm4qq/tH
hVhyQdTJSinPI03ifP0JI/Z2qyeyR3Ev2ccoKPBNJK7HP1Ty9HvMosCwCWIYRkIj
dn4id7YAjtmxrge146e91HkfO4U7+/6wocPJ1aa4BUkClBD/aY43Lv87yyfHUki7
tr9E1s08SxtkJKQqcpiqq5w4PLDw7FqNjaEkaMts8Oo7mXufWWXOpKqu3ATl61uf
zpZW/7v8C1HijRzeTL+ebRB51fvtTNpkNhC0yEdomOgBAARbqKFwYv7IvcwnXuV/
qodzuOcWKBu7r3LMwUKOJ/qFkIxlERbNngsBPlBVsDIkuwN/2co74MRnJmJUi6wo
WjXW8BZVA0hwm+K/CdIC4SnRQRTDSWGFbTbugPBF1C5xyBycMWiM9Zk5ufihx4Uz
DVA84DLHy7ijwO6MZjI8sXyUCecM899isrO6cRgFSMDgLULxzSZlmmq5D2XsqGLA
kRv3uz8EF6Z394RyvfJsigpWTfFZabQ7tSfZKqKTDsAf/ItMavTTNga59f0uA6QR
ywLUvLsdHYEX8CLCMoBSH5LxCqt9qTJgm1iXYSm76LLx+q96wgTM1UzD4l50un0O
ZGK4FEq+hqCTtaEgQSZuKRId75v+cX13196DxpsrV+c1dn9Rwe6pu74jeRdhA7BK
xhD36bgB0UmX7fIylsI0gbnVAEW+zHHXk4JO2WKlY6Pg/sI8MeL4Euwy+y2n380L
JrGEVXwKZSjiPzhEokxmF4ZsLSfOcIyQBbrWZDYFRXyu7BUyWD6qU/0F8MOvQSPi
osDsw9wD34YxGBomu7dTOJkKZIsyK9qQTdFG1dZgFB+JX9VJ2rY46sW0w6rN6gfk
ZVrnM2z0q5J8AUjC+3xW2G09t2NlfsDUSYTjtpYwWPxdoWPFnmJYIRwgaJVVs/7g
EwvGah4jJSme1AamI/7d1I4Rf83oIRVEaNEYVP3Ok7MMc5G7v6i7AWwAd2X2Dh7s
b2FOMC0b5PVMFG2RXVuUs5NpdT4HfkNY5fJoVs1I5QLdfueF9u7LyLFfrqRsPjin
4W+PQiz5LFbfolyryZFscXY6G92I0FPUIbJ1AsclpaSm0990cgqs3SYtTd1LJtEz
YrDeyXrRPjILIbBxIb3ZWL1pL3qCNuvJX5hfKusMx5yNZkTLyMpa8pNVIqNWJ1iu
60NR4dxUMSDmppmlwWb9Pwl2KaBr8s3sO/aXhLy41U8o2YWMt4sL47+uD7GjNnOa
fLYO8KpI0b/EbFUUQNRUJvj271kQFlSjS9FfpsGPnczg1qrQAnzUH5uESGbiiuAc
R4LXDYDvC4uxkMl+XCRCZGDGYEY0AuL7D4jcUFYYB4RIHe6JHaJxTYEwp3e5R/lK
l3eGneVoXNz25hxTndT7UmD40A5qwJw26CYBTD8v9mtx2iAZmQ9Pu/Fwqb+ZX3Oo
mh0TWl3L4wUjnS2Fsa+fdFSJjkGPBeLq/mzLNWEOLQWiw4ibxbyjrTu4Mxg1ppHH
SwMvmRou+BbtOuPHDn3xoQSUZzuRYxwAwOr/rAO9lDT6PEhcJteYud0RjX9T3WU2
ioffBMG9c5wOnX7lcGyqEg6Ga4cCy84UcR0o/sgKT/pL+HRhRztW6sXdVfgQSnVE
dpU2Xo+jWPuHs5UMxBOgTq7bfutcN/XUexTHmBIZ18iW71yCAn8Ve8KXterDICHn
ahMom0nKUUt/Bw1fu9EVc+GhrWYTR4iN8QkULAvSaCFmnFdi8F6W/vcB3MTPDssV
NCAAMjmQ76sZ+TVavP7PKNaLpdmqiBrub6G+Fc6ZnNtc98LZxP1dyt3GSyujLjUD
JNakH+x2Ob0KltUqy1a4ha10Ib9p5IU887dPhitsJLJcGCVcjzKLr5ch9fL8HZZ8
SjXAJ/SA0Hec2XpNp7aV+/7AoNXSmHsPLiD1DoHTZsADp2vRV9TEYmsS40Tcy/U+
yNwJzQn7vHCpcpvVkM1P6ogj2JfCpI8xG1GfZDBpNp4GYS/lOlvKkQzJVy0jpQRZ
uJnPrhFrtna/6tlg0CbtL5Ydn/D5ygvHJCyHUXqYr6X2cn6Xx8dV2IT4HEQH/YWJ
UkZHbZfTOBiRbMKmdeNYfzstO0IZKEsBeLA7K4BNyx+WcX2BLwdoCeWEw4FGMUN7
Fe8Oa4WDcuI/1ZgVScLsfgrMPfGyrfpLzM32oJIJdLIez4VYPXlAxeML1jda+Kx+
YVnRJ/OX9Lr4YKTOkKF1tXMVvIgaaXgK4+koF1pNXAcV/2OMhX5QtHkoUbpYnzSY
NmVi6l/fgQDEgaKPz9RQfLMACgfChO6O04BZSyzNQsbIPKTXvHgqBS4gebsaG4hi
2gDKPVqklOiYc5w9CJ398FyNKxB3KoyzbdKZ+neOWMJBdI3MZvBeLvlO0aK/VgqG
BN16UM7NXMmWh01kGINVx3DgusB3nisvPwcrIjguz6eN2+0h4cn3FUAgvsK0As92
P1KmDHKhkOgyQRHKZTPako7RksGsP0JfAtRhzCZiqYK/0zSskb5r7nQ/H/+uutZE
kGZ0keEInzVJJXgLNY380M4xdoorVGQQ32ZJqTVWTZ/E5YUAyHMLgadRkEqUrOZX
teRxKYvn3qPZa/cPoC1dFnvTgKjoH89dPKq1+Y/UQ067gYpiuezSyYhl5WCP3t4A
rDHj5Sr690MKClF1kTZtaHATeG5h/uV2YwtqHR9ChEp5V085dZqiK/9yJU1TcijW
G0MRGZbnZOgPlujI+13jEe+Q4iySY46tMTwmEcdE5QCZzTD9m9/VR75R32dGGUA9
mU3j/aAbUnZM/7v6wdWcvPeKcIEALsMKRmUJkqXQNuF5fI/WtRp7TcAbBxdUh5rz
JA63eba1T73YD+cxiKsSHaxb5At840KZtt2pHlnFQ08p8slCSQpMWFcvuXoDCXU+
uAtHy8U7I2Ana1UcTEGENGLTl0QCNLytrXkTZ1/B0PN3LOHf6Go5kGDTCPkd/vNt
EK5MjmqsBNxeaiqpjMsQSCgNukApxPJr34vAipyr/A4JuHQZrnzoyg53DF3hAmY6
qovmHyR5qaJgEwl2y0Sr1cRWeHc/iBkH6nP1uSjEfnz/vr0GiKNX6b6QQ3elAdEu
BA/p2lP19yNF/7dtmMXUC9xwMUxuimvjL5u5KnUIdw3kFXZnUqZAM8SJid9J3e6D
WlhqwJeKWAw1TQhzg6NWHHJF57kzHgBGHizxeF+1Xt2/Vw4aVEQe260PD2UaJ65z
7g9yMVJQ3z6pJ1rRel2n2tksYR0rwylzvA99cEOccdDnIMWcCfHYsTX5X+bS8f/O
rqI+QvKebK9pYnBOAgh16p64G7ryJ5xr/HHl3PsZnRoOTFXBArbQVaslMS8irD/q
Pp5iEbtOK+9jDVgCR7jqnDuR0SGqNNAwQ9qAQiMdY/UQudTmXsPSQUK76mSIcisB
fUYZqqzvbZzkXK3LhtzKGjp3TEquRvufW26pXxnAmWbf9yNbnzT/waJuvKkk1gbw
Lz4G3K35831CD4+1TJ6ogFRfajblK7pkEKGGJDFMolYbp93UMOHFyBsGL6I2ZNnl
d97z4c7q38h2ZUwLcxXRXM8rXVd0QjTcpAJz8Kd4mUoA6Rb6chxJVqLTFnhrRPZn
m6IBtSQkuG+phTWQDVh49D39hsP3fiVKIKoK92sBXkrUGzEnIiNVPD2Gm1JAq2vv
OYevwFznnc33UjOaHLRtHNtZ5gxLwK/Fe1MWtadOJxVh6DHDZqGgSIfl3JsUvp+e
aqFrbpi4RMwnHlb8Z/shlIKufI270Lo1Pj/fZhvIvf469aKjfnnbNbIbWcHrgmrl
2iRxku95ExvQ/XpTDlc+/VuvgWl7eXTwKYpDfLOWgHL0yEdmDhnHpg/2y0F7d/ru
OobsMsuzSanOQqfmauZHe/4fegg6rzSr9mvZjTSMGD2/DqILh7WbmXFlrQ/PKgbb
/UoVQZbNZSy2OcubcP6lzRypQsqOFL0ndbtTcY9mVihVBAImEE8K4WdWJ7Dqz1JI
W8ncYFy78wMBHgwTXqSkmJQ79abrFZ1lDvmqYpMpaQlvqPjs1ZKIzFKvqMNzJHl3
jQkGxo+pVn6NeWfARgrKFJG2FSw4f3RqoujCByagYTTNgsXQM77qXb010MElByWe
HrFBKW2P2JTQa4HDIdt0PH3JZhZBKoPMXzBbXeSFNeCMmCSrQpKB/drVO49aohX7
2JvyBhOeqchFBqz4MTSW9+D2VIPOFWzhh5KEj4WsEV2hIDoqW2xFvx4pWKXTq46s
Wd1Zji7jIOoc7f6cmtAa+d6YzArqGJ8xazvpxvYCX36HP7DNq/oKQWJHnWUWgdGs
Hke8Gbfm+1xuEMUGIPCQ3uwXZdB/6iVVmKsmkaQQR6bDmrDbp+mKZhfjh8DFcV8t
eTPyR/yZ1fQZLJOtSYjeUxvSjL1JUhcbu+N3Z1USC2oUvYp5cjXSSgkoFfj8E4RF
22bFfhdVWLkO/qaOvjTwbpbWmTxSzLCkDEggty2rHzwj1vdTpJA1bWThggYtsSZO
r86RRMBKlPdmCuMTfCq3nmqwGdUG63KTD/2eeFPh8iabPez8p5NP9iD6OgCYZuPS
azbItE5EKyoufIAqOOcx+J+JMwWNjDbfaC5Uhr+h4wM2635mRDgZEz5mtUMHb+2d
q2oqlu3PGeC9DL+r6pAqugD+hlVyqbAjPG9M19nbT6/bkDMmTgCGa1T5RWApDJSL
3yhYpSxzAzz0jPL/bq1UWuFCcnLpr7zgQ+eG2m6r0IWjq2uD8bBtjSlGM/dOLKJO
Xd6IgtaShQLmKDG2um6BBy9jaGGlg61yBPwHpnk2dN8FHRLfsZQ24zxGQQO6hwGU
2tm4+gqQrzDG7M5zw3XFnukQo3BZXrrMbwg6PQcvZSSkTHsq/ZxyxDQqJ1Sc7YdS
rkGiiymCiZVMis33sAO4QmP56Sj/D5WohzG5EW76o4y1ron7j5GDwnSdSmHc+IE2
/I6T5Nd3qvVN+pF977tnfaMPyWEfWtmlTinjdKYnpzopQ3b11/QMydEG430lxiWK
1OpF+YYp5EacsNtc8OuL8u9EKDUEPxW0bkpDGcZlDo5wQf1UoROUFBYdOKJhmecY
RQ0981gJ6KVaIm+BbZ41BFpqtG6Ylg/eFajarORFOyRkaMEANAwsCMIFCjdSYcKW
FPsOsGxTjQICdwGwG+EJbQ4PyzuPP3Hv90iplv2VodxAFanWn7h6rtNoUrl3vF87
eo4pRYeGtAFRyhd/PCIHspYTMdQFi9ZfSybwlJBmjH7ZweEHhKMyCRO3XWtZ5nmZ
8pot+wyBvamfyUiadAHJFMY+ZUneMRHU5d21TRg/WES1IGaPeLNT6Uo9Vun3LQWQ
oT/ikbiftTWhxcG40f9gmjnPsx7+pEHZ7H/JzFigkWwcwjjaHLqP8oaXqfMCHafA
N4Wf1FuI11MxnA+tiwBixy+PqQEGW+yRe6NWcGOhFZiWnMLnzEICTVo76U32onQA
NMzc9cn3bFNhXRV3hkBUQ7T5KGNfxJ8mVvmEpiPdZ9mPLHSn0cWF1rrF7heKgbr8
Dp8OdvVIz65BjlOcp8myostmcOPI/xEjFvyfGuEM+rL4VGNhcYG1Pg50I6fpBRZI
o6HGTUCJNaVOUviked9CJFU1Wk8OCppPN/Yo0XHf9ivdmLGfvIq94CniyqjbUpXR
Q1+edFwZo6nhlrJsHB91H6nahVsQGlX5kSDgDMqY0ejpsd3yeFabn+Ao72W0aaE0
E7iOkg34FseOBjI1rQ9+bx6Ux44qh0movMFYtO0HVlw9wAsR+3KfROifzBS48yVj
ik+0gm5D4GGKVeHEwHKgvnt7DHxdKOrKz3FI1ILIQmvEJwEVzphw/hqckdTDhQH5
6s+2UhoFK2j/GLCSLalBDOrmfBEQDcfIy3XR7fYoyGsbLOeh5Iv8pFnm4ICGZCyV
FRY5f5xaiHeUxcYMslbkA8HzU2pJmp9voN+aRdjX6bHqeMvUK37hPcTf+VHEezNB
Cu7tNaeN9Cw5vXCAz0YxQtY7dOSjFVTK4wuCXqyiMLmWGGjML+WWXOH8RiDv1Bnq
/g2kmzE3XNRoO7mOb2nkJPivScfcEtPLvlpnN+zVm6c0auxpPvnJkYpzlivGcVcq
XSz7WyUjnZDn7jobrRRexmusvT26eTyHug8QL/5pDAiRKNmnqJw5IA3z/189x0Vr
yKW7LTPP+tkyiSPRbszDqxy1WB7vmZglT001Az4OdirTJu1r6SckQPLUeQc7txdB
XkCtZQy8OPvD8mpWkWXwnZ4lVQSB0Yfzz1hdLmeJprTOgxC/j4eXPs1DSL//a8P9
U3E1vdoVNCI00fKeLfepfFxIZaRXTi11rAIekW7MfA6ml7edfCpiLR9TGglFCqPj
6laE3Olvay6HLMOw+SnKXoDRybnOfwfGszSjcGeO/jq0PtkQBgU+WwY2IVJTqaAU
ishpET9gO6qAQIqQI8ZLbk5hZw0h4xQYhkmboGAw8YL5quleY9rBpTpbFrMbQQUw
gZ/BhPWxyT8wy289rLxBe7JqIKONzmLOfYgRoRfiD9jLNqhVcqKChERSYcexw+Oy
0xLW1H1m1nVGXjKbzT3JJ17N6Wn9Yrgp48igf2jnlxwhJnpox2kfAgOa7oSk2Z2D
iTIcLbSEtLnkZEpmV87xyoyofszKfLpEc3Zwels3NaSO1STOtV8ijnUlTePUuobB
JZMZSLrU6+W+dXDjA3Gamelor3F2Zh3YdZCYuN1RvzQYmNa6W9hJRaSO4GRWwmKf
NNBOcfmzl2XHUkju5KRks39MYvwebfc55tC2x/bymLY+Phm4iajvmk/x/PjpmRkh
eEwPtR+zq18hW+BC4qkG3u1TU2XpaP0CkbHSI2Y8DVHuIa6SymfqjUowDrkJ8DOX
sLMMMYN10lWZVRRU0RxoO0Mj2Agz8l053pEoC2L+tGzBv8gnGgQXwvomRlytnqiI
gV+x0iHiu0lqxX+TM0vfqzoRh6+UvNwTLOlMTe2BCnqUw14cDwHfaQXZwxzDnQNK
BXR1YYTWkeaDD3WIOZlnsazz/ZBGI5ajLZSRavhF9LTYcaMReDH1wI159GcrgT6M
p5W8EZNKsB8mdybKiL/h7w2b+bAnXzujJZIVmuNDmqnPZeFfxMA/EMWWdHewz978
Oo/2ZxbnoH/WaA8VyeOJs/Jg5ugctZ1GXVykUhAttOqjSOunFs10bpeP1Y1Iz9GJ
dzi8dE0gu4RrPUJ8SWFVpa79qCO4iRw+LrCrE8A+eBJ81H9pg/uVzIug5Xk/EjPC
pmLk3/osIUtUAS8xTARBU2aWaIOYitWs0RG6gSoROQ5qIzSe8utPZs80Tl6Asei+
qBbiVutiMHsNNPNhz1voRTgl/74vzdqZM+sbCwQLB5rTwrUBl8ninOGSqz5qUlse
fFjSq6BlPb8DDLqD3+u+8r7CWOb838WOC5kaNuDnSwJSGgCZDT7BGEeKnxA3YVxp
PR7P1pM1ZjXMtUiWiBI69fj/pB2UyoEotRbT6dK9UFIfnhGwp5FfGR9YHS9mLD6v
u/pXgQpYXzUElFaBgb+yQCkaR93DJSxmP8zQhgs6GWg8uiCd5SELEJeONBm1THUw
QbYhr1wGPoydMu9EUuL9FU1TCH0vexaBlfDrYMwvVjSahFNtLrNCz4+QzS7TR5to
UVDv2Ry13xM71XN9otzIw7QebovpY4eK3rCyWvrngKsAq5seuYfdL0b4ovxnMPaZ
0gJ1bvv5X3tDMGL2cn6YrDRtb7GMOqG3qZdRwiVrkMJFzciXX0opJaIuPu5yfe00
Rqu0zJ32aqeB8Ba7xG/zLj0LU99Ow/2hq/Cf/wtA+K3HVoQoFa/WNFOdoFykqNVD
Htz5rxawHqsYucR3ycwawAwpzNuPw2/11Bbb4DTXeUVaLaP18VTi2FFh5Sa8vBSw
G8lp3iCdGYM9YSAHLvyisqKicMdb+FZpU8Q7oQIIRHjuI/kP5bcQAhWfRMr8jbJC
FCT2sDZcgzjVl/sgwbxDSaYJ2DeHnIg9g2EHgv7shHwrlRWK4PvGwOEVeGhp8nFc
G52Dri1M2QQi/HG4nXhI/pSkb6+sPEpV/i2xnVv2mo89pzwmHxSiFmQAaVQqT4ni
mAO9b3++p03LA/7vR5NqA6p1UFlZ69r3RgCtMnr3z0eiWtSznojDY5xdiqJ2UKDb
cwsoMz8z6NelqzE5cyDznIjwiyv28WvGgUi8SlzaeTXPWMf7D0KWgifTGXl/He6Q
T+pm4Qh3YtK5TuP26mHKNLtmSctrUE41J/6KbmGAk25jiOX18q8Z1VcNS1pDpkJj
dt4MMBb2tWJ2D5PqtRHbk5fJQIIuV3ZK/f/+D+/lSOdNGBENOW/sx2JYLV98lcpg
TnVydbhxouIFb+CZxmVRd1y4Cnwao4q2HI7MnG/v6PcZzBN3Gz3IAK5Njt+diW2K
HtFRtoBx6JfAki0fbkqu5nO3p+6MQpjEJLUCXQqEojlwhV1qkDNoEHnU1KTfQt3s
tFVWvQObvzQFwS+b8RNkf1u6qNNTsnfH02zF68lklpp6vCSVyn3OYaK7QRNKUtTb
BBYoyJysEi8SqG54shVLgu752tpr3ewluSwdkqg1VvQq5vYDIgWK7Fwov1Yr6SvC
VzWGZeJkLOSw8i4zqpdOnAETuAa3kADiKXI7+/6PQpJdQ9X1lfOSxVq0LQsE/FM0
7cjjbH9uXDUibrpZ+m89tcXEgof5tH5rKo0p7Rr14gdSk1H0U+UfTktzxAZMv0dA
NF7qaxi7uskFzhRbi/PSLLtlztU9syuSF7ozvS/AsvS5CP1aSVaPZ3Gk4r6abepG
0+6sRbylC7r+3mlN+NNOdrlcU5p6/zMJ9U8k+MDDHR7DAho+NMA/5QgVTwAfThW1
HWuIreOsvQCCGoih8/ZOSjWDRfqd6iAhBBbZArFCryIgACwWEgyKQdqsLm1SbuuJ
N3f1O2qy/bIywT50R5SC12i/oWoxGni0KPDpGEupLIxhG5ak50ikokIwHCMxr6pj
7Ke7GUWlmMBhG1SlC1avRPFAJXW18PSiC7/Y++3duCsdb1ExP5J8rmp5tmsfZghx
wxikhGhQBHVTZZ84+lJ2w4nyEtMEWsud6zzJ8NoS3cyjR/S1I4QH8lWxTWrcfrGP
Oj49GcMdnjYciHIPyltdBB7XWySg8Ry+VU+cZaY8MiAfLCrQG9Y4mpMW1K7qkSuw
az6oJie7rprYUQMlEUlHt+XgkwAUsTCUhTxgVlSUxnpx8ga44fxfiwzlrw2WE9Aw
ZsnzPoHHWreLDUqOVQBhqV3dr4yexdO9kJh0BhFmbZR2FZOc7xCGbE8E38tDnRAG
63kOe2Tzfg4J4ReHpQEdJ849ZlAfQDybi4NcNH94nPdaxzaQaxObi4RQGD3ROjpL
j2g3r8wzeXwZYao/BvYvLqQo87Z+IHXMuoqw6ZIULz9rTQhKqPJaXqDoTavUjeSg
ZKqVjcFvqKVjNJ/rQzQYCDDCjWbWUM6asB78ghczdLo9sN0Cuyep6SW3MMfjryQI
5B6fUJsSSnd3uWL4J7my60AUdwu22QOdqEZhlo3TnLPbnr0MCeOg+YSzBXLSQkCQ
uUhalItaUqC/GvDKphbqEGGvRGcraSwikBr/2f1kvJ7biPVTPuJCYdgg+7/OMB0I
wMk9YASCMtcfOD3vNWR2qGti9viUmnQR/4Gu8luqPZHs766nFlNpXtcHSKOrnQRN
u66f4CDbvrLeqyM5RrK6MorWjrHUaNjS3E2zgXiQZFNEHikZUgLhbJUXPscf0t3T
yJrzjQW/CsU6wDBlDmARFr9KU5DrSwucIiRWHjvnOho6AUtXohEMPN3P3xc9L+x9
knNZt6PxzZjF8PAzwqd5sKv341d46JonSJObQFlJ10SdeUqQvDpVcury/O092kaN
aWfaeQfnPzwXaoiTp7z1UbYLc2Jy7sKgcbV0H874pCPUR4RlY62w9tk+6bcezNGM
aFn0QHceH+f9ZpZxHRpF3UPbwxNtaHzRuWf2VjljnFLB2SUkeNF9NQmiSChRxG5D
RS4pTFFftEFZYeXxpOONvQwzOvGqDGDB/mIr0EgetJ3bN9vupFXGGRmgHYkiS6rm
m6U5vjdY5pmLHM+GvA1zCZt+xMyMz4WMxnZd75huJnozwkhdK68q/y3MCOe0YahR
mP6SW6uc54n6+zlB86bvKdr9J1XFPPJz5uiNKodq2ahQyz9jhPqVWV0DQUgCvbTR
ngTRuQBO0AiHGq7rTbR4xgMLnQZb9tEiojoRZR/MzoYx0I+cYKewxpld9j8d1vgy
y4iPq5P5Zy4YJ9ICGh5bTqXEwRzCr1k3gQIg3637QsQ71z5pOzeSFBqyIdATteyD
EwTHFYSWu3V7nBg3M/oDMOWJUS7KkMJVMvvbMGzCOjOFG+3HCZ3/dH+Nhj2LKMS3
DVVuZwVBeLBFm3ieLM+TQnrDeUhKM83kUEDd5chPncUTRZ5xRjHBWB0RVw5VoBT4
M2XEEVvLGutBv7vVhkX0azHcDwEczx9uRCJ9LVcFGiDFfmR0SmuBstbHQJAzRaz3
AoIVKHYX9LZEcdrb0uh8RjaUMBPCDfJU3QPXrqc+NucHERMdAmibzPu8Cx4vFWSe
3riuw3jd+vyHOtEjIoSi1m0Z0i5R1Nw5KuMXrJ2HlaisPXjY9KohAUgqXCxz4hlz
GmOA9k5EuVaHe7XV53+Dg82bvfQS7KZcGxeOVB4VtjhQTevOiDwO9cPmnEu1QeUi
IRSk4vW8xoJrEKis0tqo1PKrdiZhAWzBjTQ2fa/2IBPW237uzzBuyN4DFRMoY5Vs
NSwPFrmzURherGfV5u9oQXSl6mzk4nM1uVdWKvLtHnO7WCnIrz+526C/WrQHY5AW
mT47qmvK2yostwe0tc89+gIUWH9Id5PO7lHAZ7awIoiATUpCa7vAaGduq3rDFVfb
kmSMcJFgzdr5eDytDhI5qLKOB3jCMYrwwTaagLF5RXe6ZMjmZx4lxEhsJq09+6b7
u4qpQ1ZaEJNchGUt1iA8R/ciqooH26/z0xwj0vSpvrY2v+CAx6VZkgprpPKJ0JnC
cw9zuvn5hXWUJvjRWYHAAd0uopsylqUcWaInczRdhqAAVCKGI8pJMH3pjmfIvZVV
jM6bPe1+68N0zsgIYelyJNm+iZp1OsQ3os0fw2ZMycY1n20bNpHGL7aBjviWOJTu
5y/5iIy9nrnZWSsPvSA88y/HouOx5jWDtnpPfl2BqTrB/JcqddWLVvH9WFi7bNHg
nxWRAjUbHYB/P/T42a/coVe4cMdr5ShEbeY6Dp4qOVGk6R5biZbq6MrW624lsm5X
1FuPHh9CLyWzZDKoMWTAHv3UwDfLjKJsuiELYtT1l40q0CXUNHnUpYv2dLOjdptg
eB9F8B9cuqayH4c5c5BGU2dWJzH8Qh3jqvlEqEeBoFTXAMliaS+VeEiyA9it1yXB
RXHtynOKJlyTwXmRwpL1hgS7XTBgG+RVb0YYUP9K+95W9GpvWk9ADFsNkEYKetbV
bZmfzjhI0wHEeJLoNbo6/7kTqy3T0SGpEgg3xgtQLlgoSPGMtPPCdm6Trp9MQbUx
PaHr0xCqlCeZW5FXfJdu2bskTX720q0+Ac5k3J15IVEcOsmFyUhq/XJM/ndqoLb1
Txe70AnG65hLrN1qqJQj41PP/tSO6ffayL4cLq/unJ/b1viX6aCv7Bnt90tHDcCj
SfpsfdmseivOE2rOKO/j87/tzdI4YI65agYr9gv+Oi/re9Ts7Pp/AyJ+EF8Mfehr
PcCBEXkuELAMdNuiQarGyWphkI03+v0CI2BJSH2g0sOJeRPO/7uXy656yH8cZiYA
qWYFeq3wjt5iZUUy3i2Tsi0V9iLCBYf6sFz5fhndNL3FkYKG3yVR9xTiahz3Xtk2
1r7PjNLZxHItq/Bp3odn2toJDK2RllOvZhBp/gQosQk6ZTmPjtgW6+pRyI49AclN
vRndZHWkD6+VKKMSudAGzV5FhFAZokuGRhaQi/hhp2Hrtm9WdexYzJzdDUVwLthS
TpF/IoIIBiZ7mIIiUAhKJOVUNlWWP90el6tsmSS8XRznHecyOJoSzIRycW3+D0ur
L5BntwIMQ8G3TEkFuxrL2DjOr2SvojyKrhyHil+VzUwzE/jr+gFznO4AiuG2tbZ8
Kynzj3KrVKeWP4yMzoDrjk0Bb1DjGz13/qLVLBjjOKEZ0NYheG2XBrsl0p7Y4GyS
+PH6XVFA/6XxAiflGi5JBDBTN2uGlj0yKdZZbOjZOq/kGjmBrmVyfHub3r57LSgj
/9dryPAq/pl5LyM8Moor0tyVcChEXxON+WJ3+pLeAYB4hAQ+0LYKgva3NDc1Beoi
Rzp+VZdsY466ZN5gl98x/Cb+u0Y1+OjZmNCSFu4Aq/Op5JtrWCUXIk596xn49NMC
6tOLCHMHfDrGhFdr5AIrzJmt8eYu0zTjaLS/hJEN/wsxdAkNeA67XCBeYhuAHO6z
C1gnLOMGBNlh/WG17LPBG4y+NG2kO+w+8siU+kT9N+L6voA1fhQ3bQ1kI7Yojqaa
INU+qBjqXCnRyaBn1MibK+TL1ARub1NUKAmXLx/tl/ZXw0tVzInK4fOhv66JKfM5
u6ONdSuA4xp19hO8/DlR+KKYes4iQFx12UeMOiBkivJcVX2owBIeaIBTjFvdaHxC
DvV25KLkl0X/obPKlAdOsDZQBYZpTc8t1Y8evLdlxp85xmBTh90rOFJpiSdoQiSx
1ZbQRF2tbfjAkyLyJIHoWksO/D+b4Til09bOTkETEDZg/KHE7UlfI3ZNHSru55Rg
myPxDZN3Q7Gb6mRmvABxbeuvIAwNxlnXGQTJXzLDvFpo2xblpmuXMvZnrKAcFyMF
Tf8swx7QpZuj+llojgYyn2MFvOBlwvpzDM9cv0AYV4xtw70tPp/IMHdWKNJM6PEB
o6Yiypv+deaZ6jcuNQgDJA2bNTsqYz24gOjPKL2439Wrqykqe3THkWUCZk5QMtBN
78FC1K/jvY1ZRcrjNQqmvZGOSab/rU/oqhOa9/W9jj5Q1zAWrgNsWmwlWlu50N10
hsvPUlDziTzraqRQyqI+iTif9ThThfNEI3lfccNYa5mYmNLL2fvcgoCRY8HbGuU2
UP3cSOHZSfmSMCw3lUIyDE/xOd8aZHdcBewpIL9Ukq6Ac4tj24m2KPwJMXnu8IxH
xyqv7v5R7UZwxzlQ+DuJJPJtyWkUuZCUgpnxJ+n2XYp8Ik0LuWEpR2/YmDPQOY3V
G+duxgDugmhFjyb//F/rRlvdcJ1zMWHpRKdq3Lz7bwZDneaFqDZld+E7DHYsNwB9
s8hQZGtlE3Hskl62HobdsQr8X2qcrNMure7soH/gvdjiqgWR/9ql2gZsLr/cXbj7
Z7P5FAxC/ZS++/WzYQKf/VgTznwuIosgjo5XNhkK3Qsybte3l5oKGHTthP4uQwog
c/SJsGlQozQ7ivDIs+qKuyQbYhw+Zu/RKNihX6n7C0iE8Bc1WXAtRqV0HimAuJt2
a8mhbZ5XJ0cp3uFz4BgBEPRUKBi+JrkY2vhta4SBRQFgNG98ygk27AAq/Lbu5NQM
++pCamZwVbXQ6vDLsFE7bAgLRQdpZPrY9xGPKqdJifpA7G5SvpaCy7Q9b0bOyuWa
18FUGVY+OO0Ie8HERvYOEYsVbex1G/min/DYgKyXRvMshP3Bitb2qS/ugI8q0erR
pdGu/UQ/5tA1W95jarA/1YGYUG4cKPxjksh95xcbHBqZuW3BndX2O5hSO2ska6NG
VHPJSHbaTMnIhV/TDlLpLa31l+EPy3xMWxxZ/kuv55GGoYmxP+twftqExrb4yWvN
kW16WhFjCr6uYW1XbFqKbbmOs6ybhYiRf6vjecNzu9LOHnIH5G6YTpl3K6VPGVJO
UExIkN32HDS3PgduvaVywmlVcvpaL+2hShr+kLaWgDI2eQ7RvNnqyIjWaYftwMGm
2SQ/b7NqgXDa7gezFYvGFLy1tRjqK8BD9XBxu6X686nE4q1P8RDyQ6vOsQ8f8Emf
hktTFpHbHF9zoaTrujAGVTngorIAtr7l0GB1X01w4JsXQYrdDyOWpcxs/DDo27K0
RMWQWZCYdLoTFP82B0kWbWnKkSdFPxK/v/dl2N6yMMYmkqHxRqDuBO9SZ+hU6T0Z
TVLl3dFXpnhFKT8C51OFGNSJjfngPRflerJnPwEsB0nyEZAzh0+wedN9jGtoI6Ez
g55NNucU5nUf5EMCYeYTkAU4oMVPQ2anRGyHInHCEB9A12K1WR5AyXrclAA1U498
o9oodra0HUlzlCoRnSGFHL1FJ7sC8UqwBg3wFvdXwkYXwCir9jR887rCEFcwGoBV
iPy8+/CRW21w1FL1domDVjBuhzHHljIDPYRkp+rTBuFvWSj3b2iVwIrqX6ZfWVDd
0m2KFtiEfhdwt9th0uGJ5KhJFjRLzf2027sJOTyXKNyjZuXwxi+4V5YOp//Cme+p
41QyeGwLitOgu2hen+Rkg5B4kFRHjngZX296bVzvoHHiWGPxiv9MdkrltAPHapVG
DkMOIG9gR23V0p/6bkQUnJBQk8eYuZtxXg4yppBU3lQsK/O3/6jQNUDTcqdwQFvM
8B/B/qbUoyYWFA6wB3yTmYycB/xbmRqlrPh69z1r3d7npoPHkXRJ3Khw3ox64Gza
F4foC2mUNXLrnMr/AqnmZG27ctdbOk2kadunhISO1HrHHJ+zOFHZxaF5pnbgHAeV
V7ek/SkeN8FfjZuY9UY/4FMn4eO2Hxv591jPUZhhO7ZveGpfuLSwJ/XEF360f1tZ
QHsCBaHtfN5P0+O9j7d12IExASQBKLchgGNsBVznD7f6AdPk5KZAg8bSpAVT7K5l
3GBqH6lnpaePW6F7+prdaLSHd+1XQkim57w68MLzHas2mCmRddtU5pofwttptgcJ
OZ0vZDLXqwpFBtzVD49tMFSyCYVEJib50tqzSpgbXHIFeO2UGb6nZveoxQVYYzNf
03ZqFc4B2F0ZRrg6szz4CWESTeAjW7MK9ntB7Qh+iCrUY3F3TX8TplvHk3OHv5dW
/QZixWlaDSaSMldyZ7+YLLWyNpe2evLk2oc8qAsAAMR9zhSJhJ8ifieEU5o28M2V
fBAnqdKB4gJygIHWHteGTxKlgw/yf2flYLT4//vmR3KYM7f/41jDLrorKGgK67oE
CH19jyjBrzWFaovasJYlRdJlfwaK4JRfKphFx3niYl04mocOfFoUI3grZgo29QV4
fbCcQ99fbfL7SG5MN5Zu6oD2rMgwOzolJxkUTc4V24QKEqOyL3s9iC5iGKto/Kta
5jyTeYBFN+qidpKqfiNGDWzjO/z5Kg3879Bw9tjnUPErD/Dlb3ksNATb+6TdzquT
I6DlHAdrNs9rGkk7tZv5hUsVM3MSghnmp209rWgY/nfgCzzmYhH0sSPfdiVF/cv6
2tpww3eK0oMLocr++43lW+K796Aa1arYuyixfGGz61Q96ZvFtj1VyuGnLPBcirYY
JxwLFf9yBugRIncbtA1cMInfKxdDgYPCUO5aYdWTUCANIOBlZAcVk7/Wdxc14D4n
Xnrq9tZpqBpNKlGS7fWo1lsZY8AEKVJPi95uDQL9Mr4DNSw0IcP5w5ZdAhvrBcO9
6d5KhgUSqU49WHsjf8adLl3j4KvXRnUm+DcFZbZAUZQ6JAM0VtDlvvdj4tRNUWmq
aRaPsaOvZPkCH3zFUDxGOzpqowbUI/YfiEL3ZjdeptBYVwfp5+nXFVmQBjQKB6Wc
H6Rcs9EHioJWFvUNYfumTG9yukhD0pMlSgMYAlyPHJwGaYefidfYzeQ+4+lr/WzB
ZtDm9OHcOrfgO5+y2coByTcsHcI2yBV0PK8PDwoPqnhkXI9X7WebI5INsMOzPfn8
G2Rwid+goVY4YID0Pw5zDgbgZkTsUqds7NahFEq0sfdzjDC/dT2T0uKvheSk48bD
YVXhQGB3F5+A9peI+dILnUoDT/3PO5VgutQJzBF1jXBgTDaphqhZ4R1uOS4htom2
nrQFtkkLM9MOLv8MzbYpNOwJCCYF2kbRSYLQsNwv9N6yTKBLzcUErLmcWi6m3E4i
9lYEuaZx+MMjXlNVF/LQJIkEA7er0oZPPqKi2OXx6Ph786QBuk81vLD6uCZUcfHX
en+qBldsKkx/pKAXpbEWqOi0PB506d5Ra5yY+urBqLtuef8xHPQUrRh0uj5s8Y4K
+QaWK8MuDCySFxdoj7RNSHg4uKGUT+QIEyfE3Kqm55tRWqTOMQVPsKf3Am/KwAJP
OjLOWTQs78JoIbcBSeZcvB93jIhtooxoiRAdj1gYw33WjdqZljqgIEF1/C2jCh+w
/AH9uY9vs1VxwiB+HLL/o5gphbVJ9kb5gA3vvRPCbzY2avOKP4mLHnImtIhQ0hLE
qCdDMEtLllvqsfeiSgCydT0qcXAPS+5IrWlIyXSP8mPQu39vdK8cYB/Gt+swJjer
dNkGwYEDRG9NoQGhufDuOiMa62we0nhZoqveWepJdr4y+HS0LP36t186rW7i95bm
iQSE4zBGqvQXS/vGY99cO/+n8uVcJFXfHgFYyBHZWVTl2ecZ/ri2WWfCqemKSGTD
lHN3YWL6BD/y+mFqrtUvex6iqIHHGqNVvx9oYQmsYiuO9n5L2VNDZMOzT022p4oU
i81pc2RiGGOWolIFIrftNi2GkCRw3b9897e6DcuLZ9XgcROBbtTSVLKG9VupUvZf
Q+q+J5AzKQO1vATWRwPA9NfV8EqDY20iPP8drxq0EaOdxMyviFi/V8T6c++EWq1l
/BFKM9oj0ndssxGw0qDTy9wKzlZl1BkSX+aM69aTQuPAl75It35Ay4cBnrDQKHqr
9Tu3pSNB0uPc74ioM8aTiCBw5cFukZB1jDwoAduU23dDY49co+uMB6SMiQkDpEpn
opvQQVtXWC22YOa3WHsHFiy+tOTUyDBjIO1AktGEiIURSjadH8O6dEbknPlShM7A
tm8vWJ9M9nzE99y/2ATC/TUlZBJmNhziSK/tvDlxEOOB1BCVvC0lZS8oUSPE9QPH
RQ1NjGVCX39D1S7krfGHsrhDXhnf38kUOvZZwJUu8GhGsKSSNIKU6ewhxUN83mPp
Wwzd4+8goowIXMaXVQLypsPGDTfdfwefxoCWYoI6+Ud8dNliP53efanNy8gvGFZa
fW7Vnr4XoAmT8prZEvM3XwDJB1Xa2hjofcuSQTjZ99KcxhN8VJXD3kNg3TUlwUP2
uUatu5R/oHckG7BwK4zBVe8UpKe3Gm+GxEzbn8ooqw9+AaY8HVAjnJ23xOMNOofp
bFZkmamUp6NxD3c5hUksKkzzSl79WeIiJr1dqoU4iL7JWH1DYvhkq9q0cesU43Ge
iwyO5oE5alNr0yH7qJBgfgFgbbNqs0oaHJJMESyrZQPfLNyFuPzuYJnGY6mosYrp
MNc1VecQaRG3AXVaclixpEF2NmrSeRH/vH5LufLyJ+emEpr0J5EA8NP/5MX6zUxt
bI1eWZzcPeXNGQkEK0s/GDD85viz1VMTSgBazqwsj/jfPf1oyd4sltV6bVHWx2OV
sdlMlnb/T8/VHADa6BLudn3sxKWmIBFBnZ1lrk56lA//9WcME7WUCsOhgZJV3xJ/
0BKZlz0/q6iwqsgq6/VlBJK8wiq7Iz4xtzsy59AIwZWHYkSV9iIKNZWXYCWEnJHo
FNhAwCV5L50pIaoAeWcRync9nw4/05pN5bgXsOY9aBVPyiBrIeT57E8SEHbW+g+N
KbqLSpyZ7rZGGD5zAtYStrvcNx90pxO7YmefdaBItBEx8IP1GLsTRGMEASCY1EjQ
7hHpHbukafaDBEmf31lsnaMQoW9NTbBww4kBCYUZdoiBdcnhlx7pwFa13mvTpi35
sh6u4VX83mCrHyjE/CwzAGUXSEHtfZxJ/ZTvqZbYiZY6150ze9OLnOMO2U6+jSKc
a/UttnElJglu/sl3QOA7xP5UuyB+me2Q/VptsDnn/QZ6R+irJKtdJ/lBdrqqiHmu
nQL704hgGDmjaF+X0VleqJlAw2uCZDA8gPa4Nv7mP2YB/9P3myDlOGyi/ieih/RA
fWv4uhzcQQ5fH7+DKbWHF+rMe+I2yEt60CD0iunQpS9HaWY2YsXMTlN9J64WzXv7
trMBbLoq1+Atj688CTqviJHGTq3Mw5XlPI4ZRKtFCNTHyxD7fnMsJTQrRuX1yDj/
4VbCaqcuP+itliV0GG7j+mBF9x4HygT/3FdaMBfXZJpE6F5tuEdDREC4y24DEXO4
SPM+x22q8YxpMZsvtvO+OSilVtFQ671QbmXNfq+3aoquOnnQ1fyhwAMXnscxMW5w
IcUkE5mBxqFglwCViHtsnGfrBevp1aHt+UF4Q90OC0K+aoasXjT40xVpagM4IU+F
GDI5yGJYXD34mrOZGF9h8+25DlD/17U6X+m88Hxu4yfui+vTE2/fHkXor2kHMIM1
6UcR4dd8y1AWkDdX+qJwlQL7m5wAnpTpGVbEiuKlHdnAsdnzXq+/gbOsy6Pp6Sib
yTeILLT4DOm65qZ4IDx5q7D2BLRMxcDcahaXXZ8pKa3anNnCfoOF5IDk7DxBIVbc
L/JeKo+nUB4FoXk+Cgt5G50rpoSCdovqOLpJfQZF0s1XbRr0J1YyZiCaNdGQ8Dyb
n4S8Zg/r18JjhPH+mhXcpW41p8nEM6LObOij/42NwQe718E/XwGnD8duSfhFi/G3
HhuNJKlF0UnfkrmEQfH7biyYqO+aNVlraVllkmOE4NcYvkNNNvdSMeHuZpMNl6JW
kTWq4OfZDZow+gbKdXful5DvHwt03j6dZmB42FSGqJcsc9gwRsCVBq8/DRzUX+5D
cCEkJbuc8cX/Owx0lwEvP70qwQfl3iTPJqHBxRji/pOqCKt3mGCYDWIHsT2d1CLE
z0S7wJ/964oSesZfnaq9H1w82pKNJvCp5M4zJf5ZP2ygdOzelWITTBtDgw0+NrxJ
hm/pw6aCZx647AwPGagYmwgkc+sDkRTgQt6VSoO86b24jmNBuR2eFnX0ccVONelf
vBKDNTmFC0+ed9VlHorDY+NVaxlcGYsu70MqA/WBL7OI4+nj/BuejbJBBQSU6gcA
l21peZ1rOhZb5BWWrtO5VodWrbWjYR49E3jv+jQ0nPR9TVBMs3XakIn+J1Hn5Z27
Ebyhn7UI2FcKd+E8fh8NedTThdSogrbyJK534+4Q+SekukMFHcBUT7fpFr3eWXlH
1d9Pdc/X6JJO7OPLJwNMDlentLByDfKlsgWt+6ODcLkrtogphJmt4gGwbiTPR5yS
iBJikWVQZHKCPDcuwOzqgNBtUrbQ+1rAj/7ATiUOVcAW5mhd5pnJdmPofa8pF+JY
o5gyK3mvlWPYCh/H8x5v0NIclpTJ0HKZ3Q/RzBhJNET9SlSVhlphYiipbFSvruhq
0fP4yjQ5qhTlnd6XYQFdAY7ZLzqUZsv/J7f19Wd5Fd4DPkF/84uDNAfFQZo8oH4V
HJO/59I6j1R3HdxQ2RUYY0yVDUOc2uCuC0NJc8RqCkw9BoXwLKq8qlS4lgvLm9aO
Pcw+Kpd51ZdjeKjVc/ZyZHDZGqIDni1bSrIjpb4QYMMClaN1PcICjskTtktTQcoc
iiVnNS1bdzQ/vlKPSRe/85SazbRCW2IqnxB154/LAa/wWVUkhJLRwsi2jbiZRJ3Q
AiQShnfHTV4rrSktzDDCyp3Z9930BCkMbEMihBjbpjA=
`protect end_protected