`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
ddtXksX2+yylW5zu6QL2Lhnb2d1sD00763mmSITNX595NcHTEkwn0zB1Dry37fOW
FufOhVzEJp80NC5qZ/+F0Vk7Ik02dIR0elf3clrjeJRK85K4e3Hoo4xn7YbFUIms
l/8VZSb14+JVGURjfswrIyCUotIzlzVYZ6gzoZwDXIi5gQIBf/gI+KxNXPaKV+PQ
Ufys/12rjO6aI/pPlqSm0hCvftmBcnezN2hk1UeXgOIuKZnogjOsf0iJVX2aOOWE
6pD/psybjbnsNB6kH5uFTA5frkzIzkzl5d9+YDm9OyC+k84E83I/7/j+rk4L2dah
QJOvksSIzN867/4Qt8qYTQ==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="MvBXkzurAa5VTw+1JJ70nePUfoQXBvZOku/SMmg4TwQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
oRtzZL4VJ4iwysPsC8SXYCzXS8Fw2gtZTOskLcDV+1B9Nzn1zTyNtlo6lNICRmmK
ZRVu2BmCc2G+fmzynYlNTnSa7C0Cuel6FYpxCBlOuk3OF2tzAmLAuDyOH3Z1Yjzk
a0aHuoCdIRKv7BrZCdALt03JeUmXKPdOmIlkVGFl8yw=
`protect rights_digest_method = "sha256"
`protect end_toolblock="Jn9CQpRhJt4rnzZPRk+dOpzAubz7omckX1MrFd4p81o="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 4624 )
`protect data_block
gD6l00tciPUa6pDNTk/+t0OO0nC/UTtBwLB41d4inuAUA3i/ALrNyoJVcBnAmEQW
ptbcNp5fxEUJjnOxnedyZEuEBxWRieZFQnkRdF269oMhrZIUk16/Jjx5z37SpgvV
9Zyz9K7qeyLqpbtVHBiXFwVaDMdDfLDPL445+qWbVBujraYE2DwJ/L37TlMiXxYo
GOKj1WUkUesTq1lZSChN5U6LYYAjc/wHWrr4C9z9UjrZLMKmHcMXEDvsxdFd273C
wxyDMtboG0OjQ10sjesnQm+/fnRiHaghs0PNiAux/fV2/hulVm2XML5SYkHo51Ky
zy4I6WK+pA1ywQV1gfhuRmJFSJXDf+xA0eom2kAUvmWV3RF3K/T5FfqkT9DUyRrG
cr1dNahDvqGF8qdwFG/Yhucv0MeOZ84/3wlJVyw5mDL3yZoymGK8g4++RhT1jJJR
RCYCYJ+tkCb+CKLZOMd03gJreFi7u9GyqbBjmBruVb2K2uyLdCsrDApThNjoFmks
dSzJJm0m1OjxLvv6htRNrk29Ub4YMYdAnpowqyLnfDeoatzkSdvyDebhBaZDzmOr
aHeVFOO5o+BLyArSruXwP/iiAgs7ixQOc3S0od92HU3kfPe9oTcnbZSVTlevtylD
sTDCxcO9sLzPQuQF6Ntl5DcpYV/cZXuIlwGr/xjqNQcBR4gfmjmLOaX1DHZGWhkV
oboJaYoJV8aw0oqcKZnYtqhpwOPHeIsrdBQeQtvDF/czT/UlKga7LjkZag/TTKq2
OB5seN42Ty9nYr7nYUUeyLuGFKT13aAEtDQgouDlWFWgfknvziSWaNmxBU8XmSUS
+tbGw2PHf4+5HQCUTyZ2XZTyltxESop4wgjCvDHd55fa7lZBulN8llBmz2SI/lCY
Ju/e3bCwYzyZ/QsuE59QhFb3y3qmMNm5tOPjhcJ7aWVsnQHyUuSorHPCaTk4T1P6
PB/tvVrK0cgkqjuGbm88YEzZCSLmCKYtesFE6evielmu2dDX4etIXV7bCIhOMAu8
SJKQJ/tKFmA/Q+XI690KYo1WGTaAan9rN4hmKZrGuzXwpGhzaP/7a/T5xUZR/0mx
lrCuW7uYT6Hu0Rq461g95R6Llv/Kx/GPezwzRHz3ywNTqz9/5PZMw164sBR4Lx95
HHyZKgDp7gJDIIIbIW0HRgOBmPD10jl88krjS24Y3aWf0d2B7br7/RgBFv4rWREI
4UlGkUMGk+7fkKvjVeF0iGZLtt98/PIF/TJqDrYU404hjBq5OvaYXfz+pH10R7fQ
7Xi/xgPRyDT4w2DWWU12nUR3Kng5oiPM7MHpNm4FuGdysrKNiuOe3HcJS4naIYKb
NvhFUhvOQaEjogeT01HwXbHXjOQNggz7n28lOiCWnLe+I8DycEnr9Jkz0AO9leBs
l0adpOqwc6Zf6urmSQke2g2ypj0DAvKykHH6TPtDGHUE7dcgnHXhZx6fUK0i6B5O
UW4584RZ548iT0SVp2Fs2VO3TxEfZJhXLf/G2F2yQGcFyM71q466ZBRtxOR6Xij7
GF8clket5/gsnFWwgbMG4Y8BMMaTe6Je0H7u4LnXnqCkUHb1N5NDLYtbkqCp4qv2
QrJAYeY0Nd2YGl6WGS9haxs+rCzmu7Olq7rV+lgC6zYjTCS6n783RQlEUWkKq0fb
A0gNVzSbKwYs5n0OiPNrU82Ts4vzxWrUa+jyUjkIDac29YS7Eh0ZfcCFwRgt3h8B
nUoETanda2cf3qIK+iarZ8EXko+NbdZlxpZrYf2metFinT4OkSMn/vVud60+MHDU
CunlJiByYCi9h3dkXGIdAqAaq8fYApunjCCD0UZLokLgn+8OO3Pm4o3KM84tMPKY
fMs2P249+GdPIG+ZLJ3KU/MMbQEYkBnGcVTGT0+Dt0VDwZxLepsZhS1BbKprx45I
h/lGVLI2OrjDdzye2voja705LEE+nvW1Dvs4SNuQkND3ItOZl6iuRKq75AqqAshC
nAD8WiWtfwbpvyn65a+B3Pa0XgHgZ9qHmcYitYFFBXvfGBcpETLy2MibBeM92Mar
ORKDOYclbWbZ6cyGF0olEpLmapQC+hRrqNilE1cxlGlEnU6lmoIJwqyZH9KUkNrB
zFkQlaGuqCIOx9sVlclnJfLu1CrACpNcpTKUCVWL71ipjhZaoORnSkj7lPbfexT8
4TdwkggoyIYWWHJqxaypIy5jC2I1wjy5rvoYWJkrDzg7d9FxZyxseHuDNcORCjUN
9ltbICbFJ5BIoDxK8cnrGXQ7+zO/PjEfE6pFyV8wkdjZ1CStMCReX40l/WnEBqTe
rgDaTGIdKjdkIRsjoc+Uy1yaEW+GAmmA9w7FcqvFKP39dgoaSEtKT90B8jW9gvgL
0vHH+knp6hA73OlCF5UC2Dz+rwFJzaBAPMdogZQrzwS6YzYHdAxTRU3IFUNjk03q
Xmru79+ZOHZnhL6Wj8WCMnln1w8ivIRrm5qPGTi+rwSZ4VxqmpMg7x6hKhNgbE0p
0rS79SUgcEq8YgnnuP0PdZl6I3vGnGuH+jzPAQU+9ZzsST8k7nddyMzr9ZpSqlXa
S3xwiT1TyIKBmzQ/2IBY/hT1iNjijLMFtrTGhye0qvwnC4YU/R1fcmahNHKv9ro5
uwoySPHTDP9kXIl+mu32hsm54Nb/lUuHHHrt2BDjLZwYExfpZyq+yNR2PcBiCNVi
mX7kaQxCMX9fW3M6Ceap1sCa2/stz2QEhF19D+pUWt2DrRTzPAH6lkh/wilNXPqZ
tR95DrgalVIUUhOf2auNug9c0LkpefjQMoez+dErBIUVeR/RZJBz5MZ6neSHpqAf
WSbs8Xy+JwdRY7AgGxXF+Fn8cPzImOwm0B9FXHkSucotSgO8w2CVhbGxVWQiUcaN
qpoSvZaz5bqkr+2DohhbrVRwTYBdc28eC4UKA4iId1IsObSyvkl/gd1zWA8co/hm
x+oPuzrrlbpd3Ex4qxm5eyuB8JcnuhAo2ZqgHzpTDVb2Nrs+dO25r1sDrqOjCPCT
aojLW6/+2rhJcvENtMc6ApcrLgqA30z22O40nGXgzHeBl43oNIGD/+R4ihmbyBD4
S2VWTfD4Z6PhjEIMNnH4R94W4MPc+oMmgvKeh4P776AEhd3krZKiqSNGWY04WBDk
riFOHwChpX8/qGeSdABR8PgmCT3kiZpD94fOtj/KXlPx7JuDKBe72QtLVhEOYA6Y
hx+weFM+F0Naldq+OC8uZ5LI1+cSKfuwYPjZyPkeMpuJFYGuC7Q/yOFDgt/xI5vu
/ySP//Z7wqGUJdHuY7D1/y09+74qLmB6S2DNQGb3FFKp71ApIwffuvoy5IlJQQKN
eXP3vRrzufQ/T371f6tGQqgcVZ67Xk3DmDee7DhuZuiCtnjrvM/mAKLJKzlJmS0n
asaVft/IWK/xVcMwju9hWVkOARv73fu88gkWTHjZzqKsen0L89Kr1kipvolVyVcw
kU3DLVtswABbOTpT0gQdlS2jKTmqq37yLw779U7d2rpNoePP+SzUN1objVuAHvmJ
8ec860wOIeqvGUtoZTFRjtZbwSqXG8gFZGhK9flTzoEx4iOXBSwhHYHJG6py0ovo
NTLwQgn2cS0LwsKDCCdsT6P8720aVtaXZbCgipZ4g51dcVN/6vZWp+3q3rqY1R6M
vxt+wH00iQCQYqfSsHajOHQpfkZTfPeCOQFGO5TAZ2CABKQnll7LaG5uohiJDx5P
oZXjhrTxXJdbMGz841yy0bZdT2TATUS0DcAzLW94m0gricZJSqZmqLXvAU3RGoHQ
6f/DSCzd3UmoyEasJcHQqGLP9yn38Ycmp4sNrMurgFowAO5MkCetsRWIvJjyWDDZ
EsRILkkQeVDSxFylJisUcKVGlXm761gBQHcX1OtbzoWIp5SD7j0lFaftrRi1WwMb
qpO340f1U9jh8uI3rpslGX1fXJa3WIX8SzUxxNy2Imq9eFTEC2kzeCcei6CfDCef
3OKrzQkFtMerC8tIXTmau6Gk3c0Too4/nLJaqIfdWFs5Eb1eIfllKDFkY/L/jAaN
NxbhQVWOoNnUyrSUWKKwDB5xKpNYUaggm1O6luKgFPU5FgFQw7sJisQZI4AJfky7
Lr3Y4XMggLTQyp1pGdSslbBm4rA9L9UAvJuMW9WuxJjrLa7T2Mji9DlsmMNUOWOO
tLeam/Jq/WwpHgJdcHe87GBpZ3NVJ2HakqLIRyAnac0/7GNjRmMtl/jnoM2foD2I
h4r7iz9YyvDrIzKOdrqb+A09HBjLiXgHnIxN7QboQCJ7I1OBPo1/41yxj2UFbY6U
KfMuHuofCNz4ktv2AlIsFo3uK+kpKrpn1QCGw810+hfPNxd9td8ddl6+FEt2M/uv
FzO+/CX+rkM2G5d79+QxMTeETdTWrUyrERjuqeG8PFYkwleWcFC7b4Tjdlnt5v8X
Jgmml/Rk7AfIyTQ9iWilXkvB3iQwgpkQIokejocNhfXtJUWU5BLClkTmSi07mH/0
nTNIij33hQZQa9sM9lvylcQgqe8W4ijKwn5m3U/9AcaAXngzXjMT4dofeZ5bs6PZ
ad9Dx54twC0Zj6zyWjtPqVrtcvquybw2BsyVSa8bhPQUSmnwCH5TOCVrwn563PJw
d+fG4P5Cb5pSssag88r/LmQrSj++toTRofsDjM8ad89HTJqQPo+ZZG+ogRL+uBoy
dYKtqY9C8k51tuSWFyf6oIS2J++zm0dF/szJnGSDih+ilvg9N98vbMKfg+laR2qh
aKiL2HfoRlQizONR4+h/qFUr8WkEv6XVtsemZA/wKBIf1IpgPCT2/3vxED7fQA6D
qPcAFgC/LRdl4yGWaOJXJWEFnnESssq3aQ+KG0pE2SYtRM7sHxii2OGGg9NU7MbY
OWAg8sBO89BqudwpN3qsTEMiqE2Q/7znYofDNhJoxYgX1M8/cx/0fteqSdVwDmCF
M6aFocH5uMQS8agXjRfMON8nmoa9np3g71UQBtg6UCCxwlTbKVuYJeJn1zQ7giQf
gcrtUpI6B7UWZrjdcrRcaTRLHVnRfWTRn5Xi+4gbsQ3TbzRs90QbBaTIQOJm0myp
tRUEUzJH/L6wKlhaMKi/lznUjR/N5exF4S588TJE5Ly3VTR+GcqjIkKocK5RrG8n
r9tOYI49EdTTP8QHiYBOYfZ7qo6tXgYR4Ot2XZQelo5AlYjDknGJrOMB4xIdFu4k
2l5H8GN+EmqC5pBEF7ACzz3GMTN5fXdbKWrsxnkrZhujucIYFoiPIDSDDb+y40Ye
STHWUsiZKmoo2ucLA3SkW3LQB8quvXDFNJOO2JwRyDzqlEkMVwIF8ZSPzRu8CIGq
PuqHiCccB2+nhCPng4ek6gV5OJ73U7PEfIXeDdDXvQE0xm2kAS6fAH4yDc4tGDz4
hgNiwSmBr5GpGrD0rYfv+HKDF3sxJNzbI7HZ8CpIEGESLgq0Tv9sL8YwBkSm6ic4
FtKcL559sMGD2K/leHHqpGn/ZB4d2WkZp2CXUZrH5I46j2L/Y7pNKz3jrsFIlKcy
Q43WUa11lDCp1MtEaVS8lm4Zl8E9vGn5/bhhb+LW+fBc+fvSBBCYzqG544vKzxjK
IEvK749aVwHPY/sbfCDmldJEMJv/TX1Irdbbprz7Toj3QIqr/jiClDccq4U6N92W
DOPQ/mQ7GLR7zIWubQIyjcVjoIg2zWMwtsmMpsZjLu96aY1i233wwVMZQmJFq8Lt
jKSFL9MvyxYsQF2SVfwvVzaZygMEhDBv8Cd8WTrfNOogmJvwpqGSI2sIP/x9Wmsw
aTW1/lR+pnpTCTTr5B7559oLqxKMGta74dxHzLFJO+O1A8bfJkGCOJg/GhWgHFOJ
jeaGkr0xqEo1lpnuRF7ACvBn08kfOy5GHtk9oZ0nTBCyig5LNGxcut+S8hGPfJnt
9fMcgUVaXNIrgS/IDyjW0rlNeiO3ssn79id8DLrzlHsOz0Km9HK7ys21LXGGlU4t
fgk1WY9n597ffMtJxW6h09ENSthGyAOrtNwaFi0FDBYaBRKt8RrzvLLiDTgLEm3o
vlm15LD7nVHTGdhq101OTplrfQ39WgqLXnKiTDVXQW5KjenyyhYlUgeUjwnmfqXI
N3MiU5TB8vXT704buOcOezweV6nU4DM4CmTOXXno+xe2kx2FWE0zwC0rdCKA43Ur
Zm/ZB+uEb2aF9zMKcVKBWQ==
`protect end_protected