`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
ddtXksX2+yylW5zu6QL2Lhnb2d1sD00763mmSITNX595NcHTEkwn0zB1Dry37fOW
FufOhVzEJp80NC5qZ/+F0Vk7Ik02dIR0elf3clrjeJRK85K4e3Hoo4xn7YbFUIms
l/8VZSb14+JVGURjfswrIyCUotIzlzVYZ6gzoZwDXIi5gQIBf/gI+KxNXPaKV+PQ
Ufys/12rjO6aI/pPlqSm0hCvftmBcnezN2hk1UeXgOIuKZnogjOsf0iJVX2aOOWE
6pD/psybjbnsNB6kH5uFTA5frkzIzkzl5d9+YDm9OyC+k84E83I/7/j+rk4L2dah
QJOvksSIzN867/4Qt8qYTQ==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="MvBXkzurAa5VTw+1JJ70nePUfoQXBvZOku/SMmg4TwQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
oRtzZL4VJ4iwysPsC8SXYCzXS8Fw2gtZTOskLcDV+1B9Nzn1zTyNtlo6lNICRmmK
ZRVu2BmCc2G+fmzynYlNTnSa7C0Cuel6FYpxCBlOuk3OF2tzAmLAuDyOH3Z1Yjzk
a0aHuoCdIRKv7BrZCdALt03JeUmXKPdOmIlkVGFl8yw=
`protect rights_digest_method = "sha256"
`protect end_toolblock="Jn9CQpRhJt4rnzZPRk+dOpzAubz7omckX1MrFd4p81o="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 16496 )
`protect data_block
gD6l00tciPUa6pDNTk/+tzLxvdHE2s3DQL3/JqqujQBC/Ei+vcAB8wM3doqg5vTg
mdfn9XB1bLOis2CVSfu295W2DNwHfMSTc/8BhCDRnTlLIX0UCJs9Za0+LoM0rMrV
T7EjVWppbP+Em6PkVKCwlmIQ7JKaifJ+Y+kjw9HCGboYo5074hY+K/CBbfsBQY86
d1Td2lUTd6BUP9MUIjAL6Y/7X6Hy6OF9+gnrrC5Ruage3PJg7BvNjGhyTRwwgyMw
8HM3mQOalT0ZcoT/JjlIb3d0H+JIFfhIKhQOsSX5u2164ggywgaRomhZw1UCcpxo
YSZcsSWvue9q+o9gHYo3t1STZIjeFUXHNRIo8dSFHWPZrbKGkEnPxR7MQvBzXCjv
akmVrGWa3vIIY/MHgJhv8pZjjv7agz8N5g2HZGBoKd0j2rckKbWq8em0kTEmkE7D
iBAvGp51BUMs6JH/VJb++kg6gZsMuj6yEwUm00azgb+sN3GWH6Y44Xbgo0Oou7pm
krJlWxSYqG06J6+8Rz10RQb29/ptgpwZu5fxWT5GMLrihrvH8zWMDBXzOEy8a2g9
/p2wrk7QegtayuHvyq/6TBrMe88jHsw95MWUPklYhI8xliTN/iOghoLMBYeQnNOK
6jYt0J3n/oKKIcLkpTweMXUYrNHVPvD7Hm9QqmEITF5PyW617L2IP41uo2pgL2eW
D2gUsVPjGRx0TSzdZFb6kXGSLgSKv6fR28UOtSDNQx2oEmTASyka+e7SZlBYwhQt
vNTOyD0CfZMxSAXnWCXVY4orRdg2CMXDWONJuWMeK28Q+aA8EgaCOxWDynJurtNt
mBRxrVYHXsgE3B/MrmEsrB8WmUFRFjza1ODQzpD8avP1VE+Nq1J3TAcGu1g+R63E
OB+MaBgDg087D/IJyLNdOeRM2N5fod8WavTXxoyLMkNyky35/VT6EKoPIBnVwEhK
l+zbqpCUZcLA3qRPO69wo2ihhJiINuh0cFBXlPJQZUNdRkm2a+lEjqtgiuhGxukS
/5epeOO0lfUO5ffIsDxVuvEM6UpYWzn+yBtRKTlE4fbT0wQxfT+drXQrxxZ+pfeL
Y67FRW42JV098F/tq/k2rSySUFKRYgXxcAStAwXSxKplAgS0KjXouyZfPOcF67RY
NDNjzQBvd9k21NiX/LfI02wS5d1Tc+OpGo6YBbtZdBu73mxOZwi7ZXXPctQfURI1
97kDKjmQosmE/c+YaAP79vFPeYtfx26H6JMwkTwyHxki3TREvJ2MfpEaYwmxoicU
uy1qDXF+XLWhOveTkk9TGziyUBqP5HE0qhUKBQ3/ZUBG3mneNZ8dIwyZN/Bus0Il
RyQfNPmrFV3jTq4gWBRkelNFLuoy23Ts/ge2jnjpG2VA/QrparbyMYJSejZ5BK0l
zaLZCW46exkZ3ojV/afOKp063NDvpBveQSNOrK/a6FcRKn/pEq5Mi7ZvA5s17lL2
j1tzLqhIv1cTlVP+5I6ar+rj+ve1qiNv+Yfa3GHX0huaK6Eh56GgP9tHQOxShlag
JEBaMBPLqWO6lCmYwJqH3u4KV3Idvpa5ND98ACWe08uRuLGtjozMu0z6zkc3J1ai
huCy7FJHONxDnfc8QHdApxpNu2yrs1HPd+kcAeUkTgBrbRxzxbpqBsbY+8cheEpS
IwaFl0OZgbRJpoJHvMC23Xj5FgGwFJtBtESPrpN6goauVpBP+Z8lK8FQdgHVjtyD
Btay37x4b+k5ABb4l1svolyQFZ74q/aJxlFi1yU+xUKfPIiO2lDif46OT8Ril7A4
kLmkaHRPgj8H5YAHmu0jNadNLvsvcRFL4HKsXdALq/1+3DxIjFMMRrS9/T/1EFXd
cNTAffEYOZVyPTOqgRrVvpUPeGNuorHiBKmz8uzlhmZCi+VUxGceVp2KCXdyiE/O
bg5w10an5F5TK6nCUceogNSDRVyy3WR/eciuDN9ORSsxelqb+jO6jjpjsHHOBN2r
QimZrLot8OTE5zRUZZljJffsxzJ893SBsyAdUIJ8iJOVpR/FAkPsZSvuMna3Weo+
bMmc1pXgbmFoXWpj74D31P6nBQi1FzwxoljXi+5osQJhNn7mFiPQ0u4q6c5wwuYW
4oQhTS5SJ3okoHB2ZA6bQQljbAumGfmcVhZjVDWYoqI35SSGUkXVPwHYHmt/a9bS
LELKuBSAIyJ3YO4oWJF/pFRDTV0HF/+fcUev0v+oH1C0aC2DoOX7/XjecP1Sq66Q
T5dTVUakdYWaQaCfwQpThoVzSz9QuuveCFfjNhEmi8d5HE8yaupas40FXlSxD9PU
aTTb1BYasO9Pxz/QBx1KahUCgtz97qhGVMLDguzvnYJdZ6pH+if/e/H1wMR5cKRr
lteb2D9oxj7w1auuryjZNWOUAIQG1SFg+ha08/jRVqZO2lAevASXNVy5Ckqb6wsD
ftOvlX2JVgIfI8I8KpN/YZLhvoHKvbldqlHV2XRYCbNycJNuqP1WvfTTub0ERQ2z
tONEQcu5cXYGG9OU9vCfwnxzwZVMvNtm4kp8QAs/Q1id0ejNiYKgZ69vpzNetnS6
BPjCulhvUWFQdnRE1mpzHTjlDWwBbEJD8x6Jpl/gu3X7kgHXrEqPtxUaEySTZGTK
K7n8riPljNRqa/KDV+x+QXEk42+qDAClzdzTw7O8EouDMYSDEjoPXTP0mOK1JO0f
eTXwikajIWtqwOUbAc1QUIoYVWJgBMcaM/FukL2Dm/1g+GQchMSuVy7GyuBOPX37
91kjPDUEyyxNRvkU4yOr4yQTzanpjonPIe+Ao17QaCdlVuvQ+/FD1abA+bFvGAqk
rhkPUGX7uwn0qekiKQaeVEpEzvh01JYCo6era6LmjUAogwYaYBDPt6s24uJMNBYV
XfV0l2cSjWxU0zErZcW7ffL7q5SQkGVBnScEg/uaBNOmK22s2BmBysjv/tH6QRII
5ZCQOxEmFKjyGw2q1rUqH3JMLfX+6Uz93kGTBojP6enN0e3ok6rBYL/s75LoazMp
3EkuMEixed0EdVhaovVyPqsD9XqrgrvCFOb/2H+XqFEByBX1zMSQkg10fPQhcFW/
JDuVcjjadRfiXNdIgq89j14jLY29/M+7YiIb9tuaBCWAHVibjN1BZcSWHEnAlJzj
zrGRkvSoGTcb3xFBqzXG7qvzHxpdFNupW3FGfFU/SZWnwTObx3RQfNREHm4hzmYe
gLUuh0MlCJgjNI7gEvU3StglNnYCjtoaBiW/7ntYEI+tfSlBohD5B/RYrAmxvjyq
rUk3D7w1cWGuZYCrCRaDUAL0aUD1zNsPcllyQ8xxb6QsUMWDDt02KLj1JOi6nvwY
F0o/q0jFRkpoWAM/Drnjln+8ygdzwfgwkI+i6A/xEaiNcBXMEqXpzMHTq+X9hKhy
BL6skSXihGdGwh8X+jZJ4UiWVyvSLTNMowqIyV5p4V4/gUEocF/9jGztnKO+yiGb
oL3RuKjRNebVNsCfnQlVvfZQ3SfHpJV9JSycj9g0E+AnAiUxG9tOOjF7q2DV62t9
tanfe5yRmMHT24ApRwuXGvNlDH5N2GLhKx/c11VyVJ9rdUouUfU3Arlp9U9lywIv
PrViRjfbWqDFnrjIdIZdOLIXqDdDWkaqosXGSbGpZSZcH8bzG0rmdA5JXabmF/fM
eWilgH5xAS50V/OJUFSGkz1jeioe5zPTBkB91XHkPWdrqWBiYWeykyhsEG3OYbKo
2nv1G/3RoFvWE/AT71TkJ50ZQN/gb0Vb4u9BxFf8YZVx0jTBAhQJuQRitU56tRBo
9WJ8JT2p5nJPn4f3ryUjIhmE0wOvIuz/nWV1lYLinTiV756QzN8wpTAcDLax10ml
MCmRPYxCv/r4b/gRYrZEwPqB3Ny5WemGR+E0HCNfUivL76jBDMPiWHAzgm0nlNMI
SSEIeL5P0YMA+9YA4u7JQ9LlI2TPalgJO36rCKthPKzBpi06bJt3Marz38BpIukl
F3qxibxA7xnhTJ0HRPj5LigT2fhBIlcUcLBvByzSayosijmug3OPgLn62ksf3MfD
tKCUmHEonF2O51e1ECwfTDhT/9kEAwxGPFCSgG8xL6qjBu9fZXgkr5nfFQkspHRS
/Z3k5A85ZXXwp1wRDpvRIKVbnqLmHKOLEeQyQhbEkroj6F3urIIHJis0qMSshmgE
Ivh0k2LqNA0KHqBG1mLTY7BsBRqmdwY19iYm+L0sNAMHsuOgmcfwAHboR6H519VT
5bUCKHD4SxbrCNwAGxDpY0s5D4UI9qzSj+0tPN2skxqMjPYQuhaRMBKKOW+CH9zR
MizGPtQRs4Wj4lgAayinocGdBTjbzFYQsLMKWvO9BJw10mmZcTiqsMom32TUM1th
echu3bs9C+LSEDMxgxOH7xTZ4oX/ZywcWhXf4YqHfKuFkKVUB0EJR08tfXnuUUsl
In3iE0+2NoJcr3w5FCSGjs3BNb0hOoNZf217E7Q0IRsilIxPmlDUu1N/LlmXtJo4
wKCZLz103xGM7A7RSkD80w8fbVjl97zOej1aObJ8ZYrLTQLNI8GAbGRjB8eyhUyx
RyYhlTeT4/5BfzETWEq6zPKejd9S6lvuIzvJAt14/9MUWK0qBaUPRUQx/h3F9mMj
khEuNqLGLyGGWwN4D2p2Nop0cb5V1NY3CcXCe3rzQElW6UpLn3t17tQs/eifumCX
hYeBU+cEEcGDPNdBdqOXg2rnqE/UV21eElZ1q25BVKXH3PU2Zd/wwWC+TQFIeA2/
Fmp7zJ2HMLh7gxcrKHgI2ZYdEC98noP+6jHjQ3vui20NATdBEO2F6AZ/cS4G0bhJ
S+u+5owTicIW2OETFqROwVsvdr6SS1WOWzuLg7ZEWc4cvnKRKOwNeTT5gZObb89P
AiGa7i61e/IKtGrdnj34miNQLlhOYMumZDqK1okC7DwRikhDg31fgFFEWFjFbiyi
tlkPW5uwbVfAyXimDipjW1i6P5sgbFHC8Iy6TBqYAEPuWnnkBmTXzpzAxx0Ryo/b
1AVAGC6sXyS1ppUl4Uds2rT5QPkMF+ngs90w+8TRsznbJJXDxfdHobGq3i4PXuYO
4Sivn5wP3E7jSXvd1DGqTJS5T9xW372oqC3CGRO4OvbtJcNzrF3BbqCbYpt6xqBf
zrG4J0iCL3hmGmrobC/hKpPBHT1owFGccunUfsVrb+lr91kouV72RE4dMmny5b0t
rloagB686Km4tVWnGGhj/HKRecnG8UYKnjHgQmW5oykrGgCBF1YFd+7rMPHI9HM6
cCpAk6hLXUq2oxcATtKPWsZZjvmTOChEZtbZeIqEKM5Un+CSSc0PZbIOLTIM1KyP
EMucrVz6QPLvS6EazRkrPnJaTqTUovjhdrnIYxpADxLHlcaByvWvtY3AJKOZky7y
UGMRoin71u8ySm6lC2nWpZBrkGOod+FlyJThWdZxLC4WPS7mUsJIDzOUYDhSi0VP
zfDQpE1fiv3YxlZhHp4euMue2l9YyCOT6yXTnsHV4hnmC50htKuFpcFNcLEUf0AF
FLecAK2HBuvaOVKvIvyc8BNT15ATJnNpOJYBGNvWbdHnOfCKTG0lKt2ku/9sLrZZ
JajZ/IoSj3Gwhl8UjqIerVd4t2d2RMY22mbeO9afaTcmqrMMzfFDxUxYIus1hFQ4
2pUGnPSZDnoL8pMHtgvlu/ZL4mcFQAqK98KZh6xiW5sV7euUPa9/SmMy62BTgAeV
uHITuCMypinJJQxBMFQ2yu+HEYbArAKDandvEExXDtcLPtsvAMHON/VJTOm/pStK
BEJ0v5o74gfUnP69ngcz33I6Z5EnjOfw+CFnd4uCbUdGV1OnF7dsr74EMYGHW8Qf
G7rcy2yQ/oztA6YfF470Es+DyxafsSz3E1JzPTp39al0sCShAadfwdQ8vPZ482oZ
6NoBURirTLJbMbO6EFV7PJxSxHubV+SpZpBA80NzjrwZcx/y8m29fcSxXftIZiL7
ON4WBJW75QXn9BuGw006UY3navXmcOHNF4rHNTqUXgxG+LJJdlFfCGq6fJ/vffi3
n46QBTsCdQKowqz/VRWynHLZDPOl9SXPk67fyRJT4sdYBFuD4qR+TL9NN7h0/MvD
qIl+/aIXMmF28yCxmlKwDZfi9MP+iMepUykE2STMsqzTkmK482qeDeqBEVzYHAZG
sb/Tykjg/ouNtjpepr89tThdkl+eIjm4EFkbhrht+VBWGty2lDviAkm5gjiodbH9
EFh6MzI6i7X1mBjDSIKDO85DG4ek4ATG4mJGu3/CChA38PZcE8YGiBLPfBDH0mZU
4ro27i8CsJTRI6uY9otWnY4/XVgUkKGRbzNCleU8EuFtn35lmCmeJQs18wOsWwnM
pQJhXTsCUhZYobi/JDwO8eWoOq+orkE3Qrd6jcCqNQx3AmfaxofxOAS5gtlplSVE
ULYb0UpTs3iZwNJ6gHgTLxJ02jLVaGdMDhN+3XzNxD8Q61z5IYHbt+Lgyh6AsI59
a6xS4JASLwZ2d1yHHd/NcdoARqIb0Mtcj4eE3ckqIkaKyBdWp5m0x18sxCwWR9tr
WIjaI+8B/VJKxhUlRt38J7LmPevz32hKAw/UTEw57AUKfICOLzjsoKAM35C2A5Jk
47sCyR3ysF9nRehRUcuIU+elma6VDw17yUhbEhlscCC/3wsqIIcU3QQ/dMLWuVj4
rp8Io0hqp8qwgH6No8QjrgYoEaE1rrRd4CzhlSXEcrHFIoDtsSRmt6anUm50GNZc
EszY6XAuNShtF6mRvSUlTFov4CYrZ6G+5hLcFjkwDoLzl3JeubkG+NUWecTV0Sam
5rh46r0WcUCpnC53Owclu224JMVypkNSVfg2TgnkOsaCznkuZEzVEeJlymfxakYo
zetl/fvVTnU1PS1SeLoyKEgVKpspN3t6V6a4d9VvKCqJATSSIMgTAvPZsC/dUdD1
ZcL/apl4ApasfzaNjAR1rtk84LSyt3MBQ3FoLX//xpjhKvNGjGdtu3t1Q2B2L8fu
OyMKwsWaYa4hXI01CpCq8kYK1h9nK4r+Y/YvgPIsgk2ZvfFLQTEUOq08DhpXFG7U
Sy39Q1dvP3LC3hbR++DRrEGs8/x669j6N0hU+C73+HME6YQxQhjCnPVWspyOHGKX
RMdCBsJmf5zrDsQ61tTmzuzkVkvUlZNCj1eQaV+rfoqebSf+jmHwKU7KAKbZ6GrO
NdnFzogB1aLSSi98OPnwYn3rhbTWtv2oV6vvuPD7iswMBDyaVmQWXOGvev/Kgw/R
JHKBGNJ2Rk16NqrA7W1cugqNb5UrKlBg8UdoqaMGKWRtTfqREzbh4tqeOLOcdUpM
c1M7FBOmDVQQs+RIgqYK00ItLet3pZc6t9DZAdduiLOQZuXlpNoVoEnO9Lb9jcg+
uJZRJTor3YmxNO2onGaHf3XHNdAcKcbSwgnP2oFxrGGHMkOjB2JGvOFOhTRr05xM
nLqXRDgNdVC12hhVoNxXw1tf9cSCima2z8uwNj9XZRFG9w5iw5RoCjbvT4hM3wil
QxjsMw45QSAMC+rrmbGp9FnFkwENU/k9UegyFazUgeOVHNd/zDZ6kwBsyZUWOtrU
OlWaRUa+X0e3at+EKQlqbgr7Im/465W9RLuG7A3GdTuGQ2yobn3tfjAsaWJbQsH8
REvoD7DhhLMDo43t2RdtvY0/2vxJWYecAGHrI5Pcpahd56qSPMJL3G7AJPtHC7N2
7q+t5v5dGpjuV3w2YYQnR40O6BP4FFhBTPZklYxwniKzKSqWDxFFPWI2vHAvTKdE
IbIhHJUtmFcK/8DsWUA9PyEcEOv/L8Tj3Gphuit8hJKVV7SdFJW88setzpswEJkn
+BilT2faUCMRuKxTGlHZVNV0i6bcFP62f3Dk3TY10Wh+WS3vV5Oqp+7HsMIRby3i
JFLIYaikSWA2qaLU0Ero4ZhY7YP/wIzxyNUSZTvAXpnBw6CcvCN0JvQf5US7F9Bf
SyR8gYIMuK1RPDkKhdU1c0WiYm3bniLsUrfQugUIi2QbYWAcuryL8Pnh7olYiLHQ
x2XXVLZVWM7NA8nl5z7YD3kfkIFiOur61f/HU5npe0nWjCyUurX2+suqRjWbFc5/
HDDTS+8FgzdkGwXuiLIEHg0OllA1dk4zmYsQW9fH2jSFTTalQ1L9KeBuH3/F6TMz
6+9p8mno5QR661Nh0UOTAXGY6XZEywIv8QfEv73JY2OqHcDAHaG9RqZ3uPBMJKQs
Xd+HTwe08B3AoTC+m5FUf9LHy8rnhaeZByV5ypHL21iQBlqOJjqxopIuYndrkB7I
+ZJAFhweh/V3HEN22EPDa+ZGOR7WyjTJG4Umun5lyDTylVFcQGG5uZwUiOQ7nWWc
w5f1PKzfuu9/CvPTyurpvHAFnhZyebnpYlBs5I79M7abbKRWqz5mh71Tp/qZfXJL
d3PUnJHzraqTS6qk1xh8igXepnuX7TZ0rpFqmXn0zf+TIalg5+NcS3CoixuKsFGA
GVmfdRuA/FlZ3oXfTLbabSE6Ds56Pp10wo0rtThNNGzyCiNuW8SIzuyybKTNlXVX
C44FXBNI2LBry/vHYt5ykK7RN0jOsyvzCb/hq/6VuHVsrl5oA6yDTB/z1k3fSF2+
ilQUkqpR3kweA3e1q3pJE3Ulp7KnwS/4DNBL4n2BZHeaTAM+g5aM4ZHDbWE3g+cO
D5grbyTOnuKW4NSquLTRoHZk/21qlSnBo8Hlv7NTiPfh7L/YVHFcmcfWu+QXUixh
M5G8nq1ljFHY6X/9gdnsyjMRU9R6L/wFZSp0bnqnFfCdxnVDGEy1DAMR5q1XOGh6
UcJESfrPdgDZzkrKwlrR1tOwp2qRwIHYKfjPM/W4wdxUtdPnlxLcdb80e9MHCc6b
r/vkJruRKW8VM/5zqtYelpVV9VSodiCGYwAZ7L37jp0vc5mw2qDhNxW6ZTdpJXJh
+SomWIwN/I3UbACJZLaIHHsEFtdyB3Ll7taXdtGG9zKCvwWmzIJFYIjCtEpP0P9H
F4cxhEU2p5v8yFaVfC0TWXH7p3dqiLtyUBmZKm4pP79WlS/IDvVVNmNKPNdsEmkT
WpTVD2cD7ecHEnqBfFZdmf1Z3LvgNYmiB2TD26QmxCehAQhYPDt3vNfUk38rhwc2
m4NqcT6WQhg1jrnldPXo47XS8+v7fCQFG8rhZ4ctUImLHH0GTP4KumzDOTFXR/PF
sp6J0ee8wHKKiu3HYETx7MUDJaTPrR0X2sORGZgt9F2PfzfURt/oL/OME5ZS7PdQ
rl3L+slkg8f/Q6x7eHNcee3j4fP7kgCvf+sxy37JbwTy2Z2zZcGggJjmazIAMzqQ
2gA4zv5ktarERBy8jMMtGVnWCpknZacwMYOlAS/J0KNJmf7ZEfr+3o1yFf0yfRL1
AepJ8Ia5c/WboLmSSLBFZ6TzpgaWWt3JmI89e0ug2YK6LTWbyHV4lXdjn06UJhlx
wS5DezGepFfiDiLD6/6zHHqEN9L2weckI3kUh7JFTk+8UtcTjknxsH0R0X+cuvrx
UzMceqrpevnO2UrGAiJSyFXCRxwTjDQEq3fVJ35lLWbx3KSSbOeI5Ojp4IGfIp/w
tM044URLCasubt5b8ZFWpjZuYzWCr2n6KjL+yw30ZHVb8twTbrdhZKBd1dAFu5jY
dEOHzuhPryaUNtoGcnuGL2mej4WSg9f03l7mZZXCtURXZjS8uu5dPJAM1A9b2f2c
xO+hw8lNKwHy6jCEyLa2Cq7IvsIakZW5LmOK3tv88XhdyFvaJ0+oRSt81fXV2csN
CzWdaOoy/tBpGZ3TCqxQBHstiWbFUSfm9b1QTC2fBqKsQM6bBaBXOjkCXj5MKbNj
fYuLVmJNPWAGmhidbcxgD3daNP320gNwuu/hW40Jin4P+Nj/rGUsoeQG/VEFoKHQ
TzCIDXqY+YsOTnEB6ODdaLP5OTWfwRqFasw8tlyZevWJ5yTe58M+kV68+nsyE9MY
zwrBQZXCLqoe7wEecuemlIJVbx2hsfCsBvcrhNQxmv+xJCPNj5XLuy+FGknVJUTR
LCUuSXGUMVJGUdxZ4BCS65Y1elFuhF7nEdb6ANI32CNTIG11CYDt3wHMmZwQ/ylK
2AZasrhj2cZPN6n+rH0R5yaa4wSa2bG/nupWdmMhL3xTfUGMh3+PEFmZvsfqHRLq
y5JjzntABqPgCX4XdnrHEmexlI4S4p7rKAnfr6wcdtF0e6psTCehvB/6kpcbyusu
qC/joq9B3ir0KDttWjtFiGAm2aeaX1wGc3Yic7mWS8tA1A0ei/Li53b/+JZF7EAD
zfYE+/wPF0rDwyH63L6NELK7sKx5McrnQypPRkgR8/qNSD14XOxGJbmIej0b3sYr
PPUkrEupXuYib8LRt5+4VVFLP42E84cxESeknvBaIWHYHyB0sfR5IML/k6PYEagL
3rYqQ1PYZHpHfcSSBLTcrLFb2vekPnJf2DgFFj8JHX4ck4FkbWN8jn/ZlU6xLgFT
e4Cd/Aowsbov9CsrCvLTLGm2M4UemdBwXR6XtFSD+zhvtR8ZZ/4oMszBSA2R0MrH
K15AfSP0lILfFaMmNcIh49Vb3erYREExpQ9+AAq7OCzg3/ZAd79psakUXxoIF/KA
d+2H/VHecMZY77caNUIrndmRVazR5m1JXrzYf9TQeBuugY25jv71pibwxtMJ6snc
XjIEKgmbNxDbwDRQWeV9oVJ+NZHRkh4tfUPGG+01PZGJWAGreVJDDBCAJIcwdKe+
Hn5mCKKWH/M6AmSF4slAvFQUdfSxQVib+6TqHTneUD1raHJaYO/Ng0u/L83Xd9wC
cMd1+I6iCogPv2JdgipdowGTiKQ/4RdRA2zz7Q+iTqwb6NDoIH1vWfXJCtCKjLYl
v9KMR4LMXEG97D5ESlVUkJZ1TReqDe4RNMhdaLDZWC+Y3DnhVkD+P8i1qbmuRoqj
2UFKO0WHDMR4JZqHyI7OaCzl5zMNPm4Vkz4Hvl6I2/Ei4xxUs8O9P7lUoOYi/Udi
G+c3dxa2WPyAhpIVpCrdKrxNOUC3aInkAW5Z6QS0mU4noRbfZaW/aOAxzJKJmBh4
SDQdcrS0aMil+AAf9zIJtxK+CyWdsxkB2+nxAEL0JnzoshsEupbd7pisKDp5MmMD
GY57uhxYa5Z5nKvGkw3YEipa+qDHmOPxg6koBGxdoOfad/um1FQAR85cdMsdYncX
y/lA513i8CnoKiXiyJDHB7bm4Bq7roffJL6ScSZGF9ChxyROcav6AhGNnZEj9Odl
/BfOMvoyLLyBYtN2SVnS8EGurekV9Oau/R5XN3CsuifwdBqKkfwQbYWZYv4anqtl
TQnCiBKCthUFzMdw/syTzHm5osmfSZ8tHfSN2bD2ZLZ+VnRCmTXJGESKk2lpmps3
yugE9dgjAiFB3muZQpYh3CMHvdMQ1aBD3jDfue9mc+VRI7alIvDjxbbAQJ7i4iYG
1LFuiG6yMfw38wbewnHb9xDZhujgLy0jfQAV2pYUfOdGldItRWVFC4JMkmtV2Pme
Swsd2T445OUN4tDrQ9x+KmhAeJMQpUO7K4tMei2vSFkwBObhhzjzqW/0enLDulbK
z9FhKaoTSxyAhF/lsL20jdaoI4vvvJTomcS1o1fwhTYe7QwjV5YDLXqRMvWnkAlF
mVDQpocuyV/Djyqu9UoX7alUPCn8GQ81vwng2s3E3EYpELMsMsFPTuJVR3qNMI7/
uCmWVH9xaWx9GcxJCiSYscAxsVk86DlUFCWNZEU9qIwL3SFyUMtQ9T2YSijJutco
ijmMH9XUTdbj4GvZ4S8h3nRTxp62t2Pva6xxZ24WUZOk4VEFKafcTa2lcKutpsg6
FebG8GSi3eEsgzbkZr4nJDo80Be3OBMRRjFT2fyNvccpLQ9fc0pbYNCFQPKE7U9Y
1JajBW/LMm2FKDW/h0Hoi//KeLbjTF3ZmPwlcDfnmmBmUBXNscqWUhL05H8lDrgd
nSH6iuKFCM6Ek+KdCpCu2+fK5Olm+q36DAL2sqZfIW2Wuy3kDx/p7f426xjtn0YF
BRaK2DNGHuUXqLUjarjV2NH0SL7dHIxg/7/PfPzSlrXe5rvG47q2Bftv1y7M2Woy
Qm5iP8wfsXQgmUi9NX2lDNKpfVwW5aEr807EhnkOVCkmeBJypXrSK2iTM8gNdzci
i7CZhozVSZ3xFga4bFX3F7wvh/1gUDAiZdI/bkkyXm7Gz/OPT2zQGLmgpl2ZRXbq
w3rw8+GK9TYWkBfHTxbKLRTIOZY/983fsjPMYlU97G1Bgp4R7l/Xj4xk2x+ET4T5
fpNCc7lXhtyPebPbsclBPbUGycL8kvBA9P9xmfsFFoKf3Irv0/u6HAz2u1mzpyC/
UNQIBCavEHc8bMp0E1vpKSvaRkxpGU4lTz/RMpKPWwb2VMiM6e9PUZ+c+YNFx8MC
RPZIlEEC+0mf0MnTzCzd4OlLSfHLg5zAVfcwG1zlyRh0R0GYp8umO/FJKX6jVDno
Mo/HFCJ6HMvi8mT1NLCZP+Ei3Dk7QVI/frqdZOoddAlUnKz6Hz6abaPGBlQO9H91
ahNlhc683Ru66ncPg4OoRLh3U/uiCDRjbulRG5uLNWyZY4+t8OjQ4vGBhV/NpRKj
icxkiLb/UIS1yzmqz/r3oK59hu2+41bPFb6ImRvaLRKpKsPpFK4W3BhvqRmD1shb
6DIA7R2uUk/FMrZXH6/KotSrK7JnyJvOEpc/rsUzS43Qy3v3m3gTeqceaGkPPnlz
rDm9b+ns+MrgWfWqowAqtJXpNHzQqAEec561AbYaeVjjnl9jsusQPvt24oISn0nT
jqkR/yn4X9JGGAa/irODrGaAjXZ+CczONkpe4GxUEczwYFdz2EawQ0/zsBUuIZ2F
DsRH0/VpTCEPitPEO5i3BfdiuyPHrH4fqu9bqUm07PdP9wDoWkV4OhCaiq3c8coh
FngbVBM8Ua1shNhx0zjgMtm5CchSiYCPUBzuZiwzmiMMyX/oS1XT5FpBkR5Vsd7+
QG6zoZhvnSUvuYFBeelahdzlrmb/77o7PP2RQwGKLAIX5gEg/yflOmKphr3z6dF8
Uy41OTmTPBJQzNDXzJ3Z62WMA4Bgq/L4sXP0hWkWxwRR5bOccfT7p0QtZBNwGRfk
GDSY+jR7C+HPn7XxtwtNMUt/DEQsRTyA8Y5P+ZRTehkELgJWQUQT0NEXAYN7fz7w
pmNVSLb8sFO0cFhgQ6l6XV6BDGvTt678z9wsfv5A8hX8m7LO51/oL2mKxeJKLh5g
hFTLVkJYbjPz1YRAciyUj9KfgE7n36RVoATdKnOGPtDqybcboQc7Bxs3dFKfgL+P
ecWYZIWRiVUpfV2p7Qo8QIVDN7KvPgMzlumKgVB7XE3+JUZGps+sumRubi7+AVEE
AdO/VfaAXzU7nmUFyPPCllYENKyRev1B5ZKQ8PeiZlV7xD1m2K1xbAuzWx5Ojl6f
TO3IBTZu5jDYtOryrqQrUq+2hNfF4WWiuBQ8G8rew6wsjxdx5CJIa9wxsgif+zMg
knzX029UWM23n5SRfeBG90o7hg6B1wAhX1tGDG9SUHamUk3PLSp+loz3pGPvTU5A
Du1b5K3j92RzajXHgzY0ecCodYPYmTm4S54y2GT8xzrl8u+IrQ71qACFcyTVv7Hq
lshfjLjs/eVFQKiGOzJiTHw7mKlVXstzNh1zgmDDTBmlUqSfVXIxK9G26Q2kl2gp
im0ozxBESXj8+pfGJZNnIS6lWndS0dqDDeKeHUUJDYPgkQ7V1xK5GiXVJ1YD6w4D
g9d+TtGBFBizEsv5GPJAWNe5Dc0YFUmczV81q7MuQ2nLjhV/w44g8zi8yWnzAQuM
BoQZJ04IbF6xTNu/1b8jbHD8m/bW9y/j6obTVK4GUNuxblhbonHmae4CUZ+6WmUG
Iow3Scf1xRdAdpJqNAZCClu4tZqJguFhJWyOg270+0dJvJN07fuc3zTAGKadqO/K
CmkBlkVcMJ/aFerWeQCMXTmBIwNNk5pzF0cF/MkMig4d9XyVekNgE+5d0BZoi7am
Peq57U+LAHMwkceLUo27zg7Ll2ahf2MWhtCq4fGEv5LFUEQ/aLNa3TwOgSGoH4ij
pNeoLMmUzdkU+OwN2iyWFrveZmomGP5KnYOcydJRtbBq4w7MOOLemOiQZNCuExuR
y9gDnOIdimtzf58/WVQAAfw4kY9CUgTgo4mZ0FnQg13L84KYeULw5+l5KjNALxhL
/Z+Qu+UMk7coQmsUSV3eRBCVIawCXVK82BSMh4EN9YsQXqvv3u7zvJuEOfaTZ5yP
iugSdj0LCc2CGCs6QIHQmsY1PJOKp1jrAml3D/cVqrJo3CbKfC7olj+nMfeg8+dA
oHqYQJG5GCwR71XvO1G/LXqA3YKYip6JxnmZPSRNT8qQMM7u8I7Gf8zof/2Dwza8
1PsUVzM/+1DB78thtxdCjahVnUT10KoTOWhYrXRI2OgAES5kztH5H6H46gO2GM7l
ZaYnsmAIR0o6ZKCp3uG+J7dk0GhS5a4McMrRLEVOM9VVBnrRRuGqDubaqj/L1ynS
PzZmCUbwRrpGM6+tJMgbEUmx5ZJKu/UDVNDDQ0Z++jE0/ACW2Et5bulqp7/ltrQJ
OJGGTc40e2smrth2yProykO+X7DZB7X5Xubz4nQXChq57nmdERyQSwTcMhkAKsN0
epJIYRLMOb3gp0cgg8K1R9hUId672EQl1FVif8god+wn084b4ZIrQSnsjYCJu6xq
ruAB8fNdNNV24DN2/9uON0AkQXQY306QxqL/Ca+zEob3t6HMT3jANYmmTu9WrWVC
D5UfwPw2VaMUdJeWf8Ror80gzAwWkHOG+e2Ogx0Ezco+bFCDcNGe5JGwtmlV62Qj
dqpX+/O8Yf9c7dTht9TyTED2fVJBJdl5my+P4u92AKcKkcBadF2aqLFpQq2BqEAx
emq/evUAEK7ItHRGlHdgT4juB+HevWIJU8/dDNTIIJ6ac54QxGQsIoqv4n3+v7X0
v0RW9DpePq5twWVeCJouwsNnLvfoQUFXYaRLEf2CxRW5P4m5pYwmtVC7QD641vxH
DCKuDmHfJaHGkNSXPq+xTMqiNQ2YfSgE0o+YmdAR0kyJMOLw0FvE81iWB4zgbMXW
C9zG1VRXo6bHwgNhURfySJE4wUEgDyNXDLxFqrDT4Ki4yZDbhCHAFhjSB/vjJ+nq
1QTo/ypEs39kgGMqYkRNQfuh7HZYRWaIN+KZH1h5UOgX9GlmfiAgTymF7rfiCFaS
drKq+RdCgGnyQT/RQe7EAXoIfV82/Rbcnofcz24KM6KW1cTg2stTpcCYguNqNUNU
IXQQ6ZrsaCPgkPvNkygrJVhV7KFwlopWkceo++OFxynW6HOdEL/+HPy2MracfO2p
ct9etT+/8D8BYf5otpu/Pms5JZdkrDZd8SsU8XJewfDkkn++Yakl5OWRIa+O2IxB
NAUGTkKdpkyQqyY1Y2reGiS1zYCPLiutCe2n5pRE80oVnJPv5RqdvZgo+NFJopaf
ux1V+gYGWXACYY8oc1W3grJdhXl1HfFzyc4QrpFg53jkeMf5FoHwFSHvlaanfzor
8NkpE5XalZ+p5Wvkda31v9SnGRrD/5aX3SwRDruPGEj99x6JyHIn7FiPDWtfqxAd
OywGFT60ZtbW/SV9tqI5BMDS8QCkZSEKsk/0OWQb1pBqHnZBScFY8N0jAZR23Koj
rFWwjCh9wkO8mTHX9TShVEJvZaW+02shYedEeIunfoWuKB+2605C4JmUP6zS7xET
2l73mYl+qKJFmj9gG5XTbDcfnMIt8JZrJg+ymZrTaM70qenVGjYb+JPbghsUUT3y
QRErzh+uOAM0f06yI65VN+gPCSA3870dA7t96C7vW44YzoWqPAPX/NtpIvyjqAcD
CbWBZ8AhIDoXGXdtvSkbLuMaADcLjsHEOpO57LrpoOyUjc4QvUg3FaKvs6+WVyK+
yKvVTd74mXV/aDMMV8Fv4IOEq+aM0h0ptLN8gvBwYJfyrB5zfqyzeC53rOOyTBx9
RvUjPJbjR9qKsioWyfXk12gwMH6y4Y4wIiKmQPbOWWmft3UVOxtUAPT90obM65Xr
O82qjtmwHaKQiHMX2vSfwMrE9W5j17SWIY44kBL7gzDr6pn42F2DwVu85Sn462pS
b/KYJ4ZRjdBSz99gpUE53QlTOGkFOf6YUYXp7jWDM50/lk+ElqKmZZv+hyA5bppa
F5ScjmRFI6Vbr4kQb4Q3H6OqHpfD4YfrT4b9PJ7e8iSuEBBPqybyJRVrI5qyNnJW
nSc3si/5ewe66C9FjAkZItPRVoxJlrAWM8oiXr2eJm+kbMHis9A5ZhS4X/CNGUpI
gV5xQpZESzQ3M6z1zCi/T3jnDu2wVlUN8TQsfroTwWbwUTPgPs7v7fVU+xuRU27O
+cOTEaBM2SkT4HdeXDB/RCZ6Fe3LvF/aGWE7mPcq8xU4qLUZY0AoKv+kGHeyeRHj
f2PDkj0p4PoJ1p7ADDOmqaEbCZIHLJHByresa5oyaDHqPOIlNKBPuV3WVFvYkNTm
jBQN2Ddu4lt8THZJGYhUTSkHAKOSn/0g3HWLbax+bzBU87So2RWCrsH0YtcdTVbh
aqWWCP4+4Cz9aSl4awvNNBZa+1zl0SOLG4j6qgrlv2jhkn3a3kKChBbwBuzUonu5
MqYyAPR75AFiqF5QopY6pxv3v7/PqIimUq2d3MdfEovaEH8XEKh3bEz+ailVrDxO
+1z4/sDmjt4x52pl2GZaGo75I4LXctx6s87asBYOGGVTHS15N27T2JL9vZbbw8Cx
7i7WHl2I1V3h0Mm9kTPILbOr+VnHIvjbUAXIAbYusZpiwt8nQDdA942S1oDC6Lyw
7nr3InQGHJrM3KAPjfIT+tB4TF/+NY24X+WLBTXeXxpF6FwGNlypIocNhif/bL0i
WtFIfE5Uo4GleorKUbX065MZCRihlzy8KLQFhlQBnHIFU8SRf4bntqfyfC0iwFhb
c0Nr6deyPB5df90HZJmFBRKDa2/et/O+My+/S7jpLNz6Bihzu/WTPQLlulydKZgh
Nq4RDtUiZzgPZcK2sSWRbp6NhRuROt3vQLqPYZiWrFL9/4MWtkTH01l/5ASV7Re5
iRkITaTbmTLWD+bYQhwh8FmET+D1p8IA88c+6Vgd3iuDx0MghUOfDZZKNPmkHV83
SEyKf9a4cAf/xP/MmpGHt7/G9FfsL6pZogXpGF5ATE7VVg/KXOElyK9ML+ZCjraE
CkitCP8AYK247+nqEWfxUMtaeEV+KNqp8caoBPgTp+j1XdCzpDQHT9odQKSjHgUB
Qz/myqgU5VttZ2k2O5HirFPdB8gS2e9a9E0CIgfdoFm7RANHr9pUlf4Ij/hCuFgm
D5C8KNCgwgFqYQgmAG/oAsLht2JkgE/giKb6MNNrFD//lbzB1Gj3ZG7+yKgi/JYD
WdhCmmzc46bbfNgAme/I81OrF1iYUn97X88IJ+NAMfqGv+SYXEG1+cG1S1m8fkLG
sZhTNb32opaYkJMZya2/X5e1XVQMgb5mSq+eZqYQfiDXQPRncLcuqOP9bOZxOUG/
PkYzm856+e5K0lR0OlD15nKYiGsbjsIB2si3NG7ROnj5SfcPtCkX2ejZd2nC9BQR
77ONf0BZnYSU/Icqa6zpaWLETqfFnF2rwLMxXufCpyFuJBCAKhDaHqfRXZfawdNr
MA5PYgp8J+qMSGLrR6RC2wYmNSYtGyR8MO7rIvc7MVAF/z+RjSJ7h1CEbRSEQeQ7
Ye9cEa40ZZFuJZ3jtSrLn9Pl91YSXTuFLXbTyZoriIyl6/U/gfSQVc9zZubB7qBo
9aMZbiTkA2q53+2F44g+mY2oU8dJcvr2auYBFocl0VX5A75RMbKqzMhnK94xoimf
tEKSckpUua3A32tBNJpbGodZYILLcr1T/LtxVVWd3ljkzuJAHpW7AaOlQ4SH1dfY
dLryelcNg0C6XPhFXQoYVnw39xN3bMcOFN1YPHk3FdIFu88gZUqw2OPm0mpNyjdw
3KgB/JnJ1MxD2BuYF4G/d9QV1X7A9xQqI8997RMSC4vwj0UkDjBhYI50izPV76DK
TThyCJhyiiMc9pXOFl1qspAXKdNr4jwa9vZAnO3JNBevdWJ2Qpq4hkDySRR2jiRq
bOvbqN6Yx+cy6WZD5TgeM7puaC2eFOo/YIACDMsZO0a5rDGLtEhYOsfXYUnawN7E
6qpa/lvqMJ2Sx3RubWgqU4pU0mpcfpTjOES9tYsnU7yPoEdAMZus/kEwfCDsYMDY
jyx0Wy+yrQllSgMZo5CdLiPNpESSYr57eRiNMalTZT0sq5JX6BT/S8YvEQoMlhwj
NAM6fK9tyFFF51VgEsm4E2sSZRFtV3jbkT0iLnOgTHzot9/FYuCeD0/SCr97qW93
qQVHHgypmAuXdLsHHNMueInjZQCQhN3cqCh/Rbw9/cJSubJcx6vE+gZ1GHnfOn6L
mdY7I5KsJPM7ZL/yH5RyH2eYY/breOwXr72Fv03a884kZ6ACzB70pL/oT2CXz3Tb
g2q7EmF/JXcZPJoURxNsn6OrU3nD4K2/6kX5ZmE3rEJZJscFQdGoBny2eg3sTaK0
67ZYvDFDN/3El6QDVH+ygUOwLIJeWAr9bB4demCVSd/didDN1SJH7cj+xl67FOH0
FV0Zte96S4npqkUrHlUzGGmmIaBe12g01eJDPPftioerDY5tO4MWGhuGx7wkNxpi
XnOIy9WaituHpZWNMEy9mU8kQW8tM9RCTF5crQ44TMgq1G+qD5zPVtC3jlkRdd3B
eVakCgbiEbZ1RQD46cAl3h1Fv3/ljYAFlGuSmX/knUZlghaCNo1aybHCBOvKkCtX
nmYf1nPHWxkazzV7oZwSZPGNYutqxcd/kaN3cE2291l63xFELAORJgmNd39Kfecl
0t0G+6ysgFxOFtibbH6J2JI2v5Z7lxNUlkkrPMiXD93Jw/tnG2S77jGj8+Oj9RS0
vILpJYJH9xLtNsNeQk4d5Uds3fOu+RYNiN68C1e5VwwDri7gmfr7fRhCyzVIFjw1
ALaqt77NrMVBhCcdKj5M5y9J9dKCpS/CgyXwS9ASc2nLXK3vebM1muKCuO9e9Xo2
OeaBo6AUCu0XVkaod2OGfPReu0Sl7sfPxT2t1u329hCRVr3RJnf+4Vv0EpqtZveH
o4/lBcfFTntRrV25yNdxdwSh9uftmQMJbbKs9lUC2GgUz84OW0Ky2NF6kn58DWx+
LDHgpWB7RaFThsfdcU4Si443qXO696SBBcV3gnWAUjyQhXzrWTdKHVr2rErpcG9o
Tvq567zny1moX/KV1wOYfXNFxMOeM6rogQX/M49kYEynMcaFvYTpA+lZ0+TikUs7
uanxYgmyI2PKPRR/+ZKZOA40ZIgvvhrIs1M0bqZxutUNCnVQ9Y4K0RJSdrVmOneL
BZ3QwPrzZTOvC606gnRzlEXpNF72jcT68sBlQm+hYkpoHNf94MHAb6iNu82ljiL0
WlgUKydzMV78xQ8YohDCrHwx/6/xrDoPcEFEk8V5dlX7jQ20/zrn8rlyqWRIgj7I
kY8eeBPsIS7VuKn+xb0KKBRTkxHgA6byvZmeUygVJmkSAMKB9KHkjvZrptozCRiV
MJR14ZHnMjXTNliLcc3eJizSExVgrvzN62wMCuVu+t7njmTkb9G+L9/cxe0p4LAt
WnoNKPxoE9YkAoFMHU9QbK2XBpVF9F4ejTga3l9FZAD68DMiyz+2a0VY5Xk8hBZu
ebJmY4elTFrEKBVoBgZi3Inyw6+ACmM8IrMhrOtNTjfw1+9+o6AQqOidrnWDMoVf
8BPaj2zbVjiB3vTn1rQDsxEEzoLyXyb/Xcko1R/I4Vu4StPM3jAmHHrbD1iOfBhD
HKjQAhNCycE8xxM7kIWbN71rmR0VzISIlttNwwzwal3HNJgwzML8QlGFkNy75E3A
1YkHVfI2uwPwjH4xHtUoSYLZsx5FrhvnxO6M60tc/DPUOwBPmkUOmTV3UPNpYP5u
PK+bOpAcuRA+YZPbi5PoMMaEemnKG92JOKWdrcolZb/QPR+uj1RGFlJMb9sv7M5H
DyoAKVenWy3sGFAjBDxfIpasM5sXqSpkS9RWfzouCjxz8PAUCkevO65kxtYBlXZt
U4OKL3Q8T28/An982qoAP19h/l7yQ1oCZW2HzaDb7LrjJWui3cM2QfhR1U8mKaZ4
UpyqRiMpHwhShr/tK25hAKVap2UnoBIEax1Ub4JfAjl2csPFQ+jQKxjIodtXugF3
4SpuzKrIuYD9Q8X2RPjrjRM0kdFom7oHR67SJuj+4USCAFNEOMyvX5BBtFdK+Qo2
usY8HgaWJrV6j0ih3yp9upqdZf0QnnYmj8gA5LnrN5PWpvH8Fjhb7b6/NQH6zhxN
buem64X7eIoU6wSB2XzhBBuvb2qNW51K+xYOgt/D4X4ngvaB9nTp69cNe0HHTat3
KWuDNIPYyT/LXIMerPFc+Ap4TwrvMLZRhlN9O7ewcPje11tlU8vf5MDsSEEeejAp
aErneli82Cv9QUyL1oxqAj4q/rWYrjA/zqAUJzF5NR6AMRaGCYpNXX/i2d8YPlFX
HxFEfuZxGxBC7UvTtQsFBOSnOJFh4sjsryxlBB7R8gT4Ysr3epROhUjuDIAbGX0U
OzQh/l+2quNYbLxvV70eIB5gly7T6drr7hnvWFyxJB96jy/7LAJR9glMAIBZa3za
t/+XJtSAWqdJgGT2LQxxRBmgbGeaxuJZNVRSwYuRFFBsnGOIyHmXNc97uHbC+TVa
wVkcGsC+UjfmCANpT09twOFsn5nV8jPmJXtbqecSQBu8+pfc5bGZy83EA62XGwF1
p2pqp7xtVKlbuQoAKA/AnE29y4qTMX15V+Et+tRMZ15kY46LVFNUYBv/KqFEBV/l
iSanbaDEuEO18AfpPyZHifP72FjxZKCiRgEkJKBSP8g72RAEfuyaLsGkGzb/Rg8+
FFsJCTi2C/BlQQZ2TrkFqMi/nz9RoVURegTwIVlNieq6ZoNnMQsuW9Kw4Iyus4FJ
2WIDHkhuouhSKm8IgxxD164VSp9c+kzeAgMjML0bMzBb8KnG289OY/KBuNBxiMqC
oogZAXXXYqJxKUG5V1QHkj0lu/MvsEz2UeLkUpqdVtjsnhQ/Blqbreu7Fla6Iv9r
h9LjrMmE1DDEn4vfayIjTWaRTFoaLvEK+Oui25Q9ArZmuMHcT72J7xVLSFoReLu/
78YmZv7nfLBtYxHwEN8ImxEvWqyl6NqqwZ7kEZ/Rj/7UV2KWQGf7BUt8g6bwROsl
yiFEtIUYuUavfNWrnBf4D2SY4TyHf4wRbyBKRwP30esOkp3p2IQoVXzl9E0pKnhm
77dCwpxcOfS31f3ZfTAF06o78nudewV6Wxrh1UwovHVOFpxAL1mxUMrHMguM3fi+
qPAaycdM9SBPinnqyCtMY8fhYDAi5b9MxWUoxuQkBtZ+V79g6zRjozDlycka+Tq+
MUl9YfwGpw99xVgEo4BV8oElla/ZnLPzI0qdukZH5eExdLqyNeZrrK+dHc86tlc4
xAsIgHRSFFz1+IzYMDMMkDoVwypt+3JXlr0SoyG4OSn1a5SJBloj/okbj+yJAQSw
AZElavOOyGIiY2428W+gm0Lc7MMJqi9b2YYAtyyyOp/h8dlX0SwGfBPUE+OgshA1
Em/hR6JGTq1W3pxAX0cp+dRYtF0wsh4PtgtGOY9zh55O6MGcq2fhrOuAHpxNn6Zt
10iUqJ4r5Nhag7tsi9Ac38m0Q1dMGb3RWD8DUEmXH/6m82ZdSHQmmu/5Y3UkrSD5
6My4mjGVdRyoQrTLScXYe/uAbESUuZCpFt6AHOu3NOH4NHxAGSRmIB4s4b9ksFZE
PvZNKjQ+eeCcMJAdcU50sw5FrdgkD5BJ7WIi+nfcjhSKGlWE9GTluvJzLfFSdgFR
t4RltGpTE+ecxUocrrXg88yIEzjYYcJFmdMRstg88pYfAmL3LxbSpp9usn+0+sGg
CUexBEYINyeXM9DU6pNjabjPqpzMCsSGPfLQDiIkgeYXtbDCLODunpLbu6RHnDe/
Q434cCKUPM3RByydkBqQrI9kDjjdbTSJ7vyDbhBE/y8=
`protect end_protected