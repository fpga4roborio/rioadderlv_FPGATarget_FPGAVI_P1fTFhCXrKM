`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
ddtXksX2+yylW5zu6QL2Lhnb2d1sD00763mmSITNX595NcHTEkwn0zB1Dry37fOW
FufOhVzEJp80NC5qZ/+F0Vk7Ik02dIR0elf3clrjeJRK85K4e3Hoo4xn7YbFUIms
l/8VZSb14+JVGURjfswrIyCUotIzlzVYZ6gzoZwDXIi5gQIBf/gI+KxNXPaKV+PQ
Ufys/12rjO6aI/pPlqSm0hCvftmBcnezN2hk1UeXgOIuKZnogjOsf0iJVX2aOOWE
6pD/psybjbnsNB6kH5uFTA5frkzIzkzl5d9+YDm9OyC+k84E83I/7/j+rk4L2dah
QJOvksSIzN867/4Qt8qYTQ==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="MvBXkzurAa5VTw+1JJ70nePUfoQXBvZOku/SMmg4TwQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
oRtzZL4VJ4iwysPsC8SXYCzXS8Fw2gtZTOskLcDV+1B9Nzn1zTyNtlo6lNICRmmK
ZRVu2BmCc2G+fmzynYlNTnSa7C0Cuel6FYpxCBlOuk3OF2tzAmLAuDyOH3Z1Yjzk
a0aHuoCdIRKv7BrZCdALt03JeUmXKPdOmIlkVGFl8yw=
`protect rights_digest_method = "sha256"
`protect end_toolblock="Jn9CQpRhJt4rnzZPRk+dOpzAubz7omckX1MrFd4p81o="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 3328 )
`protect data_block
gD6l00tciPUa6pDNTk/+t0OO0nC/UTtBwLB41d4inuAUA3i/ALrNyoJVcBnAmEQW
ptbcNp5fxEUJjnOxnedyZEuEBxWRieZFQnkRdF269oObKqDENW1sCY+xU7xlgP+T
JyG8tlDf+Y2dFz1xRHI8PXlkchwxUKvtsY4JzeWQljb5gQEQES4jTdelZWu4Mjmd
rhsIe+AuuyS4Asec6atTp2XNN3NJPMUPyOkWGwVxzD396qL2iUfleuvok+iaMFD/
PbHKTIv3H7mkRTsQb6T1mTS7h+MNS6lkn2u7Qd3/SyJ9YCgQSjWMZ4xRf+AQsm//
KHlYcCC/yvdIRZJHMOIk7qStd7ATfrcWyCS5lgi46tMCA3cOhV+wseq8Bc8Yp3Hj
+JA4HLRfsMYJQLCDfQKXbQ300DdL8+rh1gFurQiJVXMcRcH15nJ3vVcqkfQ3qMoX
xG+YV2aR7Ko94w69msBkYozfskJgOIFQYm9rHZOBkzAgh8AeDZgRKL77Ke5jYqSv
Y/URXrYxpxE1jj6sjpiSUwDhgqBdGgsjl9BGhl3hi/20SxyHfZWvTujnx07Vl0HR
ggH/TptEU82kE2LK1TkidcD9rJCZI3r4+KjKSFEfHAiZZ2KZeAts2HNUOjZpUo2Z
drCMcY/QMvcw8QmVNkBV4f4eSHxdMr8S+AYJ0m5B/3Dq7YoffL7gghaa4wtkyMsu
4wO0+Q9tWfnxsEARLmwTlhOkw+zSragwGaZ1JgV/c31njGOvgCS0XlDj39ewIJKt
b6fITgfx/I+NUmCyG7wYpWWiBAMZtF8okR9+vnXIpHxShhQAY6wTkRwUgdwYCYhn
54DpHxgsaNA/spDp8bFiOaQJL/PC0FSRbeVu2dLQ1zjGGSJG1uyC3P1lXRIzH83i
wK/HsfrbdaoGHvw6YmT8O/pEJqEFn5PxXzeU4ogd+3RdCF8fTSn9UN16U6OB2By8
Oez3QjKvOKg+SIkS6Gn3CRzuWGdbLMttGqMBDHnKCjc9M9xmBtQR4AEGHCXFekMp
VlaPdtZk2qhwXhqID2vERC16Peo0qNHgsT7j8liSWKLG31oyezHLDZjGsY0FpEkS
LDaONTYuuD+pCjHJxVIx3Xqb4uLzbyoEfbATvtgC5/c2BGJTzMtEzLbXKGJez2JG
XMNtGMLSb1hZJRk5dacO5I58w8/Yx+MgTKaKSOqJkj5I/+iovI/Sd+lLhgH9H5Yh
4cRspfIjQXfe2LjUsNgUERCChzCBOW/wA/DmExzpZAEB6Tpg4BSem19ts3Q6FOao
BbZoGAM6O+CI0NCchToEC7V57lzgd5QVL16p9y2et00MJc2C2ca6sK3xP7xT0jga
dVVTNTU5HQibs5hWXTth2pGSh2Ycp0doVd/SP2EzJdyBaDjq/75pkXx8O5hIL2OD
W59cP/4y+htCiPjNBp06g3YSI7CHgLW8AwN//a/JDlpqHeabo785zVu8kg/St/Jc
+OgOCN42DwWrzi/7uxZ8Ek6hspBO4VgbrTw7fKj9kZ+opHVAIO4ydhtXkln8teI+
/BDq+uwR8ShGyy5bcUWev/UuVCZH+UNl78YZsVmZ0CHiUOq2v2Y0y+yU1DVWuMRU
QkzPd8KVp9qfo5/ahpIyHzA/RzSmCUPWMqmq/csP6eUMYLL4KcJqhze2R0WXucCg
7FGWDG2ngUDAOj+kPEC5jupZvj26oNZEPHT/vMadxQzE5vGiUMEJ6g8vW9wg/Pfs
+6Lj9uHmIgKm5N4H8VUwJy5GuWvp1FVOTEacX+R37uc1ce9gKEIe6bLWtzEEN0Jy
Yu9l8RVovGHNRBXuwuIq14XBXwazM9P/ow7xxO8FNhX8vPUzO4PIuSNJ+WzUUNyZ
s4QdF7zaitXrOsEkQbQHzNTaLC+MeAxRvmulAEIDkIcO8Wh+jzIYWjcDrFAddwV3
S8MYMeA5Vs2iSy1oXRVBBb+IBnQVsJlp42Pt0cj4IY48XxtZHpefhK4bFvecqqfR
HSo7XxFNg1W51eq7qDgn+vICebcg5IRNUitYpNxUdpq/ad0q8j7VZ+AGYpVfSNuk
T0TGy5FfhwC4AUEP33dDr6COxE4Hb0Y+X6hDm01pSN/H5K7hQoz+Edbz3IM7vmX2
kwZLOconwWjmLOSu4wzNGxZGZCTMmSO3M/da/l3GmzP+CRb+E3GQKtCt3t4AKLsJ
LTc6R9GDWxSWhagi8OYYayxVsjFo89mSuA9oU0KDWybIEUJ8FDfdq3zNjUss0/kd
2GEmrdmyw+DssVQtCtnKMJfymTXh/70OGENh59dmUq86FFz3aL16Oo1Qe/U2vKEu
lYD2mLjPEX0l/i7zerIWpVpV3JEcE96oHfLa2G4MY0PxNbpnThB9aezKmHLpejku
V738M8wRlNiIycbu4wZYulC08nE8jmsuiqE6nI2N5db6hzanjMuZDzElfXWpBwr7
NVRKiI6ThRcYucZ5Y0s9MjGIsd+F9fybLULrXLkcOsqlGYXDP6kTSrB1Sf6NkDS9
RmSYeyJEVF5jfG6/zJs0ImKsLvPrFhkInW3WQeQCSKVLtiq6/HjvkYl8HZE3PXcA
1kgiGQHXq9ak2Eatv+7KY4Is6TH1GqLSXyixJdT9A4Rv7B3J91Vhe746CRFksYDQ
Jea60AQweXjYvBYthKLOKElpUuj47Svj5ELOYs9w9Otpoa5z17DrrpXVz6z1elEy
BO+y+YHZAg8mMmBlvSI6HF1jLCAnkxtxoF9MVvv78AHlJYPLN2pA0hmwPgFE2yUF
QSc35x97r/ZniIqdZz/89IDugm9owWhgVaDBzlW/ruV7CkNHaArKa+T4Xd8VAZpK
xWc/UM3iqdHCSTPks2IDMTpxygmGs9RS590JUffjhH5q06aH5GZjsC/QGfLE4S/6
yE4m2VKQvMjPJ/h4npLLHVVxu6Ac1z7gg12pprCf3jhEcgVj4B+KZNerxOSzsFRK
93FiTsbH5Yt8GmnoDSDMyYmQlAAPbTlFoaXqUM49XQWYerq8Keh/FgBCl+i6OxY8
dXpfea45kH59vdONZXyRV2cvpjCCovAWZHoyeQD7wvuYVNIa2StH1xrBjSK0ALlc
9/UOn+tiQcYHr0sL2OMDqyNnIqzCgEbjROSuLM7lQcTOQ5SLkFqi1Pd9JEeIDluG
HtWFGRzk3sxlVMirqQd9Eo993S2upOjR6gn8Ctx52iTIueku5uP20vaEY3SzjpUR
fgR3UQN9zqXwEab5qAdI3QFTYpwFI4A8KNvjWI8ZfrBXFe6TzDksb1LL9ylIuixR
7TPAYN2RrQ6COI5EvVLKPnlzI4h889grWNYuYQgxDqkYobKi8EK9D7s/++v+l4Sp
//Y+4vrzuWrkTBas4YnpyprkqpdBlfBrEOzxIggj2MhIMAnuyK6fm+JjYAUYhDft
fgkA5CYPTCRopyuCL1tSZko+g5sSWoLahzH3jMnTtTltRWv3qRl7a3K8E8YGNM7T
hmT7OBQ4ZCOf3aypRc1U6mCU62cJelx1N9sIDWlc4S0PstrhKbt2bUIfjKsb1BQV
iNKcD3DC02h7HoMfr5FRRoPyhkO9CDq3/1IbI/ihzDEfJXv0MmKUz3ZUIoApP5/b
AC8Y3n73JKYU9c8zF6z9z3VHMzzSp6+jKTRsDAMIFV6+j1eIR7/FI/R5DQdOonSr
EoVvzwFr87mM7iVOQqwiLf9kJpr1BRXgZW/eZp82QyH0m8HabbnPN5Bz37m58kBP
rqzHDON0XXf3B5Ei3MR5x7wNpDym5gzScyldUkUl42wSt3dWki++rbCawtOmt1iM
NThHV1Dm2djx0Wqvsusp2ue0JdRpeu1I0PVOTa1TMhH7AdOvWo9c/iyEbIu/LwjP
wT9dEXu97RDc58E3hifMxwOSGSYAhr2+CV8eaJVrqbP5iGqGTt+Ed+JdbqfQzMNf
0CFGEBq8TpkQ8BhLOGYSHmu1d87zf5Jse+qv48DFFhR4mPYgqyJkOrnTJTCoxZ4J
sEu2Ean7Z6arj1mIRDEi0u/QTXWHOSmEsORqoX8XM2wuE434C2DoJi0wzCSqRKFe
5ND9gV44yK/eB2/Oc0wsTIPfRM5g6AlAVDirrdO2juE0rEDcf3Q+Zc27w6QUa6c0
S6dFVlMQ3Y7jWl+oTouR+/f4WJQhCl+5ogqqkmiesXRe7E4sUV8wHjMMqDWEjLEN
3fXnmgHGfXNC80U7vKExVnllFtDAfNWxyGYgTTdzzbLI8Oh1dtX0RKLLHyu+W03Q
VeeaBfDDVIIKw/5dNz4WaIsEZOOiToCKB4d+S2xN0R3AelvQXb2TZqlbtslMfWq6
XKuM6nIMfFgDjA6/s9fQ3hyW26BpDy/708jMStfOKaTKD5Vjq6iYpNdyCxBxlyn1
x5QGAm9SY3nJs/Kw2OPbg7euXbYbs/R2/QRgatHNhv5xpHrQAoxjiKiZYTiQ/FFe
/I0ZJfUmYyiH6JDQzbPPhg==
`protect end_protected