`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
ddtXksX2+yylW5zu6QL2Lhnb2d1sD00763mmSITNX595NcHTEkwn0zB1Dry37fOW
FufOhVzEJp80NC5qZ/+F0Vk7Ik02dIR0elf3clrjeJRK85K4e3Hoo4xn7YbFUIms
l/8VZSb14+JVGURjfswrIyCUotIzlzVYZ6gzoZwDXIi5gQIBf/gI+KxNXPaKV+PQ
Ufys/12rjO6aI/pPlqSm0hCvftmBcnezN2hk1UeXgOIuKZnogjOsf0iJVX2aOOWE
6pD/psybjbnsNB6kH5uFTA5frkzIzkzl5d9+YDm9OyC+k84E83I/7/j+rk4L2dah
QJOvksSIzN867/4Qt8qYTQ==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="MvBXkzurAa5VTw+1JJ70nePUfoQXBvZOku/SMmg4TwQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
oRtzZL4VJ4iwysPsC8SXYCzXS8Fw2gtZTOskLcDV+1B9Nzn1zTyNtlo6lNICRmmK
ZRVu2BmCc2G+fmzynYlNTnSa7C0Cuel6FYpxCBlOuk3OF2tzAmLAuDyOH3Z1Yjzk
a0aHuoCdIRKv7BrZCdALt03JeUmXKPdOmIlkVGFl8yw=
`protect rights_digest_method = "sha256"
`protect end_toolblock="Jn9CQpRhJt4rnzZPRk+dOpzAubz7omckX1MrFd4p81o="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 19488 )
`protect data_block
gD6l00tciPUa6pDNTk/+t0OO0nC/UTtBwLB41d4inuAUA3i/ALrNyoJVcBnAmEQW
ptbcNp5fxEUJjnOxnedyZEuEBxWRieZFQnkRdF269oPrzsuFB1KndM0bwPp5pxcN
fgMkqtSm7S9fOg90HIZoZRTvC+5pwJOjohEnqQFipf6rAROAMclTUQhcRnGIfqMg
gji+av07xBcWlNjqFvC8CNy7ZrWuKwV/Eu+jHlZOFb4GIUIFvQGMghYUaeSG4ul2
bxyUWEwdwOmxfYnH0W/NPer+QKkf8XJQOQ4skoH3LItcT2nkU5G/xNaAneq+FZha
UbAAxtRlIFGrYYoFqGoFyNmvtkaBbOa5X73+itRbbioGLEaKN8kXURM0gRufW242
y1hCHo/7dexZ31FmPhPaBvMwmUZpN8Oc0DwfWafKpqK9fXYihOr0aKezFWvDdhU3
gJH003U+mwcVsoR94ngCuTt3InumjiBjF7zUGtpN2m3IwSv+nxaBiCNFhz+R65zK
SUmxNPb59lRrfUW59SilGpilryRsL1rH2NDHBrzTvOCpGrlzlvhClI1WC5Kz02jU
KR0xJVWVe5lDhUATlO3UlqCsWkQ6vU1fvg916vQTMGzp/+xx5x9SGbr42YvSX+r+
FoO4dwgrAhOTc/+DpirpX2qlSfjaasRN5rP2WyTnF5yGHJAdotLWAmqUEmt3gIvl
um7Av1jikPMFvXNPjGmbTNa5zLXq4y5C4Q1Ybq1SuyQaTBXy8MlFakgLQ02R/xJT
UQGJT93dG4EYyFKTZ/jHuSQnFE9yBktMLgciv8xPGXZao5IsNzEUzbzIwMoz2/Tf
Fe8L3wXb4/Bh/Tt3Du5hytQaoceZU+dtoqbosMoVX4V1zBEVs7m1LXYta8Fao7Fb
nqRjKmWsGv/3Toika/0jV2QP1x7PSTjaSl/zDDtnQdbH6uQ0m0DWCnfJrQT/uwYt
r4er8IuJzmiaCA6vX+sIqlzADNCJ9sOM/Y8jNy6OeHRGcy4I+3cj0jLaN8VPfYGl
XMWtsy+Op6znwLVxhnr4bk9Z6iI/QSV8SbyLJ71obZUbvRHC+K/ARpUG+/3OSlgw
ZnQBM8Cs8EwPjBohFqqPAy4Th9l5u7ee7Dipr6vx8oJdsDHCdmJEWkD108GWDYo4
fp0Q4zC0NQXUQLQ5DVCdvzYOBcfiepwOZkGUKWQruoEBkZ92QlOWSTDV6Sp1RBDD
nEW/Srhypd+KarpktgMt5RHzdRJSk4njlQXvsMQ3bBBn+ws8PX8gIKcwb/17HwsG
j+97VvLoWGl/M42QZLEzNCHJ4HcXjkF2g3mOYlekiihOi57wBHOeojpE6BOl8A7r
XRTD3rZv8cAmMEPG552aufw2rxtIJ+3uYbZokKSaB3Wzzv7iTZdkikdkTprzrO5g
QvhjtQRudHevwVFUYsBWqBYA1UJCGZ+8+mtyIGygU2xKhWuyVZDBxdT8GPLbFB49
EEdQsUCIMfcpaYkLILy5qSSyVpszk2YCA6TQZfNxbjmh+cS+nsvHc7QMm1YsiLZ/
4KCRRYexadhJBBSzr97f9IFjKQKN8lOMsyXUHINFXSdyDlz+O7ZykuWRS0fNZu/+
rtAo/C76ChmAy92m7tunAPenIAgk3nXBDbxKrupQMlavngfVh5nKl3W1RzmpovAK
mGndRQ2EZnrUyi+ik7TMojHUHPw1/GKxAkL3aF8RLPWu324sX9EgJo978v3ZFdwJ
0qfodVanTaN70g5DQNQK2+CEbTVDiW9xH82MHzD3G53Iwwqf+yg7pp5mqmbrI+HB
ghwfYXKsYxsmhgEpfQB4q3lDjg4oU2UyPohkFCin6VXBBqDPoqbki36/I/YTq7Tq
sogx1tAdx144D/xh5ZRuZjgqRkAVFXnhVPkQ7nxkazJBblZumEytFrlnBbVaM2fl
cey0Bq4ZldnhzIqIq40X1Rp5uy32X8kpMPvIaZkHkuSmiA/MPY9uK3UL8II6MHx0
xK7rq/k8pX+Chb47hnSVN3/eoVFEgkT2QzvBrWk5QdZPS3pm7kDiguZnaZG5HNCT
IeDS299TRRAt6Zef6AGI39fIQ5OoBYBWOFcIN+x3N1UURRbvWadUx0lvL21kgLYp
nNmnCIPw7VqPo9lAAKmf6yljOV1VVPXtnft6G8VfW5lH2z8mPO/EbA/vnpg3eekG
TDmWmSoY7qIF2mIZ2T1DxUdTYgL5s8jC+8iLnVVc8X8BwEf15EWlHRcHgzpOgDja
JIkPDgkcbUS4q0EchmL6hSUjnm5XEQNuMVMr7dlc0B3wp4sWUMXgOkBZTda8q1gq
/DmhVhyzGo4UKSDlgs3IYyC8vt71SnYDNUYOX/O8ZVgcYOCod8PojA72CHbLNzBU
O85SP1mIh5oKIuTqCeIoUwA9X1Jc3GA6/9GayE8YFIBWKMGA8M7vH127JxOOYLtA
1ZdV5GqIT2jrid1yf8lcgVYL+XmQiJ5J86ldNa5o+lQXtssoQYSAwg67RUDadeCI
TEybR0dU/zJnelR3RKn9Jx3BUSHkXPk+4K7enANlqIuRRRhyCCYUgxZzpfL7GHY3
zTg0k2GdQ7lmXyAocbn2w+N2MH6vNLY+HAWNDCQJ8DH2yxQSFvs0xWMEzTGta1Nu
bj+QiB3Uw30NsmUU972BjrLJ9EC1jiVyNUXcRfTQZt2Cwp4OyMHtqftv9VCY4ZOi
V9VxyY/noT30D4JYllbtA/N2vUIkRFmzyTbnYSubHJ+g/pfB+c7DKvhVBfCWS3J6
IjDltQCJVn0fyueYf99hty2tX+T3+s+KwiQ2gdutWr58opy2gM7V47jg10NtchvO
KLhRmum7Rbbze7zDjT/9C6iclwqyCwOuPnDYBeda2zqr1Ig83tu10bOLM/K5++nQ
Y6fiKnTW9471hhkkSsv+OMAsl99njREcxQdTjun+rm+5Iw7V2S0NMJ97zylTUhBE
WYyy3bKPiU8eIdDbUyFO+e+sHa2x/kcHK7bDVVHu+sV6GlSFoZKnD/zrCNiAwJYl
yCFGjkx9sr8TDO6T2QwTY2esNXxRt1Y2nV0pAkFYUQ/Fm0IllBiRkT0v+GUfaejq
QCrpWMoA6OXDvgyg7BXhmgRi3wGudttSEpiNz+36UQF2LKEwqD4MgV//4gCu1H4R
qxJJReUfbuNZJMFnN2SmgjOmnlBnF1I8vg1GTeQc9bteQ1EpYdfWexwnRpBZw+LP
dbDspIVG3InzO6UDzDPg3sknZvpc2EXf/9c7HXAeuE6HI+zDqhqweetIbq5dzvC7
CHEi/ZIbgrG+tb9vZZrFkCWFUMbeOp/hjMWQzEPKHLO4mdEh4YVWO72UT6nzcmwP
YFZ5VFPnHKnaYEVWR67nRdEw4ylx8T6Zj7VPVlAn8d+u9TGspS4OI3WayU7fJNbx
B7R0sxzZ6tiMe9ddiMWz/0OxG1jEeNw0tDg4yVXka3ejW8gZ56rBNIGDZFTeQrw8
AREOpw0eqWjl3MKeLJrgRi+mDYuyddUjbvyjaa9C3Y1DLOrLSHbhFt6EMit11qCF
yOQv5wkDCaR7Hh+aP5gnXbxBGYOGdkKz2iA8gRDRiaTNRTedAmp+/ezY0CtEnmfa
GvSRjQRj8WQ8/LJ0gqSG7jCMqco6MYdfCBKKi1u1LpYBraKHebXmY227VokZ4HiJ
xcCGcdjtFi9gDu7YNAERwGtSV88IYU+D7H0yTRS97HZH0Y7OdepvKFha3x0wYWiT
txCuNUI3ONzgKIXKMD7tuaooDJ1HMm5nQYeNG/iFkHuAaHWpOSfCdGtOKLdTJJAu
jYvV4cjzANMgGUo2C8RCdGngQnf7CyctW14dncE7HHIVsPjhpmnuH0LLYpzXgCi/
TaqIg0moqkI+lA+RjVaVpSnMnyGYvuoMszm5XsJ4XOJDmwwvv5ftx0zi2l9iCK7p
L6HAnXEeSb0aGLB5JD2mwzJStN24A5zuzWHh4XtaRSvOo3dHmiD9QBIlGmjC2NAz
HIGgnpY3vV0v9zE2kKLP62+GxbcU8MQxqUzOkMAo2Lo3xZd3t1lzVDgOkBkbizIW
hOG6O+4x3caMu/qobZdG72GxtRW64HrPaCyFNGXMVJwf9tK04JrX20wvdkmx9gbK
q/EFhWmCsnWd7rbayupCR0uC4PwyaBeKiglUGvWZgs4mTaMwKToCNp61uSai3Ts4
l2b2Xm3tBdLY2uuQczJelSXXOUKTTnVmygi2YYE7lbdRM9n/U52Psvvp4m0Lp12G
n+r65BuUN6gMyeTCShjulEIbi5oP3lOxlmR4UmJJ7QYJxNztX4dqYAwWLmhJP81B
hGqifh4kZfGBQ5zQ5bemhivW4+mKRzkWnY2ovLv5dJyn4QsqQUj59fdTdvcqnqYy
5gL9oLygRR7CM5fHl5FGmh3XSAD70zDZLMnv1OjIbg8L1OMS+OK9ZVGHutV0FG+2
kRwz0JbTNn39FVMde/WUJ1BxIz+b61c6jh1KE0Lr/rRQpNZSiuUSEXozgmbrHdLZ
RDwUtj5Nl2U6xm246Vr/F46wsvWigQau/PzGFV8F27atqcgICCXTh+Qb3q08g7/z
6ilkpwh6ZX88S5SHtE0GOKz4MRdLqYY6wKk9WEzZNd15oEFRnhb7yxS/8NHmr5zU
zVoTOUqu4nJATqG9dzJLGyjWXBmIqS1wz8qwySo3yBT8oyF0kihjZNNOrMhFNLT9
TMBt8VaoYSyCf8AY3SdROdehUP+fyTEvna2PX3Ucju828C1H0qOBvct0BPEISdrw
404Uxgw9QQNbTg/CASH9p1dRSPLinsFDDcccFaosncH2h2BMnux+/4rJuDzT/2XQ
nN/5KNXsSs9m4pr4eEnxhZS5+JrwCqN2Uxx5TqcB4ifxFWObJabzl3DNquaC3klS
9SVyHGz/ySxQ8BiNPJ4ycv8RdS9mu2kaJ9kpCqC06h0NiBDTpzMBRmJtzH2rOydC
si+FfafGIDy3qHrRlWLeqdVJyQNMB+9DfP77QoDuXR5YdCJDM247rGnAEeMsEKGi
nmrSI8vZTkykwp80tD2o/hAldFn9o3udwgd+aFoMPaDJpkhL6lzpNrqIzQ2HDhHZ
b+8nZuksXFdeZsfKbkCNB1nS/zeLew/1NUlcGNTL0gHHu7V8XXsXfYNcCBHGrfUA
lnzFGCKd1jx1ax6xc0uCYcU5ku6IXFpOmyvmeUNhF5l5u9VClxkMJ7GLALW0VjUe
FzniqE5wWfO4q1b/p3rXD5YzD8IIAb9MwgJmht2CgAOivxISsnBVCUIIoVlr1gnp
8eKni+0SkGnZdWdTo6Js+myqiBMOesWMrGGrh2/AYLj5HyOUPgj2sQIDYl2Amw76
nV3pXntV0Q9gDQpp5tyN1jA9O7cTBRt0qEv2BGhpCKRAzub17qohzq+zmAH8L6ek
YxwgMi50dWmavisQlM6u6f4CFrAz1GedagIwW38bLNl7UzPrOW/3e/ooPjy1vpiB
aEmAA42ewjW6SWkCYTFJbUr/Mwb7JIsPn7Ly1Kmwh7/kHNklSoNvYtYIXmVkgBfd
jm7sGDgt2mhqiO9IFA4AQpW4NPawR3RlQ7CICOJ1c2ubBqNuaL7Pn5jaGTqCBXu4
EhLkypd/MybXGI6WY3seidU+X+YGz3s6vJb6Vone6z/5J02kQP1qb3lTwvuLV+nZ
B3gOup3ajhgG5hQ/d72jU2kou9NWlFU6CcwC18gQ5/11FYFdWmHGFv2aBRVDDliH
UjaOkBjpccRGV57X9UOidVxGZBdrrcjNIJ6hBCk8nS0dI6pCbfKvf95x5DT5mNfl
p8URpD13HEeQ+hHhasFyJTEDD7MxKcxShUBvhrVmm3kSaVUpnH78cj71yYN5oX3L
H4UBPH0O+yPb0zSufU9eCwHEpFMznRT6PH//eoJHuImyxDiVymHIlIXbMEvfWGyT
0QoAXyr4d7aGklIpfyzHuxaZln1uquXQKXje0AbhdlBiptIxy135vynRDltvNCXx
frrP8gNAQZssALlvrnCgHnAg4CgduolK53zhmDrj0/sRyMVw7G+FKl/76K+cokZ8
dNYI9vlpsCsXxUu++dFMZEL30pMZfsDF6qyCVHEdL9L3tkNd3P1iPeDLZs4eJk5w
ha2i/8r1F6O1Ux22rI3xtB9Ly3vGgM5g/9xMO+RpPppqJnl7FhM3znb5C0HGqnc1
kCQ4WK6p96kE5rJxK3iD9Y+3yN8jouQddpVL4lxahcEyBK/DOH8tYexkOg2hd1nR
GFKhEeWiYsVIOwxGUZuNQXvmdLr+wqkvhrdxKNenJ6vlWLNfsBbR7mFcxrgYweeX
3l9TCFryDQfTWNTbk7e4Cmzl4A/U5MZUplgHHJJby+RZirOPIuJJ2PGHB07K5+dy
sWuT8lKf/LLW9cK4cPfFrI276EATNQn74eRuYMj7eAV9PoH4mXC/GF0yHMM2IKtM
/72sLLRM8LzTJqZGUmMKF37QxfBA02fhD9uicvL86yfPg9vtWl63S1P6xB3vW/u3
2itsGzueprdr+VWEbwLGyrBt1DLerZ//o1D028yOEl6Nl8R7KGEGM76LzIyCZ2FE
Y5QemaDJbYm7ITfEK25MGkosQmaja7VYy7Jnv7SokUhAYJpFhPL6UkbcKvBXxQW2
eLBtDBE5uPF3SW+QTHVoEAU7E1tk5Lgmb/uZOyD+T5gqLIN0+N2vRKC4Lux18EAl
gozN/zIWDTGe2LMh1pJfDHA3AxQniBKUdgRKsSojieyb3C+CjoWj/YrTWYbIT1QI
+UyPVPMj4G6S+bK4GV/pyVPIp5pF8J/ZyK+VSni8ofkfsQhdEElNGZsc2nN9LjZG
Ez1dCfVJATZFl2ZEmCgygFT1k1fJUbxJHkXeaV7te381hAhZHBJ7gEEKmyiPArlO
q0ghUmhKtVtKVKL+/oJONeysKGv8J+XGk0Qiw0sw4gWHljUz3ubFxOikLIcfM7xp
FSuuoQZJLm06z8hATBhxVup1FZ13qLAqwhbIJG4hEiZC7tLEgpvxA8BECoUqwI/i
LV4eELsfZc9ifEd0Q1AJwhJYIxlbCU6UPVXMRr/apyR+FUklfWMl9X0MmAc/z3Ob
2j4Dv3fME59GT7d0v2n35jvHqnSuK1Z6vZw65s0+sOXhiBN8f1wu5Z75luY1yQYA
StpZvMgfEzrx49ePDEF6eQs6A/q1s5HAn+oYQmH9fx2ETB/WhLVrPJ3u4LhriW7T
Hz/MPx0IE69ZXG3lB7rbU8/ug9yvKZN//R/Wgu6XeXCdz83ufxoafCG03RhkAVuJ
tWHhP1S/zcb1A7KjIx8WJFAHdG+pyu/JHfIr4pl46xvIEyHi1jewOl8Qv8qn0jin
ApwOvDyf0Yuad9u9mZQosbIOJ4zHIdQJi13fEHVb4rsjVMdL8/dvSoJ2jO6twO+N
ZKDstoHIKpPQhWrCObYyxPsgIhW18ng0CXEgtIa4QiJYJPEAsixSdDPpXUHqHgNd
CVgI99Co4dCupl2bFIOIZtvVmQudc2qjU5CZ+DsyGcxudGSOhlS+3el1XLfEQ1ft
x0ClqSCp9/Xbc+qZYBgYAUWSlK80nZc97ivCbjr8raKH9fqQ7S6eHZSjI7SP/QVD
wrfQ4otn9ofeuL/2X+npzHUfgkZ7ExR3s8csV2B9g9IQ9BoRmlrDgtS70FEH9wkX
Ozuh4Lo1Cu4ALMqBljihhJauYpAvSu1Uiz+jHXuNAxlRIblj/dFSnus218tdshJy
hBfwkltcCHPFqN/5dp/EBHPuP+ggllOvW3oL9JHRZ7alt3MKwPBG2ooRBXoz/6IJ
uFBdYswSMtxfb4bwoqrErKwGOCskwLb5LnmK7cSvdkHc3olk8F3KzyuujvFbWNzY
7+8gruQbMizvkJJVve9aCQYT0ZRqozucbPb/SHz5Qr6y1qKk9YDpF0esuSuwfUFb
dL5TP9qFLxFivB0n20gMuU/B5OkK419OUqSh/9GMki1jEwpITkbeqCfRT80WWqer
LhX5/Q1WLs9GlFIvCWp/XSUwLubeVo2gk08XkwrdLh5qR/pcmYa4R01AcO8Vq5Qn
eMw6Kc7qAJjkLYonYXB1gp1jcYQ5crL7fGVTjm3Xl7o6MnYNDt+g0LYecw2RegSu
p4IyesiMxdjwSO26YijHFdJCHFByy85Sk2bLIZsZYeXR7mQBhUKvZRuj/ebx5Kdr
Wc9vAyFH7Nipu18yKKWtc8BFGf2N2uKAi7F/RdGS8rJBOUuDRJLXMjrNTgm9XyZo
AmL0mxnjy+CVvc7lR3VSV2BTif7OTdlJ0mnCbkJz6cnX7trqRW5H+4fUPJuGtWvr
2e+bNGiLmNXDmtwgOZONY/E+siuGrL5UejrkaaFY+yxUWXlk2h2RMqsPL9EbYBeU
pXbvuv9M7Gl6J7pa9gQne2hHFNsAVJw/z4zjPLvhZ/UWVCVi6gXPlO4L2NP96XaY
o9Fyq95qfXmqdRYk+NFZVs2nuvw1Hf08Nnd/nZNbGfgwncA5xvB+YxMkX1iXANeF
qkCR1yEI4fOcCNPz8nxee9iknjudxOR3fpclp9srMZxdTXE9DswKu/mbr13TUFuT
GVhsueBnTfO1xN9QbxpnKVnW1yBA+6pGSMOwhixgEVipkYTucuI1cKQwIqICGvN+
BdLOg2YopMhrdGSfFNrQ8kCSzLFtMA8kzfFMG28DNWg3uA1Di6AKj0WUM2nP9Omd
Iy7Nai8nywxpnvNt8Yh6rw93HLRgBftZwFQJ6OeDl/FYOad29qhMd3vZ6s8kiWJI
D5zviN0VIPC1A+feOOd9u1eoeSynnBUBAqxy6nzUlpu5dDqoMJX9T7FRIG6AY1RX
nV1qpBOysGrmnMNBLUl3bs3wN73m7QDTsnGAT3L4FRWXkcx/dcmpTZKgUlDstpCb
r1PTDX2D7655iZUJfn+XxF1EBNVxcHtYsVRK4S7skeNhKOXARG9pzvGRXtHCOcmY
pBe5cU1+NJeLGPl0LRqhmn6mR0BIckqTPzOmWUewV9M/1JSaG5c/oY06kySyGVoM
fBaYRnhbifkjuGWbnyPE10FGWm5nmrAvE6q6UmM9banCyHIX6lFMxcAd6p2RNYJO
md+qSsBIM44fx3FyLuGpNuui5JAly8KtQSIyhfni4P0oF7iByAQiZrVPEUY8EUq3
SCUjyE3r69ejJuWKRlkktI5vsDYxa9beUPlltOa5qDpW+eDOyz0M8tovwQN+ut6u
vrn2w6QuhytSRnZ6aQ0waiNqkrPM8Hp7A3fzFn0ESFcTQW4EasObnvOMNW6xO9/6
4q2m98xm96lGQuaYL9SvNOauD2fF1y5jXGubSC39jfZsomasc4zz1d7sls0GVCY9
upPDMKyOyn2PRQapS2kBqS6DQhzejkvYTHLIipRudCikfOEocI1SDSNQN+NLj4/C
EemAGfv3zdqyyEM6ZZPjxPX5QDQma8XbqgaLlcvmSvO/4tGQgxP5M3o1bLfBUWAS
7H6EL21hGyPzncFpYrSH2zTGE3Wmy4vlfg0K9MRB+621utVLVu1GxOf4VCVDBRsL
LjC4iX9hn0PKEGaYkx3vMO84azKUKNMAlml7v3OkTaOuZWHE2yyfFUBbn/Ej9FY3
NmbnhpM/rj7bdw6xukatwu6hFOKrjhYP0BmOn/PLdQdPQAui4imw1V/iXr2AncZG
ZqAPpp9KnDxmKeEIM8o3zelE4UCKUipUbBJgoWYWLg/xEeRD7b1Qp2BDX3UOjwEq
qIABChdXkvrORDzNEkejhfwUiB5x6omAwyU4lIRDm1Rg8ckr0/4ogNxDiY23LplU
5SBZU6LX9y+7ARQZMXUq7Aa/k4x0l80AtpgpGKeQKTZNBWZ/q6zJKnY+oPiFMi0j
HmH/nfF7yPUtgsAy+uNyCO0o5RSEPpaJwyUKBHDsA5uvqY9Z3l8kOvewCnYm/iCM
cMo7NwOZ1dG9iqo7mWVEocJT4JqzcK/PSlN9kzAlVKNC/GnHNgiXBNIxSOk1FuaI
VEP3O2gCoC55CP0g/1egBDAFyxtj0VIMN6Jr5eE7mA8ahVG/eMTpG6c5rgFYFfXT
05hFkJutoY9/ioz/ASiUk8EE3S3PXyzR9aKzcraJeLoemb252/DKFDB7igrql5qf
RLtJXOLQKdYP5L5Gz9IRvcvTrMGKJqcDyvXp1WDEuZ10i3RGgIHAJVPoOS1obhe+
Kt409chKwvY7E6NmRw3siEEUA6ssQ9tVgk0xT1/3dCxjRe8d+9axbsVwjCosKyKK
WuRnX9b+HX0bnI9jmi9TZVYwLKmdVZ8EgXn1ULRk7uGq3+RZSavbwbg6MdPu/Obt
YpVYSixDFYSOTg+8DYy07lSzYdoplwsXE+q718tzUAXxQNP6gT+pKFSUo591DCix
+Jt47ThTZzeISQG3bn7wkG5wvW2JKwvpT+oaYqbKRONgNwabOHVJ4D4xkCNOTD93
IBkmAa58spR4+8bi9aHJNyGwbxy5z1uwQETFgBoXQe3WGgcd7I8CGvvLddwIugyr
xTSg/LvPvd+l/fKl//fLAcjfQ4tRjMLuBmvZfr3ZdBDOxyPBVnuHxvoL6/Ye3un0
tZKmVtxW9imavYM87LA+e02jWqrbGiDsp0LIS2iy9ZIbGqnZ1MQL71BscyMsShdO
JMM+QdflquGX8W8ePKK4TZ3fjt6qmOJG8HwrRp8yVcIvLrjGu+vawmqetZMv5JgA
eQDotq++ToNZqcFZuiQFhNtnK5po7ooENd1IzBT70bK7SiXbQmo4T5WBcXLhtGKX
8hlV14IjoAfXCjE51UzJr8KA0JMqWVZKBYVzxTNM/DP4UvYcRCggUofGnRwTcBzF
DSlxzQl0z0aYV4FWOGaBuM8D6MmdBjN2c0FTnvK8p0SptfxIz2lXonJI08ByvFEA
mM7tm8vOxa8JfoloNG3InMQlw+fS3n21ipiPv8hP3gxsy0tuXzbMYA/Ua0zv6OtK
W+c00IAsLHhQWwWisTk3YVFPX/CqAZoYDcrS1iVCracejUNpVf0wlZ+gWXn4J2N/
Vh+ACUrOmp/xUcpTZhUCIb+tBzjHS0u2J/N/AZ4LjFlzTlfDzu0uiDPKtHJRhFuF
CqxIwJWiBUMTbgVCCiiekLdk39V7f8eTTJ3BtdU5kSmRrNMINSbJUwrtDfm0p0gI
AuJRpTW8fBdDm/MMG0blqQyoUv5DkWw8VhK6swHX3bbwxCTp9+lC/sQ+0ULMCfVG
I/bQ2h6sLemIJxnhpgPcdTBpMj+eMKvAeIaDuUdOq9eHu7kadEZOo6jQgydZC7nT
/aDWEwkVJy4biT6xsibCxgcR7jUsbjVj/4YbYUFQOy9fuyQNGhup5q+EQHx9xlZu
hhTCbNCnxT2huRClBvSQXb819xMwFphkw7byJOe+dlkHQVcFHs6WnXGibi5olCGD
zBdJoP7V/d2jqDEOiZC9mXB0UBMn32qiPnlx/nFR/MkBh6DiZv8szgmfKHaFCWYS
s8PJS6W4UIa1wz8bB2o7Y4itxMkteikutZkLJKFeCL3ne2cB19HJI9My2OYauFV9
a55DlHSgz9abIgLhH06bnvkH3Ej0YuunAaO59RX8kfdG+tQ8sht1oiK2aE0k1ZSS
BY92QfTDcRtqujf7NYleVcD4twQwu9UlLoh4tmG/iN+BvTzqrzPxY1r9IyXJWxyt
Ti+XTk3H/Wy9xoAqu2k5iSYgvR9jEuiwiFWe2QKRtAZM2tDnORkOaP3S6ysp3Yoc
u9RDevYM8bRJOJiucWYAtkDTGPbp14KdqGiVOYRMQ6WKDMulwJgigb3yI6BFWP4a
ovxO/piuG1WON2afR2zsXmAbGSPHdmg8maRGHJJcUop04GnTV/aBYwNUtGfusHuD
ZqrGBjaj/e3NHfOu+A3ujsVzKjRH648T1Qt+YTz8syb8SGDqZsvN9D4El4D8vPpp
1AvPMrNPZ0GyJnErKPZ+m/fQ2oi/UL3p7DvIS0wslTNUJEmrn1ZXTPsjdLpghiGa
tXUtpASoHSgwAO4XHCncHhpWVe5kwZvTa18Etfdfu78gzZE0UnfvEvD4UMM3ls6s
u2+6YMvYSOi1JzDblFqbil8s+banj+13beK2wZspVJff9/4vIgMGkIyMMZzIEGQm
OJ0KunusRoZu6fX7D3IklHccEyO2kyAZ25hNuEZ+VoFElQ7490ZBn5NUeEe7e24F
BvpM92xRSojdHIMHzaJKnHWzkayHh2wwMRhFCn4ITAnT1Wkn3D/ZWX1limuWGZRK
QTsmW+gSPmZfqaFk87HcS7zUK2lARwQ5QcyjT7DHRIjA0MDe8xiZ1c/YjYK8NbhR
yUMiuoBE6HNOIBqK3RwJ6X3wM3FDdutK7Yy/uE5ABuV74kxH8RVHPQN8Dd3EHoSk
1NGzzv1eCb+w7lrhWacqAz7KCWCGA7/qgAIfmEbJZshYpPBsTRxetpb2cxf4sGsv
Pc+g8YgYgqPAjZkav3l1qmku4Ew6Qq8PW6fNeN4bRUgaVokXDcHY8gH5iOpO0JHk
nC+bPsRvFOFpMSVzsycZUhYIn+iDR3YZ1SAWX76eypSes+GDzqpczqK28VC0IMM7
dKasua+t60si2gczEc6I0vfFc8SH48NrnAme9X7NumnzzTV3Q3d5uPBvXc6Z6JKU
rEM+1XW5t6tknmHvbGcaQF1adeOgHajXMeX7BgO9lmqbZ6+TFW/5/5j8djbIOegZ
fpo8y8bUR3Ma15QLulA7vBGYd8bx0FlZ813Oqi6esWelsdQ9oooiMlht9qOJUgo7
cS+I2aJjBn/ScNW6q2v4QAIlvJGeIdk5MNYNQCu7xeS6yPOWu4+gebggSdHd75DF
YrW+1wb8vBuhZL3tDPqVE2BXS5TKRj+eGkfLAW3BEtz1nj6ayOk5k36lEeOA/VUx
6RA/eIZ+PuqgdIg7Y0ll8xhs6mVPD3fi/cXr7Z3Lj7rjAbyK38M0NfoD0jrYfyVN
bNTiwPg2QixOliqYuG1q+Pj6mOrh1XqnDjPKlql8VcrddmcndL8DA2tTOoi3Arnc
fqg5QkjFob0nShflqJsbVxkoMXOLhH2gnFljf4ZOcuBohkI+HyOEmZ9/xMnobtC2
25TCTrlEpwA+J+ugGnrXBicfRESzuTDxl9N03PZi68tRlHvdXbD+896YZ3CzlZOi
rt7/o0W+e/TfYQ3cjZYefYFZ0a+QbJwxuzonqrILvjT/1gSviRON9Fw6/g0WIaKg
PuDab0Ak1YAs9fONFsNS0k4IgL8ArbKej0eh8ca++zUcWPM49HFA/S53n0bYbQyM
/L9TxWGT8/uc09Rlo0FlHNgpf00h1Atv/xJMsxy9zOnA0lr0J65tVRQa0y/MWodL
iR3GwSg5r78/t6IgEolxF1GlMwrbqcQoTt5QXHdIKxhglaAefNxN+xxlepbPeRu9
+p7Oraozl1dJfkMBKuiaNwofq94lmyTYq6o6q/mbX15ly19bn8GsXltVBMpWUxGb
H/YactHQtkVlNU4fjalYJpRC8Gr7BORYx0id6cbp4mkMOxqHgT9fhZeGUW/hMsmQ
BLNyXc+bfYIFsz6VLLa5nrCtgAgS4lsr/0C2j3IC9M5K5yIDDQmbSZnlfeTAaN2l
zmVTEciO5S+oBrAsMeFDDTXLDlzajJKgZqTMx5Mcm9vBnQ9MV9dCndydfUR/SqIy
vz6PE0LKkAgwqfykq9mR2yBmTiSU80hxW/r4o2Mi6Hb47crblv0AoTZuOPT0O6Aa
27vx4KvkbWb9GQXehjWVZNXI8fnLLmTNudbjknDco5L/a/FnT3/v4msbddHVVlBx
NQs/xloRCm4kexXVys6g24iSpw6CMGauTsmOJLPdSHbn2idx5StGhEeZNdM444K5
KEmyfE9kEcl5Rn0pJewR345dPr5ndVmYND5Iq/n1lRYrqmINB3sjrwYiLjGK2HWo
u7D1cB5MhvZFt6z6pQD0yBivPDOPk90+rGMr4j4cOZqZmJXhPMXf7W1Lse4sYMZK
TR7g5932feNFYhmrov6AR+/tEBxYSOM5JlfKuhKBrt2JdXTiJ4aOlBNtyEf0XU8+
Qybu9dhhG2p+L6yQmPBiIkOKNtWi7N/NnMxjgTWWVNkBO7WcAuocntcUYcOHOCJi
uk9kqj3dY5mBlEB6yiDk7d0bCbUK93ksNelwfprB02mhTtbooEdyWZ/SU0/zaUqz
uq6rPw90hIlkgMOHR/D4DRELIb1uMf5+4lF60l4e63DT4XeAQskls2AfwWl1noqI
lVGcUnh+tqkiO4p/cP5EvyzckctvtSyZFjBhcU86iH9I5gqBQBC6JoF+xD22q/KA
w0wXC5tcB2JZG4GA0QbAi4zA7RKoB0OwNGOLcs4hjtzEv/2wajJz+JgQIVJxtncy
/9OY1ojxVLMz9IfrZzY5EqBehTKFT03JPMtlPLFqw3syzi1JkvR/YypDj/NzkdZb
NI4Rok6xRS8A3RsLEuWrrUAI6dkJlwejjVUBbaa0QRJW1L99QYe1JRnsdYKWch2B
sFqKrNopvl4m3+qwYxs5qVvTDNwJOxgBzNx/2gs8t4QTPkNp4dN5wgKWQx3nudom
rm82+OD4nKKroaacm4EWNjAv4LtdN/mBUJUcl4w0/IabcSyXe40fx6K5ucE0fVE6
MX5tF6+TcvXI8qtXCYC8+8kzCIsL/bBLk8leQpWfKKtwE+TJF07b2hvCVMsi3SBA
Y9qnlwR00Rr8xwTiJgEWVz6/HzokjdRZmWiClyxW5TrS+Zot3xpJrhOLqFQBjxeW
S3RFPV2maRtxHwYnylTwRME0u6gt6puWu8SkwFV8GZS6kecx3jXK3J18DPINRD4k
ApDuRa8bxK+JH7UD0uL5KPSdI3zv9VuO9kK8NS/rqvBBk4RQnDv7/wKNW/2KrIjt
AKuNH4nAfxNEyNjg9yBX9FC/31Yztlz1fLZ+tDW7aAOQ3UPXjJKoBtC/rTq9Y8qD
GDifjQBDzQWmfchUquO76tgELpx0J4JwiRAob/YN5VHFRNmbuS6bUm1oHI2TcE5I
Xjk2wNay0hF9vmWeFjdSSZxNJbvLenTpjCU5wGlYM/FAjBGfxKD4oEhQFUEgGg6G
dghJ6Vpa9nS790yzrrSFaGZYiLsLlMP8ne9ouUGhZZARIeAdoXd9eLbS9N5Pk1ah
eiBWbUp06kMyG1OyjpFY32dcLKMOMLBE8xU7BQsiSTZ/4I4DMUSz1je5DWagQpEG
h3E1b/S+kk8bxhgyhP/NM1vemnpy4Em8thzTstE6nnZrRFtekcWZ34F+4aL082bo
trGw9MXm3kIRUpbiqydqTnfGzRxP6UxzyNZR1A/5LzKhdbSL+I1swHOi7RzUE/BN
ZwEs8fx8j6gEVXcAvPTOZf0NE6VJhVrtaHYLAvGN5EEvVu+0XYxv04gC17c/u4Lz
RXJ6c2y6Du0yVcS8Ce6c8RxOEfI17Jz5WaIrmQ4hAb2YvYfsFYS7yRU2wRc2QBag
GZEjaRNOT0L54lCwhe4e9qLPEXFW6uBD8uikCZ2NTIZAMJiaILBNPN/aPLOS0yug
MOLZTyILPR4/b97MVSRm+Q1WeIeQoOtyB8vJ1koNPh9d7+t0Iuzq9DwEjfAGP9wp
TmqzPGiYqBPHZ4XuEMXS1xxmCaLdi1uGrvd8GMqWlpAsHMKFncKDa3/c8R5QlLVy
dOoUPdPhVH50BTUp91AF6TDGUqquHw3CeTwxd4qPiTWQYixn7d7OJaf7KkUss/Sc
3wSyjaDb8iGeJLvwaPC44quv7PPobpXl6bbgs2cAmlPWfH4AHBGB7pC2K/QkbKc6
QLGv1f8zGbtXCb7M7rP47Ef0N8FXgOFARSbbMzD4RzP++IrUVJXrmZIOkJjs+y0p
L0JraxWUDWu/lOm8FOKXO7IXskNto7JyEtT90tFZvHjYlYVXT/PIGzk5J0qiSwwl
AlPrUW/pK3gaeKyvC7GI2gGiVbbGSmjZpZ65B/pSxwrSUu1wyplxeMbi9bYN5OAS
JUbUKDYgauY8A2T/2lU0nSzQ35wvnRGFGtP0gg0CcvIs6PZIEUgcsEdfJgjAHu0Q
iEw0unWCcrQU+6Wyma/fzMo5zYXgmSoASkm18lDsMG7qAUT4TmXBb2OcJESmUgUT
s8vX9CCROA4LcAdD6ZxXTd33t9et7qvBXIHXC2LhoGcE3GBP4kLuwTCmWxStIHfy
ab9mcst9YzDOla/SJQqa+IXcQzPOlERlGkcmbsFMO1y+jTu5+f2/mN7vKAAx1IX8
GmuGHtUMC9+pNjubwmlYW8eASALT3D4MAtviUl4qhvIc9o1eetVo61z8FKb8A/GL
lMfulgE68AYaOHgoGAI9u7xPdBfO00UeRd2o67Hppo7mm+RGEA4QDcSN8aBjvD0r
rhBXDQ8aZkzQ9PdPKBIvZv4hEqrrIe8Ij+HSYx9KlPjeCmttrTxtNWmNnLHdrpiG
BL7f6uBFSzvwtekvZWoNpxociEPLIGinzhJiAz0iMYJzWEOUZFuWBtwb5MoS+rOD
iBIokci4wrAJPCJGA3cwwiuIhABLA7gAniFL0jyjYwhXLJqYP+FZJ9X6hwTRUn+j
A4PhErNR63bnzwK/JR1CeUae4X1NJu5hY57Ri2gZrFjM+ZhIxqAW8d5Kz/L/n0/u
IjoSQnSSItIvg72ZUqshyN+XB3vyBnaJif6V/DuvRdXRxbqH3X5p5sG0l4zg1KcL
dxeM4dHTHMXSul/WvZwmgKgSD5oiaP4tZoAcld6JmJ04vSBg38+MUFkaQtB7HVMk
kAQOcfFi6FTH/rOhvKf6x8rq1AdXxhNLW6psXiqC9i8i4Qe/jUNbIXvU85QDgRYD
Dy0tUkS6MKt9TYeKM8R0oUSpbgcniOgNGHZO8F4s72UtkM+XSJJkP95a9IeWGBgG
UKpzQ3+j+kL631v1dHYLZ0vI8ccAUZm0lm/MAXv2mFydbAONypI6tIpmVz3522Ul
poKcGDPbo2/D3Ddm8kTKzR6//tG7s1+8yVheL5zNcItVu/l9q2lp5fjz/Iq4EdRm
oXxhGRmbBuVz28i8lrFD6ACsH4zsXuZZrclPIfDwxOUWOOV9NsohxvRP8rIC2ASg
Y+0w9B0GTAyHOBX/s3QMDAICSdnyZ83eNHye1bxANoQdS7J/OZx6RPUAcntZi24c
Vrz2Ss3SCDMTGtnrAULfoapJtDX5IkUWGqjeGT1WtzD89AV4A8om4GkKNso90yFR
I8NcwSlpMRgvdIfEvlPJ6LBPS8ZB6mZtoqR+f9ObCQyrN4pNsyBJgtklpaBri2ty
M1Z+BZOEYRcHupdMWQNguILXohpGTkjcnSHmCz0vYTBP3wtB0R5JxzrcC1PMzCUG
q5Lphsu3sskhKYB9DbBusonHjv5z1uMIi1Cu7KvYDqjLQwO1CB+HX29LLFkmaXcL
F5CaD7ItQDo1iJ6sC8YsXEz3lCMRuDlH8YemJn6dIKBxKlj8Rpr+YCgPuad66IwB
H7NdbuuIwqreT6nJU/a/yO1XOChBpQVUoo1RBHwRmpgDnVgC/T+qqt7X8o0+MYv3
WN4JBU7Lij8xHGc9471zSQLMRjOp4BQi1nmU4eiMm5h87jnGnSeOjTY7DLbq5764
dfVIpJrMr1vj/o4TqYiB6bs21T5yI+O4bGrz3m4xcQ30atxqweN7kxJ1btuhaekR
Ras6rCgVtZA6L0l33geUygxk35cA0nvNVXUCA5DrMbD1WK5nM7M0TYVE6bj0Nej0
9wiLKC0PQ4NNfvy3Meizo/crK3SkQ3T0OmV4hJ2hWkBnYeM0/VpdidFEt3p7WgTU
ZcLnAbQNp1b/zQK4WRwcQVwlKsj6NFVvb9ivJCvQQl+xkXZVReL0SS3uOJ7ZSWCH
JQZnaxPBTxuwSCZs86it9kjjmI95fcPwrELDBUaL5DF8g7RM/4PstUSJjesgbWxF
yJ9RUMljlzT36LFIjkecAE4SjRqdpqMjhDRPrz/rUxfAn3Qu/1bBLIL+vsEjsQ1G
klm6P+NQe+yd5Qw3DV7lYyoMKmhRsDOLvhZhnyF6ejpzSyOenAPiGuj3UEyxJsgs
g9bAXH24kW3ITYsZYDeYzAGadKBHyCQh7Waq80FG/WfLPbXYKz/WURkfOMUDSdrV
mDEhfqcfhGjnpXi6Xw+0As0ISYzf3iaPwDotLhk4aYQGNml4PKgXwZJ9u9FQ0xT+
FlOzEGXv2jwkvJZ29s2tGjbLf2L9flFjCLNx26hEkP/V2pMPVSaImbUBzhEyEeG5
aUUMj/IVEKBUm8P4ooPGP0pouG4ye26HVhXeX0+VvH4gtJUWPN+SF0dXz0qV2/BQ
eyikSuFPAikpZnfP29g9di90dDX0wzjIu5/xS7De90u3ifeJ6w8ylRIWXPY9Qoms
v8E01z8U0fDFkA9PND5BzbU4B9CnTGGr95oovZhSzEYRXpuvs01mEJklc/4W6cEi
IjZXvQXs4/Sp6HqfcgG1FlxIK5OMyHJEwedlzUBDii5AxSSEFdXWTW7K2lNTD8Ck
yoDMSvXHuo5X847DMKnyxfUmSoNDxVwl7EsCCUQivYWA/4o4ncGMmPpJNE5hOeVV
3bj6P3q8QAxV05Ez66u3Qqahrhd3b8NodAeCiFD9tRZnSIoaeVGYXLINOoeM5oYg
YNNHZqO7kmDLeekUKBML1TyLhD2Ic950F79yXADjyIiVFjKyrflk9eUMMq7pKzY/
XdaL97/x/v5PjP5LaMYZCZqf1kg9owhcR5RbSFmQ6O6c+/TlKnAkl6FkrpOg+AYY
QZS88DRJEGcM76TBxDZ/6RwYTvLmADD9ics8W4lA4pTychTk99w1iA4dh/LkNdjt
JZJLFcccISVS1jHDaXdSORuVEV3MDeu37T7ElUr+aljMCAUlGi5PJgS+xz5wc1kt
XwRGLfaRWn5QrjxIDMEblecaMT4G1cptBEP3W89bllpVIoLTiiv4MHEpXgTOpEET
QUcRXT/pMT0hdsODINXW6Y3BGNv2lKpoUSltrdQ9M/W8+YFWtSyVXBGV9bTD0DS4
TkMoaz/wxL/9LNwlhKKFZz8Yb2iYJODSAfl7dBPPsSov4gO3M9oTbtZjDEYwuObb
yKvfCojxOeM404NHSP+Vv5GOz9KxA1fDFa0cObFOWKlOfQKdQKsem9FgF0OkxvkX
p8ocbw99/Ss2zjpuD9Psu8GV1/5lwHedqCLWA8UaDA2zA8Zfk6JV3s4DD2qzHg2A
xsKx8nHqSPwz+fwx5ysn1jKR87FdMppj9jnTkWlLiLui7vE8j0TZNU8AcDyJJsVJ
ss3DtAOIKVSDzXf7lH2S+cwBIOfGjn25iaN7n5XCmHGJ4KyRnHl4dg2ISddG6co0
QCSYeWXbK/KveVmlm3CQG5ilMlZxdlwpa96/YzlT1C3udCt/ywQFWOagNFfBHSzS
gq3HF0y6Drif9fMCtWk43WLPmUm79HVNebvoxBioDP5ngYJH/awME2VUrOeSrvIL
jZbtW5K4pAjerh9AmwTqtKlPcARqlOS4geOrL5Chp8z0byTpOc1oW4eXJCPzA7kx
Ip7C9a/MsV0tTo2T/V6aZWyfQHr5aYAbm4pxXvwRsacUF9kNAc2rmsPZd7npIGwx
hetIaQtB2clAiwmeZpy46QPlQofTSkv4HAF/zNz5miBFmG2Mhvk7Ny69QPcjy2fI
G94VZg8jSOL4exwOJNpufLxh1/lBKT8bGTvpSeCDRbvUQvSb0pmnqzTjcbx52wIa
EWTwrQhDiNjF5HVyaa/11EtqsqxGHxi2BahsAgvGtYDcowVivu19tB3VGpQqHAiF
jqdLLAia6pckYJ/ul1gDMN9KeaMI6IgB34j0ZPaiDtUP2Xlcr3aIpGR2M5Td7h/B
vjto14XZkoTRBqis3Pk0O2G6t29Cag6K8A+uMmOR8wYl6v+3np6twsorokEgxeM4
mDwfiXZZukX2AOmYQBp/5dOArmle5eSZqde1K7kkwoNOOM3lZW4nZ7IZarGBO8Ss
8m6wW0errTDb2QnZa5pBrjMwZRJsLYtoyaywuW7lqYI9iiGLazcaGHaEv3I2eEQI
g482ADuk9KbnwosW8cjF7MCfFSBjf1nr0c48aS/AII/7Sp8uOgdcqRxulX0ajfKP
idNmu1Lm7TKXhtUo8B8tV889yl1WM5STT2zvHtqk3uyIKVlw0Kbz5ZQBGqUIr6zY
UvB1h46HeGXMZRqTWp7mOgKkKaBx1q9Rj3SayQdxkcNero5TEF+yq7OvBzhFq4Np
4smOuJYMqL2FaBOzmWI3UvG1jsoHY5CS0snfe4A+a4i7rgvMoU+OLPkVxmY6kTod
OG5b4O9UHKBCVhq1G937hh4njHGLR0Q+TkY255td36uMFdD2G0Q8hg6HegNa+g3q
fyUmpp64WnlS7cIQEzNvBL6CD7kvRDe2dT0+uk4XYxPD/zHrIc/yuvplbmBnosXR
zU6ArFRHLKv85MDhQTxhvdFnWux/k/r63tT0z/gtnvf7pOwAhuC2IF58aG4EH9D1
7j5nbvZIpmajjeX5Ba0EBAzZK/sDwyca1Kfsc2b1LWQOE1l6yZVhRaLVv+F0rL5G
f48N/u1kw9uo/2AtDweGL8dDNUDB6eo1AhalcGE+Aa4ROyEYQu/E8xkLVaR3dV8j
vi3VgUZDy0J+ug14i4uhFs1O+GIsM6eZ+Q6Gt8np7Kckb9KXZSDZEgvMKPt68Myx
jWZgKKbENu4jrEMzCkHo6pZRs5BjcTZNKPeI+DGseFjHiYus/pdXFq8fRIRO/7iq
gbD8g4GWUSVdvgm+N8iTK8emwtQWfZwQO8KnYgBqkf9EaCvJZQINi9phZz4IGuCH
HlF0toORRanVpAQ+o41LGXSQzhcgbgCvjxRMRhBgty0/hUyh0Audkb5JsI4EqkKY
hnvRqSlV9IlLpj5NYZq/RMHBcpJHaau/NMMYuVPvj1iIgFJ84OinmG4L9Z4bXptO
cSD7DWj6BWTQ3zRniorhUGACT7E5agUCmeBpAL8YW2w7oxkv0CAVzteStHo1LSfu
3OqAKHhiUyVowUHlMW/2rIil6/Y8dhiZilK7SPWetT5O/sc4MZCDJFYOlISRWsUk
U2g2OLkm3jkdfXZT/p5wN/kFnc72biTripnnkyWMSK6cJwW2n93Auy/L9j5JDzmh
rDlFm3zfILbupNSoWNjjbJPEXcXKJejhdTFgJcTnxeescwuMH/kh5RzKFs+O1w7N
aGER83lE8g7JygnfKI74jsmLVnOGR3Ux0lApZB2G4PLYZHxhRFAtQy28tfWl8PSs
HHqwK5ByoZd8FQOWgMYtMIO3abCCe0cCqNszQF3fFWRzermV0B7EwuHQfUyxUDZF
QKP1eKAtL6xsHai9kipHHanSf/YkyglrD2aXn4GaCTcom6e7bs4iRn5g1cT/rpQi
q63IznFrVtnMwFCvW400PCYTAlp9VtyxaKm+Buf5lDiw/rdL2WnqpWo3r2lV7hID
/Fl4vJZWqcSw3k7/WfyntkvzXGyDJB6CVCStn+Za4ZmgV3D+zV1ofqNuyoH263u5
j9POtYiFNF4U3tPyenQf/3+S3EvB6gZ783soMNAnEq/Qa8xZoHaf4Xaw4F+lL1fz
1soPmN67/PBEQVuXHJDGhwRZBL3v8qgcJ+KLr5XSUqqCULfv1DiBr6BantCTi1eA
ztb1IAVsWIyQWSH6EDH5BspKjvJIYgMNHKbYvm/Ej2e9Dl/kAW0DGtYNHZ0IxaPW
cSWK1HpmSI/2aoNpnV/LF7H66Q9tiLCXIOQFnBcsvKEfjgp4az7MJO5qlelqR9Yl
Dq0HD/DKLdX70OML1FWLqGInEqIncUJufoaekfewYZ6ctYbq4HLTrQ8oUrNrLv9r
VIFBJ6r3J67uuEd2KjCk+kzZSrEtEHPXIttrShZZVZ+KzjdNVYQF4Dd8Cthc/kLO
O7ryQAR+ikeFPPBI34LB4lDHmYfd5rHRHg9+r8u2EXAyjTDSD0Z2SERl/hEAAkbF
cohpB/rhkSWrj/BVwtP0NGWumT3NjKRuF7teHbX02bfojXV8fy8VlxOwkGsXEmyN
dayBABREGbcA/WidUjAj1fN/H+XcbaHl9AxkFJ9m4J3mJ5qE0beptLTY4R7BButj
4w7Esc/tGZIda3bqCVmu/MvbhPsK9DvI/bhJvLwo5RVVvWZ8u/JFku4O1X5ir1aO
ycTAWJOM4ZeBpalH+Digs8yNEIysPKMHzPc/xNxNuxVwHBo2nmxjvMY6MDl9F00t
UtT9e9TUO1ddx1pLv3RUkxOTPVn2ceLHPBlgj2cDCS87Uh6dgcvXhoN8PhNm2jxV
c0B17C9EO92G22+UZcGvo2vNcu5kLhjQTN4JGbstTMmMY5toiViOdaMcL8zwn8bX
7NzSPHSsMIuT7zhIL4uSXDtWh8Rzstexj3hPWeZL3OqCRBXJR7KjhxZwUXtZLqOS
t+UEWbRHzMiez4SykD2/7qbxfETg37FdU/jf8fnr6UADjNY7aLnptb/l1VTWmi+I
6SPCbccyhT7OAaDpICg2QekCBjx43dlq42Xuaa36MkmFwBfMJmo+G1B+chKObhS1
V9LAuxFOWUtyV9GkRULhrgJ4Ord4YtypjTGO7Rei2CVy9wn1Nk5hqjIR/R8piY4+
u8L065VSXFQohQ5+2AONDV/NIUFkpL+/h8IPxuPVoBlcdKmcWVDXi6VE0j5GTmhu
ZY3eej/k0XZf/tIjO4x+JATv+/H/Eq9cir71mALcjCBOD1bIcwe65O9MFBsJHjKC
xwddBGThOZkakss+QKNIsu2hs/AAX+kbxqFwv7D86yev5J9gtSv8udGYGeA70E4g
5GPoqkOcZF9+WMijkGHJA36Z10yxnCVbTOTX7xUrumoT8YFpGpfEwp4CylmF4XAW
PR7arzbGuBTovUxu8+yWJDif7J7k3oCYpsvqSURxIp9GuTNIYgep7wOkJ2Bhda46
B58B4Pqmth8orlbmpX6MW3zA6MCjUbC6MPtiw9LU3CvomaUzGj4jITzU2NGLXzrQ
FviZ6c+5ROkf9MjdAP/8TwJ2Y5JOo073Wp0dPn6Q3js+T8GuC6zrH0SrcCVPombp
ZNcS/biCdBA0MopP7M0gN13yVCjiTipRVrKoiNjUwBSN7tzu5+PN2nKvljf/Yg01
LGJ3MiZWfxmtt6T0hvYT6wLzDEt9WEctYinrFBglDaSjPI+VDjCnhyT2zENIRxMr
op867dboWNQP99PTFsyXtegKUp/KpHxqsCiB4sjgkZYl1arX1Y9ymxVVXT0vnWXU
R2dcUOPaA+N/rluMjLC/GToieoQPwk90qzUrCbX7+P7s5IcohAmiB974M0aAwtKj
PNakr/z15xz2yB7j0R8wvzs1fg7enmgB++YK/Xo8zOju9TwCXp+AK3ILNJYyBKoY
LLeIIRN9qf0XpzDUNu530yTFci3cbNXJ7jQfu2wB/faZhbpaXvXQjbtNUvrjqZ89
pn1r6AGeKLijCv0R1B6v8eBVl+AppF07/LMAnxOp6/yq9hwtVNBPrMb12wghIEFW
j1fbGzRaanYHyvYcCqdPQe2L5XD7RcFQxAJTT/SYE+eQDSWz0M+zym0eZuoHf7ca
sHhzXOcK3HDYuqQhVaX7mxHrpaNwkq26x67g7k/2fQOJ7iegkx+tmtHL/HHxqt21
7i3Sb308VeSUaUx2NFOE1t2U/u0wFDS/H53fpKxJ93W8kjkyLVB3oOpIP2/L9K2K
43MMrcnNMB+MpHIekIn+YdPgK85opPbgYOJMYsrcHEuJSMKuGh0i2s39QIQEz6MN
DHEKqwfXCgpJGf/59Qq6ZE/29d9oQTDHXwWc8PqO8vv3ryDBH/39LXTmb1JkfWBZ
Ln6cqWLD+wy1CydZy52PMql47gvnRpJYNk5EhL0i5SV2+72blK8nrwgapLb5cSk4
r9gzisX/colSM7BQQ12PURjAA0cDIpL/HVfOwGuNpwaWEsoIQ+lAG/QE+Mk6bIdJ
oX10fS1Hp9B8Ys8UBspIeeguYEyYlSg+C6wY0qco6CYbUkDutucIzeQwMvIX91zE
561Bx6zhccmcUma0Q0XYBmBG7bKpA1FQHHdZ1tS5qP9TANWE6xhPCnI+or51kFx6
Dfas+OLAfBewDGdQirbGqqHIrt8yxSPhBwxEtex7s/jcyGN/edqDzW01Rv51QpxY
cNM4A9zcdbm6YgC4X87ynaZwJxY5W/59knJ8JGKnBJ2t1jRyvjjxg57CP3Lkqi3M
wGeLZHjHrfbvcHXX5O/rKlZpsRIpJc5icLwSrX+43uoQM2gF15MBhEbfSSpcWbT2
LNGPIoxJZz1zkNYLoktNDMgsIWgO1op0Igvz8zZ9hlPjEhyqcjodboIpVD3FdUzv
zx0HYldbtDiLqYhWEAanQU20lWVXTfShMtahbLgRvANvipuDx7a17HfHndnsuZjM
DfB7RC1KpREN8zUBdaJCWOUNoUDT09p/UaWDlSEQN29DUbLqRyZRCis4sxf1Unzc
/k8it7unkojHTJCyYO+5IC4ws2NQ7YWokSlRTJs/N5mJIyUu3QVQc0j4XLjbYdCL
oSFVJ8f3z/rhtzyW+UN7SmTc8wcWiH+vfYl9EEjHIOG+mjyFGawbJQWL8rV7STnS
NVv0dSkJWq8VPEfkyVXUaAFPsx7TyTBT2HiPmGq4U+ALXbraE7CVW8sbx5+6ycHx
rfz4iQeJ1nm7d3uheEK5dTgPSkX0vltb9Md/aaK7XNcLtvxDSX8gz5Xn/GD0uE40
STHNSd4GtgP9vB/REjyArrytPmiaqPRur2c2wW+0Bn2oAEFi0YR7q0PxUuIRMl0Q
PLyOJpADT4VTmKgIsMm1sieu/TS1N8d4epGh9aqzlZN1rbuQbiwPVFcIhSw/kuLh
nJsLxPLt5vfIDsz9GW0DjKfYSc2s7pXadNJ4g2ydyfyqv0MW2pDdrJwf4NJotDc8
dVmM3hM/SjzYtJfD4sk/vppVhm4kvaKZMA3Y9H0CVMmxb0MRRT84Mf8YMxS4NJuQ
cieJfYz7tyBpeGItBhunbJ037bSws43RQH3DS2UGT8iyTrb5cVYmmZuITOv3bJ4V
BhNXCuWPVFNi7r9gW6YDaQre/l6DGcOfUYdSEMDnqdj/7hlkGroS3hhwLgr1SxVj
l2vszHrEKxS4M6kOUM6xbudp90adYvDsMl+Aq3Ofjn4j91T0FTIW0PFBBnufKpzV
Mb/W5uOpNT8MD+4LqnZLbfIrN/rYrY/MT8/8CrYeDIHaNmlCNhvRMPo3b5tOSqDU
JEepMbjSQM9nJphtXkpIqzspDkLGnrIHvSSAcOXQukBVrvdh6fz7SYl0uow89qeT
5t1KopbXkwsVgYZZlAl5ZWJ3JRd7jONoT/dtJ6l66hCmXpvCGURtXO9Y8mt8XBVX
Dga7X+iU9DW+49YB22e7H5MYfs62oAuC3g3WdyLWxLQ8AwrXFwUNtPB4DJkPz3MQ
qey46I3+rXzftkRABev2ogvCpHXyoqWmuaLki8YujLl759mqk2Hax7/oMx5nyz6Z
YJKtvjMethfKgYvy3rFnlLsfUpWSVFvifQQsf0OZHGXlByVoUg0m8/PY7jxTe86o
lvfgd5ZFcM0pVlVfbuZl3OO2evy3dbRIqdMDVVTmEcaIVxByR3LOdkBzgv5CoXod
I+lH+hbRI9NEqULtZW+TPKWQSDmcycknxgQ8QVdC7JSDIkgYbDkz2aWUIX+9uvbi
iOZ/Kotoct4GpAC38tjxaWBMeBxZXSzuCrSub38K0KTbQRxx/x0hIPzjIK7AeHXf
I2/7Jt8AoA9TPcQRD49vrzQZRrKNDhxiltY9wkJQCzc0lek/UKK6JN+Cs0x/pabk
fvhI99gB89o4bY5c+byBQUwe9A4cTcGl6H6zTEW2UyyNydqMRhCsHqj92WKKVZOz
2UGBD/Gbg9quqU6pNsflym+pKIWVx6QXki3QhErRmHg4mCR6eetREWiHNoAqve+z
DxsIPY/OL9jfXcgCLFRfMSvEmoqfezHAS8mtKSBa2ibDwfeYbLWcJzqVhLrqH64x
AQs27RBjOpEijJhmnMcfo0dI79oys6c9Nm0WNILGwdkbsPFEjF7sy8R76jyDGiFt
PQP35Rnnq9iH/4wMmdsZPkLYlEQVUOaNUQavKht55ab1155xs0/DOmNCjvwq2Re4
`protect end_protected