`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
ddtXksX2+yylW5zu6QL2Lhnb2d1sD00763mmSITNX595NcHTEkwn0zB1Dry37fOW
FufOhVzEJp80NC5qZ/+F0Vk7Ik02dIR0elf3clrjeJRK85K4e3Hoo4xn7YbFUIms
l/8VZSb14+JVGURjfswrIyCUotIzlzVYZ6gzoZwDXIi5gQIBf/gI+KxNXPaKV+PQ
Ufys/12rjO6aI/pPlqSm0hCvftmBcnezN2hk1UeXgOIuKZnogjOsf0iJVX2aOOWE
6pD/psybjbnsNB6kH5uFTA5frkzIzkzl5d9+YDm9OyC+k84E83I/7/j+rk4L2dah
QJOvksSIzN867/4Qt8qYTQ==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="MvBXkzurAa5VTw+1JJ70nePUfoQXBvZOku/SMmg4TwQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
oRtzZL4VJ4iwysPsC8SXYCzXS8Fw2gtZTOskLcDV+1B9Nzn1zTyNtlo6lNICRmmK
ZRVu2BmCc2G+fmzynYlNTnSa7C0Cuel6FYpxCBlOuk3OF2tzAmLAuDyOH3Z1Yjzk
a0aHuoCdIRKv7BrZCdALt03JeUmXKPdOmIlkVGFl8yw=
`protect rights_digest_method = "sha256"
`protect end_toolblock="Jn9CQpRhJt4rnzZPRk+dOpzAubz7omckX1MrFd4p81o="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 61168 )
`protect data_block
gD6l00tciPUa6pDNTk/+tzLxvdHE2s3DQL3/JqqujQBC/Ei+vcAB8wM3doqg5vTg
ERGtb9Mgk267i/4Ph+rYrB3GY3wpy8/w0aWmETZcxNujFb3uIdLOJGcr8iARkUf1
6UZX0M28i403p48sSLEYQn76p+A5XuPCoGxN1Cy9b25DMvbDJAYpidC6OEeR8h6q
pzOqOSXiwJfDuy22hQx+Aq8T6xa8VR37+pNaqJ2Nl4E2HtOaK0cUa6XMhGVjkphH
ARYsMeabDZRO/DUN2raDZa6CV20uCGkbmRL0krYie8FJtwY3O9XYlgTw59Z3ejiR
RuxOHAcFJ4NK9vlj7I1VXlnup/cMlsJDc8YbIO4XQwM4N+cHFfzkAROkwqkmgGDd
oI8G0gL76fECO3BDfDOLcyKHwEmJJh4HCl74n6yi2puloahHz3H0unHWpkU3rCGt
4vyNYUmn/0sv22iW1+pYIhqlm8af8mvZx9apb3TxjC31SMitlxlyHnMyGl140o8k
OqHN32Mc++HJZL3u3bPzzKi7xD2AHYxn9P0bLEKvoE5HpxtHR8GHDaZsq8sOJxJC
3yEF15XuTKhu6gmwrVAFHe/a5VXMB1QY8IDAELuQh12LiH2CazNhZVb87jDhoD/y
dSWSyEA3UKX+csmvTuZ1BM3YuYTODzn7jIJWKjbG+YElNC51GjyR8Vh/hJXHy1Gn
jVyXcr2MVIpdMn95xk8YVjhCN0R8vKOHMnIDZlodUYCy1kKULUhnRnTelYGENQW0
cqLyCYRd3tvkILMkJg1u8pfxa80aw05myqzZx15wHQm/CfkFIy2ULuW8vk3g6UJQ
ZuzwHSRiIh4/xPQTEGKWj8tkeqTBFq9Gv8tFvEGfvKaqQ7BBmqz6+LH3WIoCU7wG
ruIKPFJAlTI8yzxf5kSLNhB6qrHVDzl4hOmgG+wrgrYkh7t+HcGEAZT2hRXq8L5W
oDfsPLrk2xLkFXgDmcL2321i8c2tjTCAe4J3A6BZJLAJVxGYtNXz4KMW26U8kLKs
rn1hnku8Y9DNHkH6DPEiJsFFZeMK2dJLXecs+s2VUY9T7ytCuqsJ20d9xa0Q921k
Pwy2z4QYa6NCA83y3RL/cNX7gQ2L0G6fmQdyScO4tGwQP3HcjASPPn1U/CJyYjNC
wR1OmM8IlG2ivKpDgY4un5mE5MpZOKX4BJvqKGcUMbBLoNoEjNKkSf6Ja+Cep3p9
7lpg3l3DeRn5XtrzefLBgOdJxzy67miJ7yVmef7PJOTIHX/LQ035wO/WRvz53M45
uGWyZl/A7gPGYfe6JcNJSDW7jJCmhYBr6x+0wrJXY2Z1jLO9Mk72C3IgBE5z19s8
mCoJxkX4BMP7GRi7/71ne36Wucs8nAFcv0VnjyWBkNKTkZhExXp1CHfnpe/UBSYv
R+Itq18iPpWgkvL9vI+MM3EQpv7OZZi3YAPKDiUQlqdioFc2TckPvQRdTh6JYkwD
aQVdWl7Bbm3jyfY4a9VSt/qJmE17V67YAHzRyENbdMdhEOZPyqP6nSfHA6f2/t77
4q4+uuVb0FAEjYQlfMsmehNQKDGr6sTZSoemF7NXKuxIlMhU0sLPk31huZ4YJV8G
b22uJVnYg4lHZOz5F5ZhDayJx4GVZMYKySLfovJwpKZtmw/wZo+vu2rtZzis8OzP
cL2NP7nv58LH9yKQK0Y5fHEhhjpOeT/IwjjtkWPzvobtl8k/q1O0jer4Bk4XaD3J
92BiQvoKRPej/0tpnGnusqQTjmXYf2AVPVR9TrVXhwb993FFtvV2nMAkAbqKxkD0
m+YMIwVWc+3/70RELfQ8WSFO6c65RiU+ULL4kd32IGbHK3yfILJpRE9JgR82pC22
5OXmDsnOSCihxpxsoHFI0yssaZFgB7xxiGyEV+cfIMh/dj+CtFptl45469TpWfhx
fVl0D9B47Y+GsKhpq9TRpn11wDZYmSK8SfhfUGVN8gKkPZFx3HUbX89DLbUcHie/
Pz7Um4zeM+kY8UR1VKz+mFRgCuC/APCZ7RtDb/k9yuf0W6OlwJ8r+RXOTnhUgd0E
QyNRGdkpPr15RO5j11HyCW4Z1/iB9pRtyRgUfELinTdVj1P9HUjlYcHeTuOjvg0P
NdFrBE4AwalcAQUjdDt7DcOTKQwpvHDy31nplR/Nnh/N/iwtt+r/k7igihVxi+Qn
wT4IBFQ7ynns0mpc8Z7K9nfDs0K0JaR7yEbxZURVZVa0h+Nltr23+bC+Nqxi+CeW
W0yhOlt64XnCwonohwHrgYStdnmfwNUyGRS3cb3AvDjvHsdqmiyXL0Q+dnnbwDJ/
IX0t5kUXpiVCUtgR1GvgSmVhLsDvuFxk5QAjYSk6pEZPLaxgc8MwAdobLKqtDVKx
H9jDIC3I2F4J2BB/pgoHwCap2U3QdJ6ziPuhTrIIzn0bHrPRwBKxmH6slGxl5EHQ
kaRS/xYavrz6PSfjKq8TN0KSnZ5mRmdj5Ze44IFsF1VR31laFG9DDNxHtYm4OepA
5GJxwjLotMFwRYjBq48Uo27hF8oBvyhoJTC9xeKFG89+ridlJW3WyjGTxvJBSRRL
fLwDZif+SmxOfIDQKS90Qe7FENdqIPVMqiUoGuEwVanlp5/jru87OYxRPL0rAaeY
a++ipMDMgOervJnaXO7cU4LGna+GdSoD7Bzjnz5PiDskVhIlDRerkO4vKDf0XF6z
aAdxV8gilJpCwEwkqTqeGlmrINEipYss1Z7brT2NLAsBCDZoLQbhw8XYsufzeIVN
W8NcHt4Oj0/0oRd9YMkmngXZBrhJlPJ/lNxv5SBCBDuVJ4Wk7GFtqCeqEkcrSZbI
yhz3UfbM9od+mhPO60+22sJ7HwQinylsxUTfDNoMt68N2Id3eoCJ95MyLgDsGvF0
QjChdaKJPj+EFAAR3XJN/ShmfdwBRlm02JvctH6uD5RAUo+RKghiCvhKgEVYud+x
Mhg1BCAss2hW1K/+acFVq+gfnklYCGYbGxaEHVkwsu0EkSAUEVVHTvyYGTC4Lchb
gcv9HlvzSJC9ho+CmJchmiFOdKg0j1HHyKzLfRhjx0P8+b8jITWd3WtJIcpmF6Ro
keb05P2OZTIeThxkYfOqjtSjBv3XEr9xgeWOgh/Eq0/GL2gmmoA8EYCZQ0zS8key
0MIMP9xJEaJABNaB9Rpeny9YBmsSncrvsQVQ4EC4NJcJP1zIyd7hgVee2zCah7+J
h+Q80+Rjal7qNT3/Dq5deTeQnvns2sTReAlneRVkyk8V9nXD6y/1gT92C2a38H7B
cGg60sS7fevt/sYjkrNC/t8R7PsAp+ezBkk4I8vxCN7nr7A2bQkaj6YOYA8VLMQN
/rgv/21EQS2XGIzoxNhskXuA7HF7jqdyJfjR1Xdw9VKtvxv13kB4C55nXZnXz4Ah
VTIKYuSehMjMcQ72R5KViuQ9BWK+7YjpGcAKnSGOKkKSUfgOO/vUz/rZwgy1QwuO
wflemHZrcuvxZV0pAwkcJfAxH6EBlecHthHAArg182ELtKTJPGFVLR9hsT2r86cb
1deYVAVUFovIg04nEbR0GujJP/5EZ5raFWVXMk5ewBWqE0etDUVTiDIIRByuW3Zr
u6Fx4sarS8P72HS3BvwL/RkNWyDBFdzoby16ec7/ux0f9Po3Jxyeyvu7/wJj27uC
QybEEM/9+pmL0jnotD93qKj01EEq8N0ne9A4G2dhOK1JqB7OWtbrKJX8wC3ANCIN
8XS9t+/Mejy/+ZB+zrlMiT8KXDOo9s9O/8Z1V+5I6DWL4qiywZ9sCPrDQ1ex4e6g
eg69KektGIVQqNEo+BSy/7LQhGSnQz4Mn7EmbYgSGEeB7OVM7bLkZ2MGWSe/6Njy
mPRsOarU6aP9mdQLxypV3RbyncwLfCnCo0dfSCwETGZr4lhBIBYI9UEFbNvbIEs2
XlxHiZi7Q953T9EBQ9N1J01RI9jIrglClED1A6+ULeEJUOMcjBKam1m9vcnmTNUm
NbxHBxiA9iZXZqhUZCX0cP3CHjEkuT1lnO5p/2MxbLQ4Plyatk4DJufygaLv8lGa
Eou3ou7FGKCFj0OqYtmWs7V2D1YbnFZFiVL42Ne6Hw2+ckBIW9ir1dF94KF7acdB
E7mJ+TYRsAiMWudfM0UUW2j8oNYxOvVPfra9N+u7Oz64J2kAc9YcwuSsWu9LGpSZ
SW9eM1XLezHzy9d21b5ACaTVeeL+sC8BXYy8q6EnqSs8H0+IeVMgDpCe60d6TLxl
mG58LudHbpaDlJZyPZav8xEWD1xiABYpEyBkP+ikb8/8UJRa4Az+A1yD6vuKZt4v
W2bMDW53usO3ekI0XwCWBOP/Klb78rG1JjtcQ+V2SlkdflHk5PD55U+/nnhid5mQ
op3vB9tGyBR/ir3b1HIAjVnx0lQ4fFIO9PVtJTNaWD/cx0eNeWlTAnnnq/ZG6Nd0
BYZWKBa8U/leEf7GL+7oI08yysG5E/PNDSwHA/Y5XI6ofuBcOfCtlnj/E0j8QMu4
378gE2ML7XH7VNk0IALkEL9C87HRdscbi+zmBa3MctdDJUHMBuvQvFUHnddqw0eQ
/HC1GnfGGR6iYPkZKzPvDFSD0TU+8pCdCXTrIdEbRBDB/rorHqfKsTmv3s1Gagz2
CBoXzMVIkl2Iuo/WNQwG8YfO+srN56LXJhiJ8rQedEcugfnRMj5j1oz1RG3B9fhS
xmkxBBlXJRkddXfudyARt1EALlIw9Co9JtdC+0qCCqfo7/H4wkv85EZlfrkvcLeE
5ui05JAXectJ78V/z0JWeGtuoLJsETbNW4a8WaLtGZu/jPAOYBfzbc42qIufaHmY
IQFa996rxXZE3cpjLVb8/D7W1HOdWR1jPilS5Hk0BP0RENl0zbsje8fGHsIT3Wor
zxtaLx6NdSPVcURPBeeLvs4S64JI8enXrVNxIOxkPQ9gtAXERWwPfTEtrpdDTr4C
vpISs02ZmYeD+k2BsbWSfUEUXZIquLNZRFuCbPG1jIk7LhXhvZzU4yUDsYNk4TMX
ZkeaIsOascJQ+dJglolsAG7iXtOxjVOc/OUYood2BcDoq62XKn3V1AlWJI1Aa2bR
VQH+xDHpgSaIZQOpINbpUUYCY/MMLz9Gh3LIQWca/74DRI2UhuH/Y9gJt1tnrZMX
HLDXdju4q8lEsHThHYBDNjxdCks9z0SWCNhtwLFRqrlTUzfsWZOyTi+K0i4UyavJ
pdYH6ael9IXYZ1kGNnkvl5a+PuJTaBtSP4+Dpwc/WvC1vlpEuK3TmcyEXR+C9fQ2
0uISWTBoYW1rxTp3yAagBSYOI6xQNjn7jdh7Rs9E3HmU+LFXV432I6b8tXUSTCgc
H5/k0gwHxKUBqy4ruM+l6qyaFjrxj68Z2lqSVlNe4QY4AOhOhuHylB4I1YkbRkf6
4JetjeKRyhuh5dYiNk1GYobvtHqFfEl5FkrvSeJtiBOTruQdG7ypzdEuGy1dULY/
J8dz80Q9suqa9OB2J7sUz68uqCghOloxP4j4mozbFbr2rfGrH5oEuZ6OvXfSVxMG
Q43X4tM+pUCFSkiGCoGagbtLALhxtJfTBZ2kiib6pSxlbSSId/zbgePzH1geVunH
kAwToJYz4jPsVkfLHvhEs3UZfVHyUOmfyfHGvkdRzz4/qy6m1nJICCaCWK6OMUCW
7Uc8Zoa9A2dTN6VaQkeHZiwmbKOcTBbhGJ9Qm5S5B2N/f/7PgFH9gBz5IZb+/XM0
nyb69tm/tUc+cp3HDmT48W47HNbuTwluBlAAiJwDFH4zFqHap6IeZ2J3Uos6sPfR
X1HAvfodVlpbJoB2jGwEgkXjxjuXP8rL44SNcODxAPZoEsEDr1PsVicP7VO+lVOp
4ogp0aYBSXJRA8J081fq4yqdJdGgAIuPrR41B5HPm/2HeCSP1Za7xsKg1xzA8ACd
puNLLj2oEkhe9aFezUVcCCg3Nbzn6qiyyZeTe8kuCS89ng+j0Z644tHC2B9vOOTh
Sfn6kVVODI1mk6fQ1Ld3iYZZbTx1qjaja3RJBZUT96yqTriF+Wy++uKdpZzmVNd0
5gR8y+yPg+DyrQq9Q5xo+OChrndi17JaSfQPKHOo+PkBTDFHrv3kpQRA9185mY7K
8tvBJYWBhRuwWIOG6QqMLHvM9rvoEzsaa2MsnGt8g8rs9BqQE5UrGHIgu6fxtNkj
4+MLHB6M8u0H1a2QKukoizGwuhBNeXLPnTgAd194AJj15z1QQCfeACpvIcmXuFom
7hTOqSIRNn/iNUcF+MdEq29Cmf0xELbcjNtRM9eMvxPjM3THi4oeuLXnj3HA5Ai4
JXP5OntUnE4kEA9DaTo5Ql31AWDUyFeLRmWTLDkKPIJOyH3rQ3N/pFpLL0WChcJt
ZYD+E4BB5WXpBcJHb6yxs+TsuDubHmYYs1qeYj5VpkYzKWWjodG2J+UKVPYFZJrz
uvd+OMcZ9OqagkdVwZbP1lHiPlh0CPOSiozVf69YgFM3ykgY6wPzF2PXitg2BUrh
TzBn4dYFk+OCm01PnOlnSpTKimv9+UiB/ccLeZsOWUBKsr9OGT5VeaD4MZ6P9pK7
t9fr/jJ8RVtlV/N1wbkgIQio/lJIg4dsJYOj1J1WbGiJvMP5KTyNwwdq2064+4e/
LxatKG407vRlNpSWY9o9cgntnInWTlIhxvhxqZbda12gJ9iZOL1weL/0arAC7sPA
NBAD4aQbPEgZcg/9uf0fM9pFvVOaALNSgz8bo/XSGLKC4urnrsnySksgS5SKuq/8
nZrnWZSLjl/Gr3tLGcGHhvSr0oJ5xkX8Lnu4qGYKcQj+fzvInbsr6euiPv6VY0g2
k0w79wnU2iyn7zBFjtSEFhTy2h/dN62s/EEWdlcZG7ubtljugSsnSVZkMWy0TJQd
FYYtRetZwfjx3No1FhV9ibFz0emJI2EfkixJhVPZtphcsAR8KHiZp55BLYtt/YUc
LScSzwMyT80NKhXzywCZIpwKsD3AFoBfl8bGH/ogkMcHUAukuxgA7KTGZs+nxjq2
zVElQfpvmIBKRHFEdPXUS0MFj2uzouNidXWA1+5M0f/X5g5ZDMG3oeUfYznt87WD
bvQ36uBI4EEH9qAj0bYbWR2pfeH9QD/KJUF1AlsC3M2O0Z0o1hTF8hrkb5nXfABV
esFBznnRvMW06g0Q14Vz94YTMO7UuXHauzNukRMEbiEYuQPGMkqvSMALt3GFklUx
7qZie61dx1suFugLhKe8pqvNzyZNENClDJ13iQv8DnQSDd9BTYsulJjFnGrkjUZP
8Oa0xXG4ZEbB1+G/u34xLK8yhc529BYzWgeTHUkgUYqEGDj5KzFW7sgmsTiLfwHS
LlzsmI7+G3BWloIDA7GABNt1Ff6yRZ3oKCqOERphRYb6tBm/V067YJ2MG+hZWWc7
cl26aQY4I4MFctEeVKp1YFWHQzJKQEcp0IDYGpXQsg7qNzFXx6qv3cBvJimJTE2/
gXB3NlUi+Iela9JKaVEwf25CcncKF60udqzjhWNtouxCpdDePdSGK26HP6XB56a7
hgFo13OCesvwCP3RjECaz35bMbRiP+S4V/U1VRhydHUzONrYXswRJRfCBjv+0n9R
uLlQ9kSph4dxcJGJN74a3bf/ZrZ6+jIGrkNllw5jS9AFi7Qz4cSHwmK+fcsedG/w
G7AvarhPXQM+4QQpRS+Rr05YyfLxPLaJ8RXz+AfkYr2S9Nkl/RL+6KM+CtPcTedp
Jx9UuL2L5q6VoBlv2Ru7X0u7N1Z4tXLO13S0VALzyxy7TTy8OjeUoJxEBkV/Fzn1
2La/UJngdIwM0NjctWN5e7lVzxnFMe5NwiWDkJ5qd6jxl9pEKx6g9ZcuhwNIJ+/s
Zu50iYgF/Ni/9AyuBoWzChEXM6uQHz3PMAmQibLb3O2bCBSjTossTR/Ln/o7d8Jp
3D4cCdelCutp67E+re0Oat0MUDGDyCY+fBPQlrRyxHqe2k1JHFb7WM7eD22jElSd
aAh1q1z5w5EIGOS/hmI63nW6VxD0kD7PguuGvtENmP5fAPPOJa36U3cmPe9kZH0w
h/dvS6PUyixhSS1BC9dN4N4neer2TROUGvnJ2sxTsyPTJUDsZ7S0DQYkBN13Ydzm
6e4KHMZDUF9e8pRcE/at00z85Ml1NCZ68DTuwYoS28nMHHipMllhz0+hHLExFzAT
Pf/t2EpQbFc/UJzv0AtOXcvoDDhwOUzUZfjvThFdVb6MIgPjjQoFbR5YOrwK7CYF
SKqNLKr/z2vyo2fAywH9YK3+IdJhFziUsP7wAh4aFbKkf/lbg93sbkHHzFVlX8ky
TeipsoB2dvpsr8pUDbfss699FUuUv9fo3BzgWURY0HQKxdO3Ui55JveRWqQsqdOe
BZW9dLbAhP6Q/tFmCuniIBe75R+7SX9GUPDAEkypEhbjBTVl07GolKI1y5eJPCPp
gZuFa2hP1iNPvz58HQPRnvYN3fUYoXhD+Ls3a4s8MYkZGe5OgVAhZ+Hyd+Wz3J07
MOghxcsS0kQSFOMN2L0x55YpUyXR5pTU/FMogFDHVua+bJwlk4pgZ6oDsOVtLp/Z
nDKgXTM33Lx2OcMkEmU6dXY+WA2LenL+8wSKXcVX/3W6c/e70pvqnRsLwyNofIl4
UzC4tGT2ImLgSrCEZ+XXJgaK8LGVZ5EpmYcwpmyNfjd8y+KP0ESW4vOJ5+tsq4nY
PcicT8kwMoTFSNUI8P5YuQQ1G0wkycrhGpaRK/o+9UtvaoAN+bQRaiRQa7GHvyH4
LaioxZl6cEjs8AHd9Tt/kZksXYGy0/5RGmFR6ay3wYpxHW8vbAQMtaRlMuxyG/Ae
ARzf2rV6+QplZLAS9fP/S55lbUwi/dOvHDad7hj0l8zZdZ7v5covACHeKr4ZvIhH
+IL+D9A4sY+ZAruzSadqpIQioIHV3lU6hP8Aoi1wXm3UXAP9XNRhdgpEasXnA+0V
snx89le1+hYYcQEOK56jRbPVTsTOSMYE+vhePryAoUiKENg8gQXcXauODolyCbbs
g0mzzo8fTQKzWRHvdTKbmK5cVYpXQi3A18VIdov7ferhhcgLZrsp6siOdg4qCkSa
XyVpHIM/mo+gcOtl43Y/QtZ1Hw+LzJfBwwDI77FyXqi0f8VhBPXWersnYNL6D00K
/3GQ9P9L6rkRAsPNigweciCKI52ITduPuXCpcuQ7IFgdqofYzqsHmwGGQbf1Dl6m
9sVMgBzmoZNUDP5yXcRkIfcuzDTEDewkR9L+ihimq3vQKGbH8tw4GvURL2Q2xEDI
fWRdKrddM/Igk7aM6H6P2+NKqLKzWED45Md7u0PrtT9FeICXHmKsHo0gaTUQdoFv
KBc5f4L369V48erRA6X4a4HlcxWv6GE1J6ncH92Y6P1TlPCPgQShb15091h9XnaN
JqIK15Wv4NdA1L5Mk1L5oHkCgk3A/4feSgIh5945yC8BdTPmHEim9HT01c+fyzc5
hQsbFD6EsSlVJea+vUlyYEZIbQRGfmAJyR1zW0JDKAmjydc/8KZ0+9vsNRf8g88B
VtOW1kKM+Yvb2Gjuk9j2R7YV85Z1tuKYjMyxpftTspsf73jlSXH742HYMS43NGgT
r5u5Eq/Jd/7vBE1clNFQDFdEo1FCktX7C1bmEAlBfxdDlC84RsNE4atJBHl+Ju26
X2JeRrHLaQ+6xr25fJ5vTfDRt8vXPNf4Rdx82HbuB01Rx1NwWQ8MMBu8x3W6pKPJ
uS51TkvL93/KDOHnq6wYB5+mGkyjkS0oNiSEVWZVHMqCHOOLyNVsUkbAhmbaa+If
Np40GrN9gmmPe65v/bRP9hlrBbEqavF3SBHNkUPCyWxTZzlrE3Yqi8aG6lreB/2J
QAbtAqEdVgKkjVA20Ifcb/Vd4I+Sm5SAEkWd+KxvhTLmSF2JQvk7CljS78JqXIUG
4JRLGmF9TplgexxEvo0Irf4PghjAKMSrxk/8i37emVba8UlZf4+zYgkqESmGQlQV
CDMkiuGU5iWHisNu5SvCROrbPS8hwS5tbQXSLhI6wv+1JeEBFm4NZAk+Reydglau
/yAQg59bHgawjisARxYr8DQyGJrUwmiLvCPqmvcRlMvIryy4OM9NhH5EGE5RQn7W
F5CTDhv0DtCKnSjPoXmKkesdvmjfVuKUGMQxQlUUIhdQBE1R7W1na9Yi3wHh86CZ
ELmZrRRCJXPvdX/e2SDQYwKKgtLti1LryTgAtu6gg4850Fg62S3e4TZw711O69Ub
A/ngEbzOA92k+MNnLvIjZum5HsTUs4O19SOJfpmZsjUxnBrJt8gf1jNwO9kMAJTg
+WMza0OcqStnnEiD2OOvIX8P8JsKG5YDN4KsBrmwwM5RJSfHSbOz9yTRq6VPTunV
+273Up1vXlB9VEx3TLj7tm3RWsmtyEUVPqNT1Az2sFYaaYtU0rzssiS5sh9/xZf0
bTUOkk3xclA+wZB90kw501GYopO+1/r8Hl0i7GcUavMNTLxfuipCCkVsA+LZ2aBo
UDPfjPChNXZk7e73LVprqkrlqLOVSJGpeO7UZHpZLcPWML0o2dft5V12s75nQaZr
tv2amb77hY8ujhT9f1av5gX9LjOvRsK77jU0eoaidM2rhM+TXOUkrXAHX1lOyXh9
7Y8DYoKyglwx1CGnqjRw/gigRvT0Of1DCgl4bmsCBjtm6W/K1kKWm8qgG1q9rUdQ
a2W2G6+VZU4yGbSi2XygZz81fzRHPRBDMwYIkD6UnR6ySJzn+MOlMtv0uiYS5SFm
isTx8KeYLJSAMi2Qa6FVlBLB4/J2zvZxaJyJRIkz02U6Mcp4LXr5e8SbtrXy0vPA
8w8NKWPSfG+WGLzAlfI50kUe7PvDNRSh2KVdISzgjwfBrHaaxwLIz63cEMhcaruz
A6qJB9oXirw0Wy6pZ4hjjt1dCmnX6Q0xEQXW+vLnjMhTXEQ+rIPMbdZzv3f+YYSk
8E9QB3W4AcEf6Uq10FoZNpVf8flvz0cyUjPDX9LomYXpApsGSv8tSaJaR3BbvFsE
nvTOfMDC0CqWpBuBaFhVGA3ZJAV+R0M/T+ess53d9r7BA1TqMvE22j8GVTnZaUQl
ry3Z+pPeiBlNZDsQglTh78CGRIcpnayOUbf2JDAX5exPGOreanPaOJgM7nULgK7/
arTEZYLdVV74RBQxLrryE5uxRndupC0uJlqXrpj8mP25W2nYIrtQ8vBz5goIVHvP
7c0rQpGrek6FNFiAU26sT+/MN6xpx/lbBN5p5KpgFg1vVbXOalKSln2vfk4BULpJ
uvef3SN5jMF76XilNTro4ujhwujbl9WeiHX0HEX16tlamlNEtioXBRkDi50yvsWJ
uQCuAHMyKiy0pMCL34j+SqLTi0pjNFSHW6xU2OLg3yPL3GSowYOITb7utLDAGZdB
flkTRmeAwJOgafOLENN1axHLG6EDyEnKHV5vVk6p0hfwi/lrWIqYBrIXR0UiyY5f
gOha29CPoVNpgG2GOryTQwDqxr8389uVokTtp0xU+QLJ/pisBXj1Uvr0PynzRJIE
z8zS5VXSX6jFhKNYEOGBHV2L6Nm6sB9zIZPKiv0I6v+C51VJ4ktq0oPbZDNfVaBL
5+2GHZZkQkFujWO4ipJXBYOfj08bkil9y0TCVC9EyteBr95W9rs9pQmhuHy9jEqo
PI/iThLgD/dbT+A2vzbj4RTSFT988HbyxxgAHRG11M0RsmVl19a3rnDoLXPleKS7
Q37lrN2jVXNsnUJO86sdZ1aO6x7OOnbiapW2yty4FFrs4veKeeNdR99OMXv3ArIk
dDFHhqW6kbUnVg3+ClZM4NHWUqh4wa7tUlGPC42LgXWbQDlZlPSVjQmBELiGoBjp
jacLG35lBZIk44e+vkZ4X10VgGGeoEOqdNotONfrJ5QEZ94aGjuQRHlMGUOOBf55
EcaO5KNUgZQkKNkroQ3wT2U+uJEUK6is8YPTYjYmXDq4cPO1cVCboMDAx6nHeesR
MdPAQj73t+CtsaNJXHyRo2LPbfElAjfSv0w+uTVLlLudoIfaI/j4xoPOOu+n8Bqo
Hkt2yRi8y8ZcrhjnScIQfzn5tlqm6FkLz3M0AIhqwcdpMlKpxCdYaDWa8QcOh2H8
84o+UQNrVIeoFyEb5lJ41a6WtL6ZG9q44BAq2SBOi3C74h1aT36EL2J+9iywkAHr
3Ct2lB2iCFleXBGWwVDuZun5m3olGCny/I1reeaFCq57gqhAbhyAzfZaWzqHhNKe
sh9sX4cxu7iu74tV6Ko79MMXslulyPfv+emk38UEyrIgr4AGPJ9SUQUMuZS4H3F9
ACwSIZmmsyogj9NrpfKEWHdkwZhHjWu4QzpXN/5kQdTOm3llkgEX2LiKT5tN9Xcg
QSQdrPGlTlvnj88o71sqcXNNF1xlOh6vwJ4hIcMgoM9aEeM3QFYg+Uka30YBan1g
Xq8YW1DDizfIi82NTyqhyq0w+1KcmCdG4orxF3B3PI2XjvpbKQD6S1P6kDSnauQR
7TPc7Yzu+++VfQcGHZzUJy8zjNBAOm9vgQ207oXT9wGiIboiZr7u0liO/pWpBCGQ
a7bgGPXTtOcZQr+Boih40+rJGC3VKxEr1/9MpU+EZm1/Cbu1cmV/G4PbEc0G5NFC
8RoxXShPsVOmwaHCsBkP2q2BQPzuqJeCZHbob0bH9Mxq/Z3N6IUkMS1Fmj23+uQ8
a0+Oe9yoespWNID8eHGB57/YqOWyzwm6ZX/AVbtYXRaMkircDh4y4vBiGLkrkSSk
TKxTbVoWk784x83KvI/yOMiLbho8Af/tZ3GG9sV2AqUF8N8FcSCyL5pURzw+d4Wr
6YJKXWbNVnLsBldlq8iejVCQRGPg7sDx7kaFobLPpDEORlHRMP6Prl4LthjkGj+5
TnFZ3efH1Qn920M+Nc9d104E0YdfhC0Miti4K2enGQLQmjRMkrJwZqkiyFwRyn0a
sfFSz1Pmo67Oxi5DU3Vthc/rXWGFZ2ij1UkQ4t/714n5+O+sroOGrwWPVsamsjcf
DFWfL4qMM4qPkgtdSBFWtE6iYrxQd+Yz/5rdTogISHuLoWKY2YQj1xTEmgogel26
gNZ9ltM23DsyuOiA6R8f8hTjkUCTC5MJi7AEOJygTHjj3pzRLCpF4ds7sHhZwAmE
5sT7qBUlL+u7RR/NUYFPB2CAJZcrQ3EQ/9glHV9pvMzFCnb7tnPEzHI+M6OqSVmO
pkR6h15g3uMlCN+vYosBNpgwPLomxIFV59XHGOse5mr7toHHh3B1vjm2Bw/C1q4d
CUuA7laidc727ZHgeXlC7LofzgUHA4h+Ji/UmGGG7SGWPE8SEo3evBQ1AU0jQOv3
5nyNzDcKqom/WHfFwLVmHPBqUIjG06xfIqeuk1TYdWe+89HGWgts/1HG63VoxOv0
VPfdLWoRndJW1OGZ6mFmCl++tSJRoR3Oo0MuJmY5KOkmICSDcal1PQZhoyvhcluQ
XUV0ROl7HFg3yLSfKcnnA5MDpBymTMDsAdAvxe1hafiVWDcnX8ubNhjHo1P0AaMC
uKOVvOHWAb/c4DfaukxaxnqJzEQ3bGUwIY1M9HUhM9bEgBdxYAhL3tU94y7Y4trj
zi5a+aH6Q8sLKdZaE7WNoiyNCNpAdg6yraRAOdSbFuq8/UmXtqTWImIAgwFUdRFF
/NnJICbP300EUX6FAXs2pmapfFIU8Yg+S1D7ho9AilqbemiagB9kBtgOGnU9uSOC
tGP4o0Skdy6qRCrkOzZmSvdT0rEjVWCnSRdh7utS+6b7xbHv7XM3eguoVkb4y3o7
c4FYQUoGPqOKJ+aLwqcNiLpDwC4o0ngQOud59inR43BY74RVS3cZmutPvTfeiI68
9+PuBtOdwCE8FY8RRs2BSlnXOaRBT1HiksYPo6GdtvvGk6SWV0MjL7gEkM/TU2+J
NB/hB233EslXcjf7ew6EeL5ph8UoiYbY/a7LPP9tmWz1yGsfS6D5XlPXWk5YE8WQ
yIupxLO5fGMXiq6rI6Q1SICzoAmyet2R9B46Hy6kaZt/uOSkb+mWVfnmIIwKaNqG
hyPr4bS8WzJzbym+GcK4rRjKClU4x83XCQuAnkr69vRly8TdHwqWr2crTLwrFas9
tTfoRlsWKU0yNh+DJNFwvU359raKxuFExIManEL88NzI8xls8IxM/xv9pvBYwWCU
gLFUnybQOf5nw5C3WjI+FxA8KmrwJDhFsFpOIvUm5ZTjrlh2MsVKqIR+ujnWysVF
iV1keP5bHPtVsaxUnoD/OohhA9V3sAjw+lwZi97sUvmwiyknoPBfocxDwd4A76x5
dyVeiQjc0ZqBl240Eg1+R7smdh+9/X56BtOm4XejjLKR0w1vzHY2AjbDeWuJvawi
WOiyEQDAolfw4Qqb+mo+NRKzH9mepgo0YZthXPIOL+1cq/3fxg/dymAIDbfoz26R
HG1RRID2uQcW+XLF4MZyy2VbhW1jd38NY0Ty7ETAoNWryg8/vdW5M7KAhOx/Uz+5
CdvzmCKFJ3reO/e4hBo96jx6zAQbuhOuwBB3iCIkz8biUkDTQqGcyq1SpAFOlDYK
aeyh0PHQLifLBtcrRBG8eIy864sWuzRaebOa3k4T8EI2tfVUUE/6ZuAg+jnxNUmF
zNtqCCrkvPc9JTysbM4hhQWVwjPN1tal6meQDsqmizt2XABIo2p05X3zsYO+S72p
K47Hw+OK+nFwHqFI1Vu9/m2gyHYXt2ETsJZ6Dl9s8+EtAdj9MvRu1yvhMDh7xUNC
KCWYvDD0O+EIP4BE3UhhNhsewxg6h1IBPSxONeva1ni1XUdnLD2mWgQYrq1AvYeZ
78JrjfkicwXi+IlAA1Sp/oFPS+t2j+8Mz/XYRBzlWB44RNBDd5wPAXoMFGjquc4u
KO5X/RttUZCiLvjKR40E6sECElqKf9kUElBV6F0B6XdN4ociuY9tP4voD3v+R/XK
tR+PnbhjGuonN3GRuDpsy/7MmW26eV3iI9+zhTer5KBIk2ONfnUH1aIkogf9w/sz
fAPICjVJMcGrTpeKeU6LXTxnJiewjsy04+uldhyKOSVecThwijWxA4iCwLx9HcF/
dK0YqTXRh6Udc6iPgfGrWzbGKeHClbtefgUqll1w581dtjVM/5ec0axZUqrQMePs
jWBVtp6fxPTJkBv+ej8vhsm8XC6RmpMUHZfUBA+8TR4vMMLptoU157/KMlUP6qGs
4TxHcmAxDfLM7YOkZITFczBWg2JB+epfQbQztYr6qgIlTRAJORgt/AngrMw9hLSd
G55xKJ11tbhGdEiwcUa5rxUCvO0TDkNEqsHrt/hgVUahTDiqJQJMUUxedH35HYNn
12Q3z7OdqWuWoznuluZ1sFX8ByDlYkqzQybQCrgYBZUu//hdWId6XsseI1pmiU+5
mYE2KP7b4dU6wgexHXMxu+qYR559zAs+JFChZ9/yELhqPeqCHsEHqpyx9bRH321z
PEAaN9+oohKxOz9YGx8DdKfD+FxOZZ2DLMb1efokQ16/sA2Rt5prFAtRJDzPbXZn
ibmqro32dRDnwsUKPu46t2yXWX6oVfaj/1xTb32UwouVOFV15lPGzF/xa5m6vARX
XE6Gy5/WcL0xmHr2p1IZ/Xt8wcqSNoYP1ryvTbIgD+S7Dk7RsySJ9BP30YLLxXDP
EWxB0dXm9H8kGYpcm+k2vzVrJeRPOUmYNks26k4qzOswWO7bbztpJ2v2WBvyyeot
lRONELNZxIJIdRjOZdFwXHGTPuU6dRtQ3nJLrUIBY8aZb7wr2wiDuSF/T50m+qCv
0UYWLF3w+U2hgQYH7b022NGBruWIklVs0YtSICW/elNZSDjFO8WhMaCq+k//bHeO
bOD1L334/Zp3zfIG1ud1w3NBi28FlmGoIKE7bDZXt686TvNHeORblhVFDxPeGXfb
k2lMWgUbJ2oJtF9JHK02Rkvc2Hens9i5xEpFm1nW4Kwtnm0wHrv1jKaLo+EVW+Vw
O7aqLCBqqegWJaztEC0+ob2TQT/2wBnmFPfHhtzXxXhHKeQIlpeMhc6R8sHG0i1w
faNcj4BF0Xl46cmBZWd8yxC7QZluwTEtInOmiGIW0xpV1Kc/XHdTsLlgcmNWg+Fg
Mhb+KBExHo5RA+4Frx6UKrYpLAajh4sbufzWgOE9V9+IAQZQjBa742nlaiNu7Xh2
IuFgfH8jI17avlp04bh37GEn2yCkhlLjkrIRg7l53/BIgtMw9WI3lYqMqcLcLia2
hgEiCw3DaPiZCOYfkUlYJC1Ej2LX3WKbn6m0SW9vgheM4k4pXBntC48lCyjvFBeI
ib11Zaf7Fy/zCJdcSv31HCg6YJ6c/IT0z3crRpU6+iNfLl9JAFaLV2UfjAbubkZz
3eQIM78+tnekF1s4+RG05jUb8yknFeJXUtQdmJjp3V8vOEP0OdblVNIpqTPbN8Gc
bkHG/QxsKzUXQ1XS75j+tqu+VTnveOpvmfJe/IcXV5YH/wc5yF1OiHk0uUQyrBWT
NAT+RbPCDG4paZOpYQ6o41RDz1DLAU+zm2ut1C3QQ3Q/6J87RJfYKV6rK5DGfxdH
dqKq0lidmo0NC+Fh/IJDjXPqIjJLHSYOJfwsIHslms1IzVOUtdtlOzAiOMiAIJ8r
gP+bV8VmB3/Zb4/FTxEBoCeP5BJV9Y1C31ddt7GAPfqBBi9ppD5EArcZQQInMZBE
VbEPpeYjirZixZhq0vsd3BiG2pu4D0tUDHvSLjM+/NAaZzojbxnTx0NbjklQM0WC
JPvHU3wAlTlAi/pG0c2GzuaoNfgOWkJ4A2Gw7n7auPTc6x9+9N98Ruu1WB4Y1cNB
bv+QFjUGtvQ9qclWzBZEsW4POr1nsmTUI0F0NJOmfIKJlkmCwt+312RPTplmmYWm
lWer0y66ABOYY3JwuLIgoYp1F4mpEiru0a+UzLbDM5tc+PFtaamHl45+YrgsI2x9
0ADSiZDOXfWvUyvmHgaby5m8dPTXPRI3h5sbbxEuWku4NlOlK/Y0zkqBt9Zo6qqi
oWJkX+0w6TWmV3mAoxkj3pJRe6+pIix5ehesAkj2EEM2NPFiAHLC6QWKHVLSKw1G
vuqD3XTfyh4U5BS3aHdHwE4w2kEYqHk5GFLrxazQ4/F97ooCFuc2gWk4G/eopaBC
325muZQPsnwsX67JbsXRoSyaZzMjCO/cCYyZfbQAPnxEIWcNZmPbz82WktfiGZxV
G4mhylBtsgui0BM07RG4JKH+7TR+bD17ZuYACBqktloT93d4TzazAX33J7N9c1qM
ZY1paStS8X+Sv2E3m3cfoFcdyriY+A+yBWSCNO2lqQqwwtTMqehbxX4QpoR/miQ1
crY3UMQfDI2ZheXGIHxMFtAejYTWKBAmF6P70kEhH9IJHp9cUR2yBShJj4qhIMTR
BQ2nSKBWVwv2gjL1NDHMrNAvvBN/NbYn07RyDcUsLp4DuQUzm2xEvDawNJEWDYmQ
jhSlSahYO2Fa+xVLvFWIVZM8echRzoxcL5dV1VtIb0stXBt7E2BT2c4SAwzlbqRD
7GePh0W17Ofhy1RAS5N+yHOlkWPB8cTQkB2vmqLoct566ksasY1AuV8xlVcV6gJQ
4WRCbYNzDTuE36p15jMrd2kajf8D6D1LI8cSx0iMCafetgkNs8BlTd9SEfjjFiWl
SpOK+m5aBb5nnZPqVScBuDTrKaWPlj7Pjg8Kojftyju60U5fxseBHXlbU66LA7Pv
dFExL/73WTmE5+68qd0ZjAqR1a8jp2Jz/hXV/GRK237OjYAGgeDhvFpZAHYKisod
l5ZA22gK3GiHf7ldpG9XLT8wvQ5/v+1Le1T2xqWlQnAgizdF7Q8/Q1MSWR0hlOWd
ygFZqGbiMk8Nvx9wRIzPzTzxYVrl8cWMOQsIP0x679flNZ1GJnaQK71p7xwWDZAp
nDLF9mopsojzuU7+Hz3B9zxbiHWvJB0vOCdRirh1viOaf/3aAtzbhbp6rqShWgp9
2cNCt2iJyNz7P8blTOz4jUUUYEmUDh2W2GuM7uY5fgfHcKD/kTqJNZHFzY0ruoi3
ym7z7E757zD4iA/DVOWnVtZ24y03QF0VUHoCpXKs8M/gRlkdk8VyXgQMoi8hV3Am
kZuF0DWHJIOiNZi0ro4KcomU4Q/HiLxlVvPdCos5u4nq4iFInNNAh9/R7IVGOXEd
hTCEvWS1VCzpOVnoHencastAEau9Hvx1ya+JD9xswLxiqitRC1mj6HjPWaMBCnrR
A5PvIKQFQqdfkndR8vwvyz0XzAGVbPlZ8VZUCqxuyqflipb95kTnsz/B/cbp5wC5
HL5EgsdlFteLyRwFBOqyitGbzEx2ZMYnjT7kLxvNKlasbmVUx1hmAd9ixSQO5H4c
F2sBmDlQWoRQw2/b8pfuHB/VuZ4k7FMXRSW/aj3rVJv1IC3aB6h4XRWni4WzYwQ6
smcNF2f3j/gpSRq0afZUtU5JFhEVQcVjJJAzkAnPW7tdAzS5FlkEpxguLdtvvKE6
sO/AQFJ21w6E8f6+0n1QNVOkMpF+X1hRCHCx4dRu9W5hcCYCDR6dM7CgK1mBDen5
2q6kT5mCejdIRXx9DJ6Esljfh5FHI0wWP1+VnTFfnSKucTox4cQJYkNnkWmeCANF
hHV3C7OOLSBNNFV17h1qlEAkJcuXlqVy2+HshafASONXpFoA/uT+bIEAoXxqTVb0
cudphPTpenVl2kEUaRqj3BvI5TYDW8ukJhVwFPaaqKiFH/5YEXDjLaSVV/ZDZIK/
Yxtx8tp+JpiO/6ld6ZNDE7btrsGaMrhqgUy6ECqHmiKGyLOU7tS9nEEldZlT0JEV
IcrM59IK9dFb1xiDKMnZHGywtEzJTwDjNHEQX9S4vaXTRmMaimBInQhMoVImfwxv
A2RjXcl3Rz6KoHt4Aj8TAHidfXyF8k2n9n9I2yf0l97JooT1f5QgD9xlGlvYyOon
eXQn+hqx6e2SCo+IGTA5902ibgJz46ooVLT9ToyFNf3vzoaVWmd8ZEebgZqZoW59
vzjGg73/3Fx/3SHz+IeUuB/Fmnbs9kzMtecF6alJeLrG5Q49/C2Zi7kiQJ/aOwDt
BtcPH4jD+aBWgaOrAfiE1hEkBW6TfqI0tr7a+yoptGTHeZIO4itZNqTON4LNqy2a
x+rldGXX/4QvdU+tI8Z0LdZHqPdTFz0i8UugkGdga2qDrQmgR6NN1rwtQzQFUA1V
88sQToTjw42jChoIJG6kC8AFXUrmaK4Br6H+K2HP2/7yXEmthzYHluQNh5ikrafL
6Kgf7I6+c91fTp6XsFO4211NESgb6ATD0j3f30RFf9LjtzPaMRFLs6arvWBIcI3w
kFVjwp2mblXxSbq89ZM0rtjzYRFeev4eNfeO+GMgPeanXyfbmCkzLC7yZIGuNUu/
dxaH6s9aUoNB3tvY6tHnngAsMC9nsWLCea7d8CRO3C4CuTCz4/cHuh1upSxFMDgC
XW9vsP5S+7h//Xo9CAmby+ZDyll2YA+C7iJo8fLkA6jgWJWIM98fOwDB1nzxlbsM
PWWW2YfvVVPqnyh9u7v4YhcrkDboMCHoLzN2aW7aaHkkpNclLrOJ7PJpfVSuonl3
tW7jIE0qeWfshdkuW4b1roRS45PK7r5MpSneQMwh8n4mo+4oIZnQBTtP9PUvwXaQ
zsan6vDeDXvLv5/517cfB3wQuTT6jQ6jzr3IovF+4MremVqDPS2735Tl+Re8pe+x
sky/SjZWWN/meN4OavRq5aZt1f0ugy6VnDYqLI3vOE8al4r1xEnNkNHb+pn36mSA
4tH4bR9JqY1cwdJuU+fw/rHoh3vx4lVyiCHZGgWa2oAEFqwSM9QKQUl1eQFY5sED
P0Oh8Hxzt8VAg0d4Ht1nWz8ARygHvE8uh14PBwkmmKyGdCbW2bfYDaSemmIUlbMU
uS/eLe9M0YRetKHUWlWS5Ai/Ym/QHg3XR0mEJgcyB+c6GmFxFFJTPYG8vne9soSb
sco7bRAbOPs5h3tqygeSp8AoBilec0xNknBrGP8HhFicMTv6Ho3jBGRGAI5y5nwj
VW9U6ZanKHYLlzhn0l0ZJ/eigMb4ZoumFrks8D3auuGdby/GxsiWnUy6bdl3tzDi
udHi3W98HAx9OUZTiRTAjgGxa49gqksxXkyBxbDYFTciXm2CKSGAxcYmNqMdGPUH
HFoHkEaWP5W6GHmQHt9ETDxTiv+g5YC8BOy4nixpzWcf7l47Hk+VAWuyyiWvlfW9
dUzScOzQe45ddBXGeKtw9p0uYhoFgIbcRC12Hb1zRvNdaeVGdGLj0IVhMS5e74sb
8D8VJ8SvAeFKcr6zbU4rTUfTFPc1k3ecsDrTeYhHzv/+Cm5yis78SdOhofmwxyW9
Xgb9/9Lxk7GVb3wQXb/BLs9YPoHDnWPa81Y6wdlyCXGyLo4lzrCjdUG5Eee+X3Jy
pj0iHDLnu/+Uv3MBZVlnhWOig3s/mHqp04cS/DrDu3Cxm3mBuErz87l1L3d37pOG
iOjzGe7fV40znCHu6CLuKZzbG+4OP2J6Qa4q3oa4XAeBZUznBjF63ymd41iXsQvw
phYYK691vl1GOxw8KwWa9zqTTk2E4AcloBaUi4v7IckXPDYXbXbL+6AETwwGYHsU
R21a3njKWVfVYl+t34R76EkkdhrWBn7ACl4ORtzk9HZIIWNVdyPesn7an9xVc6HL
PUe7exyjMexelr/x2BHfOXTBey8INeoh4yqzzz8c+9vWwX/f80yi/7WDyaT9pWbN
X/42AG0GmX7AVaKWmk2O7QvysuCW4rpgCC7VXTQi1RRd1Lh6Ol3WNS5wwCVhMUT3
xNTytT+ZQjUwRn/6DRi8BzS8Yu7dZTkJRTrl1k00zwoUTpFRP+YLdYY9rphJBO07
JkINapJGGxWHiQ2W05/K3olp2RBrMK1nPRKWcoiHyjsXOg+82jaUL2wzkX8qeExk
V1uN91rdIAuHXCqf79vGIJobcmC8r96X8rzj0VxHy16e2TKV6SDjkF0nzHBxf/jt
DrMrh38Lhhbag4oy9Q+t/OtjaksAvkHSKrgiZ63q/yg4lCZo0iYm4QYKUXQvThJV
NlpozHUsF6mvsD9gAdmKYSE0wNajv8tfVBlIY9rqlavBxrjuZvguhTv4uxS+WO/R
yDmbEK8dcPtyQWiTK0we3Es1pUopXnvi7z/pQQA7TjeMSEjItVvRrkN1bzrz1vk0
aw2hl1zaBhjgH7tgWmxvIBi44g6ScXQL9DQqG7gUywBQdF70MhcDOvvhd0jgTqUz
fZ3PkADJHhjxtPct/v7K719QDwNCWEBIZ01tportogjEielY10c7qpWbk6PPcGoA
HQTDLvZa7CtolOBrDAQREaR5XDuGYZQpgKZ+MCaXgdmJkmxS4j6jfxjX9vm8lJOX
2KUSPFRSw6g9uayN2ENU2x3N307iHs498zGzgixzNCdOlh8bTx9AhXclAYAzWDYb
usIdkadYKzFKuh3oPBWZCXoE+oYBuGb19UbfSfLrNoSwHO0R+aC8iaLGXjoF1TI5
29aOyZBmiaSVqBeuL/dio4X3pduSHXb6vkV4yTj1ooJwCSY2wmNKJvYUWm82V7BP
cyG8Unhfdh58TZk8JGlo9gNVSGG1d53JDxcL3KKZqjPLgRdo86vzRb3ijAPC9u1t
6cgrqWNtMf8YSE9ulTihvjsHLdi09gPAQ8eDg2b+z4QverJNbUK7v2kv9lVFFgyX
RVXE2jcCHJIE6nIj3EDzyWVudrngDzswZO5UiXXjz+i/CaIjdq74G9JHd0vwmNt2
8TG9MGBfBnKZMiHZDwQTkq5V+Qd5CPOXk4MPivxdiEBp+4cWI1ILtK1MsVlSJDqV
w7U7Xyog+SzmI1CoT1aRbq4weLAtAHQq/+9ZnlSgJlmTDUYM/sY6BwqnRPnO0DGM
oy3tFCPB3AO+b7PHIzXXXItVpIf2/bE5fQNaeEmYqJ3dvha6adl+hOWojU76s6EX
8JYLWxueX+/CaRoSrikrOO9WGkK5BBhbZ503iOhlnqTw3OYae2s1VHH1L+arXVOW
P4ha1WRhG0XmSw1/1B4LPY+w1TvGEvnQqKWL4TScyhzkpp92Nqhwe0xtYUHIiWkT
cYOOgOol88grq8Rrjp4+BkK5DQ5M2D7x6st1gtfqjwkkuae0Jqxo3Od7iTwXijmA
PYoYGVo08rRavrgy6qKSzoA97RnEZS4v+uYXYZel+/0aBFcBKklMNpDFySkNH/4u
o81hFAxSIXAbgNkyxgMF88EI8rvzL5bGhsDe9G5Y6n2tT4XDEGUjKtm/BqJHthAw
XFCZdl+nNhLnXJ4VkWNlsZJvkh8Zc++91/+amGfJb1lb/H65M8fIEQaAPtWtbAlf
Czd9daTNPAy7YFto0FEsg8UnLxaNO+EpQydVQv1JeANtGmkB2Ur38USm/OmwUrPu
nzkXas+W79hU1sJYo6/nZ+Qc6zzJhWnOXRxQQI5DCEcbmRAWFGIevtTiNT65OEsE
zYe16UabqXvnxd6zKABTB0Uac1H8R/4Ul0lQlHCOzOWxcKhTNkTgtVDgs4XGKcm1
PwTqHSuVsuCTgEwKWaW2GHB/XytCulb8efT6L1qlDz61hWoMx6UNHdqnu/p9DcKm
uE7NifhGb704hujFfqG2r87rvS7rlHjRwJ2kWcIwQJNf5F95oD2MN3PjuWpRwLUg
vtvZ7q/XCNmnHsHtsSEU3NT/fSKnth1Uor7bEq5iIPXGxIl4w5kanNmGpj6EC+O/
MbRWizVG/9ulmKPZQjfhQ7Y1KTMc83mySznKE1B2QnZqi5QiNqXT719zmAvR9J5z
PqENA91JjXO0ns41USW9oLxdkPDo33IBAyOwkARVs8kUbKR5+/a4QT8rfsZLhel/
hSPc7QcjrZNes6Kb/6r0kZ+Ze22P4J9FZxaWEVFgn2AxcE+J/kzBW7CWMV4d9muL
h58b7gwAiqanCjrgTWKrlkFbt4SpjCSBDVhji2LtkI4Ek+SinKDIl4zwFF50WgnF
dikil8pNLTwopbZwGcn/5b8qDPuSglfxk+vwGeg/XXjwvFLCRAaUIoZ4tZ/pLJmZ
qnq+LxBB50WKV3OIzvziPnVfCn3LAIbKnmX+IAntxla+uaXv4xV1g7Q0jfxg+4HH
I4+4s2dIgcikXF+YZALkQ5TNnCyIEMgB76iSSPoQyZwFUjwUIwVSDo5OqD6Ps0S3
iYc4Po+baJgto03Sr+w2ywaVtR5pr9HITBUS1uodOY657A5lkeyzwmv1SlYAgCjV
BxmLmsWi9Hp6GJsuc2lwS20PZQP+wOdYGS/NBXKJpIhJkKGOx1lAL6M7rMXCh/Ey
mSY9FgOFJyx/rjKWzqu6huROBDC0VaSkI1piD2sAcmdQNHfCvFwBHmOmjzUgDlJX
khd1nnNzdiP/l4kYCHrCCiNgjGBAJsl8J+9Olc8c5hS4a78nZLq/eQjtkCu6v/m+
1RAriyjm59hSCNq9GsTqJ1XGbPLHfrjDLbiBDSSg8t2Jgwy1oB16RdVLBrZhCbi+
5bKx7kOACHf9BK+jrUBj2CZ0I57IYPWY3DDz/g0fCu9GYw86h4QOAgVK01dIGbMP
u9l8tX/gQ3+b0XuVNiL28HV93kP1EL3VUkmydyPDtpwciUtgQhCgD6mYmuYCzFho
oHiNmNayiiZbOR9eMUrZEJ9Uz8KvDgCcj8mtdil+B9jk42/UqFEcPfV06ANLtPXU
ehdl+DTgWVfMdJrHA5Huj+cce+L4JUQ9RIYmjIHWJYSDzN5Jn0QkYxTH/aFmrTOA
7Nt5fIu0oR7uGL2mSi8V0vh6A8Jo+lZp9x/dLcOxvvFup2F77CQsmWcAMVNVg1AL
g7yeAwlJzczmyQAX8LUU5wcBhUtWuOiIuI5lTfBa5fxUtIXZrg7mlhYShLnOqyn4
Db/CXOVbvNjhFlvV10FKxvyE7MiOLsg3uLLJWXm97XdABsW+wLlVnKNnFD3/vfGD
HFI/V0DXzGxRERWpz21R9Rdw4yR1kPYFObYA9OPt5dz+f1j6FHH4SlIpMthZTcJq
RKd1OBREzx+GsAIMiPK3tzTW8aKkfbM5DeKx7npSMM+/i585puyLA0yazEpC5EhJ
RU1/A+Mk+slkHQbVrQvBDiLX2kr5XQC6fZtuQ8kVV0Br4aBYyVzh0ezFL972ChbT
wUnvrIIclW8ypwPRRD3bv7Ntl+bOfUtIy6xIuH94TYeEwEcThrNMU8N+LyoMkuae
x2N4CabnNsVAgLmhHqSvXDjBYPzxXJN1gbFw8UaoTu4GbcBJwQMScJZRiPOXo8+3
0yIrD52kZEc5ZQ9sZB62KmuSCuG7+3BePfNf+H/b84PZ5eOllHTnRueqo+o7WE5B
W9Vr41LDW5DZAeXJE5wKyBfv8z9r1xeGJ/pbk5yzJuy0JvCv8wk88Vwjtty2Yuvk
VByb4QZaoz9CPSbo174eH63aZmVvX00kDBMMoKP506fDcVAL7mgWPAdVnL9jKor4
E15YHnRdQoWccF5avcSS6DdOV5v2hdC+U9fa+NAQJzPsurGbOdmcwK7F6njh8qQO
uED88tYSclZ4eJRVPIFJFvQIufkQJC9AumjxwYkMrrWa7oELM3erm+uoNelE1puq
9kjluyLfkc3ZAWlO0blw98/FMCln208xy3oWsR/SPgmBozOXQs0QgWZENOLu+0hS
x/yqbsaophV6UDJ4tWmr7+1ICdC6bxvboiIaBnmAEYpuGMc4Tuy6qXVGKgHsljmb
bIAepCxVSoKsrX5XtJPz/J7xEgVmz3EI0xSpl3p2R2KGXPS77Q3voMJS/s3B3Rdn
RMycdbvcawpVpDenTEXo7nTVn9noTGsYQV2MmiIsUVYFB41tVxqNqNhEkoUlzHph
JMVFmql+BQ+g/r/IWD6504EV+g3YYfDwczx9xQX1sA8a9cUT+nQZeD44RIYwFYGW
N+cuRODkxZxAGWqd93rs8Wh7j3kehrcjwG4vtdaJutxhEjfVNahTQiSxNG/3zFSh
exCKXF/hj9I012L1v8OFocs9gvQBGNcnrUP4rbHsb9079nlHx9Vw18hpvqAPJhSv
Y2gCYhsm4+0bWs7RtD/8qWbvRlBaYQf/SUmOksuKdjaq6MELvrONiEtsEsbTJ2Rq
XgsL4woUkVbXxjv72zS1ORGEAzIdxUrQzbAw7zPPGpwT08BlY7pkJbrOehBTo3oM
8+Bww/JfNZwVIsYCSFIdBCpCjUUAzh0Z5T+6VOoeGMe182Vk03tHPF+ECwY9GpMm
yaOP4lwzasIyvZtP/7JtmP1kkWIiT4Q8SxRwuxjnwGJYl1rb0jlBE4Vu/EFb/wr0
yk516FIME6x6akJLyetkSX03DzU8eYXzRFXho58p78u24L5AO+Lu2dWC+EDUGx6M
MASuAnLPFPkBiFGbDvtvEAkyHPmEl3upu7MBZ2CJ84vSCTkAPXE2e0Loe7oCej7t
lKV+DvdNfP3q7f7+3ElLAO4W0ovtqmIjraeU7lMy3G94TTWQnVROtn+GRE5ztbtq
znApY1GAc6JIyNtvcgyfyVWPpsm8Q7VeW4qTa8ssEzm0zOsS3yFYjpfInk+gx/tn
8pnNVmLtQAhPYdGCG/KP8yCWwdM75bFDEeAa2g0mXDl3uWBTgBLej+caw+JCnfGQ
uscyfRa9Qd21miOQZV7SsFXnsmioBBnhF6IW50WrM9cS3GhF67sl8sUb2wulk8bT
SUMLhWBl8IhGdW4kCvwwk42d881uZFrVJBrIZafLPRUBPgAGzh/vnrqxXUPExkQo
jKGxm13QeOROsqm8QFGa9CI9hkUgRHSAgumgqOycSAkO4ne5NDjhldiE1G6juSlD
9doJs4zJxy9qrZLTRtwm1/8e0KOh94TV9fJ6SLhoKM4TErSVgzIFZypG5u+ngUce
KjNObs5qfwRlKyLhI4SDMEbzaioQCsF42D8L9xNHy/U2lai1/AwlmsyCA3NK/fO5
NC06qNSvHs4w2SHegIpCwiTcoPEMblgEeeHbEP55K4a+wRFufeJcsCSZYTAxKeYh
5bCg+MZKXII0Awe8TMETdlHyzZ7Q4Ut4n06qeY8D9O8A9h54IasKdkHJBDsO7K80
22jDlTSIAu80HJgUKj4H5/PByaI8YamFcTeN2qEDF6vhJC/qWM6yqYyLQVIfUxGd
OlRl53YmJst28k8uJRpheg2eMhkarmG+x8Okow4UHZIU7ZB1mTnY5dIYSXDITgL7
z2MVp58l07BEmxZ6RDaz3XUw9+QMv7nvdqaCPeWkZRj2W/FTdAa52mDWz8lq0wBQ
6vZrBS7DtwtprZcR0p8mmrkeBpo9pT/beHett8SX4tr9uoK+BlWf17kvjT08KqZO
z3H24WIoSoB1qwdB7juHqmWQHbf89wrqK7nNpY6KlQLLZHglo+vjYN0rsb8CQwty
+26J4XDT6M8N9IwP5u+HoTEgDyMDN/HSAokbXp+sNEAfPRTeyu7HNXBqmcJHWcJc
GLzUVazH9ToLHyyKnLWP+4FvwZtLUW4WXTFXGgFI/dgCndUZuVabS3PRkhEyG4T7
ZoxNvXhobpcwAxSJ/DRYP15JI6EMXIBWsMlGbMY4ijLIiEe72nnnq97LUyQsBUGa
AcXL7b5rYJAJmuAKrSzTS3WirICA07D5fxO6upYZa348ncrcu44vlobCM3KdgF+i
BH6ryU0Uk2aX9T/h/j5Jkm/gYy/BP1EMpmWS3dhrrMreJA63IeGNxIYhknrJXUQ4
Vocwefclfzhag9zmGc8NqyPvN+1Y2z82vYmTqUEHTRbIQTJK3mm2PVMYfcs5Akeo
IFqmI6mnqxbcT5HFQKVTY42dMVmIXDSpXhwgJaKNbU+U0TlddT0+tbz7dogjWMz/
gWVFGvG+zGqnZTqoGsCSl22pGe1M1BQTnQhdpGpu00cN5HRz9HBIgx5XImE6LYcd
/hJXHa52jaixYSIDUp2qZOZ2g1hjGF87R4Da7kAa2PX81hQgmMIOIGWPvENB4uLY
BrYTmWTHZhqY4583aRltLUqcWuiOBRbFDRw8BmWVf6B1Ea4JOF79dUJ3IZQVbVUp
XU/srBiXpZckYHumKj6S9HcihBSTSJ67yzNQDcPsmOmu76YXXXi0fYdCkEpsFAsf
atX3ovRRYV357kqYwyYpDuvWwgFnPeu/AJoU/lksQRGvkVFbvNWra9gxhNLDFng6
KdpO7HJ41l8Y8sSjGubPf7+W4yJaoLOs4htPAgjGE4YH35yFmq8K1N1cmCiMuZGD
f+PcLHOsCcptrJKwAAcncCbNkHU/60CIv8qQuGh1B429iv4F/2MHWPoly+TIJGf4
a1Ip0yc7YQvngPO4vIMMgtRjFUuuPXyCNEkSORronIVxBEFMnx6r5vCq+2LQOtZF
A7WmTKhA1T6vktsxhly18i5ez0mVSAAmCXPXCW1I9jLHxCBKR+GCdPrW/tdYu530
2R6dKl7QtIWdb/NjlrppB8XQbyVmndWZP5aeYKKR98M0imazbhS0PlRDUovbzbC9
ksUNrRaqrvPcUOAK/u8qHXqhRpOpuOSoANg9rspysyC2oC8glyPYS3ieNR4afSKO
JPFRyGJQKFw+pYYfeMiykA/Nt7KUjTQqpTQKNS+LHE5Tnvgw/9Ni/yxB1frlCxxH
Knd3YJNlWHsXBUkhVMvxkQVd/5bcTA39+MhgKWmkEtRl49jyafi95W3Z4CKL1OXK
5xLN6IAkBIxydrnRDBKN0IkNcxzn86Rlv6SW1IFtL6VTZBKYsiRfwPvA/tIH8jYX
YfOILwtn5BiGlXhBBnS9QG6+jKWvs5BHoT93OSeWecB8HQz1Hr4WTSva2kGj6BZG
r43PTfcwNXcUUohZqk5OXlTUzY7oZptrl4dGcJU2mGzqOGoyh+5EKRJ3VR6ksGOy
LZrwEpKfn9grONBbjRgK2N7jVPJF1Jih79vqzqLAn1mVGsblMH9G1u6xd8Svih4Z
FtTWofhNNvP3Q1Jqj8bk5anmnCF4jy5GbR99vAWhfUx0980O1G+DO/ZqVryVwpQ7
w6llxWZFZEr+Rj+TTtv+cHRVaWEFkj0yECbBwW9lsQZ0EXvwCmsvoUa/szNPYFeT
J9CuDlkyIq1+UDYDCODs3IyFD1lSOBo4F96D9Zsi0Vxf2Pu+xnoLHyGMSC542uch
vWNY8/FqNbC3orNvnitMlw/lVqqzwA22s/vyoCC7w9XJZ9VkCkuaTYyiwT6B+ff1
ko/b7viv9PDaZ1cdyyGPi3PC3Egv5ZBmHmfnw6vrZi0q5Fj6R8lDXti715gmys24
35eoceWZHDi5cVxduhiIH5mk0BP3kTnBRg+HuyjjDXL8/IMXuDdNvlTwS70AS1pD
hkD0udkBNDZ2nVF45gdI+JMfrGmAc6Js5+dqxePOMLMO3sN2WtFYWHCwM59nd1XP
OwvTk3PiqX6/65xwJyp/hlLMEIwS/jn5h+sNS3bDwUwwCRKPaA0oHvAaEOUkaPQd
JHXA30RASzbfxNywfyAoq4+fkU1sE6OJPBjdlIxwy4/BdM8avwOFGkrtiLIDqCwh
UnBjNGtK32DMAckbaZxAk3YyVtS2tDMCBAmS4OgB1jR850KPY8t1jxfLziwTjWLE
2uAs328psST1bmZRbGCIhh+Lk0z6VPvbdPe/oYoMZUC+Eeqf09k3iO1/AojbfCtE
BD3RRXk43QgcKrdx+sz4JI4eFw9NGZOo/auih+mjQCwVkZCmT/gZ8mymkUWP+yOV
E/B8KYsvpfs/rRXnk65fk/rR7tJaBDv5GzVDFAyWX4TgAIaMKMMmqhJ6iBxmK96L
DNyn66U2mDrqDisZtCi2vF54oLhQlCOgTsXMVO3mmRSpuTaTtOSL6MC9fqwfBlBO
aP6BhUflPs1FCrvWX0MuthlNLLJfGvS7EcdFBQ2rC8h99sKzF0q3YLA2+MX8to4k
7afQAaREU2tU6X1SdApOt/mxnAAQpAmmLskbenLDYKP49uj79zpe3O7RaUTkeSQp
nwPyoBCElHyyZSDtcDy0YIEJmgmBz2Y0lOBHObGfus3cdouUcN6w123VC49hNlq8
P4jfmoBoPnaJLvfsHqqKdqQgGIdK5QxedV24UZ235bIIMtFr5Fz0O01KNjG7RUX9
5auOTj291/oU/Ojs3IMfCEBYJqjsN0pU7G6a/8SrS48ehGqIx/jGQMEzW40q48SD
mjzciI2WUZKp+Xi15OfFRQirJ+yjtOe8IQQGL0HHHOEkb4v+dWkv4M/1YJVX59tO
sx6P9Ehv9whJ373p1SvobmZLwq9IDncp3ztpm8AxK3RvfVmh2oJaCNteqWKucBxd
Mrr0JOJ4Orra213lqsFkfLPvrIAmtJ5S+0BdzCPjCW2ymoTg4aKHWewKPTMlDI+m
IKzXJdfYsm+XBzD/Sh54u6m4HTN59RF5GYQ3hoPwSBR/f2QOZYxzXKl6WrfMXS6d
L6BUr/K/hkbFpsyS0um8DmkTl99EULXlriouPwda42IjxtiIQ1uxIKWtbuP2Yh9D
A1XVXGFwyQcfK9lnHeQSfU8Hvu7EaOxigSqszim4b7RaWVveIAHdito9qVLizUac
Rg6APXOkRRqnHYDYD8EOJsMFcktpvPfyXl3nrk559jzMUC+oYx2ehXorHQkXQ0TQ
0Y/5MIFFe991wkeI3OIREqiqgLiotquznv0tmMRdB2y39VFnaYFkDqFOspLiRmLz
8b8R53YcYELWdcQwYcZBsrsRgHZpqjskstTXLQNKjEYI8QrS45V+aj683cI3CX5f
uBxaSUifxiLmICbWxv3cfbbt6Z7QGih583VSqu0gWbJOq01UNPSD9EkeRzBJUSNa
T57irS3rPlShwKwmkoXJqMFgLxOf+MSnWvGEtK4aCK3l1Vb9mD5FiKC2Cm80go6Q
DN4geG+ahLwdCthxLlz9tSD2We5ZxZSTk7BHiBZ+JPnltqamztjb8/AIM1A8oweN
41UW8/uiep87D1e5kcKkEUhcgzH2E9BMZfJMafCITT3vTn5EhfbZhkZEIiaN9qUg
wfrok8vvOgP3bnuQYr646MNXtGK0K3DJqXGqQzxdPlpqpR2wVf29/RITgCL5yqI4
fblIt8Sx/hyOOgM4Zb/65EHmjAeCuMQ0gwz1QVeOf7yk+qktGLppNr9RgZvLKm2D
E/GZfsD5H3WABqdtSXoubnkmKnhKm5DSfNw87sniYlUGyomxJ0x2ZM09ySko2u0H
SZjWGNJgZqDrSq/q3ieQwtpDgmVZZ3Gb8jnpCNHmbWZ1AQJ/UJAm6khSH9FDhOCq
JbWzqaIX9XRopYnnujy5bzqq02ODDgOwWnWUUB1hrCow9WE440QOCYvtnCOnmBDf
4m8frRQXe0Kt3BEjGxLzsrg8WLXTetTykV7T0loGpVEqNEDGPQdbQlb8YXlze48F
O41CTefq0+l5FHAPwh5sPvXwRtQOH38c7x01+zUT7wwRul1P4WvM9YhlX2aewMwB
CaRx9hgt3z4JrLt4tDlApIqqnxpTmhJuHAj5+5dh4oSrneYOU3W3E+lHK9wifKZD
EASmp21S/btV+CnMzH6jtsGFP5qyKts+LzHNiDlFRsWNjmUT7bhGP+6m9g9p8YK5
G8W+rKWlr0RJ/vA9ZlulRs81e1t7vXMCXMsnRuTRvnEin1oB3UC06e0pBa+m83zs
+jC36+PoafjRU8+TOjf5U14Hq6g6Fkg7Kk9hm64tlhbFBAy1w7mxfSxhWd/NoWhC
ubv0FHncAFN4LduZuoiMpAH6GlGkeozrUfLxx18ES98hvEOM7VJiT5GD3j2WPyhz
9fduNt0zk/3m0IQDmY5I2udWKDi+OwwS2ubDGSfphvIKDCTXmr1SHmaAthIozTlO
HyIrQsxyrlygUqNedGIck60rcb563cs1yAEtFXq0kROZ6qud0UBVQ577BvmgMZfj
0Vfsf6qj/nM/CH4KFL2OKiKDfXm0CR5Zg6M5g4J1BHOH/YMV1snnRpy/+cBVfVYb
mBWBypTMXu3QcgqVkWQx925Y5WsJt5P/mCAdqynYDlp2LTR5ikG8JvBBYH+aHhH1
VFP0le5qemrqy+fKrqZSY5HjvH4h0If58Xl25PdW8FUYomnuQ7HAhmvShJNIxsyT
Rf+cCJ2p0O8qdavsfiImFLV2yGFBL4v73FUyt4amnyN8S3nh2iHwPfIEmjkl6lmq
lEPwhvCz7BEEAYYkRjhnTSDSpq4JDKppTUKQZorjYyhKI3JFJvIqiC2avCO/RM81
4ziZa5f1N8sGB0RcfkP8BLHYjvaHV9gGp8t07GNRff2UAmy7z4fr5toCgOE8dIQx
FV/+KRmRe+3wmxPdNTWbLDnfv16Gyaqj5hzygpd2rb2RBVsIiYWys2KNx+hNshVY
UY6o9NAoIomcBPJYEtK0AFmN9pStS5jLIZJA9M9ETnquah/o3XdZey/dtHTxo7PY
8qL45y3JoqQ4Nix+Bz1PxXUATnfp7RU563WsTz98HUUx3g196VKSHnUUHuLEnKUv
sq+qP4FqZ2mafI2XAq0r+4iQ0mVCmm5LQvHGJ3rhswcWq24+OvcUQhWeDARaOBl5
cXAPmFgWzxhppI86g7y9SAJLuZukOnL0innXXO+dxLea76XRMxp6Me5cdV+m50tW
cMV3jNibQPmT87CSOmd5TTGHnjYy4k3SSBEmvH2623Xd38SbgZ2xGX/B2IH9+jKC
zcuoqNr/fua/e86pmaeSYISJ6V101XdmenDelPPT4SuC5XMYT57yG8FfvvdR1w1D
ajH5oXnC4J6ImMxqTJIF/UU0ccJm5ichHbTA0PvoqLJ9arD9Rgh52sJaiGp5wj1m
k5ZwH89+FEg6BFD75lqioQs1OoaUrDJGpZEDzkkwNX7ZnJAsFCtWIuzaVRr7mKHy
+Oeul7fpZUoSlExWpki3QgENamICqQ7PqzIVfvQMVtzEsGI57j/42+caSYE1zqG+
SHYNE1MpEYo5rcNXf0U9y7marRL2qVf3E6b2SiaguKTNLZRFILui3NqzRJtnErIF
p8XJ0HHndcWrW6mVFmsdq+C7M5l0WPh70Yx7cAMYZRELNHaflnt3KOdPsqvKaJuJ
nraoV5GZdD5jShX/Y4+KD8DRG73PtluTpYXqXaw2IPN7gOZ1BEfnpP31SHT3t0uw
Wv9DC/D3H7aj5FmBoONjUNW1GqhpPW4XsNAMM071zkV5oDNLZ++FExXtWAPw7+8b
q+i1ZMGDTckOSwuB5QdkPHi8NqKVHLyaYWPTBTQxfSVnDMghZpHWVw+lvurFBd6p
GFhpRJ47xcbCXhXTUA2Ru29KpRpqEo481PpjGkWUoCQc+XjNB6CQJuEPjoKtaGWJ
CMrmP3x8Xx0UUxpmwxyyun/PpHEhyFzjk7WZKT+hb5fRBfag/8YnT15cXYPop8+w
tei+R/OWJ28MSGCsYGEQjHLVTlp/prmauUg0o17EEdVW9hFFyI8DY6/shIYTLipV
dWCXW42poiE5bFVmOBJ8YmmmpPo/F0PyxVWTda++kfz6OqU6TqJ3A/Y0ae0kzRpC
c9x4YPdMuv/mTpYaYQl6+Yw2Wmd03Ua/DjNHs4Pz987W3avJRkUiQYuUcZ3wXiAF
XyBpyX2jmKVJkX7LYpbdnIA9zAQdyBkKi16MEPixmD04pS7F0yUFgxDGdcceupZX
vqnTRSwhTNRioMEmkOApl9bM6w0LwsiFowhEsEW9z1Pn2LANH6Cw/G4fG9OJ5yKb
RS4qoUcy17l4NzJHvUi5cK8eMcq4OIlqh8q3uBgeYUOZmVH0oOKpncZMNPbcaAeJ
B5tvVzHwcDUPH7Ys7ujugMTzF+6j0DVSHPp/NJq+2AXDUWr4vZmjkhpIBFBScNeO
7M4l3imIOWmNRwjgGsLDLRIw7c5yVgSCtNNCErynfGUDxA7mga3EjNFwr61TbNVZ
5Rp2/kpkmU/QkYMs9nyaw+TbucY3oQvbzLBmyVOqUBWGsfnegA+L+K7EmYuGYc+M
4B4KfsnGrcHQsZJiR2AHhTjOvW+DESYi2N93Cu6X+Q0oppmAsQSkcWImo9UHPm/Y
0aomd3feKBxfFKu1f7W5aL+PyF9r8kZ9puOL5mlF/6kfhp8w8LiMbEzzen9DDPK0
Gj/cWe9Gpxs7j9meNTv2y9m7cDyU2dLvcsNQ/XdeY5DdYeR5Ge2BAaahyDo5vJ3T
khXTSSkPklW7Oi3mYRGGujJa8B2E7C3rLJF1uH6KeYtfEPXl8vnWUL93LLa5eRze
YdCjuw8vMG5DEpXk+8u1koN1JYCWpxzH/BL18gWQQOtvIm/LmPvpkpzPSdqAM8F6
qeooS8m/w5RZ1CtDAJ+1HweCfqGfkaPuY94WTr/TWPq9QhzhIYsn1Htp4xObT8sR
78WC6kxvc92Cxm2AhgIk1a9JOPzfpBoZgGFDtl5shEXX+BYY0+/Pce8Xt/NlKK3h
NB0e/MYfn8LFX+GJr8uW1eHMNje8JNW/U7BU9lia3LMs4Y47+XbgNv+bI9L+thBK
054BTVnvZlbG49HNmuRQJ0MtyzrNObFaGKTgzYuc8bXRGZMhgJF+yBc0uSwKSy49
ZLEV4qS3nWSs86Rxt00hYfWqC+yvn5ebTRF8P9xLkAE3wbWm5hpOWvYsgzgGg/SW
lc7Zo7sLTM8IAdNYw8eVTLUKrWJiZ+WtUASlNT2AQhHGW2gyTTvuvwlkITw3crjB
5I9u6rI7jkHhMOm2KVeEHmJOntk/SR8S5eJdYXi8fuHuN5/8E5QPuKLkuUwsChib
KzL5OsZgJ+l617t1EP37tlSEbIZxViU5St8CBTKBFEq+46OfkjZAVqHiWMUedPiy
Ah0Egp5PkpRMDykHMYN2GYkswlLjptz+ZaGQlH1URxFIY/P2iYbsXXpAnIJevh+A
RHjUwcjaJGJKb1Ec+gvD0c5OPlSb+mJh0Q4dbg/GdzqxqGUTC/ksZ5qgE1djcVMa
m5WKfepvt5wKXT27WyBjJFiIs4JI/ZFsYKrTYxEhSuRzuzoXTxP9c+4tRwzncp6x
oNwKhLFKpbOvPrGdJmPyU7WTKvFMq/jaeegHo48j5u7pYbUHE8yOPZ9M/3Nvc3TU
SQEIYttKP6tP4bmBNE3XbVQ9hWeOv8L3HXyHsifH/Mp5qgPrU6uY3cyW8gTOIaNI
n6N7m5hTowXJ9QA9b17jfyN18tPH1rNEFsI89ji9t78KYz4Kf5Fpc6KOZygUDuyo
zut3J/3G+mcprTgCxr9qm5/wchofk0ZiEBHWMBhD/RRoQi5Gr3BY+/wwna8iHg8L
JwhkJYF76PBfTyMJqb+ZyjaO0VfFex7x0NHa8cWYyhO9CNTu03O0/ZV6dlJgHehJ
h+qpHNIXaHgiu4VauVOTlgOLWAJWBbQWn8b2KxiQLW1BQvk6jy9F08q7FnNumN86
j/S0syh+ViXR8zwaoPBaUIPeNVPuxSm+1SeKilIaGnBP3bXZjAdbE2zeDaliAVSD
Eia9LtAFU9T0wMbznu2xb7ZUzgd3uX45Jgu0kdZYXMgCJzbkYfo7MLMCvHCgE43I
/FsCcqCNsdBNY+aPbw+t9ZafDWTdgjq8LYC6SfqCGPI8GR2drlgMYqBkQGuIIM3l
zh4bJm8oIJ5+W+l0Cj5GJi5gX3pJVAjYL0A5XrsuGMDyeJ6OoZVZFeWEqKFPO8eS
TKM+zOsDL7MA4Ok0ocDLCbtPH1m97Cwz+6sG8lzl6zwdXg0vMTl5dTo9A3v/GQpH
xlBi0N0U/GVF2pVZd7+NekxiRNlgCaONqhX5VRyXbYNTEfvRvJurBzBIirff7imB
kHFKtiZ4jDDyuhNiJje78Ra6xkvaZqsF6KCJbxdvPmazt+gYMAO1ZQIEsMJMqLA1
wLCwPJOTDsJetFvFDvR9qEnZ3OX80TPvtuWOW+ialOCzCwocrI4mNyVE+Y0Cy2/E
CtVQ0ZuCV2cgAaCs1z8YPs0CVgNbQ4QmGqKuAK8uPotwptNOXrwXQ4YQ99SFbH9y
mu8KNR44ix4m6IZxr0+8497dUqbnCHJAxBScXLotntFeYQtKav+v+mGC4K2icvBc
VJFz+kKYmvzopKXut1OdV0srjVWJnWwvSlqDihPUYh5ln273W5E2M3YrX8h/sCm9
sdFw1mWSWnEjRo2dS9Hi9fRfBTB/GTbAv6gbFOOWkGeXjUhArdaAIXUwVvE2R0ze
BW9TaqHRzdM7w3Mk7jgExMcBg4fT0dTOLl31IJIWDdcp6y+T8Aob/moI4Xm5p3yo
xtlxLu+4/oL88wpMuls0KEUHlzLvDGySmqJonU7+sj9jzb0zoI0RmgMkHFHJbqtY
RCOMVc9CLrPV75Cm+w6LOVCr5pRL3mww5pjY/7xfrt8ywFyMwmQ3dLFuP/wpUQW5
2MwW7AbUzXZgVjflHnUE81lnMOldeCGiKBzJBaDXUa+JUx295gtzMiOk6TIPGXak
NC9BJxMRszDwQzWN05OeFshhgvQzRwzq9t+IPoIMqnwTP+t1OUduqWwyl+8LGh5J
eXoVlZXdDCjRxBpic64gaL6rfvbUsLnveHHtnEA6066VRTwm7n7Luw7e4rhWtK7T
CBlxhWuy26XNGv8+bCv1xCcDQ0WeIdEQCzyEnbyjq5oqBp8AyrJ6S1MecjRVKUM3
G3384D8T1EfwbmVlJGBuwRxad9tA4T6+DYt+vtUa7YQjx6yQteszcBkNmWHrZmf2
anYa01uqf7ERDeanJaUTwG0RgVdOYv8OvRrpbns2KocfHg94HIYCsunptJUy3iAe
0GiaVpM8AtgGTYO10ivMd4Wc6gQgshBo+HVpd70Jn1lRIq34xoVsOl5vDKbMmXw7
q2YGUcCqSn8VcHLGs4sCjiRBATPkFdf3+0ea6h0KcaWlawjfo7PcjfogY9jZH+/q
DzW1Jvs7ctQ8TqaoL2xNbyIhRrXDu1kPP+HEx3GeSKnGh+zpi/DVKnCpaoV/kOb/
XWREmtZj3U6HS8X6KyXEZcU8aPP/ThntaMy//+Ew4G5BLfCX0280yJbWH4yIxdya
oOz89VxUendXKSyW0Pynrst819vWWz+aN087K7Egn1wetGacStW876NrZvRx+HbO
qeefJrLBtNn2wMHnDYv1r6UuR6TJPvrHQPOuRHQ6X2Vu7GCtCbhejvgxxTv30qN/
wg8kEtTKxsh7qHek5GLIZ+5hj7S4UNTu/roSWO3neLUNFwDGtT0G3QFbQmJAuAn/
6FQj5/OH/ra5wqutCLnRUlK6cqXQRSqpwDmtP+uszrKeMoBrNnIXM4wrhusIwFWy
wKoXw14g7lBBU98AaYMKg1wUlRf1N6ikdjU5CDGreBZ+nG49ksaiqMg+0u2Qctqn
Yz80S9jFJtV1VlyetJuhvshqLVLWfHx1/SAmDTqUoJxx1NnoiC++kaTpjFYv6HI1
aZbXEpDwIAsX5dY+pghOzp89mP2y+NsuB10j4fppYkPj5CjzIeLWgvo4EXvYzajY
z9+xT8jfwhsjRskSQPZN0IyNSDUqfZHPHGgDCXpsDiIu+iyetoBR1mPYgX2y9tbh
ZXsmrWjn3Wrico9w8dgxharW739eEc0mLyyjEgzRxMLR7NHhnHV6N/uVjOXVYw5D
Yf5Nb9hUq1Fg2IEfnmp/VmoJbpX2+Ml8iNWzR50/YhwkPwky3QS6UAN6CHWqSfE0
Q4dz0fY4gzXTpoD4U++cBKJRSKC3A7ugFti/Ph5bRSoGaewQ7q8XPyAcBGQDPXT0
cUe6gamRItMYO84DYlAzS+wYIaZ458sr0+//fM31iJLREByq/ywdtuRpi2o7+lI7
U+Xb5NIpyuu+5cpuVE2+Kge3vmrMXP9LsXrlI4Y5w+5wtDigOST2kFXySMKC41vG
tnDf/HcMZB25k4bk5F9tv7dSyjjIjj/zFNwMHSibuwzTwuuMv+gecXKjuj2+tLJI
3zKyOHC5721Qp2+hOLdqscpC0nGdDlEvFfstfFACbmuXQQAgz+vO7MnEng0ObWtO
UnjBARSO+qLsE+FqwMzm5ual04JS4cL64Zo84g6PwCyX4RACAU/mh2ugzOCLEVEf
IIOSp/b/yo9riK4/VdgegOQUmiGNQki0Yj555A3abnlnQJaTFRiBdQjJvhYMsDy3
buLj9AEwCMVX8/EKvF13oFXaXUpvuZYpA7qXRfzAolH90yHZqVvBrjQ0+V5c+AcZ
Wcmo5HVtLrd34H7WUc/87X8NVhKGT+bCE6gwZyE5vSX1QJU6ftMn+jUv7jloa8YJ
Oa8xqiJwTQGSMwNQVemtjkossPQjAIlrqPqstFu/Tante5TEUk1nF6gnoNSxZQJc
8KdTWGvxPGz/3Lb1cJ4/q69XhYK78KD+/utuKZDSye+I8tkiDIFVHImD0fh67lA0
WwrNRJsrBUtzsZpLgqnqMP2aajl5xhVi3IlNcW7TnIqT2avsDBNst41L0dWTTPzG
Ez9w+cuSnLaKYYpVEH7gzDSsWWNvPJORCiiNB6hGwcZOLqcUdMrEh1y+nVGSn5NI
4VU9k0xSWaRUSJSLIJU9tfhnqEsRIV6Ox6eI1BsgGdn3riWfJQ8uRjEx+v87UhuO
lsjdh5ogDgrmCUXfQh8XNKuVChYDqrpegjn4mwis9TpZW8Pk1JfPpsNzxtii3vyG
7RVK3uXikpXnAM53dX0CP96cKvObSxae0UsC16p1b1LWj5+h40VOEp1mIM2lAoSt
gQNF+uGn9j5IElOef7x1hVNM81mB4ZdOsa9uxGgOH/ScriPBlJMyiSYxnj8DKj8a
dJZv3Ri8Lz19fJi+OcCt72MbUupn07Z71nD5ZtvMhdH9SUIWLuB9pEfudolywAIV
l3eJJL/70iCe/SbQWiWFJvK3tdB1IW81CtVrJsBXLiZMpK4L9MaTwJ949qpEXy0k
jyCSBjGRLWEGJvUomQOX7LH9ijyVFjFOygutGp0r44dxxJUKE3GxEKC7teCSC3m0
O5BkURZh5vsmXRkmjlahtnVp8jNrqtIp94AyEqZKGCECtrWA3RDRgx50IFFqoeY/
RzEx4BejeQLYZXsvRCBnD5ddnZv3i/KOqm97SxKMMUreMGWwdO9iLs8REXsw8I/E
2/W1iEOnB4Kkq31aMg6tncTOieNYSLzsCLmvn/GRAC/Kz1PKDCZBXXSEO8t1gemu
yffxeh7A/Qw1N3kJFv3SX44kqwvcK60s/aR3D4j5kXdCxNbz3mZn+dxOwFEm5qrC
2yrmrmoy9TynoCp4suBXIhLFwFgxglH/roaK/viOkR9lzvWj5eLCtirywwQjUJEK
RZvh3YtZwj7hIQxNY5Mus2bIVB3A2xXMBf/wkUFIz354w4EzcBBzd4LsWtxQum/W
KGJst+0VFFRGMU6kSlt/htJxTijJRBXd4mpjm1Si34i8CfVXs95sGHhYS8ckGKd0
esu68qgAMBCaRhK3pZ7OSiYl6NRYeNXvzS3BnJX14/G+Fjk70Xbwt5xTocz/H2k0
/dso7C+srlfZSfAQrAD3Q2j71VZ8SHeHwn5GKdG4ZDTDL9p8YF9D7YISdvM9XFgv
mKHf9CIQtuhrSHZMns0UN34N0c9zek9IAfyjTmpVDh+6VXK2MnQpa0/b2FGGDoxS
T6qRtpn46VVGrEL0sM4ZobvgkHSkLILGqnWsR56FDiB2CpF8QjUOM/x52D6E22UP
TXTzgljSVBdrdiGnEo/AtkHqqWGDsiAdmI9byQfxGu1Wi2BOP50uyCgKOzl4y53c
H3J0R87/9jsIwgCq+mzgOkkyN4uslVVk760a/NrghcTnxg6/1MX5vnK7RODrWzXC
VqAXpE4CehUm6GDhsGhIcC1peZaYrNEeUX1qHpygV5KoPgDMNWf4iE7JSI9/YL8B
ENSEmWMVKSaEjCPFVouj6QR+To4rbYjgdlXB38Eo+NLAHCdGpx3YKm7zWVLyR2HP
21cedDiywc+hrdLVrs3xkzqBKxKhWuMZmJDCN12Z0cYEL9s/qmUpJQAjWoifeBEr
/7gkqQJDP73lnkIfZ3Pu1kmY9j5RoejZNB6khwCDG7ONow0H9ybi47FtjebKq8VC
5A4/GteDCHN8BY8UGy83PKi7Uy+MKmRq6CqgcLC8Fi9YCoD+vY+vZ9rKMMbwxH8A
lWZWu8rTnEwZ9RtxGQx40icKqZ3shuSV6qiG5NIbNanoH6BnS3t+VChQqXfD5pwO
WKYNxjhh7QP+TF5fUa3je88StApVKcY5d00rL+FMh2Zl80y8wLsFQHtJdp6opKJ8
JAKrZ9o0w2M1+mjprlpBPFFh1cEjAt7X6zsg6f6K/y6fEaJjp89RGKKK9SB3tiaV
M86gMrhGhXkT4Tbcq3KZO023TFcEVaqkAWKrxbkinLDeS7vq+1hA9yG1zttXieix
vkmT9OsJrQJfkKM5mcHbVuobcOFpmY+noeTLMZQ+sn4m+4SBqRlcOfhen2nRpWhX
nYN6zxq1hDt7L5rDojxWVsEbZJP4kP39Cfj/P3kCeKKiy8BuQiVVxswwvE0DsW0L
Yc5rO948Ug0dT3mWHZwDZ58hSrmz941YHtTGVNcZSXvp+F+ZYnOOQS7XLldZE4zP
9ckIPEKPbQso/wgHCyZ1ra3qjWo3pHDw+YJ/wQ8IxmNE7r0OJSgg6UD3jb9z6I6U
prZc4wvt3DOILqzMY8mQLjlo7dxacvuCV7t2fNmtUMZxyLJ7ZIa0Cw8AdbzhdL5x
w13xtIKwQNFsKRlFLymW+EFBGOrLbLeG2fLmNdO/RGWqC9nFto2/UEj5s0cZT2xM
dEQ1ZNmhJN6Xuxe/e04l+Y/e1c81oqRNEqznbzrqyiWGxpJhvyR1CZbgzLyME8uT
1JofXDJ+pnHD1hr3IR1fd+OixZCT5BUPeRlqIERGZWQppKnZd7pwLayDcCgUiU1U
35SxlaQlKzMJGDcNOO+ns12pqJgljiP8vKRL588R0bEN+4LS5BcFJ9iw7VnzNOhV
6j2kvJkzVRLrohB1lQ5gAHFn1OIYRH+tXeRq7zoBXyS7G+UmzemfztUHMpCEFoSl
c0w/CeFkziydQ5JizGauvH4LJQIQ+ryB8frbFmDZh5Vt6NlEIDgBHHQ4KmQTFh9o
Mpxj+IrxbCHZcGonFcaB4ryJOp3Ge0UNGOTUKaqKG0U/+qhU9Bt3ZIF933TauBv4
+R+Xedo9RbAQfxx0C2IVNeGBk4DDWjzCxZtNnE2e+It/QIA9eKPMlrxI3h/5RPuF
YhD6dnX56Kq491joS0QvU80mex07RTTu8LOuKMxu6gxrVh8ZRqYMUC6aYZD5fd70
FWUo8kgPxGVTBa7yKmiyyTHwxDoqSQkopVDnLL4ZL0u6vURBskUY3bsdjUW/S7KV
KyOivwtiFiK/S6ln4DmMIFS1EUwxjpx3fEb2ePaTMIrV+YfLN6/rgWKgvUZ2AL65
4Tw3y315S2uwZ0/naafWS+wJhVIv5pNLdcqVAAkM0chiRkAWsUZss3rLa7ytlp8M
uQ4se6+XM5JFiAbYfBt/JXnZBh8UpNFxAd1TMDZ/4zKDN5QdFLC6BV91NwnGffdv
++Ug3HGUIK5OJxs6gJaWRvYV+ReiZTneQ8Qt/YU88iCErdXMHEipvt8Gkhpwn1Ws
7KRrxSlRm7sl31PmxS5t/E8RKXYXtYV8bJ5N7M9Ensz7F9etvPe+7mdl630JvXoU
Ey5stucHGsFEkM2awTAVmHLlIEq7V+yOUle3tGW17kUTJY7eceUmWkCJWuTl6qJw
+o2PSaC+rf29A8pD+ZrNCw+qYanvK92+lRubTxzttscqqCwxWNyNZpeJr0zQE8OA
BX0xIOfDZNkwZN6Ba9Q2yZ5ZoumkZAZE4LbNgvWIPUJW0svtikGq4BMe8gZtvOOp
q9Bryut1Mql29erD2Ks+8e5yiidctCYcJHz0qrWSUPksfJ1ce/Q7EoK5UlyhCRrc
TKQ+jJvHwckm1KEjstxSO4FKJoEgS9rgJ2Ed5yN2uRS47QrfK57eOB3gzxLVQVFx
Q9BqJyF74lbR8REREDM2NPONUcX++hTu5Iz64BTabsemg6zTKfsAZXaeom9WuIDG
++aZGLEQTxb/YhAW2qPUczUlpV8/NLnKL/XmOmgQAD6HMRL/7Mv64u1b2DnLIr18
G1A5RbLY3y24BCf8SOCjSbIgtNBk/SALAIxDag0hkqkTnfu70PtGo60mDIM7H/e0
QAep0/u745hwljiBLN6kICl1N9DycQhmb+Q6aBBF2OHZVr/0AyyWtyee3+fkwmix
4AOUtdSJqz1HRL5ksVkjdS0/sUuRVlUI1hRH0XYiELwtLTx8efxqtgc07rKktVYZ
qnSIX84jkyOjVJ8qcq0WB21hgrD3MbOolyNoeJDOr6bhtpAj1txCh2oAu7jIglzH
NnrVCInuUg+wwdW+p+Ng6rOwlYNfLoFCQNuCAsn9zhVAAAZZT36mDpu0xXUoBOCR
uEgpulKDV5pHV+1HNBSXg9TmXwvzdvFtrmDKJH+lSeJkBcvYdmwRRcwn2HZGS2/U
ZYAdhMnjV27Wcgt0iRrAbj+Y6XWXt/5BerNoeCwZImtNWfedEqkNxNz5Z3bjwO3W
5WKLcU4Jc2Ze3AvPk1e9s8t4UP+PG9wmdSEI4BwKW4j9OPsA+oNL9W+cAD1ex5CM
+wqCeDlqY1xZUTyrDctpVPiAJPXxvTUgFENLo6zfbuK9Kqrf7k2iYcioIfjfgxFG
nw9h/Mm6/b4ftavevtirvGgtQc+eLwxNEQgCibA9mI2zXqoEBD/FcO2PnjCZ+94F
63ehEnnRA06wkg+O9LeNjYmjqTUJ/enWt+Tke3SYcCdikNJmJTPDVFsZQST2DQvS
Tg9AfD5EBJnqeFBYvQ9NJP01ToPXa5y5p2dZuvSvbF6Q3Ktctz+qb85XlW+6T7Nz
PCrAy/xMN1XsWYFrN2y5oK2GFbZhGRNkuXyv0G/escE9DhoKt2kn1aAW8ZbvNXc/
0L6c4Nyz76VhsPFrISQQwS99sT4i4YznhIOk2LOKJHfdo8Z2sg9Ph0a5pYpFA6Ia
GhU88OVUo0s8Xqk3g8kZj48Mx+gk5zgEeXQR5GVFdofz2zzU0d5sTNxqFNVn4bC4
JymKcyfq2kHPw2qUoc91smF8je5niavWhg8kmfvjOclAkpbSj4kxD9FvHqguhlsi
ufcYf3joBRVTEBA+09GVMwzbjbxQT0lSrqkW8j8u+zDNKecGC6ed9zfloDUoNteJ
HyZ/jZG+j6LT1l4bwjRS5QifyET5eWmZTlauUyNYmcM2irY4kXE+YnO+0UmhTbJ2
yX77bpEb1W65LWXl0pcV5cojICZEpe1WKEW/gMoWQgx6bqaOqFebadUIkUnjcOJq
rcL2GA7wpKOzYWp9GDqwMu8d8y4nB9EcI24QJHxYotAm1chf6jheaaHqeKsxrng3
f4mi384eM5j5CfsFt/DjklBgAqM9uMP4w+atNNXWz8iAb3TGt9wwvj49ykr0Teo6
t0mKVJQs2YPBFT+XnTC/7LD3hyVMLhqvQ1fxGjXRygGttL6yebZBJWRANfNN+q1P
ITknOyUjlsGKI3rOhtXbCReLenF5SzE8JXmbKL1qJhDpvEwK72ZXdHkN7tNd/2A3
Tw8eSmt1Gg6xu9MYBAKk49O7PbCWTGYkd1Auy/A2Uk0yonNb3+cs5Y2WD0Cdqofa
WRtWYh73dCsUiCnDHuFDRZ6oN/3XlRl3o1EKT0nlyJaNH8Pi890bSq2OwMNVUebr
0WqSx9Ywu85KS/TYzDJMJDmMpMemcwTz15Ubt2gh4UJ2j+mh8mVAuvbW1AmLr+V3
J0nG2AACBxv//1Vk+WGSfHsajkFgOeauMVqkm4Sb5CPqbufLmN9ln8wosC+Kci24
VQla9r2TDMDxVPygOrUj8TrhIKkR4Yvk/TIp/G6WDSgtbA4CwzQA4oBr+sfdUc58
xTCC7O+9VefkcyD/qDbDUtJTG8KHqXbx/V0uJ2NIQxuuHoX9jCIL9LHcpsJ1jZP1
6jbQLcXIHjOVNGslXrK6ZWBNdWE/O3fN2jQU/kAHQ31gpjDJIvBxu3Pfp7XLlOWs
lKdzwDB+ZXXJjjoL7wlGmvcykZCtRViyReIN7PYXnANj/RmTqlPKBrWf0zyr+j1+
FS/qry1jK4L5k2LKueIrNLln+Kphuog72oam3SLe97MaTjjb3lceFBAoDuGF/9FE
p+GTQXDEAez9RrXKiEkXDix70sS9HTaOqVyNR0kGk4VGlMrTviiFqvBpQKJIOuzU
Y6KhzEUkaiC9YR+zio9NFhlhlk+hKvXBMdSLMIWoTdVx0RTsmG+wbIGsSqxOfZcb
FCvQGoNIeuTQBZXBWYD458yGuzIqWfYR8jnp7cloJRKT1Z6i9t2hLfug/qQ5Z9YF
3LaY6a/1A/LAXJmEyY8DpBZvc4bur0dfviA8+BPQjZeA3lGAQqVYvwB5xwyagiDy
Q0ayPwtzfJCLXeWv2hF+f4Gxo7eokSYX2oJ70CCHhF70mlE2ppjogOiwhM+iGm+0
QsW3KL0/b0pm9sPRveb2sXRvuoQqTtK34tFw32/V0f1E5cMAZgI83DU8CNYh+LIK
gh+sl6yivixOKLd0NBjNf/8UEfy321Xi9SDrKFwoH8C6djSBWmz40DdfeAc7SGIa
6yXYX0soUYxtblBKzV+Wdl3dVEZCbtql87AijBu5MjLH5HOv8PpWgwe2Ziokv+Cw
fHI+dL6nN5b2PYYID91oClOgMhtFxWdlrtpsD/42a7roNzKqirFgleKtjNt9v2og
KiLd/FzClT2AfvHlMENY5IR2Pp1EXewQIxJrGLfFOWPgjOce4c4WJGu0TATgtW7X
jMt96kP0n2gXSoRhU7OxNADexrYAuq06cioSGiQtEiZ9SZf19ExLvd23XRMl6ck8
NAAmTlTYD4nOWq4+hgrllVQX017BRgxUF+gqIs8Eczc5gOUQbmkOO6jUwMzBA0Y0
ZPwCa2deaFhPXYouKxG1bORgnVRPw4qdtrbsqsQEFl4B8H0ZcYJkST+4b0AlhX21
CCfz5HvVz6O/fEPngVf5OY+zkL7mImdA3WGDYZzbi1/YzwwdlNcqykncg1zil9BL
SBrXUEm8+ebEcUZ4xtJgHu9M4MSQsCvPRPSLTEbanX+L/HSUTPvcBREZbX8HrCWn
LJ/34VZv2uoAweRRvAYuazCEPwJYt8+qBS5f+OGQ0puoMBAlhAdILBlCX45/+GhV
akR3169nEz5P6OsWpjHC9m+fIZDY0l/zJv7Hk2yaRBw+a+eSJ/EguGhkckQkfBgE
mQjw+CZp3TRMIBVzOQhr5oY4NwU5DPhcyjjsc6+NWLVzcBtLVARWqwBYX50quEoY
hfsfm/GBSOzBzbWbLViODI7TO1GR83lylghWUg49gHsQTybz7UJSnfpeEcB9aNtr
ZGYmq4BIpho9tfYqKMMIssgE+I5IJrK1a4KfV279fTgtkjKv52WeCPhOd7JidHcz
Shy5Lbg/y18yVYzFDRI4rNI3D4BPsUd38cBeLgnjONHw77muEnHbHsrtaI0u4Z8Q
67vrH+jlmfKQtsgZGEFDKZulnOKfRUOwnrDlOxm03ReGE8LO7lyVNNN07a+Bc1HN
y0v90YPwyp/BHarRw/NQ3/LUVc2wkjhfNQEXxW6Yc4ZHrmSj/fL4MAVbBMvPPKmp
78gXbtQ36aM2pgUF4twH2rtvVXz9Efe5TRkcYGt8EGKeFyH7W8vg+onVnL+xPnR2
2MFRe5vwqkLO8ZE+YWjmnQRb+L+msj1wVsyGKKQaFIUHcf2N6X8uoNkjyIO1Hfwk
KMwCZxJsu4SCSeOS/ALSqKQl4IsJFDkjzD9tkuqgPcf3W9nSPrm4xTII+yOt6U0y
GLZJD1d6hS+Et345agAVlozZCTwz0ZuV/eh9g5lja45ihUNnoFElNIN3eUxFeq30
JupvIq+nfHTsv4IG9Sp6O6SAyVw9bdkx67uZ9v0XOqrlevdhGAN4v24EbHgDVN7z
nf7j6oUV5YY1balfvc9hti1gnALbTE0tuC+w4tckY0vssX9wZcFKH3VNMp8Fi0lv
W4A4MrNGBhPr+yBg1/MsXOaZqiDisg4w0foHOj03TY82yfXxH7cHZFbsfcTuHqxf
tEGXpU/Q65jBkOEHkL4Gqj09weyJkkWBQgkzqAY2RJa1S5iZygYbxp4+BfRT2ljU
BPUc0GobCLHEvSaBN+hSyKc0zUdQiWn/7kRZGOLcZDPy3S32bMNi9g+hwgorctlT
K201/DfgF2KRXWQu7OiSElm5DlUwCu/0pvILcZ2bovTFpvibOXX3jweUIyZoCHcu
PblEY+q61ho5ylkw9i6jhRf+P4YriOcuRZ/GE0X4E0p4hyM3Ed7R3EPb5BxECExn
8Nr4tNpS/OTMG+/u0f/CVRLu3HBpgNReNRWK6wdMqJq1n+TK28NmE6lTztGj2Cr6
/Igz5FichO0LrIv99uzS4BR0ciMi8qZDtqj9v6dY/Avc4qBHk7L0aztnTnzM2k4T
H5E2HIf8jYSRe3CPSvkM4v96H2Ds5eOznrMRYXo+mIM3Bp9nOtnWQx1+F2CN/TmS
WrRmC0HGggXFNMGYu8zTU/EwFBhOWxRXzwF7Tkm5/6MjL5rbJHmRMCO55Yiy9rQ7
W/hgdgqXIw0r6yu1wn7AHyk8IubIXK2Pk1V3LyOCujh/SiIrH1EhuapF2S30BMQ7
pvc7Vjj+cQX9gG4RZfatTkBqSEA14GtcPCIxEs244+lUg6MxUyZfN87GbjX6U1xF
4K8FqPuxJ5caXKkAnuJsywKkteugwNPW6IHhCLOMI1Hz2CfEd+KP4mvHjCaPZ8xH
px7lOsz8DZKGv7QVc/JGa82Vszpg6TcOm7fTq4KCrWsoHEPg+LDNvDEe/eJj5xpS
WM6u1fy7alA1wJS8d4q/vHzTL36nR3vZ/w/+KyWQAGzoiniOAsbg3i9QETiMx25L
xQSJKwy4Um5tdzef3YLl84tzE7xZ5Z4p4Q+m0GOUwSqpSPGpDjvwynNktm4BCjXE
K5aprEzaw4iw7rpILvRDntMSM+qBGBPq6/CSSjjP8xOeUJRHe/258EVn0So3RYMF
aHHh7ZLpHY/NnyW/El3wXlaWGoX6nm1qBw+VbRI+ISry/krvE/yBeQS3mXRX7Nru
AX8cADYWfeYMVdVLCpYWH0N6z6RtyEEPK6fBfj5vu7Ip0qDVw2hPVdsc1ehyMKJr
/m2GvAc63RAqjl7Z8OvKVfKXyhS8Yk+Z5cjHqEpHyNdNX90ucrM6Bn4T+Bsb11iM
tEbfrmTUhoPhjyZm1EMTsanQ0mAqtz7iGImLJS/51a0WS7z76sDoQdPNRJQi71HG
s3Jq4bRGp9MrZbIHay24U2q49GcLAoHxqG5UHKkiEWk9mPpU7VA6SbDgetFiSlP3
5/Bh6eSH7+6MjJO9LGHz5TjswrmhQyX6Kb08oH8qIVnK9QXJgOFjgp1H4aRLLpOf
OprKPFXII04Uen3KVzHDy+LOUiIeQaVD2mIeyi7SNO48T3B98PmpKpDpsnrRJnlv
I/heuv/BY4tVg2Wsd59xJwAHoJP7zJm1s0x51k1bQrs5/t8w60GoX+IAK3Gg3LAe
lBfZAD1kXl8P6Gjm+F8atjkr4pgc4NCRePuUFE8Ir3gI46oHSrKhZYHDcfvtylxh
mOc7xj87bUE+OKRnkQj3yfpBf3hKECzfBQbRFB2Lqx0dxW5ULDScVyTe5uf37TDp
5hOUNFjLIg12HEagqmOGwxEiHQQzpv8rom1IsrkYInPmx+66ZvvTa7UAM9AiPd0S
nAmBRurd0Q6KnmcZLR+8mzhYdKC/zFWfetHjW7LkZCwJdQcDeIFGBEenfRHHRhCU
qkcE+E9iBOcBh3sk0Agp3bUF3+l6aAECc6+k7bOcrIEX9ISUIAQChWoD8IyNslaS
30tn+Jgy+x+E0ZYp/OnYLfx5js02Z/L4LDOHBIbVaK0KpfRRBF8tbO9X/k+GfmA9
meEP+5QTy3cjHEgaGwycwt10ZY3wkUvddD5Q3yCBQOstokfYWsh/yvlzvW0X7POx
W466zalxFBYFSFFvaPKkajE1orct3y0CUJVfKlPzsJWnBe8/ReynvfwHj5261O0o
TMuYwcX5pHw3G+TFid15hkXD6Vkv9SimJO9j95Jnp4pUME+xA8Vbf4SHecjr1Of/
ipLdCMN/n+XrW8CNDXi89JuI8d4Y6tLve/SkU5+J3ABy0NAMgtioMu5ewXJOaRYY
rhGIeYOB4hiGr+xlQcvPS33t8ROvNavaeNxSrdv08kecW/XkCnDC6vwfBOfLezOr
98IEs6rjIjywWrDSmv3n+NyS+I96bTUd2ys9sQ8DR6FkH5CvZpvJJLCXq7S3kxES
Y1B5KwffOUAdbKrxEASjrvk5FWh5F9SHUzmv9XiuVongcuhiMjESESEijI/CUkXi
dLzzztBkK8zI558NJAodFh0t/ARdrmPpxSkw/5m0NZ9yo+Kvjyj/9gVGKIAX+/v/
/5xxnrcmHJKzdKtJyHNgezaoPSD2rdl42ol5NGWU95OAvAjidoGKS7M84x6e5auF
9s5ysxci+ot+lZxO51+V+YGAdmB7hzOZf8D57PODBHJQE/frzgcTXojD4d6V7Ieo
lmqMieJCusImwVWsIj2PFYhyFwIvUgxcr7K7sFGn5j6o9e7XOZ7YF03QHJ0rtZxk
sV148Tj+53d4cQX0piXgXbKqJxDgsKv7tQjyHSBCUb81GhScyFT+zH7BkH1sgAF1
udapv1RocmA8RWbv0kiyqesMqaX8ZAmI+We8HuOrPjlFvYRReCl4K2eB3B4cpKRs
bWSo4cHmaA4aJL1aWdq9+QmSjVWO7vZ9VPCo0NKethZBvXx+wI93Lj+W2Mj/bKII
BTlmohL6NytH1PaQUrA+ZA08w51jz1vXpgHu+pXUa3+z4LDlDcRN6IRWwv2bFXSj
K2UgJW9wuAZ3mqi2kENmtLqseOWyEW16+fQkOclK0YrZBagFRZC8dQr3wTBmn7MC
n4wj4lnct67FZ132BjrArarGBaJevK5PzdsRNw1Cfa1m08ZjI3Jop1R2ksmDRkL4
ehP7AfX9cwL1GcbduodrbEFZeXMQN2xQy6CR1TYtl2JYGQi36OnYNOti4k2ODjAY
OdPL8YY0IREP8PaQDtu8nhYhcXr7tCqWG2HYj9WTcjZ0Aj3q8aAnhTtoenYMoQpP
jayzlZXJpWuNZqiEqkezu5cehCfQYVOADOet/+0mqmXSiFDiFfSPxCKk2ZdTSeTY
NyvkoXMbKS7CwGLO/6gFDRAyxsa4v8LUGF/MXioefV7YjCR9d9LpdHPp1AXdOcjb
yM8gvGaL/rnD/qjmwDNnBKiTbiAaaPgED8m047ExtVubcuuV3N2Mmgo+mUDW6d1v
6O78QmfmEvbbCsa2fI6RyOoGcwy0ctnHInN0gw+XA0uwDmsmO9z5bIVIfMGLklMj
2051MJpN7poUEw8ZBHJlb0PQy6MyhsPnORPKAl3mt/CHh3u/OsHocCsdD9o6elpv
npIUFDYkZ260lLd166u/nNHMqAiESAu+Znow5ih/fcG4kqwcxFyJXcUU3qZz9WoW
nBUJuCKxZtlt6ZYwahDcNLpsm1gbIlNOLFF4rmkNQ4URLZfCOr4H/Ro9+YV0f2pu
rbBBMg1mdJx0VK3O9YTyQw1qwY9biRoPG8igcbNqjYzsuit+BZzZ7MjhOoLZT8M4
11qhqnq1hBpH61NVl4P/rDXkofRAwJXl4tSfpPH7d+F5D2KNWmCTzIOPB+XQsAX6
KWq0qmDFJk5Ix2wFduQU4FbVwjq5J4Z1JnTrMa8UBpIJ3FuYQ6673AbFM8vZb4RS
YbhpGU10bjqUjg7NMbpn1jWWiRinCIMvWvXN0SJ0CVx4ur9+sDmd7t/ue5bw87bm
g5COOgqFAjfUUuPURIVUasN5uliknL40Fe8egnpJk6ZWoVuUm5Uo9YOofPiXQvs9
lmjFhoYPpFuaqYZy4jTs3e+JZuT9HFGOM70cqXdRG0KHldfP23aZUEc8IlJlGDQq
RM5zasdQlP6WTscsnnsi4E4J9jUoS1aZDcRnfmjsqLcbX98037VmFylz/zf6OvaC
tl+dQbqw71hd77svLo4aZlY5xRAXa+kjAp1zP3pxiJ0xcYKjE0v0gu6YRjwI6MCm
t+/Wda7s2HQx+tWZ24JYJ6EG7d+bkFkA49lEoqw4ENte0Q5fYhn2hTbKDWJeCKA/
emXmKx+8Zy2/XAHGzL+9NnwHRLerTywuiRv5WEtwvj8WBxEpTp9RXvo49Y1lUBTy
IojmdbvuLHsphECT2Uth/ily5cHI4qw0g17x20Hbh344KN7HAD7mHA/AtLmOg3te
yt8hsAjXMBAgCcgw2MBwYzmVnc0K1EVvZd0zJ9h5XFZyJKEgzXhELnXcOgLK9W2H
e1macXdMLZT3SNcHrn5iI1NF4VFKt7GAg027f13bGkAaXzuemxbETtQ+l7cpMqrt
XlwEtDzBID4B/bRdog35bS423540sq17a4MsWg94Obmncrw44xKmxXDhwNFYd58J
s2WsAbkT1kazJmvYqJV+0LyQ1j49UtPUQ/lR4nM20q5+8vD2yLZXI1B2WmeoWb68
eYG3yZ4XiCNUxgPfIEECHonP9mnk8hwGbN3NQZvGRjYycBfeGJWQO7jUVY12/ACQ
W31E4ou7Vlxwv3P9EQejCeetYn5P7w1whE+gWoXcljZbEah2DMp0NnTM2omEzEIc
+OQveKReN5jQsYeb/D8fyXBrSoyqg6bR+0Hfdv/X8Oo6sb+kIq5OwdAysufz3lr6
oQBb34c0BmypH/4I9yoqa6cy7L+T9Z2/Ny7b+qEpY2sUXmkGeLO4KB4LrtbwBD8w
58o9Whr2hA4FOx8CqLSpGkyKrHUNfkCIoqGnP3rn1SlRJp90us5PuSiRIr6CzwYf
9L8v4CN3TOB4RGCzIffSRENS5PT6h/g/Kzq6stBiv7bpDpaEW0JmxbN7XyLKcR7J
bYcH5ZJqWW2AAodzfMDcXOBHhgvutQgjXjWbSX/ZcKquv+asUMXKyVS2SxsU9WlA
cfd6l4lXH8OsK214WJfa1WyK0fcqOBb2hAlgKx5IEZQm7UXTMySPL3VJEE2ZOpUO
p+1cm2vtSAJwRAFaB6dLDuWT7MykQaVCJn3jEFj4qvgQYmfGE3+PN1DJyX23h+w3
MaYFwdj5mIydjJah7v2g7Q8dCXGp7SXhNpIh/t+b8Bk3dV5gZIynqSg+IfB5VoQx
UTr6pRGkCcsONIt+HnYKDJu0MyZvUnk62P2kz/8WbuucGmsitWJ93m3zVIwDts47
JEazT9S7v+uNUkBYc0Yy5/v1rFVbJWj1MwfqmML+XGszJcmo/I5uJa1CiUiOLyvT
ad1d1LE16FXMttrPu+9OV3fDWgAIE9E0aiLsjto8mLjWwwTmqCSptzANzbZLSwu+
uCXedKRNVTQ7A3AVIiLm9E7HGmv72h+1r4uInTexg8NuWTNA2Oh0hXEwVex5ncoN
Qt2LHXiNHdeIAdFBkmRAymcOhvyqxaN7FUBcpb9MGcgSm5tdokXZGbIWmY5i/Si7
3/mUqpXAiyiHo/BkiAmeB+qKxqyUZJEU7qUyyrXW9EfuNwPfnohhoS5R5W5XDGml
OJFIru7kKzKmYLXrAzp3JWnXl0rAbv4/xzZb9ioCZQeucr8eT8H9ZcMcKkfMPaa0
/l98TkPKvTakAdIQppFO/O0RSYT7qxjk7YwvrNkmbybe8PUI3MqE4EfKUOUX2JCY
kdvxVOuetJsXv99PdFxG5zzpQy0Ee5YgLNj5ecOeobnNo6OOYT6mtrnvZZdDeKV6
c+MypsvNeBMR2PdH3TOrMFHkOiYIOLgQtW0P1prYOo4A6s9QcYWfuW1ag75eCc/J
lngPzr6/1bjqAaxi7v52j8Iu0nLtM24wrhwD/puv63PeJGZZvkYzrAvbPq/wFxha
IP/0doSXXlQSCsahB6hGWOljhZlsdBjjv5G1GrwVrM8p2MIEd8JStX+m9d4o2/yT
Wa+eMgxJ3QQl7KY4E7/euR+193N26FuDoIwTqdt+bcYnqZKQ23GoYx6aJDE4XU+j
p/1mQIJFpO7kkJJeZ/OkAU4YDg32OwVdUldZ2ug1LGrUtymkF3KlnISPeUBL1RNd
TDbTwCfIIe1v1QTSFCUrkIr/dd2liwb/XvGGFMPWnTz4u5FrzPABgc1RxWQDdFbS
IAx8lWVl0y5z/0/gCDGYl8OSaETeLh9a9DapXXiZX52r3On6WlKghotcrGcsJM5d
o4DGXeK9u9dMaf4QF2tAL9qWYcoqbwHsfZPXCULWqdawZNKIC2i/Z9R3rbL3ps/Y
pS9uU+ANQHKJMe2xzLCMnOo1ERZ87vYpe3uvHLspQ8+/pdsBALMdJxO1+gKxgNus
s8xohlb5YwW76+aryF8JseF3kDhKJMMAHPbDl82OwVC3inQgtnF8D3xUnEujlbV0
hbvxJxkA0gu9Mspxl9XdrMbjozioWkOjhdDfWpgO1a7m2GCI0TSbXRskAXZG/K70
R8Hh9DKsu1hLVbD/7jlOKUc598cMaNwAIlbYb0sOD9plIZxSElC3x/2sBuUBe4ep
jZorsADxXSKJMJQOfqRzX60+Xh5EiJzlb+VMW+KME4OrNeiYPF3AnhnbSrgNRAgU
DRZKwYRFfHeELe5nhBhe9FmyQwX1Kgk/zZx7rh6SUKlnnFXmU2c1+pi+ZLOUPlkY
OVLs5AUtrlaNr9yNITVrkFDSD+flDArOGwBxa0J8GzJ/Jc+8rMKniaH4eCemgFnp
QACCJ0yMeUFmT9k8zTzsWUznSprjcgeM+suUM7eNgw6hJY/x9pgO6gnNO/xdc8ZQ
X1Zk4hfYB1wQqId5BAXIas+SUz1XKDva8ueY9gUbNZLVJn08RtQEX4zBNsry05rW
wtC05liKRXzkE0OIICwajj8kxB++PNIEuEIzuAhNbiEheYhIu3PxQzcANV4UJmpK
NIHcyMwZHK2jezfKcMKg0NGMz18gXdqfyPB2Hr7/bVt2MR50yueJEyEvq3lXAaXj
/RQ7nUUXotcf9tJckEsXX6ohQ/ZqLrwPphqW/ochMxc9bPkDSDVKTOQpQqqfLrEy
2CHq7fAn+oXICZ5hnHt7ZidEf7cMEo2DYQzHi10el4djzc+b7hgq95WZlCAwciXS
kd/d/U52u2qh/anjpFMPe9ot+9ZCeeC3FPQ9i90ih/1fLAdVbZ1gWfDJh6SjFMmL
O79sE37hac0rinxkb3Ef5VgWlXYYx2/pgSTOdwSbqMChNizIKeWO6HF6F+gaU2dB
SwaegTCltXCzX0/2dkBj8/CJlC2MKCK2Ga+HNOVp4THImH5dQtayoVg0Kv/m30hF
kJhopH2q7u2fR7eMUrSKTLPF2k3AUQcoVY7zKSUrKtuhkfNo4zDG2NlByoB5xtuh
hwFg7suO3ojR1FwFYMhxkyR34rEHq2PrT/j6N0xVYl4IzYgYTUGy055d52dmVxRr
lZoW7VTKkGMePnwIYKyazP6u/s9VeaWmlru4QH+fBu85mmMsN+2BkGSTuegDvwP2
DTxiFie0tFM8NDGt/HsA0FnqPhULDCXLXqbLPUzkP13Cw2/JWG+k4MzGI8E6n5WK
nbqibswO5uRpPlbCxZJIiEp+pFvbUX084mCKVDBOha/hdsemVf13W+n0cdfzAcco
3pByWHmggJwNCZDlA1uLgUa/ZqE6A9ZU19C0l4n62bQXh+iOBNF9tqGJS/1pmMBG
tOag4nuEu86aYiWXcpe0AyQWTfMHeklptB0oLWEcmUa1rSOuMA/6908zKYLG+66Q
HfqFoeS5OWfaHYbObhirS2SzQaUhpoQRYoSs2FiV+J+1KJUJrr9WE1dEphsAAKzx
CvDlPtiwR4rnN76PjrbxOj3ccCr5UKO6h464p/NgtBA1YJTlG6v3bFh/nQaZegNM
uNoniu+WUQ5TbwbHKtTsf7ntX0Jz+CU2dycsVVlkTRFmYvGup4kfUql/N/1zfogU
q7oVLFPxWZRi9tJaOgZms0Ypl/rngAkbZXeurq6SD4WQV1fYfOlpZygnmySKJjfG
f3kmUwMvguEzn2EdOiM0qCFzPJ/K7n9bpjb6Z/sKilFUx2G6HZAX3bgjQR2tgRJn
Gi2J/yahfd56g6fF/8YZxxap7onJotl/dx5I7WJGJa154mkCt4Cpt/fP3J0B6pnR
VSLFafj6AhDO4RlDKelgvlxpAQ1a5GncBjYR9h5PDFMCPNsWWWrmpv+BG0NPjKDW
ThRaWmCqTGWQzT8DZz6V+0Ic3X1dXlhop2jrDiu5keTtA7pxQvTiWBvN+1RQDTTG
zorcyhTSQ13uidm6IJWN85FTWM6iArAYb0IwlWhCKHZrXXLjzzbTEz510+lofC3B
riE7pXBVe01y+FPXpYGE6aAKpjjRQdXBqxQUaV5qd0o6d2Vt9GMC9828hYgXmBi0
YO+aEMTZyMm9m4x8UeCt4tBybE0mH+BxMVBdxIvegDvKxokNSi1nHR5UdAUEzYAc
4p0hxoX2CSf7Hd3CZkzhOnEi/tzh3arYtDPxaGblYUg8ccdQ69U37se7JRjneAna
a+C0aTm+lw2BBtnG4tOuaeFgtHqUm8UVTH9KtDFyM/I3rdZbPuqKHEoXMw/VQfep
h6/QSYLw2kkWccXUf+yhz8mpCQAN7GVH5n9ii9Ri1MP0jVa4pGSPsW8L7d+fGcVM
ufirMWnJ6x4JMgEFO/HhbnlQip2gK9UhXPnFtdbA+BbY3hxPS0yKdChMFs+QeNCl
bK/jk4CODPS1m3o5/A4SEhN5Or2uP4ukeksFkvIqeV8ghNGCiAK36YVoQV+vjh4O
RRn9vkYpjbk+Z2o9fl9E+p/6GF77PfllErf70jPisJ5UIh44nwtyadqo7F9MBqvX
T90Fkv7ro1Xtt8RLCAZlAeWZ1HF63EqOxz6ons74D96PiA7UP2rvfkYEQbJ00Dga
qdHjIwynrPrBPMmxbIikJG+/LsmT6gUrEAxtVlJ3ZTJY0yZbId6m7DFM1JUQNU+O
NuturkZQwaf/ailzsMeh15/OrBi+wRcULPPnFHNRMPpXPckyDufbZuwTOCzht5oK
tVjY+FP1c7Ve1Xyg6JDJjwCYvMUfZb2mGefunq1YJVOPy5Jv+OFlTbt+n5G2BPew
aec21UiqXE/fuEQnWep5LwH9BvE7PPmTS+nP5zRUdktbjKCq05/AUxC0cvfFQLkm
yW5u4wSdjzlx/aTMImV4RjFN3pE6CUM/9uy4OyyYOrAWu3LbdgqDsqjZ+JUjy+tX
raJWHffirlmYgdlZWgoF9Kw4WC/C8O9lzP1OciJyKju+pi+Jl+PWN1SX1DSCHZsh
BBrHXiznd1cbEEtDJIPGMk2a5i59E2xLnZEQfMSMrm3djY4vez76v39GS/szzJK4
N5N6Z/9AjIlEOvnAVKWHePGA8lA+2ydJHCXM9eZKm3ERB53bokdthwNjpFAnjdn3
HyHoEN/3HfrxkT03wfAy2e6urGufm6HrnCeUm49vn3KT+RCZGMJcGyHE1mD7PnSm
PL2Eo4SbdC2J8mpJrG4ASKliaKnLa7dsE5dr1sr0m7QxmYPTx6ojxrketbWyiNk0
k/nh977u4iLS0y0TiZEUtwg4zGSG/lx66SjT8zozIGEAmdM5yQvN6H+LFVmsC32E
wJDMLdyI+SEYMWGA6XA+udrDJpFNWt1bgCaWTCtlZY0O+GMajfwHrAMqBZn5ZEtY
YulL+AG+VGqMnUx4ri3ci+0U9gmncS9c5daFQCRaUOtxHFhnijnjHjRIU6sp2Mbe
al4ILR+b92TcggEbMOT4bVYdgvemR7ucpOzthaXr9Y6z2lkv6lN3J0g9tRXcTIB/
1o4xvamIhZUu7wpOd2uaUWXeAnbGG8S9iK7ED+Ftk5vi9qyMco60PB8d//nKoEw4
L8rnm5+vVq/VBcs6rjhVTSZQcOV879gkB38rs5LfMJOePUAWK9bX8VYa3pP4l0Rs
ZN03FmTrU8mO8SkiUT4MtLyKJvw7XISmgcOcOcsTcgOl10cWtSycmNPlEvseGyiY
YFL/q+rWb/hG6Oh0P1RuIiY4oYBvNJnS2WJ5s7CRz+tn+8Qbxeb+nc3qiYi0dHFq
r2REFzu9OJgWYli4J0JtrkWKye/K/O9/5iDoACa6KXIM8OLYaXgzcvFhP98a7RmW
sr5aKZaxn67CBgLK2tR5r9GlxhzxELGCqgMIdtDzDrK5I9dCpsN/2YRfH+EGczYV
64JwGIvkXsKsxXmrh7ZYv5L6gjZQmTi/7OqXSmBCTomfXZKuNeV6RyMkY6CCZohQ
wrrKJsWWjROL/mjGY8ZOCF5vFOSh4ZOO00Ym3dUoIju+EKD5oZ/QGLjDNfsiz+4q
D8tMP9wDDWBgkozD0zMYzR0LHkoL2RPUTJxKEim/2L0cOVFzqwBw7dFHYoMuwVK8
aD9jhrZQDdZxCURv85Y9EqqzTfsoprT8O9T5H73iWSOJfDOhCybonEM65EnroIvh
vbufXeAJNiLWEOLdq0V+uKdH6TCPvuGg7qAJm2TZ0MYl3up0Tjjr4OHV0KKKEV9M
OCvqG7lqBBJ34ngcbDY8CzcMZ+KbDMUSfJDLgAIKd39mxzx3tetrZravP18adL8O
iHJhVImItW4SXxSLuzoCxAbb1WtwnCPJAdFe0Y01PriGneRZ6wDLMQEcw01nW/KA
bkaBvpc+tYe9TG906eS4BvIOiPAALArAXqUiP+tJywDJE49Eyt/KMYa2a58vPrB+
h5EWzw3YhCh20umfkwXeEUbv/4KJv4kKgakUZgyyGfO/edcaDwBjKXkexhXsPRG0
RBb0zBevLCqIw9gytJYjxAc68dg72n+uaGVwFYSl8VB8LjTt7bLL7itsUJe3pWmh
BYs+jmWmF3r5pJSE/YO4n/2SaggYyiWzNTj6UDbeZASndwZbRjPQYLnoAS3bxtfC
wUt1/hkU9YkKqkJlnchPNapo3LjzEaLeGjU9ZLKc6yIUKkUmIp5DA5baMUY1Gd0E
AFBQYphLLTLH8N+FDUUce0lSVgs7nbn2V+Abe280bkB1fok8bHHpLmmDrP1rbVUU
4HNCp59CwGZKSZU6KQZ2qbbRwPWeNF+pHcMeZyaRyjX+bXbUlzMweXsqz6GKncHW
sNWEEVqWC5S+RoGu18MA5EIdy9a3tbA1ftpszE/po0sIaBaRa3q4c0GKhLXh6MH0
40GvkCFLpjhCdZv8nRU1AI/0bZbt+JoxyZ+SfPQuFI84ehLKSJwCXSkUy8vJUZ89
CuLa79DgV79HDYyaiwSt1bGGaNDd8IJVUu00310YrDs0eKoYcWdC+CqRLQtjMKxe
v/toUeg/iP84xX9OkZVtHC4hYpv90OXAYrfdATx1zLPCSQk+oIxw0jFJk9oXfzKy
KFBfDMgGSss/PsfROz3akyzq9Wo4pUv89e126HlcpvETiFMRCwwR9hHITQ6HaLeh
eBj+Z0MbRlDDQeZ6HPFG2av8epzwq5gpMk221uusCEPzqBvht5RN4kh40vkbcrew
i/ff9fo/qrVde9ZQ+XThd7s6VKZWFN2VbiZlbI/QX1S9VBfTX9uG1u2HV54+oJ6b
WaTiSvqjJD/GIg9DpgcbEMwguXQeIwaI6NidpevDbktwl9PWrprVRH0mepGR2ga7
nxZ4cS6xkWQG/Yh3VfcjYfa591M6k7Oia03bBIeLrEkaHqLETlQW50DeyzFq5+Wi
NnL9IVNgpa3PhZRWyzhEiejgYHGge3chGZboJlrMHGunuAZeIeEBnWJ+Y9iNce2g
mj38+rO/62IAVN8QKqwUKjnAU/6raVT8zGulsiXxo/Z91UidpNZJ5vJQLIatM6DC
4hBgj/XDCUS4/DhyUZo1XAPI6YsP/tz4PFEKWZZFtaEhPQxTjppPWxaCxIrFeYga
HlVKtW5CzTWc9ekrmzr+CuZ48faf9PclT2q79KjWUE8w5Fw/UibvhywgF50wu0Kw
K9DE/MHW3KxbKw7/hyxKBQLxzQnlA7VV1Uv5Gi2OXtTfYVUevJWoRXEn2x3fcHI8
7ckcHpaOwEEUFcxCiIga4rEwcwNCc5+R/D0Jj1w201bQy/wMg6qHYh0V3N8USwjB
RiQKsNpuDoLsPCj1DAeq0T2l8WSTIokvH36apfIN47KmL+MvtoRLsUdOnqi5Basl
UNSBQDxyF8Lyl33AwcB4jtXeDGZ+Z/daR+29Zv0ooEgZBvZRAnANNMBfooCShiWw
k/am1gGEvrhcAvFfvpU7BABQssMCsgE8kt4q+V3d8H/pV/IkmWKyAUmoaXTeQIqh
Seo0efFbRME9ibgSdxgNHVWDI8Z/nAicNeA4v1YLWkVhW3QXWA5xP6J75TXKMvXu
bEh9TVuGgrLrodgSDH/aPDhZFGB0KWXT+bwWXu2+RUsFmnf9E2hBtnspXWQon62S
TsXMy+pNro5wdGtWNWYXt1YXyG9C5d1TpjhpzmKbR3+Sqx3AHjY+PmtOMHGskKTV
b8+AXIouBo1Fl+YULZ1fsPnhzEFWGdkl8M1iQU6l33SRTbTbAm4M1hwLSjG3d7O7
jM4CNwxkWi/uu3N1fBR/soyOgz0SJE1gsErfayZ6sQodKo5FBbFtW76C9hq8gRRh
ALA7K+bMlqfKqVUIKPc6WBqCsLLoFj1A2NM27XRmNSd64sbAmHrLHVFFUHrdyhVv
Bcg9ZrpgzS6ovUTvdPQOffMg9lW+MVhwefoSluUfxxzeaBZhZbCJTHluomSzpGc/
DzphXX+1r23IIygnxv9gUqrgkP9FUMj+Y8SEvJdrNOhUYqRUOj9yB4vh0Ld8aH3T
ezNqn44RhVHI9+HjuWvzL1TBeNEISYFmGVOWbwm5nk5YX8anZTJq444MwFulNW7o
rKSF1teg+3BkVUhMBo52raknz3qNx2vF0BuYq5BvXnCUvgffxbn5uhB9r+KOhDfy
3rx+JrWQe2lbFKxsXL1tbglIb1RSKzZtwyx/uAmsBuYDGJXsr8o1Ff13lAUMax1q
5QHzt/0g5Nos6rDWyiQJQPM64bUpYcWwtLSXVaJM7BXAaLUMJ/mS1zXrXgYa7f7E
Kzznp3qoJIX/T0HSz5Byb4kv/SrSpxEeRtGTmt+59GcSXhhgoYflV1wXYWb4zdEJ
uHaAW4KlCkg4c0CyJMK4KH/ghPZhZjYgsW/8rWWcIyQdc92jkYD5+rwG1k28Kif1
RG1TtN5aFLu0JQE4qCiMpSTUGSgCKTDlqRzJz3/gv0WkpnMXpolLIMrjrdiov4Ka
R8XHvgvYcV7UsReV2mSL27weuzdNWwR0EiDFuR9eVwoMOJxUOUlq0HsUHkcSTcov
HT8V4JSwXLMKk4QCak8n6ELJ14BO8IegGQh2p8r04LQ9JJekhLNx1XkSOpPDJY2P
XTt/WFiBQzN9hIOjfiQweP+pTDgabRARudbdAt3j/yiBvStIt5Ksh1xEa5QZfims
rhb+AAshUjp1Ek5vFUYp3Dyk5fdhoqs0ukG8nPkkZ8GQjpJ0ojLccN2xzlpcHizB
+H1LSSNNxYFRPO/6qPIR7c/8Hw9X3WOGVU7ZxgzMZv2BlvLyd2EX9RaHFwX3Dwpi
yg1birm5NqJ9w4fgEP4g6QyyGDeklLM5NqKUUWOW5CYp6ZHs/Q7ztZtY+zhloKl0
0RsTFaWJQV/HL2Gi5y1oHBCvvjg0AkwI5kIXOwFFyY3ITkwgFcinK2H6BL/SdV8z
z3PUM/k9TJUubG6X+2f7zftX9eF1C778qRz3DdnbDFH98fA19E987rMXTLY/jCHk
+IQIx+TPeQXYHT0QZh95wzzhgxubpx/0nIBDuDn9fzeFfMvADuEueuuDp8nPw5gg
HcsDHN5L5nj3X0MJtuPpkmFM/qzkviu/HPKhigvRZ+Y8+dWu3LSunt4LSmW4jFY0
zqlfq3WOHGt/Jt/FwnTHHm8voMTNIf36gYBxwDV/d2pN00PBDggGYYM/+91n93Lj
LrREDx0i9gFRv1L3VelUXYWI+T/Lzc7vMiQ1RlMf/l3fr+lexEd9UPNdsTyHMpXR
j8GtDshO0OlpJlXdkWw+H4ujLu1cooAESkLslzGvdgd2M2MJ4cBcT9tjmYNc+ILv
sftZF6A/4fkKcQrMuz3sR5QqnsingOMv22D5Qes1MIiwq+lO45Wv3GyYecWMo3NA
ZHWWEo0fwagbXr20BQUQujtrRZ3gOet61CBrPuXhfGTfuz6pXw6X4kcEr8Gy8rAD
VNFeBAdCd1KBq7TjpIRLpvWqM4mMHNK58tuArOuw9xay6QjQH1uCBTuKYJnAxgUU
MD5l7ysEGGDz35r8Y2y5POyWN5/Z5OXv4eiDr5GzpqL1CCJOn3AljmkRjBCVrziF
CqZQDFWWI+AeBUr66gixbvMAiOp7fDFDqd4NxcIbZnDVpuK3Xz5nzO+BtcIq0jr5
aZ54bT74FQhIuJXIvXsWmhBAx2NRlKD+nUay+U4b8XCP/f2cX0W34ZQkCmPfsCu9
aW4aPO2vlKIIpTr4kVdxiNBPUzh46FDTAHcJqra08UD+2yMnvMJ/LVRkT6uMw9xX
0yeHoZ28fCWYjJ/2+aEqwQS78JG8+XpbHyH4VmaOmVpbHhMTo0QC4mExoi6WkllW
uUfNXiM6gNYObf9WuhqrWoOGC2TQCnke9XEUyDzZHLIf9xLRGN8f9xWxcWaWEi1x
75cEbk8rpZEoAqLMbzkBdTxTkdX083sj8REsy7Xpr8OQbITHiC+z78YBomvnikRk
QcD7sCjBhVbY92ZY+yUnO7QOIs51tfJPRopV9c9zEHhKZxJZ2nhjXysOe1EPdgFX
/L/zA9rivSEDhXQrtmwmWqDzq7OqmZWuYT22Jt9xm6Dd+WYEcSD3T3/fsTnqmd30
Crck373rIrETXb+Ryzu7W6BSwcyAIFZoN/oKiLDEeHPGkuKqhjrOModSL4z5lSdS
xPBTAMLR4fNMPUuEn0AuBplptTayGgcnkW+bDVZTWqhEWRcbt3AZaXiJ+TqWm9nS
n3qatvgREb8sUjGVn7gu/kLPEGXI7iEyW74PI2nLeGIu8L2lFrde/QmCZ4w6DcI+
Ncv8lL9q2VYzML2ALXm9LHSyMlT+GvQ0XqMzKNIgIrxtQLI5kZWG/Zf7qT/w1QTw
f+RKfjof8/xsVJlKEUJJhoOQNWzzGb9RPn+ALdgMrKGQiMuLtUThc4r2j0IHW5tt
YZGgItaCxDATomhvegyoPZeEWfG1bsICvvErsMqW5fj2S6Kdfy1DITthoZJ7sTaB
ixdX0LUFWgswI8VP4Mg/bFdTpnnbQ0F0ZwzMtzL/Nr0tYWFFq1SnzpXFC/puWAh6
I9E/oDUIhxSi3MjjF//fBm9zsN7oQuHNivAT9lrDvPEwZrUjm4dv+qSAjMbyj+ny
sLmrzAI22EWggIrI2z4BTNh3gyTpFge1lnluE/koXY0rPY+RTe4tKu/5wNvpSwMi
Ydr9xDAec30q6ebqyv4NRNGfVT3UydC+Aysdk8VULHpAZwsRMoXkAy+27Er0nZNM
V+yTymWKxyI0k1zddxZoOtI9bxN9DDEEg/CJ6bfOjBAjP6+d+j3u4pdCfnJJtk9y
8YUmhiF0+25/JYWDNf1ZRHnuZxRQrIXR9FSuYEU7M6RRvseN38T36np1LZNwgU0g
KFTbFq4oI6tDKHzU21scZCG3ctsoK5zf+rvOUEcVe2oFUkw7vpfMGDADBIFhNWnv
Yn4ZFm3aVM2FZPgESji/1f+n7Ptr9j09dKfBOIrN4MMLMvVHKW8Mpgql83ZOtsJp
JlEDlWPyXYZmewvo87nEw59aojVoRqzu8XS4BGFzCZkUDamcuYWOlXrNTjMJzWYE
yt8IKr0e1BqSq0s/0osXzfakJIz/MIvnc9MUcoYREdg0GUEUFujAFzUo5mWqW2Kp
nn9pHA2oEIXdq0EnS/aFvS3uZsQCS7PRw+NtbF9GtMpfRHPlymJJiB5Je8zOjLDt
qj4+Do8wwrN0fbtiNaeSupc0W/HbXayCVk2KG/MvvJTafeTYVvP+RvJx8p/AbgaB
D+oYbGSlsQ89kTygQqIH6iXiVFiyEKGyia8Ea94wboZhlgtD4Dpnn43q1xai99Ah
HtnMkJ6Gc9GajjbGUJEOS+5EbRV6SXmmBbsV1symv4qr6QRmwf2vSM4eq5KqmD2Y
byn6Emc0bu+kS28gS2KielOKM6wG2Mn19euZ1CDTnq8SbK4lmlTJ2O9O9ECTObwS
QUZedXcW/C0NdaFhiVDo0zyJkrfz00oWkYTyTmdM5cOjJCgvWmP9VgPzF5jEug2O
A4ivstl4jJ9fN2rJk0ozz9H6E1K+gvE8yk76Yqezxifmom/wl0GOrJVi5dqTZPCe
LA+PzeLMR1EV/g7IKo23C8f5ijeX1SK/UUWmZSia3sCWZXIv1ccaq8UkyLmENzB5
TnB+Y+CmxH0cqgRA7+nLfQU0HmCaOew+4xSzi5HwbVLn9e9kRRPMgPVw2vhicpWA
l/+gv2cKsePGkiFCDeyQXYb5PwEO1Nz0Y0GJJoWBDr0hPlFbNw7Mo/Vm8AACR6Ci
z0QxMWHhuxkNyODn8RwztvNjPJOtOGO/xNqnhN8MzFtV8GcIKDGSxcDrApWfu+UD
bh8PUNFFZEuK/BFB/G8DCEZPdRl3y/gfIM6xHO+NTbC8pdS3tmYU+JbGoTv9Worq
GrvQrTyYWlBLF2kMSflNMkreEdMONRowdyMqYNSxnNWjkhV2Nj0mYkNN3UoccSK8
pxTbXUtEq2du3BoQ3+ZoX6qCC24WQU0vQOjNRdiRqJN8hg1g42/0Wlsv7VAtjFdp
rRO0NRClGEyL4mH+9LU/nl3RaRcKExqei/QRcCWtRBgJy3MmMsm1I/00K+kUiV0q
ok8wfbKvOcsEgrPRe86JWAU9PdiH7TPcfbXCnlQAJZB8xA0Nu5dvxz20gHE1i3lt
WysNVKqk1bzCsqsodWVs3G3wrp7Y922IhxmLOVWdTB+Ee9R2kZaAx3KtUmzYaqpW
92RNrv7zNiiW9QaqhTpuJWJ4X18GQ9QVU8UFV5qNm5HH8TVhYCntewcHMOi4gfVR
Z9Fud6U6BI74WUR7UfrBM03Ssv8LOuLFHsM+LCCkAJYaEPI96MsFWI6XBAMAgcTG
tr8cnwMCKFZNGKZCzYbMzOR/52zM0XwhYkwSdST11bgOg1KWBoPENYHfFboWPkqf
K+Yp1uWFa3co+2frijQDS+8rEWK8SC8Mp+iK/6/71dRhRhefaz6BvQNfVMG2G1EF
WdexR6N7KFY81WAG2POWakJHUPLxvMy9FvS6FO6X6m48UhK5POB8474kQ+pKSq1q
1CSmi8GW5DM4rRaxAjUITepJ/1X1olIBCoodtTFEjcachVuhiJwH/rhacAcc+LgU
uTCeLfKj0aXA64qqMYvC4TJezYdzDpbKmeddE/LoUsuZkaJEb40twCa0S1EMOkI7
5zkA+YUlhYgIY7TxyDDmTQR32SPKB2rFyZNtv+//PyQCFeqVhIQyWKq5bF/6L24j
QkUKH8eOJw0xlKMkRdyY8MjWMeOzeQ5o2duer9zzzxkZYc0jbqVHGWXo7xUnJ42Z
/F+IpBypj9Ly7vnnAcfZtM9nJXeo9rTxcmm8w9l2Cw/tcNP7ormtDg3nBKK119u+
+wMvJ8YbneoHlUEHhI7CDp5W5dyV8/wNIPfjxmSd7l0DyIldGFUuy3Bi7kWJyRzm
PIZSbBLyKuQerqaUzI8y3ls1Wee2jaEing/sd5VjM2469obdtYnz6sOAkaM+h5dc
hhv9FZ2DT8tSkC/qO2+jHlPDiaBXh3yAL29rVgxS8Sd7eZHJYiWREEYIM6CJHWhr
xzVr+os95s2NwqQ+Y9WW1A4tYVcRB7vYaU04OdrUDFxSWF5F9a8D0CmbVp/wFT0j
m6UqR+hKZv4/83FivXrs2YFsV81OR1mootWsNfO/yzrnssi1FjAyDXR5vpg5SU/z
Rbl8XL6XUS+9vnR0yLe1Gks1Eahjog5Wirj9g16qM6dnLRaobpDq8dCb15UCwqYP
DB57w3OsEBKRX7LnhBzJU9bnxILTBS0Qu+eowq0yUiXxk0SThfre8vNa2VM4/uaj
PWQynyZK6jSHMJ0ZIreh27BP5YPGPrida/ptnG4x+ESv5oF/5ZmOwmE18EXoAsC/
/zxcZ8QRqUqi5MbUdh65mE4ZxTkcjaUcd1FEhdPuOjyBa0gH/H76gtGVVXLUWAy1
PuJyLtXIJ9oxgUzDx4qdb+XW8SAJxaCbZKBogToidI9x5g2nLL7j0jpwsZeD0YJX
YMqwg1UIdRtB8jXZKK2yzcMzbtSMHbxEpGam3BaTlP6+Xbqqsy2jqUdIxtpdOM0L
+cP3CLIISvbcJGknX+g45vqv49xBV/jQY/o1hmhNiMOroYiXz5ivsrXDUeneOZxJ
4IQ8ue1F/WGQsx50ApEZ3v4yfMNPKnNDRVBjd2UDnKEw+s29pYu4UrcL8se7dhZ2
uvA59pXK8nP2ex0+8OcBpuQDEXL9lp2/sASS/xR+ZC8c3leGw9/77ErQJA3bMSQU
hWM8GzUdBBzCiBVY2dDWeBOwCetnJVbgA1ryZ3X7mPNb3zACRStZwSNOxC9RLOCA
gJ9HTb/i4VznAn6cqHcF/a0/3tfhqNNHb/6vLXZ31uS8Nd1dy+IywjbaYE9lhcLU
iJ0je5GkipIb7kc3AAgoP2D/iVQgICFH9vfMdjqt5coDPJ0F1WX1W8kkLJSiwDBt
WXKWrI4C/2BhsAqrMn81NLVQQxMaNP+mtYHK9JI9Oy88AQ0XBU7hp+rwR6sCJJLW
S+Asks4xh59cVVkOzLgrXnltymRk0/ORz6NdFc6blQAIzx66HmJYHq4iUR6uGYTz
K9Fi2lmcW0LICSKfESzFZwbkjA3mxF54uKvhC6wheWrk5F7q1C1uWW5hIE63r/UY
WOvvHcEoOVz9Ju+zKP+VywYRXvbWwCAVm0ns4mPZ9OuHK2f8v7VEk16wMVpRgykV
QifwUz4KxFKhEvs0k3wdJ053dZQub0iSjzpafDJ8fHE2yl9PTe6W6H1FpNX2yBnT
IvG7CaAmO9Hz1/B1k9p6dAdxw9J/oTtypFs98aBFVdbf89psX6OEPtjyzx7MHwhf
Yk0ib6ld6fjbQqhkqnBJ+3i80Bly3bH3kAJwlXRoJG0b95yFKJtwvMuphhkAH4BL
dbjZDmDulI1DIXywiMjPvk1iTD2FkRF00U9+AJef1no9IFPrIFKXZyHpwZ422hTB
/HDxtixrIVWJGLz9PvjN7tcf9URv/qb6jDziRvNibXiPWZ9gPElqFIiOsUN8YR+Q
VSt7Lml/oSmH83HrNj2fbcbMuc6e4zMHpS7/nMs5zUb+XUQzeQ6TL/46+8Dr/7Ni
Co+88e14uCI9ysK9kNdgXM6cb1myi7cKH84GgHqoJ/SARdSpW6sQnuNpQfPRpFNO
F6sPz0ZbQsCQcBvu1Ac4grgU6Kew596BX/MIQq2DYv1dJ2PdiJ3ZDAkkaS4JAs0I
BT0YfXiAOLLGmC0/N2jZoN57pKDNCZ2r8UTp323hNK1yTaru8d0YFXK3AO2JG/I+
Vs/EaVd3R8j7VqGvnt0WaHA9iNl0Nfqh3MJTiuczli1OUluW+JFOR4BjhAA6xjc2
Y7/J+ZXKeX+NpDraf5kMsViuz0y72TbYDWEYY8NTlNUQ+tLwrddJkXwRA1hhkyKC
zNUcJ6H7v5mwF3L3gzEia/zLY6fuALaf2YQzvxbTXDe6fG6kAy5ZpxnMYbWZQTG8
3NM+tlwmxg98HcxwUFoN6vGMsuEr5iwnvYaW7TP9GL71k1yId5D18SJNZ4IK9Imo
2UKbQ0FwNLgSHl1CTxdx8O8h1OpJH2CCz6GrXxfWasF50f/zU4+Yg1P2xvc/7mQn
h3WEmC44EZKSlGjVA8TnFxSmJ3bjrGp4Ct/f2UuYX2IxXJ4vCLYuHwTcGc+JcvrM
J3xKQ4RdJQy1Ezk48MAUslOtrJElsqHnyRdoyiAWzp63ngH3riEGJhS2rmzeqIp9
VFDyRv3mYpNN+wagqVnmq9OwIyRJTE4UbcVUO0vBXvF/HjHrJJ4KX/q2HbZ1nxDV
T19pgz3OqeHP2Q8yFrYv/kZp7yZ/gIwsX2fWBQajxnSZls3Q+DvMn0WevYStvUWL
SVSac/Ad5H+iIr/ObXy/OKHWhBRLGCmHMwNRwrAb60DQxlOaw/kIr1keQgwQMS1U
8xuGJFf8YpvkKpOXzapzaQVAH/6xXMokELyQAKcpZStuET4Q23PPMjXqWbxxs32y
qZ/h4I7Z4/XUYVuM/BrBuo/Zpb8O9Vuo3UcydIaP2O2VgwydTf/HNu+9dR6Q7/P0
Bbe59OmvSIXG+Ng/13aWHRUr5pHcm7mEpSEP3qXwXEhMv5GHJI54Y0w1FarlKTjC
5tTKUumh5S5hkFV5CJkh0axnd5HfCUuy0bAw22SrGY2qF5Fusu4R3CnElA0ruMQV
Q1faHJG1GUqyJxy4E4wpM+jvlRpw/uq36Lqjr51d1Hf0TFb3KWcy33fZaSbo5idF
fOK5p/FC3L9pV1MfNMIn1iouUgcTHCtgz8MQi09BiwTpNtDXa3Fq5frE3L+KlSWs
ivr/uCojTXsk6TF8NrAXONArFTfAguK7NjVDB866AGeY3A/59s/Nwna7NeE/mtR4
WanOY4bO2t6GIJO/XZK4rcNsX6oTrU6wO1mXHcyVUSEamoUtHTVyrux4fmmuhsVe
dRWJYkYjnF7Zde6Mlr/DLP2XujEECyj0c8IyFUiNJQ4BhC31e4fn4+GZ95DbkbYt
SJxKc3l/S3PRjIGdCLG0/jV8QtBG6QtEWkqIn4F6nh7zB4TpVJTQwlu7jONcHna8
xlpisAnFphJnQlTATFU4lKw+cFPU1Fe7h9vDbFHAPli6abeYC50cKS5YMUKKYDh1
4bBtKL+ENJev9hT9fO6IblAXLR5LUQg4pPpX+M+vl37mLMi3ezGW0WzKZQIdQ7pM
n48NXCBwFGW7ElzUfnSV1q8vwtTXjpGcSKm5cATTyqwGY2/3xIZlNrtIDAgzbjy8
095nrSjmLfMRIRC7LNBOwT+2bpRYRivF8k2Eab9znp3zfPMEOVX+GEsMps57luDM
w3RzKTVGqaFuz0J03X27XPYCGq6dm4TJjGrJxkNoEv8Z5pKwRuJom9PT2LIS6fW8
D4EBW0rFQtbtxUcFyJUNJhaG9YDGWANNJzFoMU0hNyg9mQZM06hl144I1HE8FMl0
WNH+t4DHNNrrbjP5VfJ5Ls6u+RDPCwHCh+2YBTRpf0kRIxToUM5Uy/BOGTw4u5UM
pc7fj7dXv8eeEK4ZGfstNvzL6ur68dMQsjZkNZ4BpqJ1LcT5BFLelDY1GA1DYOML
VoL1SosQ77BvLFD6wA9E4RI0yEDjkWY7MOrxf2ZBW35NWKpSWPN6QmT0s2hfr93c
8vMXeUxp3GKzIYbzEMmHIsmvYmw8W8f5v6wekS+v/KMbARnoYEW2I8Tws46OZAcC
xtNBZ9Uyg2q8ocm1A/w5DmLAM756FKVH/ASE+jMajJqaZ8UkomVJ0nM4Rx4OHjM3
+mncINAyN9hWc6v4ukX93OnF7WFhpYqFWBtGi8USYepCNhFycLeDip8ACTAPSV+U
/0fhJtThN2ucT14ec13aRYPG/024FpP80O1Eu1/fMG8FAKkgPxBSd2Tbcp3kTtAr
ThMKRqbFTwb6QDhuXGdUJmSB6Sf3X87GJ0IkY6snRkusrCO+hOR6rIiQvYWOm72e
G9YxzQO9H7/TF7w1JLKWQcpJ+BDgG/2uPcezlTeq46pu6A10LO7R9n72bCOaKla5
R5azm3COV3fO5cFB43+Ko75w5Y7vzQnnfN3F+3IWLCJF6A2QQjruitp1+I93Y3BW
WjuebYbf/3xPwH+llObS5hL1VpC77mQUeTrgQIdSzbSyRaRPX0AVYjaw3ShtBUWM
tFpUU/wSKY40DBUIqHk9LUbEF5rl5qdwhxdN8Kqv7z+vDNmzB4m1cQWktqv3Dnsi
sAGS6fPbHCMPAodyUlKiz9M67XjaPo3nRAY89T6xk9Ly+BGpv2fCmufTarS5G1zk
Ne6ZSP7igimOCNDGPuflinT0e5T2B62aytPh3nv9KrPPisIT4JdJl6taDGD66/Lb
VWFz0TfiObWtxT33fS3d7PAjPL/NaqjfKbdCAbi/3elhZgGL3SpxbeqLThqrdtuX
BakXcr7IP/GO040nnx1MIiQhuiJa4KJkp0EmgdroGg+iH+dUzzOpqpZy0AaaROWX
hgkt6wybufyTwmBuQvKT99YLfQMuWSkp5kUvvUaK/B8lBNOWCYJK0KEcb4or7ycs
/3MadhAF4+6gCnXqdXJfFcGl+TymWrTZWSFRGAVISpkqb68PhvpHJw4oJ+Y/uQ+y
8FyknOA02zUk61yTIXmqghH4MpSpbVO9yTWtipeDAnnNRUSwo6U+MIYNpKqK+Dmj
Lz4d8xh4hQBEsvpUqAFBjZSSQHr7K6ai5wWkSZ1jWxTPdQPjKHl6jd1nu8UoL3jj
CZ0JG3OSOhFueLKPznKsFfESxr3N9ICb/SGKVVN8LcYQlv1VveXk8N+H3RkqEmbs
ez26Mgv84pKWm83XOrs3k9ttIuWxm2ick/ca4gicdEL3fS/KWrqveoexs7FtWYJ/
7/c55HSQa/5/amDS+lIh9WxqIjp8ltulxKkaZHrvCMYgsA0QLHGMuf6MbZe4T6rl
fwnEghA9rXpZf92u/VlGfKUXWbwZpbS7Dd/weVE93Jh2N+hGSqwSHpk2eX7x0NNw
OKksrYR2QMSccHNzgFCPMtNsIUwHNf7bG6ui98Pk+tzrMo+j0udq5GnyQc02+8FQ
aUoSPHxSBH4RP6GbpgIQ8NscdmDQmJt5FWHBZSW8lyTyJpVvEM6gc8/gziXXCL7y
DdbLyO+l6S3orJb1RASPijnIb8ubejUHFcG4lEZ8uPsw+5SlOxTqtBMZVMD8qNjX
yjHc85lSoED3KoY0XQknF08M6yWMoJbDQoo86MYZl4Fi073I/1awx+BBpw94sU12
/pyTnK/dUzX8TLPu2l6+VmuGNN44SxQyHa/ZK9/AJFy1CRAaNF2rkzryjIwkC2sZ
pNRgneeeNUS1RWb+9HDxc+ZSatjyAGDANYkTVQVeS4160dRzzGft350nWpBHRpaU
d9X0ZHMPk7lqwUCqPIu6jbnslTeSaJxwsTs7Nd/rbm7JcPk3I5X0LC46subaMkBd
5n+EC+xd0XgX8hZ3JKfbTZYoA7li8GpbHNnwmdZyVTVExXccSgpOogEtvH3RhX6R
kIePFXPzeza1iDlG65N91NMyGnh5ZRtjrUAMyzERPN5icQbcQ0jKiWHhf/Ubyxee
Bp84EnC37lzoxbZnp/D127Dnu3MugeBM1UxvjlPkwzaphOJnhlQipXQ2lp1MwG6r
A/osL6wHNSWrHkAREnGnaKyDMs6uxKd6by7p/u1kAf/pynzyG7q9e05sJmS+/Ktn
5pHIs0AieFNilF/Hts/7msps1o6ToSf4gTVSRYHPcH2bnY6NCXvMwBaQyNoFMJjz
XvNpZJwTk+Hez3r/Ja6sB0k0pXHEifPpbRN5/pDBMgQh8GQqLNd0VX4XEE5StM79
vCot7agUEXdaO+4D2XWzdZCdHNyazwf9wrCw8FDbX1D7d7JYfgMud1DMf3AkjEnE
EYQtTFPjBhO1kkuMfepIxjPqNl1I9J0fs5eRppX+UH41UUSi0Mw5kiNsV7mi/Q+P
TdAJaNziTfOOEUW+ZO3jsDMEk4VSmhANZDUaSsFurLrBATvApFbMExZMFEmpNj04
rs4whl+Qok96gUk1Us+NXz2hHCI9K8t1Bwr9hIi3VV33Eik2pkgF0pc/EnZaiZlg
Ebrhpj0CDnpEFvZOua7yS/ISdEmiYd/Y456i2w7CMGI2gP6Xo4+Y+mTuJY7kcFFO
DnoLj3STIYmwZGpxmcl2hNwe5iBg/QvOOgBFmoS0uNIy1YH/jNR5EZjSY4p09ynW
C1NUCnWUQ61a1AYT/PTGwpiy0OtbNeuElOhNDNbYfqcM7mVsVo6eGVEOOttttRoJ
Aqyypct6Ol0ybdrfne0hPZ3wTocJtaHkBEjrRHC3qpncYuQxVWe4ToeRSOYO6UJk
yXREU1oJad1qiNnFXmEml2ulGV382Y0W5FMdHbDUTy2ICHBaDR1ELO/tm6NZq+0s
sCzumfUnRu0sRa+fyDyohCGKTMdwqhTC3KmoBGfGg4jveqj5sBX7BWSMKoxyoJgb
IRlRAE0GXlDIepDXW7XZCIwJVlrOYxEIwJF3mOZed7aLPKwdcxhv7AFTxkGFpoqA
M+h/gGw/EUxlbU7L4FXXWicA8f27UHJ4nSYlvyrROx4QYGoTZnhYTFjN7XkRztDN
dOsY4f3CCfTBbX2u9k4k3Nt+EZd2PEBpMO1T9CzI1BmBFu/8xXjtllV76NenGPXB
P7Fl3QSZ+6IJh+tN0rnpfme5s2mS1PAgY/gGVA3AMv+RCdartFYH7maW0uiiUqtP
OIHG29AxNuabHh0yKevlylHSCUH8S2VhFQp2yEISmUO3eHI1GBF3It4KVwa7oiGd
BEIQ7n0XkST3tPbKyhck1zfLRioKbHdz6GJCMws/teSNewszn+RBXyTwsqP+ch4i
uo4v8QiKBLLE2svdnB3M6lC4dWlt23Hs6Gf4GOxRWWdXjrXB8tu47zc0UwpoDD+K
wlP4P5zqx/F83x6t8wdHu1PZj2qAqAx2G/hGhsS4mfxH2HYWNLWz1dSVrBh1BOvZ
7O2MqMfRRvhSAlh7qdAwqkAYBw1Xi5b80WdkiJyU40JhNjewhJdsU0dyjGRdFmUo
KDIuCpKdUoVP3qc26mxpDDpl2ODpDH96hXE6QXNUXT446izl4OqDX7k0hCWEcEk/
eSISJ9mb13wHttoYnBO6NNbRjfsn3EsUCaa1E9Ys8CkHbxAyqOKz0MoWjAPJ8gmU
RpRm19S1sdOG9/q43uTgdxf+SBwsrSGTUvttGXPIxR45bnQuv1ho+FVJjD9cpDfz
bujiC6yFo/TyCIQmaUxwxSFXmZVdNirfmhqfSHWhDzf6V7k7F4N3VlkqYVbuGp/m
sFcRiJ62AQBI18Xb/MRpkhPzfp9ySd3PeMSY9GwMMswOTqTI6EgZkWERIqcH4Nhj
m6txSqSTYHdTEr8F+dHCCTxEsuulnxOHbqVKNSc85F+sLtVuVm63ealvewKLNSH3
msvYUWRnkH/ynJP9RoR1sRXlUiCoResCS5dcoS24mf2vvpFe1+VPy/vHL2+SFpFA
9mjZQT1JCtix0sMPnO7KIZ1cr/n1DBcpfUG61phXfZVTaO3jj4vPxjeDiJ1iUOMY
cTW5U/UDUq5EWFUPJ/YlzHcxTJsaZF+BTdGrxRGN/ro7AAlywxfIEGXGIHqNhJFp
yB466CQask+M5seOu1r+ohCtSUk8zSowaxIBxHBlMlHokUZSxQN8JGXdawB3/FqD
59LEV1gbrHXOgthRfJqV9Y54gxmYo8a4Z2DsB6jd6TXpB893IGi4LDAHoKjkcuhH
OlUKU995FBC/VKopNYibEOYRN8bfnILp9XiE45cj8nX6+QJh01t+GYm5+7V9FrGN
OfT9YcVMYB5lZqyyKDKxcVKsXVDg1sp9hEYrFfhQRUlfHDFpL3VexDlu5Tpbbs7d
khMH8/7HcvKI0Opfrt7vBlfKJa6qBljEXtylwkrAZGBOrjkMDI0OtZFBW+9t0s22
6tI+lve9Db7QzlQFZS9hzzlLGOrUHNH/JLFS8rctFNFVyVo2Vu0JXArg0sGfo74M
9a1n6EiZ464IKd9Xc6DCTJ5idVEGc9lNEa1qlHZXQmveicMqJTAxH5Dd84paNmoi
hFgnwMlmbLf7mL/SPIPHDigmsUPzl3nsu8xIevaSrWsEKPiKr1ujHXqtoE4goOv3
ewIV1vyi0oaqPjWVdxGg8TGV6wxvHmnq+UAUmljX5atoTO+YLMjm6N/Xl/gx9HEt
a4pvBtB/KjhkSGODPH+0eC/5D8UBjUDR7oOBjbYqSZC+Ao6RdsnxFDAyJqqqfrUa
1SrHC6k87Qm3SwvQrSNHRrgn12L+P5m7aIGpW7wHp3uVMDwDaPQDBI8SVu1IbI+9
RPT9Csj1CxKt/jk+iBHqzUnnOwnCv6VKvkllYUvOHt7JAdnq+iLkfGkyctZNuqBu
OJJEhv/FaQ+V6wApmBEeUQk0N24/wgJQHEfyAvtpl0gXcHGDNBwdCEc04VpmN7Zw
MZY0taxpB4eDRWvghhVpkB8eblY2VJNqgVyJZr/Ly3FhyoL2jsoOz1RXTFSeRNUL
nVEBG+w32hd0893CgBjoJ3r0cqEW2fJqjNsV244Id+X4AACrjm69i7zxCxcrLQDb
3rFbbdWhZ9fDNoeA351g4O5WjD94JgS0vTKhYxsggekKrTfG383w9h+QGinnA3FA
z2iLoTm3dNbyLO7hswVprOabH7F6E+LXFO98x7DZeVhpLsBZyvD/LEQPi9g/kgZT
gdxrmhKJPVsGixGMFlniaOQ85WLcQpTpxb7SzDzmF2XbUE1613kC3QR+cWzrOl/S
gi68O5mXTgvsG6bCaEGA4LBWn9DU3th97AH0XFPoO/ETmohN6vPcAJR+cLUbII6r
ttnKR4Rwv1KsEq/8dVri3sctNN1opWK0Bn55TSudX78VJb9eZjQB36BItYOddvJk
IHRLxAIRDwMSWOY75vq6ofxkuHpUdutGtWZmnKycpYvjTNi8grb/MT+kPgXYIqLX
NVNwILLx60+KLmER6HRYuB15suoxzY8sA1DHf29BCiCLxmIBuvcy/EvCfv23OHxX
34qLHM/5EyHEd25zCaH3sTB7LFEOkyMQqApfmpvISNPkcOBH+dknfiKqtm7p2Vhf
jco0UtH2Adk6pEDAzkx7vGqW7cV5Pp/JR1B8q1UIwqM6z88w7OEO2rdsoATiINW/
aKD/V6yb2ER1AdG4IURA3yO0pmbeGOxqsRfUB5VwPFPDbURG2G2vJnBLg7cUlq2R
fqD5bpZ3slIcJFuFVfQFdr15VI0AEBYDbvsADDu0OC62z6DLf/KUPQEIdRGgi8gG
cwSCIl1/GESrjw05cTGHimZqHACLCiUuulHqqPSus/UVxzYcCR0aX9J84vxMgSxT
rEzXWvl859mttY4i1iHxI2yYowAK5aTHl4jQ/UWNRYrgoBJp+Smk9VaMtjhWRAIj
p23W9gw+sUVlpuD6JoxwVVGWcAtV/2VTLgjztk8yE+XNsCZBfHvk3s5A0L5qYRNP
rllKiATFlbqXPH2iLhvPhFTrYWec9GYosGDjxxUwQ/70CXBP/whxDeICnLBFhi76
koz9WpTyVFy62OqE2l1D89FrdvdDyghSfBLEpZIbIhhNNvwhCMomjZF19V/amkpY
SpUhZ1p+DnUvfrY+cl/iYxgkF3zebfBI0MgWShqYlooagnW2U5ubAl9K1qbBeA+S
HtqWezAEGD4XqjBkDn9hpCa58EkWb3QBHCoN/4ktgX0UKdI6ClnhK9PHuOwy7mbr
JQU60cpvvMlnst5C9+pOL1rGvyHk7f/gUzV0aw8O0w+VeDOy1jVw5/1fjwzeqq7J
uGO9NbMrdnpS9xceSeTIX9/vBUoP9UTffg9HINTFBBh+jKiWwdO5TZ8HLbydvqcI
sGQDsUN6XWy9CQMtwbty3RU+rvKgiRrnpWCCSpXsaclfQ77aGxexcNZLdf32szhX
cQzgEBHRII/Z88Ntu9HokUFyHR36C8Zrj79lpjlUz9yekp5a3/jtuqkCDlUhWSMZ
gYt4klICkiLR3VQLVbjq9KjWHasoH26lYT7jBFTRoljukvZrG/0gDLOfwsQdUN3S
Chi++uTo3tVben1dV01y2haPxTiJhnKs76/AGRmPs/T3Yqj05JQWcqMqMjmZiuLy
uqx+CBaRvnn/GVeIpAAf3KSsf1kEWUg652BPlE/Icd/fLGvaWLVN0F9yXvcOxMrU
c1cFZwNBpNN15c9SeZ4/sjf8yFd+u4nX4JeNQIg2gUUUQiUNePRw3fAvjDUIdaC2
yKRTPMMlsO4leXezUZC+s8KeILG9q5IkvugV/k1me49exIyL45XG8IdyAb6XJ4i0
ec11fM9OLF/smbEXYgmBbFr1xB+RBNT+fG4NMXlA+7flcDvZks9Z8XpktS1l/830
Z7PBHmKIyzOx5G9vby/3K2qiyn+avtzMoVWp9C3aexULlpVF0YM3nBCurmipjscL
Toa+muORusMriNpVBX4nQXIhO1mwwcMj3CVk+LIg/6EMX+iBZ4CWqTrUuUCx7eWM
0CNO54Tn7Q8xUMCao8vf48iZgHxvomEcBbaRIacTHZ9nJ1PE8k4vuxy9zSHEr0va
i/ybjZEpHnTUWjr4nsGtfiqU80HJbJ5I2OemF/pu2UsG/Ouea+yJs+IxgtpdKGR/
sfW/PbTSuBFbU3Y9XV9fnQSnXSlcp0PhswXRbMY6aMp6APYmQzdhB5q0LXJGIimR
qujjyUzpgwmHjk6DUadEitSskR7rsgfwhwWLf7kAU9/uWdc3QQ08mnyV3NAoI8MV
ZpScCL/QAz4tqwnlBFAaA+0JZQXJjg5bqCECmUI8ZaAHHDWlsDBEClkpUUcoivLH
lLKPk6WaM430Cpn3TXFWchjMKR5lCocDke4Ng0v7pKgBhOznUmDhYpLyAPMU0PsM
1qqx4FXhKAHthSIXaW/HbU3nVxN5uoeWL4wJchJKWM6SpnhJ9D+D5edUoxv+l7KV
T+5nofug8R8WNbg1YnKgELh4N05E3P2uKY6YWaFRAPst1X6Te295d329ePzp635e
64GkT+ytamFB163qo8bgmS53DlR7x4cx4d8vrUSI0XWrlVkMrcMK856fpdclJm7c
oRqp5+h+FdtLPxXMs4RXsB+SqsBj9sn8+p/eXZduHjpNN/raenpc0KAyUKdZ0T4S
cTEKd0EzddbzGcOkt1KvIjqVZdvapKhNTqnXslPbuEAd+qvXFafeOHnhCwbUsFa0
ZWZsO8nVjBte+jRqUEXjfJVU7XS/CqwcsbWNOvUQD3LXIg3clmbj35boLNFcGF9K
3N2LDJPTuuTViMCb2DPn/MP/lBgkokr+McH9+B2mI5YbQvS9vG5iM3pxhcOC8AtR
5bf6ccU0JHyi95D7vr+B5633QjrFWJn+XFubpURuoExNtCT2CKoFdXlIsvdWxKKD
P5FcO0NpuUXBCIvAaTnyi22PVIZmcr8xxnzzcmDuQ6Mq+17OP7R+ebocRvRL+Toc
Q6dE29U4LKj8txG2pNfZLX3zgoGVWCXhbd6ltTVoGt3g+Sx3EGFX3/TvQKqjZCpx
/j9NA2lyi6ANgYG81XpwdK9v7/DGn/ggVeBj5XAp0iWmotehQ8NrsOhi5t4VXRJV
MxUkFhL1LigmYoaOHqMFnnPJvAqB7XVJblFwTloEQfVKbBg60kEGEP4Nvb0jtJ9C
SAlkWQiBjzPqXS97DViY0oi9C58xdtEGxcdtIfVNe7pQ/3QzlkP7QOnvYVc9O5R7
KH5fF1SL6e/Kmu6j4AynOR7+f5w3C6B4du4s8Tf21ZjOeiNYiqw6Him4xYDdNoCH
ImboK0/rtuHzGK6J7ASroOdzUFuEEdnXvc7qe8gD8ztK7rHf5LRWEKTlV6BiJdjN
SdCy7zOU1pBXUyJXBbUPiIMLfR5eB0ckfrC4L8DCMWR6jPZoYBIT1wLrLzxwiE+v
9gheBIavTJKR26IgZalUfDFQMXHst1eiuv92W2LjZ3tlyquT8DmduY8N7P/6J09Z
E6GQR/+H6QTllpSs3UkrmAKIm14Y4HXSAkgLHO45Xl6DxE2juQC8sbZUIUOKS1LL
oRzMss1p3sNZtPGEf3F1O74kL+6MXOR6y0T6TwGfjLTzeeleED2jgkdyo+H2S6+C
vRmD4zChp76ni4g5ehAPDXcjBYBBo8ml3mND6Vk58SzAK/92Sicszo01UHoNh3+G
FhcbJzVwrOGfPYFNCzqHaKner/QM33gN1VhPiI3MnFayBw4tZ+5nQ3xB1tUt7DDj
5XA+zjDCGaQ77Tq8KrQxTyQC0BYYRj7RpJgw3tWIQetZY646FE17D7ZFPK6olYIp
H0DDXTm06ptKq4bxQFAnyAMEUG3FYqKWZq0oQrH1fXuvsn4MJDUPckJJ7Nnwd7VW
9lyIvvs7eRN/LaACt8SOt9WePoF4PTel2sQo4o/eiDisSqVEWCWsZxnm2MWAFXSg
D6x6PnNWGAo1femWV84pxO9dfFfELMWd9U+6XRA/Ew9KVJIwjyyd5zG7AShVaxSy
dpWw/DwBEVndIneFWrnZBxrSWeUJXi7y6yGkInHDT18D0VqAukeoMBAFKWovxE4M
f9NXI5mHnqn5O+o+GG9mDCoUZpKmVhBZN+sJ0I6POPB0EPAp6wRcKUfgDCQS3+Hv
SffpzbOwJfjKh6bCV089QlvnMYZiVW/mP6TAPLxD2pOCEI9Tpfz+Oy3fE9JRQtZm
Oos7P7UU+KciWs8C2HFoZHhPh/Uediq7jCelMnr1SGZP3gbHYFdxMrISZ7pbZ2F6
PwjXP40EM7mFVdzkodgJgqqazpDRXouVHd7tIla94cFeaBLYJlnY8lJGIyjzS6fM
z0uj29LoME0bmFLTefheLDVJ5Phn9mSoeocE/LuEUNY1rBJoafUB1udn3c5V4oOd
+pje64UQU/Z9Grtkih+oCtz9deT63CD8t2UIrRvuw8KbZif0e0M/bsuzetYYqSUT
Os417hmh+Mk3dIaNL43w3nLvFvTeGXT27DEX4eBC/KSHkwcz/8zSoXmai5mFn9gd
/flaOQ0PTWUfyF1ISBCnfrUWMid2imeHMqC49mIODdlPT4HzpUBYR195cVWbboVv
efnfwltv/uBhXSp0fGign5T1d0frOQ022vjDCU9dCbbHun5qRJiw2vKWQCyr3zna
zecjAUu3PFvEax4zlyBUxPbF/f0MnAr00iXYcfwobxxizU0NiPdqU/Rlg6bKTfPy
oQAxwI+zPWuWw2Az7+VHxfUwkDwWt1p5L/EwUB5K4lG1B2ytVmYRAkxsJNeVopKi
Vk1Juytxw5upfbfBwYyBLCTajB2fq0/Ncn/Qwrzcax8fRdqYswJfKWAMDMJPxZnM
b1iIhh/wvTbXRaoKtrW1rzPN8nfyf6MDoIt1YwEsluBvmKgm6qLg77anowJZXnyy
fass6w6GCT4beijoYcwESQze05pzpnxG1ZMzCTjdNL/aYPbfPX9pa5MtnYasgCsp
t2OKV9vWD52OpgK9LPEGz5xlYCAMPEsQnaYgUGDGwj6MvAp64x4pkIMTu5iKY5Hj
l82NRd+QyRCOxmkY2cmv8qT45T91OL6TOq+fu8jRqY7bU9kYs8eGKaN+6rkChbDT
BCEQTL7TdEKiPYAvQI9917PrFhAPZoy8mOGes1fhg7qc5reGBe2UfHFJors2K3nL
lO8Q2xCA7jkh+enNPFVkEUffAJ6B6hEqhcvR2L6T9Qvk5SlIreYkh+omRUzc18U/
P0yQtlFAIB68FsAh1uK7chrxtykl+DNEso8B5uCh//mD7BhfzT7Ch6Re6qlHfT7O
WSI0XjSxf2xCPUZUwPP052IK4+NrsJA/87so1bpS0QGPKtEFEJmETF0WykYDt0We
6UVgArDm+g90BEptVytA7ul1GHCwvvQ1x3SZrx24Ok1Nnc+/nk3Ct0MVAZAFT+2b
tJ4K4gDLDAHy0zDJh+p0eGq3c6z54XN97ypDMfaXxOt9AwaStEx9PGmlS6uPm7TV
3v1XLIXDRKna5P0CX1RJ+0hxEjxkhUl7TW5isWf+2gfeVjBJEEjs3Ms61kxauiy6
RdDMPv7BsSu1UMbHfg0+szmHqyk45HWSatK7/hKMa/0GA+g2mLFyILA3chdQtuYR
feucgKZawsqqa2BWc/DqW77LVZCFCZbLAdV153N8VzkA5NJUhbuWEvF4ypa80VPN
NLoZdW2t3MHHznjskqWX3FMN0HYqR2W8pS2a0Wg+VfGFoHbYnL19hDP/WKKu3vQX
lz1TYdIEkd1UcJhosKHng5qV6t3OL8pjRpJOViPEYBzd56+BvrtW34HLmRnmspuI
qkvP+jtSBkWZYjwtXm1ziwj3lF5OP1+8N6VTQXViGswZnIcMGIwO0at25pwBHx70
usya0Oo/i9/CgAkt2NhysQymwQ4D5/JpO4/rd55YIIH/dIzVDFO7UQkV3krU1xgN
JfHvALj+nz9VqfLXEzLV1RPOryXjrkUCqJMEZQX5XUJ58BAqZae4r4i4LjGxX7yf
I9GbIojbiy+OXdtOJSIMjw9JvyFaYsJW9XDM/D6FZyAbGUUyCUgAOC8AHkDcTj3j
eNDSvGjKXgS5wSJ687E4YsaODIB740jgIOkB6miI/QRLkLjyHWJfJuq7IS1hRwu5
0Cl49bOzPwgAWGU4VuIn+INUKmKBqAReTPlifo23GvmxZiZjlLjSeMw7I1EDmO9U
9wueJe3Xi61+Bc8swWS5uSMx1rq1+3v4RkfdmU97uLjYMxcQtjA0I2TeJ0YYaKEy
d4sodqGkb5uCgwN2h8b0tfD7EBlFqdIFuvbQtOX/h6+3f69F5l48wMdFJqGIutOE
T3ILUZPlAS90tfZ7HFxzb6R519AkmQq39BsMqdYEsz8eo00mc0N0wYjJbAFdLLWM
lzEIMRnKdDgZVaV61pzUTnQfjvtTCuo0S9LFtsC3akIQkdT7ujNAZHeogREnIuNU
SZ4EkTsvXUFVzjOxTt4+HaBnBqLNtzAJDGN1X9MewvKCEtlquHLwR0KlZLR8t+TB
x6LSG5TIQaepzTI9agqHE4k2nL1K6OwPXm91Cmu5RbwDEOnzSItZhI6SOnLbE6gy
4HmZgv+Oa64bcnRspofX2VsDlbJRtxk1HnIEVKZl417Q4oRmNWj2hT+I4XkT/M9B
qxSFrethdV5fs7siRYbepqz64hdHOJ8Cti6gq6mTCM1X9MH4QVza8ShVphjRTQve
Dvr+VeER6xCN0JveLDpU0Q41tvGZULjO1dLnoSjeDP763AndrrrTp26UB7syglXN
fKL9EUFfQyANctRjLgnr3c5hoFOuhuOoQZlWsvglK1OatWgC/hBo5VIAtsWW3On6
sDb0c3YK/WHdP/nII0Lgptoz6r29FHlCbP2J1ntPwESGbrbloSm9i547KdhZ8Diw
8Z1bfOyD+8e0vFLaUSHRs+TuogVvOwZOXl3Yf9uWoTuOW8OserW9n3PBYXUBM0nc
qIXQ/Y9/8k4ZzmBksu5h6zHLpTia200k0ZDUNc0XrdZyhyL9/PereJrGt0P66p+x
WnVj41Jd0L0H+E9ZRtMf3myBCm5FffvlCGFZSycVAMAOkKsTmnuX0GMUqedd0PhY
cIyBxC+5lxdR+dvVDksTdVKEDfXaUA0/MxxvDEg3M4154PZSZCZWlN916YM1fqnu
E+6GdezCBmNN4hWIjd5ki008SzOTIHkI3RzxCStNqsUW+R+PS6sVAAdVRCzZSV/d
WUyf05fZhbV3ER0wpL/GcrmU3yOGj5iKjt2G5RkoX1g/Po/pp/B3nZJdqSp9V6EP
Mx7dqjc52QFNX/KtFPpJE1t+mrL1z3uSlUKWzETM0e9/DcZB8mnBKUK1u9cICFWr
B8AUWuy4I4gkJcw4m+lUPEcuLamjc/xDf2207yIFmMEQu3NgKjNCLEDVFDpYrA82
8888PArX8Grb1NkfCp6i/Spn9eSHla/DwNDZ21SxdBOYn6jdJB0Tf2YGKXNFpJtb
cU57yXunwpbrzMffWAmHtG3LvTxa5fRjpL77RRFCElxfQ98L87szbRdugBI1cn9p
88eQwg45SNBmKBseteu74sIbt5iDJ1SrMRZ+eLJ7+p/XI95L0BCy2YiTY033zhm9
ySYe4+03DbWhLSzBftTWzdjs5lLIbN7vhe4hzLfxF7ZUm7Ojx5XCk5QaKTkD8rlO
PQw8fJOfLT9Ug0Po0sPyUzVtxd0YZ8O8vzI7+pYBJI82uSKcrDY5oTndXsTO1NC9
lhlJXl9Hr6nOjXY59gdTYfDNmHRDqHDjONnOyHc0UuUcF6+Kv9G1yitaGl35g1/f
82TgCowX4bE5TlLwAM7VbKcynHWimb0JA2rpYzT/N+RatLX8UdIeGtTK3dlLSRFt
B7K0Bwe3ppbMRIfJc/tSh948NyJ0y7nPEzLz+BZPfGeqtI1O42ixVgsEfrL8vW3K
agRwvltKwjUwIaaxobWED3K9tCOkNshmFZ8yQbZvPgK0m+x13b/zRG3vG3+ZZVKe
pf2czw/Vu88/MXkUA54IaCzr5xi5f6FVuky5G+CZwYFHGU/T/VYEmXaxrcaIhdqI
k5wiXvtNcDUbZstmJybQD5zYSFbPCqgMX0S6kFijAGtUinH7HGhRI685RGIgUl1w
twBqYk2lQ5CRMGhIeMdOP6Kaa+KvJS0H3fOSsKLbMCY6tf5QYdkiHKUGZfNEQUIP
rRyU2IbCAzGoyti8Lkll5MByFi89QTBhG+XmNXOCc0ESkGtK4XmUUL1k0s8djqQn
gGFhqr1QqmgScu3ekvJ0FYzvIjzjHRF8a/EuGbcQ1QGrA2C67oGgbZuxuoWjS59j
cNAy5+Muku5qHV592s04Zl7LWcUOrNllJ+sAH4zy/lMoBVDqRhtnWdusBzLi1Z+w
k6r4Fc5mu1KNO0Z7QaXzIX3c0EzZLcDOmUrujmJoBKxZPAgDhJXH4RMOO/q8TLyW
Bulu67zoOWkHNXED5k321y+RwW6ahEBB2VsKfavfj44WGldrAiOEOBhsqU6Gru1o
/lr2HIf/tDmGh5EdNTyZ4WKOWbea4dCLfGyFC2CxyZ8/k6rVMi8BW6xCMX/awzor
ypz+X1LNa1tAO+wpDYMCJhU+XfFKud1x1aZzKGPhhMNwEu5J/lgzfhXtiDStVjHw
Ur4G4qMCgMrb08OHS47zSFbpcXwGjHW3K3MSAC8rYmDbim1IAR6cYnJDof0x37JE
aD3Erdk2G/ddAlVF44hqvHH/ihiEoou+5wLxvTrOLh/7e5n2VzvNEO4ZojR8rEAS
wlAE5jGXVVZDaUTolOwkhTGc6ybaPwcEkZkb6i3gZbA4lzYWoSiaQj72RLEVpvlH
Y4wQN/AenaNEw14hQgCKISDzD7wVfEchryOD0/CHYs6Jp9VMQSA4vb2iINhIVRNb
Kg/kSrz9QV9JkPbD7zlcyMNfyqjybK8Or/Qcy04/35Q2z26Qq5/OtK5dS41DHaOs
FQDZM57sKZipumO4pIAZ3QeUHe7hzobHo3w20bt+mAFZbigm4VQN7L5AD1nX8YRl
wKx4I4n1GmkghHL2cxss2R4Yl06DK27UPM3iUM0IZkfqcNPcevwxBVtHkcI1bw1b
5WfSRNk1H9hG0bzuCaOa9JXxugSWydMDzLCFY6gva2boLX3RBwZaCCsbltJACMD7
YxwRXlI9i5JuO/6ldFAtvP3zlDjStKvB5lVg6ah9BEgsNlzjpf1TCJNL/7y0rnvU
TzvM0twX73sU7zvVrAgwW9Qbr7C3j2b0ivMzyKfhEBufpkGypSUMt9xQckRURigE
f+STPg7QkQDvmEI3KqtU2Yh8n2qfa+YxbC1okWdaLV+hB85fHSj5T90jnCbo6xC0
Xlp6YyVNv1U+Q5SyeDKeNiheUvbc62tDRSZORBtcvehPXaV3/NtyrMyjkT2TReyk
nUW8yr69fhfF2XA9xWahMxySojw9xPg4X2XSLNjEF0JdJXla58Uxxqe7YQBCZjJu
JJHduq+DrjQQcLgsLcgo+wriiujz0naUv+AZbKPcr8UYj2hIuLlhFDHxnA5yIxm4
vW9ID92qROlXN7TCvh/zizgmrvp7O4MIM/3AWzLLEABWYr+Jv9yzEwnBp5leVjkK
CEBOCfWCLWP2yDPv/F8v4ZzzcO00Ic1gRHGzXJO2jxyk+LWFUz+dt0e4m3KaHQPq
jIguV9YOll64qiIIu6BXyK8ihheMBcKjxsyJsV2ofU5EAS5ihZjZbCtvmVCg+E8Z
DTTiYcg47hDlTIov5V9HMIBitgYiE0EBzrnQ0SY/MFsces+qTtlc4HZ2zXsBsbbt
h2obeM3FucxI1KSt2qXNSeEw9PDFZiSo+I4+pazWE9fNGg/gRIx1LTszV6MetX+k
KvUn72WXLcGxIGFQ2XaqHa7CtlLVZEv/iHrgXovd1nygqH2Vn0rMzdp3W33wJjAO
ur0kSPQ25WcakTKJBg30nFyo6X+ZIsOJGdVH6CyVwQp64cNTZL6ni9/viiWN1CaE
oBlgOL93oPACJSqSaEbKhfMBBkTfRSgTJgWqc4kQMtmOTWb2fFZA+E/M3JUfbZpS
3D3lFqmXRGK9eF78PRXuJ+Fb9DsLuumsPiUQTfiE5V0xRRktdwIc/FGHNJVcBvgf
HcxB6/UgLui0gQ3IXBbRdxVMmImteG9NvJr9eMLRmCVPRgl9wxN8NYZt89WCha3z
bB6Kz1Ikjv8HpI9JeyLhW9AqH+31BcHKcBNfjWEoxi+9gmSCwqc4eK7E8CjCLZpG
Jan3vBHA13h8RBFPfyunT+/jLF2ygFNghvQJVzAXSHDFspSS1ND1V6oieOmgd5au
PVxgXwHqeUkOD1e6MVH2BbdfEufY1Ru1oC5NenCVoaEzneo6lTMMb1Ls82KRcQII
56KA34+XoYJVrq9EMWwiDlJtIA0QLITZgv7KB92nORA02n7jVWAuOMHFVVKrP5/N
lD7ibwC67066XTIWCTlCs/zo78Y0K8gSS4qcXwO8cWN1kwHh+luoXlxJg6olm7TK
ItYu8NbvhH6hJpDOoOQG7IV+Zx1nB139OD4CvgFIqFCAn5ifCRyDmuAydliREAHn
zjAO/4DZ5HlkrvCQ47L0OJbwgkfDzP99v1ki0HDT2EbARKsNP2lPeNLoIEzwqHh9
FUXJ9jd0bkm/46dO99qVg6AddE0pJXhU/OiaLIOv3Szrjs2ZSFoMQ+cSzTJ0gzY7
dsxk9Gbq+32zP2HxbxTrFQ==
`protect end_protected