`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
ddtXksX2+yylW5zu6QL2Lhnb2d1sD00763mmSITNX595NcHTEkwn0zB1Dry37fOW
FufOhVzEJp80NC5qZ/+F0Vk7Ik02dIR0elf3clrjeJRK85K4e3Hoo4xn7YbFUIms
l/8VZSb14+JVGURjfswrIyCUotIzlzVYZ6gzoZwDXIi5gQIBf/gI+KxNXPaKV+PQ
Ufys/12rjO6aI/pPlqSm0hCvftmBcnezN2hk1UeXgOIuKZnogjOsf0iJVX2aOOWE
6pD/psybjbnsNB6kH5uFTA5frkzIzkzl5d9+YDm9OyC+k84E83I/7/j+rk4L2dah
QJOvksSIzN867/4Qt8qYTQ==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="MvBXkzurAa5VTw+1JJ70nePUfoQXBvZOku/SMmg4TwQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
oRtzZL4VJ4iwysPsC8SXYCzXS8Fw2gtZTOskLcDV+1B9Nzn1zTyNtlo6lNICRmmK
ZRVu2BmCc2G+fmzynYlNTnSa7C0Cuel6FYpxCBlOuk3OF2tzAmLAuDyOH3Z1Yjzk
a0aHuoCdIRKv7BrZCdALt03JeUmXKPdOmIlkVGFl8yw=
`protect rights_digest_method = "sha256"
`protect end_toolblock="Jn9CQpRhJt4rnzZPRk+dOpzAubz7omckX1MrFd4p81o="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 25184 )
`protect data_block
gD6l00tciPUa6pDNTk/+t0OO0nC/UTtBwLB41d4inuAUA3i/ALrNyoJVcBnAmEQW
ptbcNp5fxEUJjnOxnedyZEuEBxWRieZFQnkRdF269oPqD2T2UnI5wIbfyuxMU7Xd
gcTKD90ByBUjHuBTCB+sQrtEgJrvA5Qv5VN93tRJyGY34D4R5ZQ2M1hQJQ2IbMff
gDsHxyLZlnmrAoEH8wDOCUrH3RS5VcL8A0RYnUPlRqdzR1rXRi86GrScYLXA+Uho
lSkyxsdyRimYqujB/OJ7XHGA/qjAP3OMohUVgkaeVykNa5l17y6myiFnZIqmvf9U
MBi+LXytlxF9Ck3m2b6Xm5E8TBQAT3mBHDCabbchqiDITc01yb1zCH8xERRHPaAq
DrlIgPMBPK55SRFQrHzTEtDS17TByjLUj2A3G1N1ijBTal5rCAiDyyRrUzg3c7OO
2AzglLJodQpTrW1rRUnXC5reFdDGE75ktK93wsF6e/XTh85rh7AumX3WhP0R2PA5
FAZz9VOFNcytvQpos8riufKBCQF82UD+b2iP2f8HZkppoJc2wejofLKs86HD69AO
+A9KRKW4O9dOIHTTrh9LKDDn5jRhn1RDX3meQWjs4j3gCBMXSRJS44EbVUteo1JE
39o7ptPVSjU/SJTyFwzjWMUYmSwEob+S0alMX6tZEVryFTUJ6xadQZycN9ZVuJqx
Mou/5mnG7XFOk60nqB6CjH9DSldfP5OmSiLqPUnAxXPZuZP+Kf4k7Nb6SLVgJA4K
ktaLgaLN9aqJLW3gynYlITuKNtvj/iYXGKCiyZbtFCHg2F+XS1QzV1AkXR74CV5H
IBnyBOZ9pZNp9HFfms9BPEPfnLFgf7d8hmv7J4X8cckAmCTlQoCIbWz8wepTyN2c
rj+UP6x7PowBFk/qSAwCovEHw3ZqSWLVHSr7ICu2jD33mXLRuTi4h12qCqq43EbO
5E+WC7eyfJ3ewDss0xyZ3zfpSP/nErSf9NySk80Ox4JGKC4paCePgdUm1QaxPV16
jwUFk1ziTSRGK3UAzML2eMpM5b1fuTRwfypBpo8GvN3XX4V6OeOWBT9F4P5CCUy2
Mkly/KqtiiAvyaf0ILd0e9rImEc9QG8PsVrR4uR/MLDg44TSaAegqJ8Qoj8pVS6v
FgQuh74F1vCu25swRyQedskc8qrYr65xo4egZwDOZ5iEhLJ9YK+zdG3ff5AqWVz+
97N9qLlGc317QAwjw6HkQTK9d6xGMunKvhXM6MmOjsRbdulkfeXnQlPKu5CIUJC2
7101a2Kk5pzDrqunwbcwFzMh/Jyf2yKbuVOJ6P1qM/7EPScdI9JNoUeu0xRYITY4
Rq4EmBjV7a8Yh/qma7AdYF6VLcGnjchiIV2lrIhgZfq8QvWu2HNcbIXDol/WvZIV
WVPZDcOGzeM0HZ6H/kGFMexqJn1AshdZHLJfwRe5K2f+He/m87P/pkiifuvzlqCz
9Xbou3iie5EVMBsfDQan+jLdK8b6EHN/veKFutCZe/wXShYxQDXE8JKQ27lCpuv9
/qTUa3RaJ2m9XK8bibTu8v3gX2c5XSpgtFw9vdSbDjoEjaZmPzSWyl+DsdVSQnXC
uDe+pGUiPJGXCJrd3XvG5Zv+UzB1GZRa8dGJVSZXoV1ZEpPsge69VUJIlhfTiKRK
N3ZuNeenXMhx4XWhaGcS6JY2kAB37YqrDHDsMfoOjtMi+CNmFhm7SmMJJM5cCWtj
f6eGzse3oU48CG3WmeTG+hlovZB2Ccys7zaa+6CgpIuEXBDSzdRGqSTMUIOruJAy
o0dVZX4fzrBIkEqu3Ga2V26i/wtkSjTROyP8OIH9imtuwSshY9AEmCcworRoxeGU
4w0Xr5xXK44jzf48HveS1o7ziz+WyZq/EqBQxgCz0zt1423KNzaZsakoInWfYGCP
WyrnhoIYmvUOe/9h9bI2u1NcqOkEz8yS53K6vcXUEN0sThajHzqbqBhHpkZm2EIF
Ed8mGCV2JtYfgLwHfSbty8Af/7KqIOvSUj9LxBh7gFmlJdhOeo9yWniNXAc6+6tu
9BblUegKd9DmrqM0gIKclwofdSmVJB4XF4L6LfhP4D3OdOs13w5hTs+TU3z/DsqR
WrWjvDO6ukPUdonxEB+Vg24OHvx5E9kVewgVM6rxEPC78SPCGl3ELp5qGmg5BGEY
gYtzHmkL8TsaDqLjBsYcmX1Jq6Ik1Y7ny7il6N4/0CXS0dEeL9DyBQXZDWNGRgTn
nu2DkObYLftV2acX7/CFA7Mrpqt+2vRvw2vJDtHjf/5KLRAZsUCd4fowcEHknRvo
Pm9P1lqMCR5skBCHl0XmTbWepiJhgj0Rt39iJX5VklKIXRjLTEBF4AwqBf4ad5sc
2jF/vaR1dlQhVAA4POr1t5fu1En+l0On2vXu3s97y50Fa7LyDwHlyEMyx4kevyOC
OOXIv0WjGqgoByu54WjoLk3sLg7Wo8fapFWD7uYt/5geoO3cpYubfiqccx09PIoX
kPtxe1qxlMQ1vmsd7IakkpaX3hVnjsGneHiwiKl2YiuLMpCaL1b1vOMH5hbwoAfU
9MM7QTZBdtqzeQed6KxkOWYprUkBJ8Py/uPWS/QG8//DtXtwUI/a6s1AO0rI7cMX
3vWx+IRUYK7SEQ7wHs8NeedoSB7nXMJuHgw28CCTbzXvDZQ7TvCYHV+oZ/6Tzoae
Vivg1oYs7B5V5RSfQuJVTON68RsKSXdF/zV8l75R+S9nMfOQpTKl+XVsLVlJ5dYb
yBxulolEN2T+hb457n0zsMVEcgUmpXSoe/xk80RmYvEKvI1pojC5gAgxxsAsbyMO
RgxyayNYxYyiyKbKq3Ju78vsMFSjS9GuMGqTs4diYkht/0OXijv47GbvrN91jXb+
2hFMXYc0VFmXZGWchIFH+AVZHHWJq+iDofzxSkmRv+GMZlMRigUcrxEL9wDEKvMe
qHhHYOm+6KcTAoRqMFIlP1nyPEIppLXGv3rjTslKZzOQsWv48xLze+WbgxoO3YN0
VNdV6fqPLqHgdeEVYkm9yIagb9xtcjvJRaXzKfcwJW7ddiXYM27ed8rKB6pv4BI2
yYI1Upsv9XxRfX5jLfgwjTpSVl14BMV0QeYMI2YFd0t917Rc3RV2kfJpWGAEoKLJ
/qp3XU5CrEc/An/Vd+hUq20SXh9XOF/5ewnYN0pdn12Isdeqg0CNM5Ur8g9nA+9V
nC6/2GzVFno1doXtCDPqWeBhq2n5Z05za0ZUnMw8fwfDreW4JNvBrHfNw+S/NocM
mJQVoDdB0qTr4NimLNW58h25DNtkI0o2gaPjiOEzkwYhWByd78BDDDdHZqIwmPta
fk3yizOiDmL3n1mIbdtbF9bJ4hZzdlIl+vCcfg79rG6HLRb+83HHW/ifmXUvZjQ7
Fi9Py7S3bW4SrRxKPBU2bo1WOa3l6nhhSt1iqZ4+xZG0p+OS95c4Wn/VgGDG4S3C
ARPe7fxSx8ksmMw4gfmvcgRyW9je2kLNpWs1/wU2WyvDcprceUxxQSmYchJVvXY+
5yE4pHnwJ4FLfk9uL3RWCQGFrQw8N4LBYdMZa83HyQa076HLkuwtMy+xvC0VTpGM
mMjNXifMTk3TJEfo6FZYSAbAfgO8wZtGsKOiRDo5eeVxWkxT5l9CFYkDQMNDAEH6
x+H46BNdzkrYNkQXN8S2PRWL8AwY0eRpJT3oGMndVZG/T83rwlCPpLsR3uLiFHPK
qQRbfwhj6jrlXYb2oD/zdC30IVmOpmr89aMH52zKivMK4n/Vl5jjv91sZI2cBPZ3
f1NnlFv31+GGHIwLJQFMkdJnhbL9KrezS/cxHRLNC0H3q7OWbuOnpNGNDOBQQGfS
TCEutTSmwGV0qBA0R5V8OJ/VDzRWaPwZW+TiZtVBJ5o1eqv9ljDnEz5oGIea30rJ
98hDtrthdFwuOpaFbnwdlWg41XbtBoRmM76ZYaYF/t9j5PIvJuXk1LzkBcsMPo7k
CqJXdrYUGIGKLN4h3zF6x8TXarVhmutOe5kjNJ9vq0M9nKVwIKUHV6v256OSJ5L9
AdutinKOIExP0lr4ubaa+tccm6Ka7LjKRarzibPYuxUPLuGRh2qu+QEC5iLrYnWk
9fEL4AFJUxAKnuLsZzstBuYtrrK5gptraL/jCUJ6To0QHTDs8UXtInFkPGEmaFmj
zrWm/AHUIQL9CN52MipCbTL1dW17YL2Vx1P7Q98uMwJHfd3WxX26fOinrhQCgQgZ
KMDjpDxrut6NdLKTez1nvTHau+ZfIDajGWoqDXngmQE4utvnIvY3cPix3GNdAcrf
oRpCvRhnCvM2GT0rQ4OCz/y3j5RRCh6stjQ+tFOwGwPXkhjbzLVktrysm8UnXq2K
C0tZe/g2aL84FnnTNy1WZd3Lly76+laNbXkOMHRiAw6X2a0x8I67lefCy8xlIRR7
NxhvP1po5/FSyMlm1swsEpZrbZEH6msvo6mkLOFnYzKZ1rMm9PLSOxxubTIy25U/
LHqTlqVp9CAQzpr52kbzkuLQgJQ1/qDTSOWy9W2QmE+vZl9KpCZ5EtsWYV85CyCi
Kd743oBzOVpOpiyo0xG0CR/p6CI5VcmkVJe4tmAYJ4F/EKRkjlk27ke2vebtDmUM
KvecLPWkNPkfzZ2YFLBO96S4bp1WpFeiu+rwfe+Vm+qjt5r7829pSZHzsWpeP3kw
2e8GS0QePOM9PCwNrGhsDtLvb75m/Jaho2Nkz+iCPQTGEnrt8DS5AVPvdYEAq2po
sYS1kcda9jOJIDnYNNrLN1DNRh5PHM3sre0WhuW1f7f0gjV73+Bj5COc/T+XXPI0
/HcTprwhoJZEqU4NHD2r4/yf/5jIp3jLgnFXNOBsGcIFCO89mK4p5eN8VJH81/Of
gXqm688SHdUwkcm7vQyJJgtnn7VDK1OxVFe7sJDWYowvBkWlgQlcMgL2rsqe6R0S
G7aqv8OR5/9FujYtMRNE3ZQMs2pMLRSbW6MmzSz4zbJ4KRSvRWgAONqwoQr9ONRx
OhVnuNKBsHiTHGhb8BbRu4x3O5mcvvi9aedpuPspzxYH6nj+BnTORd3kSKd+S46D
6j0GLHz64bMCV13qRvaEI61E/eZ5k+7DfQRYOOrVPv4aSrLEihCux/9mqP3gICPU
5LY21cOuN0ZrLMdXex2CX7BRv71Cf5tsJmiom8H2SZ0WKDFzhdtwXZd1APUHUcCM
b7rlk9N3neYyU0rf5aZJAxRXcWSfvc4JmtM57DolOX3CVbDsincqtYNyWNMp00yp
o0hCFoqEHVtRxs7GKXgeLNT4zbbYTNxf+0V4dGxbByP5tkGe0wKRjyqnY5s3StFm
0nD759ggLxfsjdthwQ2pQhGULHNK732EVCXQ4N9DSf0PQBalw05k2zRySnlg9vhH
1+lvCQ8uwsn85ov+PJUvTwijEy69bclLxrCzlBaNPBPfFEjc0Xubh+eod3l1AT3O
hNSAccD5p+bpVVSd8x1V78JqfApeABNzuOER/GCA5ZvhuYH+b00gzrrikDlR0ef1
U0noJeplATgmlDm2x13pNmjhLRz7PNwHTGNWUOwaa55Dj1ckEPDQGVNZw1eddoyQ
bU9cG4eoFRBqhsh4yQAR+pPWF/I3/rDsHBnkTMcO1UUGtYhlfTdjMn8ZAA0UUS5H
wv6KY+fMM+R4YRbEc9nn3sGN4mDU6AAKa3hjmC8XTjkPN8nxM4RjBxrUzxU9uoVl
+0phWrPPxjbByQRwi4T0X+zR8dWcdyKsA2xMMS4pIXuRn7bdMPl3BhTB++35nW4O
Mflv8BCnxIp47skfIT7wpFVUJT3f3RBfhsEkZY1OD5KfxTHhh5HvUTQAbcDWQn3r
f8P4Rc1nJ2mD2OwtD+KkOHLdLilQCNB5ZB4xC5pzmXaCc0+fhCPJz2eZnc7/Ggvb
u9Ax1KgVNFZPc+yfXwxNb+vZTBKiRwbomLhBN6SygZGEJzmE+lhcWaAp2rzC8TWK
RvygQpqsUiPvIfsXsNOwl3r7pCdq50weIs2fCzpj8GNIdIt9BnqwAdcFtyNxCnW8
J4o0H6eah7JYXr/lnjg7Qtv38Glha4rmGZTPIApz3XJpX44ZlFQSPsAY6W3xEaas
2d1qTq7aQ452wc7BpzTbEiyjIAM5I6Nv4Xd1LRywSEJ3wZ7yBtMEZ73osyWr1iSx
/fQHHtmRGOFrLq5aPorABVeYvyVKVt4dh6m/GN1gYLnKA43b89/yRhdLwVlPskdD
2Ixq3EETcfLcFOJ5X8xLj2ZZvQVlH7IbD88C9OAgyw5vBZnYPeBAtV5g83SPlK9Y
e5aQ/805GKvl96CAkypRqpuwipn4T+HJVKuZJqksICIK/3xXrlepeAfZbhoXGADZ
PLdINuLq91Zr18bHMgICqWPhx0W4S8zwP62+28CNlGUjud1z7feTRFfJInTkFM0z
IbQGATiiv8BDT8WK9OOLTjUSpAdV27jjl6ziN81C6DwNqs5ajRrlbhCA5s+fV0er
oujI/5LSAHq4tyvhO8BJGi7ywm4Scwl/Le/OwlBp6tthvpKp+2T3qz6abJKxrYZL
f601Lj0WIoenwp0lBm7mu3ImAoWxkoR/upoD+9XDMyyj09TeM3H6BOny6FAwqp+X
CluXxMjDVhFrDDvFc0l0+sqoo3SIk2ZTP6tTgpvQ/j+cJYaRQh6LzGAQG0zvC+CH
ULx0wnKHAEykjIfLWq/I/uZ9cGeLXn1zyMEy729QW3wONJh/cNfpBUlt3YwFE2ef
OhqYrl+SbmzzlOj7fyEzHHs9e52AScD80QZAMIfXz2obhW9v/2Qk38QXjn1hsksh
oUHUhewGH8sIfTO5dsnqKphYwG31ve6Cvq8UMLr9QVnhKhEopkxmPLJf7HD01eev
EsQt2XZCa/VIQjynGTy8GPmFqXzBs2j9NEh+2InQM0EvBTjtTugwoA5jCMxCeKKm
ZK6ahmpkFu/aLkaqIaxe2TKgJzzeT4v/jZf2abzFEVnbY+GKgaBlqT30P9yhVoDg
HQumh7HnlLhK8fhotDwS3U+nkc4HGKVfnEwzXObeVr7Po/fJ9sLQzT47iWTnSyoP
NMKgWPR+B9dKZdu7ZkLIWPs3U8MQsR7e1f/Ncb0siuMJqJ041a6MlOjiv73Dr9Mc
gJEPrtu3QpyZEoE6kMFpjtLnP+SEzHWcotR0ifrzhRFevzv9ALPGhze/D8n36ClA
M7WgtMewLlF+7J1jxKob28QAcfR0d+FKJtrJNbBMwFSnyUhC2G3NFBQDy8H1FjNq
Sgqa9yo3JNQHKocRT7Tk7I9yTMlCWipEW3FAXq2cbAwaCO/mWts2hXh5PsUX5ebi
p36Tn8r+2WQRHe2nknHBETgkb4ibSEQQbY4UFEOTyOBTArX6vNsGJZQHoZeJY5ye
j99rC59sM1KFRwSkt0oUfluqf+zJjf/rzwZ1salEx5LcoaobA8jEIl7RiWVQ6a9P
o+YCT/KxCVmyWZ+a/rRw5Veevsb4W94xqv3YcMGBKqz/19dAD773Kmd9oWUHpmy7
u1olrPQ2L8udMEmRhY5el5D5zgLz36M2Dm3EKvX2b/sObzYQ3BfpLieuQWKXuJnr
Yp18E/tlz5js0JLz0G4pNFTHrPBb2JzVh9Kbod7N+mOxVhkLysAhLEF/kkesQQlB
M9VS9+EEooqsCUyHqvSvDbuREkHDoNRsKBeoQ1KpT05rQmK51dEOpfk9mFFPYSoA
gwdSto/qV/IlZL6XJy2mLJ8B7QUJ1PDRSkYqHEZL9Cm39DVdYQdzxdLchqopseRO
+PShXDe3p3gJPh26yvsUTE3IBsCnDrzNW5Tl4eXNXcUStvYAlY0txm4g8MqTZzOP
r5LuUHeUL7OIdEVC+l/5u0hbYebUV+AE7QLDJxX5WDy70SdPHt0Mu60ipVajfGgX
LOzxGH/VDc1rqiLmUfutcSY4gDK7/bRcI0Byss08jNWwe4aZbYjJuRsxnoAO4h8U
AvPELULS5oeo44Scxcbspeq4APyvdscNvl23BSgebz70uQRNK5PhHdFehJGyHTMV
D0T/1F/+lVHkEM44DAMqETwfMZnnekFkca+/RyZtrq+6mfmUoqUu22DANYeUhyiJ
Ht+GsWc/thaTKa3It9xJa1zMyUvWia4Co5znKzZPtG2M+AhQHHqqKPe0QbQwvSFu
Zwldwe9OWmbKIW60vvfKHta/5v76rvC4VpuVBZxPgC49/j/WEZrQ0CSDQOwLQ9uz
PrI33JPgDffniwbKCysK3RERbnOGYgjFpHk1ueb4uWgp3b80EzeHWq+Mt5aXRqYL
WaVXDnThN9+QlyQ1zVBWrqRzCrOGmZs6yk7gpY8sLEi6oWEfZEtn89PVSObjCyvT
Sqpm5fDsYApAYrkX/hV9hk8bXllzNCa+3euETEezQ/qYU60SZoBswStDG6IXu6cz
z1kCY1KqFiERHng1aVbgnMPO2+Ai+WCrg/ygoy/YDcBfN/CgrcGcxAJJ9iqRGFx3
1dfiWgpOKXmbMghD4+1YpOcEZ0Z1+61WL4snu2qaf4RXuD5SMHPo2bkABjrQ4Ht9
IqBOgtf2ofsLS3NMkgd0KHJFAbjlSuq+Rt7lM41qCsK0BVV9fVDHq0k1wrVGXIxM
DJ/UfsTEYMr5VgQ00e9cplMv6YdvD0ERA+EqVX5vMMWSI+ebnt/uGZqxEMdDV9J4
EkV+/fgyHSSjH/hYEaXcGCxtNW1x9ob4xL9TbNtH4yQPoQsTAOfb01hcJgrEgUvP
TNwvw0Z0+nbVkFFLUBdI0yCnUN4EJyZdHAJmPxFkwsonEAa/zdNBHNcw2ZHVdCga
qEM5Swchh+IN6ueo1Uf+DaU5yrPs6KrztdWRFWbpbqSXtIV9RsBDQrCQ7MhUW1+u
YTnmDvgI/SJ9ztfarifX50Fchqz4GsicUOdHS+vjriQYBYIqo7N74nElnp/vMjPg
TaSn8C/i1vHzwK815lGhkFbn4scOnQgjx9Uz8VIeQZ/OryGPZIGuv4O/IbFo694A
hNfEg1A7bNlFhaSe3Pms3axXp2Nw4A4MWReq63f8YyibZHcwrd1sVuKT+tuglV2N
e4curQG7MO2uVBSE+ZP6qu0QMRmsLvGXhSBmr1cSQpi0kQ1nOFn/j1WCH1XXxDww
anYyZ8E5KJ6Y/+OEV2je70j47H9okVjHqU17MjPAw1+qXsjYN2B0gbmRjfPP5nyW
/owe0avp3w1BcyhYQauCkr7UuEM+IC2Mnsuv3xqBstjXKfcYqYbRyPatT7bRhr2z
giOvABFQUjR3CElo851spuj/HyOL2R/o1UYyLdF37D/HrpX7MIiDkztriURmPJjJ
lxNEB84Gzn6PX8tRKnhUqOO6IfNlCU1ILCF+6aKSLFqIQqTasIEsfA+rbqb1yQRe
mG0SuwYScr7LikjbuUh5WfRyXCyvpmZzMNK2pE+L7EgrsNvuJyKeEzHZLnwJC8CR
HtwK80QDEDf5B52bNa3pidWFQVu6XFcOLp2tFEdJYagvBp7AjV7xEV/2/Ie+ed4l
TtXkS/40JD7aItAk4G7cWbZGcyzpBa9kFzvtJ0vCBl1IaBBNfH9+hu40ichHlOGF
B/YLxzypl+RsG2puSG7+q7rS/1dXEWMFbygwfzdMmxpqJoQxUYbqMomOwSDbNQEh
TX3NryNdb8Oyl2Pd7HwDBkFoggwuRiKfghL5MIDy9PYySbWuQqbQa7U8TdnZ+Xn4
r1UhTCBHqmVJzlcZqh9Ytf6PcnuxZ+A1CMYN3e6wE0HHDvTTDRfP54Ixl4N4jz7q
Dve/SsMwyshFUYLNNVErUzhWWxX55ggrm5wpjZR6IWCsNaiXVA77W2vuiuirEmjG
7/VkrzFg4+QI4uOK1nGVSacfe5QGH8XAYEWWJ0v2vqxePMEdBs8YaCPLJMSenGAC
643q1LUXbdw8vIPhqXrTvitv4WCXhp3KY4FB2c7k2fF4TFR70HRN99alcPOPzdCa
q1/GzHPZ9ftlkUVA5CP4OKdthz707igtdqYMimMOdvlqPeWjQOYiICNT8vNYxGRn
3UwhXx6zNi9YK9NVANWClwQ0KWEweqf8omtnbEiecxhDT7853scH7XIohCfQYvwu
DE+zLNyrRAdG50KrRaiFjHDYuhaovzl2ZJ2DuiPMhJ+UoH0Q9E4Hen3tL7KquS+c
/vhlDfOwQ26TjVUahsPFNZK8l/oJ8+iSxRPke5W0soenTlEw/bPO8ZIL60LS4OXw
B/4rFFOVX/p5ZTEoJoD/MKtXA4TCtG4h1uLEGZ+cs6zQbG7Vdxpeq6jtOUBtplJB
3zZ9XuWx0JBYq4e5aFbp7Qid5n4fDtJxzNnR0mxuJlavu+kQlwtNU8jsA0wPq7M7
DLCTho8Oejtw3WbP2Xx5oT3UOLmmZcq4Brhi+GsedmrU5xdu942gIS3gMclCYX+/
/eOj9ylv2J2cFL3hOGnA6MYa91ZnoC5D391if9/em/Utct9XcyR/rcZxvOt84hU5
u7G+rCE+2NVBMVnIbNv5r/Jhg7BGOLeUaR8ep7zvP3hMTLM46jCYrtZo+A/0QfDC
Lk1OqUYrllCGA/l/DniYWBtyQ78UfQDRBbB8WMSJ7bzAj7LgyjaIBTHHTy7STQYd
25el3SZzoKx8FZIh+9oL2aPcXD0hNfKGo13kt97su+88fcTDXIlgtx4MX5HkLawl
zUHqKF48ny/OVP4vtUSWZ5BX6npi0ffOlLlFVxG6QrdvO7rXWHXAd5eEHLIagswB
chVzUybCVlmZnJt6S6M6/t1tfRJJhJsUNZNepIJgF8eOIEUVQuX2fp9Q3bg0GsC1
nf6nSCX8TD+Ba/QKXyI7jGcTr9NEt3/Qay+8RWhFJJ8ny2fbiJWvd2ULaOykQLDU
vqNtp2H/8MB1hwTBjEO0NJi8jqWeH0XEP+jaLjnpA27AqDn+rQet/0iX9xD1dbIj
3TW5xdVmHHi31W3EJ6vXPkGUZTiM2nZ0h5mNIa2jusY9rioMhRJgBsBfL/rNXpy0
SKCYHU70VlbOGnFe2VF1z4H5gR/HXgQ/SxPydXXYk1GNor/5+rgEwr5K1haHs8kN
dnSww+SRrLxsrM4VSCqrzQT9AGCJAPnfoIscg4QytCpT9/SoP+cyxV9+792a/mzL
HtQVa6WwU8EYH0p8JkKUae7LhWsv77g3ZwMu5QZBEW4gPGr1ngPINl5FgQ1vpSaC
SJT94nq5ooP2sepMlzqI76C/9tfqnrkfdADojYQnsmZNBDpQDtw/BKbiJmeTzrL8
IAwjAenx4T1vxjJY31F/KDLkC+4m7PT+kQZm+uqzBZHizW6ylioPOsxAxckkxZB7
ERaw6lkRZ3q4dwilgXzjzB+HU/KMZwKF9BwarkgMtnRzm6pI0623xYtq5hEve2ZZ
eJMisxRscLyRUPzUsXMn+ReVA4CkY9WKbvI08sj+w3Y1ARjhhReTBMsdcEFvb08v
RCvLIxkOE8Kf85w68dTOYwfmdu2O8B6m2hGnP2h/WmX5UaYQpkNvsiW5XUbl4HL6
QjL3Eb3lQf7sdTjVk3urHf6CQ+zVy6+uA0NZMUpdxd1xgZLsYHGzkNzCuM30zoy2
p3GSXS23/ohm2AMjSO2hyjh6KHUgCiwZM4inggLONGGl/z7t8qDxhFYxPrbM3opD
qTw+UHx8/g7JmSp2m8zN2O8CJwhtjAERQKdKYOhI73kk4iMoUOzj8KTvZoefknq2
QBKP1xeF5Cy7iuQBo84mTNsYjxWUljYIw3Mx3aiyrosVV1UaAF36J9YmsfEBQqdX
ZRAX1qAiHYXuWFbxvacWOcht2k5hn8s7FEocf1bR6C8qNoWjmrzYdDKqTLYTW1Eo
/I89kP/MyYHre0xmRWFaYsXJNorrLg5/WpqB2VuEZM2oqmeTA57W/laoye4c4EP0
9rRHYrf4zfd1wvMJ38fiPGjy4vzF9BFKNUqQxr0YYwby+NHFFnAJU/J9lnSPX1wF
5JbWnrYt/MWGEYRlByi+bjANObbf/kW+zCrV0PpALjqyx2jXVW4lKUeoSH/oCIi/
1zMCCQr7FFcuDsXrjrINq+PbYBS/KshZUJjNYm9kCicGPdGf6Gz4lxA5suzzufLQ
gX+WZ7Vijh7eueWAR7DTYR0vfbgML+oYDTahGlhVaRche6zy3XtyJviK1+lDK9KM
fXX8MYJPIgNPHB7O7LY3Jn97UQP6MowpZa/YxmXsFlpjUoJLnRTA0ZR2TxS4MtUe
G3EO77sO7qNRzV+KPVuzC6j5Bf6i7b3pVyTq9gbeSaOtjOyPmolMozqRMQsvCA/L
YeDwSiFcGDBuAVRyHsLKrdZEiDq3rLb6lYjXt7opydLeSzXuzxWj+YneAPp3oU81
Areg9LJ1JmldcL6FMG1i2x9tSbhgWVvukAzj6Xgkqpn2NfZ5yf56GUz32QTLlRt/
956WqaqyFpc0EQFoPMR1x2/zP9M0spm0ufgp+WPmEwR9yulC4a0DrVvV1NIUCnEE
0iPO/14IP9/EaqpIWHSxyTx65HdtIjMJv2XSgQ3tumu0rgKNqB0cZ4EIi410fdN8
wUeA81FpiFrQ1Y1BfVH+s+L1gyio6oLrQDEnAkA2FFRtz6jPgZtremXis+OM/mEu
xGDwSaYsVR+UP3h/cZ9NsrGhaCEHA7nkcJBUoHiFJNdZmguiuFfrOryBhyudRig1
sMfAkzSeGeoAmcf0SsFNnEhVbKjOb3QTuvZHpTnhsMyDIzQE/kLXglRBZh7mKUbN
UkpTvrX3OA55OWB0NQxmo9ybCv3BpqKvXfTyij6ZZLr50Yv8oys05KQ7qO3ffNVR
oQEAZX8GtJ3l/2YURoA1wYx3K0ImW79ZS8FAce36I9jqyOzXhDsAjN3rpasuxiUx
4h9cmNCJo9vWwUahUwfKF2BwIuzwv7JFjTug86o/NheYtsfJjC475ztjHFrBBM4e
kgeLeblqc+DKDhEW7nSfbyyix4eejEy2eKw+NcQ/n+hzGhlUOG3UIknkD4UlwUHe
kmjPn5GWpUbiQadTtHLmHcWn32ruSqgxlBTho1I0rANyP8Rq26Qrn7Dd4gnVDNLj
mBOmVgoanN4YgLZBJgshmZPGuqhaG8cUTm/rS7YTrJVPzCBhOP8k/8BZUE3ohDc6
8acJCPFcMZeeJZjURkcvnl9w+MEwYpjzbwt3xp+i9fsycJSi0Q8RI50fIouK7Xqs
Ap1WJdugqjf1JuGHd+SVvtlbki7RUZ/Ul+MPbVYHOk+gvWHfxH9hdDALbGyIVKDV
DoFIJesRfMsL2ctPvKQGaKu+6RS7aUrG5cLDumMrahnf2cwyII0mZ1W+okdCk1+3
yN0iHZjcsOL/JVqpEF7tLrWEKJMUpbwbuqXNYybQ2+vHdfJVocGAsMNbiHr5AJi+
N6gagao+m8KQDafL7Uupbgh+ENGIG2n4zfBwAK3OhzgvdChXhrHZIc9IGFpGaVgb
W99q20yOOvDwm0YgeEfRgssWGPzvHOccvuGNwbi80wTd0FeSgCfCRvNqfKFsrMDt
Wh0+21DSTDe2vi9tZPk6uAPSecTb6/A+1Hb3CBmkRyXOJoJf25TyeKjH/YsLhs/c
zU88rDKnDMPZSchgKx4vu0jLe9po6ypf7gmQ9ZMwt51FVMewHHfXJNIa/oIr61Vz
uLlxetQNOoSzKhYFQgmtr9FvK9H5u0ADc9QV2RR1KYcVAWwlZvR63GFrUmL13/p4
ud34sbVxsjm0GnxV2wi9Ma6UNgKBetVfP/+C7Kop22ujoLwy3RTU9nc0WOsT6Kf7
VVMxqwH0bQNYo2oDDwPsS+kRqnnluT0FqKsVI0CBd9rbt1lOc8HlA2G5qyKj6P4n
ScwZHa/ovcvjC/GfNLoYpyKZCzkmPOUmPKTvnPyxaI0ZqBawhWzSqQF4nMDyerOi
TvA2p436yaPI0XhBpNVFYMkO1+QcEA/hZ6DwntOu7+xY6env71h+9dSykMG/FJAO
YfrgoOnI28WVk+CdQKexkrQqKWdbnAZr1O6fG3thHJCJC25dTayPgf+JEBqWwBo2
PGYfzGlcF8cJ393St3kCSli76g2aULwfW+WeyxIXMaVpZb0AVUq+4EfSI+dVsbpm
R8AVOiFT/LintesJQ07z7Sf6kkHvN4plD5T51WTreUh0t0YRWffHG1vspBFNxjJv
6TOT0eKYddEX4UvO69YBYwZtI2Pb9YenfQKdjYVxIjE4HYGA4sxDMKTqAHYNLgoV
UAztg1pPC9NCHqjvmYnTem1ZtXZO+Bpdm079Zqc6XGnzzDpjrfsF588I+qX8XKlM
SfaoSuP0Nf4P/C+7W2HVD4PC1DUIeSyo0lSjnUBIzVmXev75JB7gceC2qNUbthKM
LnMTLqnw8R+C7F/axGJuk6UEA7oZLqXgW8LIysMPhsGKNQ8FMxY9N3tSsqhCeXaF
c3HC3/Hmqx9yWONQud0m4bunThs5dB30LLkRBBWjwqsODl6/JbW0vl+6qmKtniN8
j+MNWy96K7P2Yor5k/Q2/qalEHzz3H5j7ufwzD7SByoffx0I1x47BG3tHo+It3Qa
ZXsxst5GqQFZxmXOvxDZGAduISqa0hWfjGoqAQP7poTw5vMJ9JJK7HmEcaRlixOD
WZZcsM4EqtSjyL5Ay2QO5VkrvqJj5Dg4dhjhc9g0sAMnnBaVJ7DR/T8gnZk4TYLs
eDNoxWRtNNVHjisg6jTnets79udlYW8ud0H+P4iDhCCWlFSgPdbSDbePtDYiZ4pH
F+NtRk17ul/M3r+XdjAjF0azNAPq1bhyELSWZuckwpzzt5HNS28KRouoo+BEIBHM
K1UD8J75zv16ZXkRcxqU2OkLphtOWl190KnHZ7wXOBL81TaT6ATZ6rL3VeF5TZul
I/jEoN1briaXlb9LhCH/IqhhBAMBouWCoaIQJ/gb8juRav0EUZ/vj2ey1sry5fJh
SznMffnrUrTgVQSkIe9YpseIEfzhKZJcagEoM+egcLXLa+zmZjuGacBwcqS5QnC9
sAVrG4f4r1LHg2NwAet9Zbx0NIzGkDpRPHLnEo7NOkZorrFoci9aKWDhC3FVO5k6
PHpAIhslAtgqX5kUx6E/Bejz154CfvD87mxbbtv2essMBe+167eHdGUzLG8ukNGQ
lAJSwpNXM8Ne+s38PR4gUd8WrQTIxOVXropDkMU+3LumRTD8vXqr4jf9ZZ6bHwxC
mEc9hGsNfVmYIs7B/F8LkzAbWB8x3xzJ+BJgm7t2K99xq3boInvxhHTKogzC5aBC
M8++fkHInhwXOAD47rmOjTnD6T3zcPOqJUnL7aN5+98J5kc6vQjOrSUt6rON5Lu3
x2kjKpgy+mASiT4BTdVT2ale1+VqPQFIgw0xaS5rJes+cQS1oACBybx0zb+4S8BH
1CTNPLe6BUXbzUKRVBYOcDFim9tdQtZXdkykUlizArDeRq/FrMJ4QmQcLWdMpjE3
yFreCwtePDYUq3KNIqlwYAzoynXOZeqcb7KIbL4MAFmAcaRfgVvhWK7avMgycBgw
lK5k3qJICMK/js/5nLu7567SdpQZsuMoVahTXfT/cziY6/X7og/8uY2po4I3PQKx
i+W8uHs8De/Pt50WyMEUtC7A98oXT17/dJMDGkG5ubtx6kJ0TXJhcbiWVlSPYKHP
H68vxoVadVgwQtlffjXqEp9WNY0goJxH8sD9/gDjak+M92HVL2ZfNNj8nwDUziSH
T8M+C4Nx/NkRcSybAvHb6DMI33Mq3NfNn3MuS05fSgbpd8ts9eMp0+JyznkHQ1X2
qkeTEjse45HEGufGzy2o9UQrbh0XacFUAVcOesBi5TQ7HDcQbGk6FdkqcHWfQAvg
M9XzijbG54+OwpUiGUTR6Kk5A4F2r84nIyOXH6F5XzkdfjG3F/jOomMTxMFnbghT
9VSi1dk2bg5rQ/c35PL3/X7lLIttK5iUFGOemVJTd+N6cTvWX9Etjj0XhsVHIVvL
2vO9/hhk1ei0EkbCPnxJNKSStrNNzuUhPn3P9/f7OWelk17OUwsNXEH1OH8GKBPI
/kOsqZHHSMbrZfmUU7CFncLiaQORA9SgCSujTpwycdsezZ52/IuC2mk/Fix4073R
Jy85YP/OIyag+ZhNBXGAoLQ/AmR7USA0oQiTU5R4HTxyw3fe3MbCoSSu6mrJC9uQ
33jXFF6sZSd9jf/zek9yNANz0UfbTSYrWe03fiT4WIas52uffICDE2omJedamF4A
WCmAGHfNCdZbvb+q9qXWrj/bpu9WaX+d+vn+vJb86KxAsgJxERNIuUTDhpmeb29a
IEvK3DrOwbgGLdx84Uf5LZxju5Kv93v1OATBj8iRnXf7lrBcqXVPo1RlJRMqvbwv
wVMRexbBoNBqYl8pVLoh+hUgYB0QQgiGcDZJBjeocBmtLHN92NfYY66iEveN/lK8
jN9GicLFIMMJJupb+oVprCp1xZ1t7akC/JReq0HBeNIOob+OjbfvSY95ZXMKf5eO
kgDGJCOJny4dc0B5xTP5+xBCYiUJ2pIFqTlgEdCL85OAfyGlaWbOPWy8OA5oLbna
HCjQs5neXRCTzx4cWfmueOkLHL9AqLGPg3u4CPO8VIE/f7t/KWSuO6x0wES1swBf
Qx7BO+HB9ETb72SDWC7M95WLOQ5VZDmHyxnLhrTm4dKRZElF+NMlY3xh2ReTrOXV
x6c5jK395aOztFxXNZHUNOmXVZYzlQWOYN3Ljz2rMisWazchoH5rXMyfdubpkoPa
Jt2Cc0yJggPSY2rZMjY8COBbSvXv5EKTTHQXV5ifIyduVRJBwxK803ko9NP2j/eV
JsoTfz+ufVx5pswMFxoujZdGGS42SAPpvU+86SYqwRWL+wzUerULDERviqU3QvXB
zl+YYbmwel0a1uhGjST8akSn1mHcQOI3ZwFN6HhbtBNafBO1DYoIBgol1Y9gL3Hq
ubjYFDhNxLCr1fLw1XG3J4Y7o21JB/0CtWArpyHaa1c0O5zzoJRTljw56oPGrnUn
IMSohSvkFoCuyvfc3lTI4tZOnKaCwOQClLiEhtqCJWc2EEzGDBfLVUcWIq2Ddmnm
FBbJUKaEyGJ9J2cTbIDOMGPuy83Xn5TxKMrOPzmKwE3pI5UJjTsyu49eYCKBD8XG
Pk5kp4Ip2pwsBCVZEeY8t7t6BhziRDZgF6MsJ96pwEb1d9SafdGmN8HbVu4LZwQ/
GaxMtJFeZw4T8ynlRJf0OHomyt5AcIXU2XaxRXG2FOMtTnNR3noDAwLrZholbCbq
LBdn9FDcovdyDwnD/Bu++kfk4+G13Bup82WGAEOwSDeuX3vCci5fcqxZUaNo0dgN
aiX2Wbjd8xPsJ3448biN/j1dRWmC+4DUqEvqhMgR9DsXbztIxyvtDHFo6YIkspRC
8jKtVqah3qaCIkq2PZGjg4PEJhsH7bERLkusjZXnmxcCT16yyZ1prDfCw6XPTSvm
NORxuL6j3XL+db0ISe1gddoUc3dVMHC47d9oOZBGyBkW5LL8ijNSAuPSR0fVYgpb
wYjBNJX0+PW41uXjwFrsCoqPRTxsglMS7tX+08yctxVg7dYNo8gjdqGq1UCV1hyO
k4H2/LdYI05TEmkxAxvMhOa7Rowa3xzHBAq2WSsmNRH5xJxZQgp1HNOFhGztPf4M
YeZGaPVWsXCgguquVLrLnFo14pvzMU8cPMyzAz2vvU4OU4inZ1l+KFY50Wtd/93E
5RSRsypkwOO3LHKSwUb0zpe1PPNjX1Wl87dm3rYdb+LUgHkk4KS7pXtPp3Pdd3HH
pBEaBkH9TH+sQyiTGP8bilDHJEwJkq+djW6q+4FqfcPOpjmAWgvwmIFuQHo3AmSl
+Hrh2i9MieAJ/+/BrAPSzZFiG/1BLXjtgyaUJxJjRj0wxpmh2SB7Y/QMBv3XkLE8
7GvPft7xy3lnZ3cBsTMzLhN+Mb9Tiyq650g21jdmE0FL2BzcH6BDAieXUyVr9XBb
Gdegwzss/0JB5a1NjbALJjmbnfKmwxaI1NJhkOyj12Bz0lgEtqGwemgAIBG2fs3m
FsG7Acr/+mM4gDzXw9ajs/U7g7PmcQZgkaRRIiEf72OJhpb2nm2dRvhAXYBVvxYI
LdUqe4+THTfszfa5X7+ZDZEgfwvlENjjyUVoMvRpzMMFwkXsrhNUA4ANviDh6prj
tPiSRv5bEl31WKOAZut/wEBMzIOpQNpsUPA2FgE84lfJcnMWf2BrLeKzE3NIWOjb
4rd9VUIESIM1Ct6ksW8aiE9EtdkccfXs7HdvLov4OZSNpq61KWHklenCSyGSKoy2
gXLg3ooCRfE3DGRgetkEmKreGShPqtISdrfQqZ1StvPd1edMJwphSxXi7zN3E6eH
ncz6GQSMUNa9OcNaLV9yigDPtC3ki1Z5awgnBElXTm1TRIUx9nv+BNlZ5yW+rLzE
k7vzLTm+pdcXwz5uaSHJ2MNBX6kWInb541ek9ObOZztG66e/Bv6gcZZ2IZAnDqvy
Kgdp2rhmvZHuIfPFCboYd/v+iEHkROqr9ekZqnsYBZW2vk7TlEwQBKGb8eu4a/D1
fXNuo2H3HM3vM1db8BC4BLl6O2IUhGpyshxM4VphMkIs9TAKE2fcsU96Ar1S61TX
R48/deTNtls5l4FKQdsDTdXzrYQrZrZ/ztHk/t+jwPeiNnJVJN4QbRZGLFu3QMCA
fjDEDcdoobv/x+zSB0OTjzV8FvO4ekptDFcuTWRV/qFfF7lfRCv9KNRoXog2XoIj
0o7aX5UK+G0aT0pQHKgi4T31MWeLLX/lI/uvqXI7iQpnsPPMByi5FfVuIueaAkLg
i5R3sya6yFUaAw9emyXKKEd6i4a6ks1pUUNuuastSuSAz6COu1Oic5L4NriG7Yaf
PV4Sw4yRZIEgjOvMYXpKWsEQu065fa6AShNOTKu58lyLTj9azs98kw3+cDvOPbn1
WGaHNXtYxIWZwGZpIzo614A7cSU7KVptLbfWTwB5ACPKMqlDeEUOicvI4dIIG4lm
qEXFjRJ3NXGp4U1yE+i4pA7OBJ67iBkceC8/aU2tannTzIEWAx+aSCu3+hqXJRjG
VoWpUcfCaO5UWLR0yUiJfIBVON7M70UrBONAxfht4n3ymrX6tptPzX2aG05rVWHr
fD3Wan0/Kuhlubtyyn3hOYGzmpEygfQK56yfgJ/+W5WGZoy6hfPE1RSikomgnb7w
JTcN3A6y4r5Vlswes3mnM69k0VRbwmXo3kfvFhLCdYyzY8kP60OMJHWAuSxfeCdH
gOIDEfNi020+TfMChpqZmNY5A+2oRDjzL5vBY7fSNlNX1GaW+GfJ+g6JzPcVS6W5
m58TOSxd+psNeTvx8zraX2/tcD1ezoQVf4170GtPveiKupb4Cp94ls9tiou7CINJ
FstdsLNePRxk2JPBGk+Ly6Z46ER3YLfQyXP9LLLhz6hZO/Hyuo7cX1CXzweYLSxj
TrKDl/+PKx++lKtrGeoXxgOp4CLIXClO6TIIU3bioXbAouEdaQYV0kXU3q/lx0fw
PQCaolEqyI55seDpnxTk+gRDhhERkVwjJI7HE862f/p2d8OYB8EB94Js351pa5XK
sGTfAfQFcufQSGfas24WT1eNXPD9DO5JlOCVOJWAiYD4FrQWhl+n2dzPC5nzsyCe
1H65KrtJugjRCF/EI8LDHyNYD5im6XIWP6+7Fj8CEYyiJ+p/dbNv/t2gKm2lzCYO
eNik75XbMocLV38l6tNFy5WbH+u/XzJuJhYBk5b4WQg6eo9IikQQhllXkEW8/NTB
oknznaXmMUcfSZ+dP7GJEMPxlEMLlUlQHUjpGobk1OU/Silstmdlpf8ofJfriy7B
SIN/iRHTmgWZCC3tqVs3/gSqgI0LUPPGfkkx1SlVEG3JUAWShmb6+jRzaDZh+Yk+
NvFGLfM74Wfzjd7J9+VZLSyBSedFPxrT1zxHpR3c/f7ln5XIk/Xmq7/NvvHvJ6Yq
momqK14G1CgOpGcNWkIqPI9cjzkDy1B0u82zNVng/nqGr60xcE1u344mJ7lFNuxs
wkGfs70AJR2ElU/cl6qLW66YOxWe7rEUfFsW18JIUK/D38V43wnaBJ/8J6wmi5LH
+eZFHlmgQjhQg08uzgn3gI3IWPrgMUFe258BICXRS3sRGuc8/IMvfS8trg0QiSgY
823JJrYriqpEBp3eBRr+lvSjfqw51iJCP82y2Ms60YKjp+WWpkDSTiU0relUu4lr
dhRFJWBN3aDCVaNp5ACIO+DhaDXbkkjNmLsB2FYbW/zTh4IEQuNK9JwaeJg/fGey
kdmVI/dTG/+JUVWoeRJGvpPC9hC66rV8tNwc7LTKNuuzs+oQulqCOD8kiCRyWx76
2Ngic3gDBNmqWa9q+yzhy6PXzsBBxKortsR3McHtoAMpx3uplPzawirYzl1EsUdV
nrjXq4EFnweFa7InamFWwPaiyvbqGElozKtFNh4VIkHTFX0Q7MrO5Fz/P9dsgdG8
hP/FsNP+igsMXC5b+7NybdnF3TWROEJMymo7Y6h5xmfPsVVN1fg13Ryo1HAx6KJV
xQHlXRGr+EzfZNKgsCeZLAhJHhnN1mJ/1RNXK8vcaWfV4TyYKmFc2dhHcHymlAHk
hL+9ZZbpzg+AwwiLnBUstX0YxnYwGSgsNIxTA2qW3zx36/ePshkLxvqP8WzVIDF2
zkaItqQ8vWxk85X59vu40iMCyIS+yK9YSMU5ZT8nJO/8xKWbHTwCeVPiByCt5auL
xy7BwDn/cvgRrYaIkgJJAARONK4IQ5P/VMOJ6ynpmyK3LJI+2IKjfWjNXg1JGJ9U
a+oUqmNMwkvN1ms9xLRTYlIlPNzA0gjut3FptfFQFVMtm8ltvPVHNUdGTGFRUfQb
gkAW138iMH9Yx2lzgSFlXhcy7i+J8g+2lq6bRq8yyDEpNADzCeoSV5GlWaMfIryc
7PUo0goqm5xzMxST4SLfmbijSFjxBhKg4kBsSsHP1fo9U67Rt0TpwGxfA+4QwyYH
m+vwWdU9ellgJ3NwejpMVAB17wDxhR1RH3QwgwC246suKUizw8EAqwV0BxE/u3E9
Ect5PDrjot7RT3FaUgoqUkh3Gt5KTtLZc5/uDalLIWiMwr59gye/Q0okq3Q1FAbf
1qgTuA9ag1BueqGq9I0Wz1xxMPE9/SMyUEoVm80oN2p2HQePgGiGCVSzUbYBui3q
rWeUFsHEDoI6nGecjTC4wZ2im+P9fBBgT1M5pqdg55b0WivHiYOcXglUxcAk6ifF
saYEiw2NYHBa+0gI+dR2tBNvnCXgoROq4KZYanitPRcpUujUiIm/J6grWQxvF6Qe
jSJk0iyg25tzqBeBRBBvVCIeclUp9f9aiVMg4KsuyS3xmIlWc689F1zEhgUniib0
kbIVKqljsfzzRssTZP9NDK0WND9qCP+pz9pnIuzyM5an5iFab8p3cNOUNSeO4N2X
AsOG719kEISmKicJYM0Qx/T51+okvSgvt0y5xoOkHwIQ+1eu8veOPmS60KI16qN0
uAMyulT6vQXbTmZFI1u8BxLszJM84pv+H14z7n77/Vu1kV/eR0Jn+3rCGlakBvEz
H7BhcEoI/MBYLlbEyXwLvxK4bT/Y6zUalrUp9tdSkZjo5Bo/zIOegoH8bliZ9TAz
HSf/dUXlLDxw9ozmKnm5/P69L01rCVYD685WT6Ldv2bUD7c/RFtuChCgrDMGLvdH
OtmpJJjOuFl2AnMHdAIag+BvGUOPEJWZrPqoV6CxACqTorh033cQXzdrNiKVesRZ
UQo3tJOudb0GTN7p2JWEIVTYKEWoa7r3DbalUlh7GAh3iqZVTqWh4z+9J/jPuVTC
Yat8EPOVfSNfQ4A+zeA8Tltnt7gEmj/q39pEFZVZZ6QHzOLzWwnY6iX8iQ4qFxEd
6pBTRSb5OtpfKX6JEt4ebc4NtniwMdKewbYxFk4PW5yn4tMNVZrWeHFe8bX2+KrT
QWWBlsDy4Fxrb7MLEYgmNoLgDkdzF6bUlXoMmjXlAX1p3Rmj7loVm6Vq6I7U7h+h
/MXt7cr7u7kIJfayEFdhsKf8vY/bBR1CzeqNpUSYX3cVipHvdtpNJmtCk0tH/mlP
w2QZ0JD8cz5WGAD2ApJlmd/HBViZ9DoPnxmNShuLpjPe1MjfbhZ8An6mD88P3TuQ
vqmJsR/WsF/0BrhZ2rGuAZAbvrGmwNYjLWbEP1DgscE1GFOiFLuDZFifmSiSMbEg
a+KNCf4IUJbIiMylT3yidbZan28GNQaHlbs5otxPrToRl3SojUlWnpRFglh5rDeL
tgmRlpBl6WmmKGxjLzQ+M8HgQWDla99qSwjBuQ4XDANSI//i+TZsvbjOjKkoKpKv
LiEycQmiOR27JUqEi0MG/aDr3vpEP2zfKciAHG3ErvT3UOHIkuRrHlqZGN3TYop6
xMPqeEWT+O+VL2ViQt8w8zojsB7wEHhEKZ0y2MqdTXGFBkdoxs3rriDxJ36lx9oo
RdhJ5ypfJIYonirol0Ys+91tDVQ+P7rO8f4Zy/ivAwQJVo2ACMElzey1LRMoLIXC
rkFi8SoLu5EjIteOcln9ynktTvCIIt+qLllOxcCbLxOF2wmOJodW/c8mtEXHNsMO
quTf2Z6BmWQIy1E/yChR9y3dxDh3aU6anzTCN8hIa+DoSxFiT0uTtYaZyHCwNkzv
KHJ9YDlxln2TeXmuutM6PTrFzVFl+YJ/dMCw3/jYgyN5R+d0rrs2kgIs6TmlwBRj
F0/vnci8mz5BtAhWkhfCDAiEikfmGP37MGKbCgDogoX35V2EpL/PtMzs1ygZrgGY
wKpCMEFAA1em8DOMOvpY+yKZ2ackr7mTVsIZajmAh/hi5xbcYzGaxWpk3bJpvzAB
CJmBHUN1Dk8mLxjwEh1vfnptmpo5/N/fC1GewGQQGqfi7ei6rLRtluPM5FzRiVl1
2IhCB5/b7byMd7nwDvkk8Dft0dc93tGRBreeyofY2RElYxgENOsCKJXz4OrGnz3W
5aw3IaL28ocWqSuOwr0eIVNdLoxIoednYN/QaxKD/waYvE5gmfzRTMWVyPZTtRL3
eWEQ7YAkptppLywnLZ2gjytgdpop/hGTag7YDXAhCXivOW6tsGkZRnKEXr9ipkyY
DMf8CiauOZra9EZB3O8D0Z4vSm5qeF6/4HJ3CpjL7hp7fxmKO18UjwIm5rBhNDuf
KVOx9JelgJZkUlCW7+8FXT4+hS96GtGnCweXUs8VNA3QdZKfyfJTglwwKIj4g8OH
Btrtkm8+yCl+8ddAfjeM4dgpT4pspPCgeanpV6YeiEzs7UgQ0sCK0YB3AEFjhZc6
9002V63n412srcwnlIEgctDIfNT1pJn7bPjS0kcRdW2hU9q1ADIZBJZnEB07UNh8
77x4gcbTDJ71poz4oLeqJWWTdYzplZq0EcAGhpsW01SOch6z5PhGKc53brEvALS9
E/3UrDaW57tO/9cpHu1d1ChzIgJPRNvQ0HuTMcQAwkBtK1YQNVTqxNWdrwUPC994
1AmhOhLLhb0w9B5Hco+gpLbMdHA0db3qJ4Hv3Y3Wd4NEhB1LHsdeubUjfE1iIoGh
shRj0Ag/Wgd1K/uSGwBveSikFOvMJnd+6EY3osD2caMiJhi7+I+0GOICymK15xm1
t/PzVmpim20u/vrMFHKrwp0Opj+cBfkYG2Pwr5Eu2EddYupcqzAgrUyDo1+uUxWo
7iVKYBAHGnmj+vdW8X5e8Kpiy7SuiuPCpGcpW1WABBva5vvRqMAQ5KnfwhApNFpk
qpE3G8FIZQMvWOi1+1k4bD3Qr4ZwePikU/59NhyL1BWvasnFq66MNmVV2HIbJGzC
hxTy/AzUC+iKuvX1vHACsQmIvAtvH0RM/yjZalmM1fxnhdHIFAbjGd8lG5YnbUvf
e3rDtv5XOq6PAqKSfRtWL/UmDaG9Lo6mwn4fZo/cdkEdoWpTAd4iRxOaZboh7KaH
V8aH7kMKKHlaYL9x9SVKOWQ+NSlNp9hSA/b+sHmJkXtiSZKXeV3KhnLWHlkFCErl
pJuu8UgyfkCgyy/q6HPLa4H1aEx/qZ42H4fxAn3jyjQGeVtgF0f45AxcLNTBnEL1
T2B5TTzCZ6YQVi8shz1PGszRTQUgT9upejpmH9/nL9k4UxvVxSHFqVGzhKKrvItk
UA9UybAjGwXFUv6udlZewsNRBDUBu6eZIqAIPNd3gAJaE+qxseE1e7DIJMPeynsL
/8Nt3Elik+jW+yEwgY1J2Z6b0ZllCGWiuuAALK5DUVD+QoXhgi7EcGtaRza58NBr
9zeneMQPctbf/JwNuh7T0l1inpUlmdPuDsceFPstS29KJTK8NkbOCgBRozleIg3D
PbbyfxYlWTsifzTS4oaKTWjJuUUY9k0YOyBqSG8Z6rDHKb+KpbBhHo1SIk5+Tt7o
aNyOiJK/XuW8ZDat5pbevxI5ZSG1FkPrX9rWbF3k4k/ORKuCv5sLePDWu7K7bJHB
TclxKGbLdI7xgNcp1U9CugXNEhijTdVRybzDi6O424TogTfRFCL5ZU67VrzQNYbl
Mm+eIEM1KbodSMn7ctXkgBYHtcKH6mlZnwDWi8LBNjClV9aYUuMCPTk71DkuQhBo
EUmbkpISVgT9Rkz+OGrar7N4MYa8Flu+ybHbIqX2XegN2fxt2RhxzEf0o0fuALbp
wcif5/d6LCv/mynfMirMMcTbcWZ5W7zaIhEPGvR/gwAxd3MoSJN/Px4XbXhr92ON
q38UHy/XIid3+o7i1mH6OZmBsXACDluEGgPe2eHqaS/MwZ9oRR1C+ByPCAd0f2x+
Dx0PrcKlQt+gcoFh/qtyhjMLVI3YEluVvhByr/LMCrJxblm4uYuwHe/NErrkQWgY
qfl3zVmcCqFNuhlL+u9vYe11LpxcNzledSm9zlF3jDsfd206zo2olzQ7cF2facgB
6DeBcWrt976i39NZFLiOwt7s6HMmd8gbmwJ9ahb5mxtp9AigS8S280mK8RhAqjTX
9ClyKTliNMwEWOqoiP0y+fN485o3gaX/N5gKT2NdsCZ3LjvPlHxcK2QDE056gNpm
LCsq4wCFnJT5IVYAKz8ahCzx4mt2SDglLl78iUW0VM1H2ZDlheiUkV20D1EMOIK7
6P8S1hU5eFrK+PPIrqtcL9lM3Lg40By878bAfio7Cq8OE7ftyx2BT3bzctyiU9r2
eMSIo5jSKzLQSQQpzVO3C7FZvoRun5unGbRGbnMdUmEreaoUimpYsz2gftI8n+yG
bRWS/NHY3N+mUVeR5PneL6MX/12N4jSiKEKcSUx7RX/QqlodDD1s+bWFmayoLEAS
5FRy09fdWhnpQgi7ZXGItOfU2KqjYQRQamuuo1yuBuqX7hKvdNrFbWAvVu47rFXP
NVUgJpkKtOfE7g5apL74wQrP1BWpZqU4Gpe6Mo71maHVYJLYh7Udo0VSR+Ey/ZYV
Xy0Co/n6CULuTd5LhqjQLkO4gLGvElYAXBK9RbJqO/HrMA3KLV04nY2mznibAkw7
5Rhs+l8hPLP+6CdNb4+rmf84Bieo8i7m8hEWLwxoyLaPgbivdRTVwCQtAnCJTNYj
4fqsj1PmjfbIRCSGrZSEU7zFsToositmN5NcdXlbI4uZNUPagXIbulTuYSCg3HMh
P/oTflkpzxVr8uUTr2hOy6/rQKj34Z9tXyTeowgU3wuz4CFRQE13Tjcpiv2D2nq+
wW7ZkuGfUe1AnQEi3yhF92S/qGakL3Abc4ezS981TcgPu+ybn3UzBeT5UGS80cLg
32TjI054hlAw6pcpfkVJelj7DKNsn9ffCzVbvDlSJ2vWssLjNsCTAKTvAvaBYw/6
Bdj6dyStAxbvB7HcuDJrE9dtQdZMEDLcU2ixisuo03FkCx/UOTOKZ2N4F7wRPZtp
4Ww9K7kAuaRbA5MwAo72xyYTbxdpO56sgo49f4z6UqufamZNHygg0yhQicS8KE8U
6IUvp8Oou/issUaPKl0hc9Ln9Olvy0JMHCJTi7Kscm3tfum1mG1N+36oF6UXtr0J
slYwxc2VK34lZly5VV3Ts+XhFCKs4lWfUesyuPnRhuwklM1YIkmGmCfU1AvSXAQz
vt9uVrU4q2Dk5GruDKmX1Dm8ZFBl2o9XLayGj/dHzD61lABpn59ITvLrtH6yuc0z
Hv1VdU96bLmXeG8sF81IWsMtjFwJkvV+KJCdy/K0hLITnUkjCKDwheb7kMgDdCsh
FUX0F6IMV2ZM3JrRVX4TX9zsAgj/itJrRGLGQjWXNUO+zYtw9SR2HWcrddZZWAdW
Qk7mOXxGGn2GZNMoG+kTS9sm4LZc9hhnw2OTtU9RmFPNQrajBcWRRNjZuUKmG7l6
Vs+NSrgVZN8iO29LZT1ZL6ajKSIv+lSi82GG0iKGq432h3+/u6Wuw8iXeTWGJf9c
m4Pw7zUjgaivkjqeeOlofaa5SOE+UUnUtrbdmr5uCEU+dg06rI9SygJVc8CqN3ED
/cxZTtv/TKkOtAXoyeAjcXMvJZtTrmRUfqlCijTjSEe52/ZAWBnELB38grCD+W3s
/frSvHwuA1e3X47whTL5hZrMbqSl0zpOrBOeU4B3SIstrjdMaiWJt4/9LmG3r9Mt
fl4hrJQ4FBywsUm4c4Dx8FzYqEr4iPHdhxwVVAOVgWUrxDLLgT+36WAXWV8bGj45
0BC7ExLqX5M/dLTZUUWS6LImmWyPkWNCgUrI0qp7SBm2GhO5B90mVXK7LMJsaaPU
SVnNqdNVwrQVV5UNfG9/LvuMSLbJJHm+BQUxO7AvyClamSBCezZn8G+fBXqQxeRr
S/nSaRkvC+KEPG+BOGVTtp/p8Cn1muzQmHPKCTnMdNg+Y/lIxV/eh1coxUU06xeD
EDLSvHHkhQOQRdb79ZNbs9Kq9KQa8wV14POUxBS1XYrvCQTtaSdGoy5yay9/1CHE
IW5O+Ssdryfy2RglMUAvk/s5/2+8obflXYjqYqPE1VzGHRYsEjfcQgpzx3+6qSGa
aT6Q7Rp68tDtstsD+s/VUXL/QFdxzj3NCz/7GQufPEiEQDJeGkevsw8ycTVVe0/A
ztqiJLxEncFbQ2mSVRnRKL9l/3AajtUoCpAAo2hYqGxhcbJRNjodHPBS6v9NMI1o
ox0Pzi9FDy2wqZ2P1lFtVT+9YZMGAtq8LxOZ7XZWk2/99hQBtmGEt8o/kV2nFEGu
OSe/TcQMZJ77i1S8JCoUI1KTNyyLKTA13MtwH1Ap40ocTjzKXTg6U4pqdm8KlLf9
zZUCYfWRhzM2GlO5YVvu+5LGq6Ke/MGwUNFzFbPOw8xaIzbcErd062cGfTBv3iEv
XxqxQhhGmty+4C1hlEfHx2Q7q/SpgAu7uTcnN8N//tiaHnDkxNz1TKOrN4ywSnwU
gxQenzqGaE68GWpED3yxyjsWv6qjQgt0Cog6LoSF0GPgclGatvTMNqF2HJpSxVFr
yvr07eDLNoJirqo3wKj1Upl8JRNpBfwO7Wm954NheCHu/RG/LzkyPdbtE/MuYKdN
R4EptgooxQFfOo8dCJAmmHMBxlLcyORjJQqSsuo6fqzL7tuL6lZ2yPDCbe/YMTcw
vp2icN1D4GERAtpdLwh8j1foVOy2HVfeC9iJrduErVgD7c9+3ehajKRQDvsGWQai
cW4PA7eQUwbbjFiMzvOWyva8A4T64ZpGxmCf3x10QBnvzxikDGBnEERn6Eujdspo
gDj0vH04+LP8hiZzj9m3yFx5KNTF0QtCOXK62Ii82VNFaJKCVv+Q4ybtlZTulQoi
I8J+g3p85SXXOZ7fnBjmITp5YN6Dvd74r8WpCtMFMT6ymAWWQIKyGlg726b467KP
1dWnEu+eAUJnRta5yHu0n1L2KRLysObvAwfhK4//jjoZc8ZuXXz+n6hPnrvsUuhy
IIeKMqv6cLeNsaHz/Rhak/pGqmogBzxKTMsS0SDjPOPGuBdmo+/r3kPoiJ3a6rNN
oCKm0udTEc3wURXG7g9m1QYD7KF30KD4daH6Y1eMWsRwCf3GW4FmtJKvbOwJa/ap
LKm7+L3ZQQrXPJJciqIc7Y3VcqCNtz7YzEKiYGaFJAgBq2FTKZgz+MOBj6qExgpz
bD4bTsyc0DlgCe+Ysk9OEGHu/eawqfhScrL4n02OoWTN2WxFFEh7o2HCGIKXe+G1
sDJKH/j3ZqMacvv8u5W2i9PaLHFAhHYEALEUiIarGRKko/Aoig1WQ5yzXKU0HjoY
kmNT57A9nGt/cn9TTFsVGp4gxrxqb0sf2nXNuK1kCofvqhXJOwbzbSzacw6qFcNk
XhFrJg7gA9tzb3QCqedIoFWWgEQL11vdp+q0pb+KWeqs9aIdapdNgRq1SbV5nkq5
YJTnARo0zd9BhZIsdNepcd5uHZAKYEwxyUSLd6rzKnqB/YuI2CjyD+lgNb+bp8lX
4M1bLPpynJPfDxm4Q4l3jsXWOyUqfhjZHUUPCBJZUPQEkpPCxqadHlOu8949d5OS
tOo7sSOPfstxJaQCD9CmKfWuxcPiLMxmpVKi8s6Kub2viOBCQzOnIg6OkgulSmsv
2wiCskKo/X1gvkhommEoulzatJO/T6CeM3TQswEhAskTv5Wmkpzqi4cLH4ON5yyh
EmNfEKDpjCKJjtIJ7lpN/sCXPl5wdLUUQq3IjiyyMecXP7Rtp+XGBwXfcqW3k5sE
YAp1lNT9zLxkOAbtmrjpAbMy2IGkzIJamDwE2JE63BzK5h5KUKeY4MEfHrkLbWXL
mS5QuB5j1pMeOeZM5Vzi3PicY1uMjVNwvjWAg8Q2TBy3kP452dEtDBHCLEZYT7QU
WDjIapFxgVUvsIxXqIsD+NgFz/Xa7HyNEFyP5CkdZp0pgs7va7e3kC0msVQyqhnb
ZaUnuJ8yPP1gqZqh1jdoFHRNeM2uAKGOrp8BKb5xtbEhd5eOECvhCGpXxSae+ClY
soGkHdi+hC+ovO71c+5OZCYYlYVxoU5XmeNdXxBiRoL15ZhKruW0bUuDaMNVKtFx
o7T0HxfF5VncNhezSj6uN2ju1RHDfztZfXaeOAj3BUwjW8zlocFFpvDyvJbE98d4
S3EDdO9uVvdyST73qE9t0ozTrCK+uyMJx92E7GFXaQl87ynF08a6ZMn2+fQZiPz6
6dg2vMceUCCKnAG1wIXMjoOA81TOPNk/+Mxtnpyp4E1tTfdbbN/eunkkflP8vofJ
Rsc/lE76YXhNwmKKQMLrfZ14PgIkZiwJZY0GusPi6yYzPO067BfCkcWB2ZOvoBKE
jgR2Hdq8HB7r60Sb2V+iWY3Ty6gJmIjtOrqMizXU4EVVaMWAaxgaaFmB0tZ4/SgE
e6hIp/gCrYVifsiuJHVzFHrqFSir4uf3R4Z5sPUNM+Wp3N2H6zEGt80ufGMTwZGR
CQzMR3BtT/6PZQdsH5NmlXQFniOzAt8cdREZhW1LfSYtyX2kXZKsEHZyJd8nOO5q
LGevjZfQbfneeqCe7onzOd223UIP3VVf4QIaQCUhDEtqw2SzSZ41J7zKoaViJ1G7
qIOmYN64CYmNSEGq2Aq562Ryhg6cJ0+eXdF6g7vFcLPomRgRR1st+UBNRAnoiwbp
2X2PIjp1bHBes8zOmEf12R2sTw0PY0ONeUj/QgXUxCN6eZ1qNurSx13AemYKOPCI
pKQaDhlLHoxSLPhVgB7iFcGNdBEpiLIW2wZRFkL1je/12VT860RwITSMI9JRadMH
805jJLRVn0MDLA5Kr1EKjilaUbSrNgH4o5fujPW7uRca7cu8CWSZp9swhIWnFL8k
1NF4CECZZKbYiHTveKrGXQztLNQl5gk7HbguiCcc1o1ApRf/Ma6YXcfQx4lcRpK4
pHdxhbAwFNeP3hvJ7un3zBBci1Ip0rIGUzQpzrTiDXRfMJLsYHOAfcAZsDE50Soc
pWeU3GxqdH9TFMADYMcEtQxXZeUlQOXn78KWzpLAOrqtU6mvGNfPRwRs6YAsymX7
tqQXZfmR2HU0OuXsC6PjLdOfIaPgeXMAkB62NWBJpVCp5TxO/MZ1w1kxoqRQY4gP
rYefwQhA6HK0hWZOBKtWmOuprp+aiAPO1hB6uKrShTzuNIXbU0qMT8n4eG2Fe4/B
oppyCQroEBq2yuwC0dHx64f/9uOgONuHGEylHaf8V/onUo0nGxcS9HkjLj41V1pg
2i8rt3frm9kG/PDmxCC2zQ8ECIRHvsR0vi5IJLHaaF6HTGjAlCVh/yhq8D5JuFjh
AxN6OdnfG3cKFnmkpj2+QG4Dac8chLhBWdzKm2+RP1QJxDmnpH1AM45EdhxGsxQq
DSUDgEMlHRdeHlv+JJrkDbd4smLSEtUrZZcMh+U/FiLaCRELcVZ1+CIkwmBKhWI+
eZ4q6bpgu0W96J5nCjswyL4THFBjl0gVRopofVoE73U8azd39ye+iifG1RRMm2ee
Kb4FI08eGm8wUTPrvQgCNUabek600+C1mCmYtGhJ80z9B+e33bYKXdTVubvLjZBt
xj1EnFt4NxkaFNi012qQ4oo08XOhIBnSj8HpI+H7RDrB4mCK1V/R+MhoogdAIbjf
vQtWsHue6gx7bSUl84g9/r+ywaeQBvy0Tzjqm1ZiSJEvjZSyQ2BdjLpsB5IGGWoi
UT613a8c6obpDNSruWWlrdcRJ78S1zG47IJ7iVcPYv4Ux1sGBGr8S+4ozSsANMEf
7RlTGHxL94O/dPD6GL2wob+EAkVVmcMgDieu/8UbzFy635Gs07Q1UvxutdcujcWo
mrOFcfaEsjAYCBw58TLdoIw7ZkppXHu7lBvfycM2ZABPtqSIBVPSd9IkvZKHv0Is
fBr2qpnlgiiuX2XWJIbZF58crcirgCMsxZTGOpKHMlnpX8MkzujwQyN47I0Yx0PQ
mcj9V4BN1YV6ChsW1QILNuacX+f/FCA3Q3O05HYslzHvVCkkR6z8+2laATHdoJxl
w7NLKq7QQd2W509yrVE5fAO3Egk+0PX5flnhCfcNc8B2wWYWE8duZjQDIoawaSgh
gqOJHH+XFnkJ7wxT6xMw6l1HlIA00UHlLtPAk4Fn4XJN2Y7qHP8t1tj8Wpa7mDZJ
mWFSx2KakiaDJ+VV9valauuiUcjhsmnpOiS5RnBXEGR8x/gEzw7ovboXWswm/i3M
BG4YHgEtfLR5m1DHbiYYAe6XCo0HNd9XjUOXsUMFkkl9LVF99zXxRJXmwWqNTkcw
4TO3GiHCT3bOViRBUhVJp37WIgCqoDrw1cd/bSdpR0e5rMfgK5jgMstFMg/LbzyI
UACLHN4dbKYrKS+6STNntLpkqnLYyw6HfHO1kOI7lxw4rKS5b0R5CvP4+SivGn8c
5SJJ1+mVNO0FMsfrxi7wCnaOfY1Da19xZxUuQDbH1AikfXKfzaRxQl9h8M7B+HJW
sKhmyjLeQmOcIIbAYeP9QBFwmWpS4j/LRRM2y1YdxXAY5FbmVHpkxgFVtY0MqSnP
gbuc165HaPTgj2B693VqGQzwg4QODpBqdLsQLcSIaa37sMiKu3yZGWygYkmCtoVn
rdnY0kv2ALObvFwL/BZHrA1Wn/XmEWWPYW15079iuZw/xQaf+wIyPE2e1mi+54rI
6UvstgagKFWYwepLlaopppjZKrOazDbMpjhuYw1nlbETgKCJrR5SWvQ3FymJxa+2
Ty4yd6QCta8k/oUeritpPsKJbuKK/i7aJOsQoCntZGKWmhYZ0l8la9v40QpXpPiO
T6k02XoBn9mknLSIHhPpP496/bsand4cEmzox54Hg9PFOEAHaifFq704L8LNOtgI
wtM646G6ziX5aDrLmn8yNfgMy0zk4b6p2bZLFLe9F5Khj2B5npbsfopgTnMlo5ab
RyA+ZHsNrmlfmbXzW1VuccrhPwUgdv20pL65VQjbsAfgYOdYzs40urcTc+GZPElj
munHDOXV8pzJfrEnbYffhsW9Vu5PluGHeEz7p6CPovhAZGu6ymUc0eDpzpP16ZYR
QjFM+hCodERUJ6ygLb2V6lSrEDfpQJe6baA/OcLNbUMDJMJX+VBiSIKduP2JgZ2e
lLrdVGSxcVrzIKQiwogniHjYPRMQ5cm8ox0TvE7LxbQp48aMnE1EFa8XIxqWWXGr
RdMV/x+qRa2Uo5NCWiZf5qcd55jiHuayCvYsKb/388+lSKA+W2SwR3SQxoJ6x9xZ
p6q8IbbY7cu+aMDne6wHddlSCyuxLFu6pFFVIC6sd7Nfdhsq2h9fofA2BDtiBfU3
fjf61+tZmg/T1iIuX0yijZOErCFeqkwEh0CkchOGpfI3oC4G+EoxF672LHn+/8lD
BYNJWkfLGCB4/Tj+lKFnyIQOpnyYbsuelMD7WeQhH33ZYmewcw0Wi7Zk85E7qbP4
OhcE39KNH+LPC/npOjlZNe6d7l5xKcYhyvAn+4m3VYDTU483j26D9bpaOKx4yIu6
z2RvRcJT+OMdbFkxISm2TAKbFC+P808ShZnQb5huiNIoLtz1fr96k/pnxTdFRQTO
gMfCrJe9RKx9mzPBr+np7h5ADkejGonNMcobai5lVaQ6ScqzeQquVpSaTvDJ8NeD
pgVyQaHUc3uUuW5831V4IC44ankTJ6Tp/DleZQiaxbw3iy+cRJ6abRkvCBBZ61Wl
OWRQKHC+vbMwQMg0ptmZ1ry6SdVPnGCe6EXHWEqmoAMepFqeB5DxaCpqoir3xIKp
eh/2ao1FNkKqmRCEmalvUCHW8fxyjh3RmOz81jr0Hlj5IKAjltoq/DWzUjDxgL/f
OFbx57hFcDLrg2+JBAIxVW51ZmZRVPzdW+VZKXF7g4BlsdTy8hv1ZV9r7puGge9b
J6aLn0MylEKXGJCtvweV9k9Inn95xhsAqybLa2h0/jP68lrTPtHxdA9aAUPZbZmX
U2xtTY13VvyNk3F54ULuaUleMgJSPCubojVowkcBtLgPXAXfAZGT4Xp4vEErT8k8
IIQVA+geK3PqZdxxnWQ6rj4XVo4AfZVBMMT3646OWFvc/rO0dB5c+L/aIv/KDmqd
gouo3krEEs5xIxsUOKuJu+C0Les8gBMspqfNmYcHgV0KxZlbi9XILKT6K/tuc/OH
MxP/as7eFpcMdYUjlJ2hrMQX6yhCyfnuuj79bOxszjTphypOvJr1FOlBuoLaONlD
N4dTQZEyjS0x8j8tKeiU6b6EB/SnUGhINjICD/cYwAWP5pOq4on7q4F2R/G1AznN
XrNmQDa6L5TByFfeh9JVORg5x4LLRRyMLfQW7qtCuTcnh7p4eREAqiOHy7dtTtk0
s1tOUqZIIx4aanuuXLRDTvzjLUUPNFbL8T7pRpZ4HsCbvL9DiKtH4b/Ivy0XO31d
RjDWBJHhkcCpKIzOdptsYAV0RDho4m6AvxZ2CzAMH1frGolCRdPFxYmSowIW7KOs
+3GaZpQkw9hDjVXk7pObsFx0hmod6TDRTDps24uKU9lJuBqsvOrtHaGdC4+B+noI
PNBA+TK8K6xa3J0gkgHaLmS0DPfEyYSWE92eenXCm/rUwizLC5oN4ibrgQ+omRLd
OSReimpLGcp3HK6vRmQ2Jw4iFdSdEHpzNn+L9ABv/uuDWWit5+FUvIxWoEmQlHY+
Wi94oTEU1xUYyMBBDGU3lXwivhx56wmdjQu7g0fFRrjBz3EbDODC0kkyZgX18BaS
wpccSHLpZa/k2W98fG1YiggJBdQ834YHf5PuSaSWiWxtUWEUO9FzsneMsJitK2Ei
hHOqgiqHPpmHaIM3ZrD3YaRn+Uo3vD20giKxFQS0d8ceThOtI2T0Wo9fNtYxPlO0
G32EKgDrEn4XJtIJ1O7fb0B+TO1Aa30QaAZw1r1Ikzk=
`protect end_protected