`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
ddtXksX2+yylW5zu6QL2Lhnb2d1sD00763mmSITNX595NcHTEkwn0zB1Dry37fOW
FufOhVzEJp80NC5qZ/+F0Vk7Ik02dIR0elf3clrjeJRK85K4e3Hoo4xn7YbFUIms
l/8VZSb14+JVGURjfswrIyCUotIzlzVYZ6gzoZwDXIi5gQIBf/gI+KxNXPaKV+PQ
Ufys/12rjO6aI/pPlqSm0hCvftmBcnezN2hk1UeXgOIuKZnogjOsf0iJVX2aOOWE
6pD/psybjbnsNB6kH5uFTA5frkzIzkzl5d9+YDm9OyC+k84E83I/7/j+rk4L2dah
QJOvksSIzN867/4Qt8qYTQ==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="MvBXkzurAa5VTw+1JJ70nePUfoQXBvZOku/SMmg4TwQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
oRtzZL4VJ4iwysPsC8SXYCzXS8Fw2gtZTOskLcDV+1B9Nzn1zTyNtlo6lNICRmmK
ZRVu2BmCc2G+fmzynYlNTnSa7C0Cuel6FYpxCBlOuk3OF2tzAmLAuDyOH3Z1Yjzk
a0aHuoCdIRKv7BrZCdALt03JeUmXKPdOmIlkVGFl8yw=
`protect rights_digest_method = "sha256"
`protect end_toolblock="Jn9CQpRhJt4rnzZPRk+dOpzAubz7omckX1MrFd4p81o="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 20272 )
`protect data_block
gD6l00tciPUa6pDNTk/+tzLxvdHE2s3DQL3/JqqujQBC/Ei+vcAB8wM3doqg5vTg
mdfn9XB1bLOis2CVSfu295W2DNwHfMSTc/8BhCDRnTlLIX0UCJs9Za0+LoM0rMrV
T7EjVWppbP+Em6PkVKCwlmIQ7JKaifJ+Y+kjw9HCGboYo5074hY+K/CBbfsBQY86
AyoN0MKhsIx+eViNgnWjAyHsRz0TWGT+ds00nGNUf02PkhmCLnrE36m2NBI+6bSE
tNkxD4M9U8hHpCtBnYYOwhkffljIXDcSX0QYYswLtWC3oSKmyRvsPzH5MHW8ZlUt
54d3NBUSF/zjYAlce0Vxxo73SqF5IThRhLxasVgIrn55zRseVEOqa3NRsJjc3ppn
l85nuE5S5H8oIbuph6KYmMqYIGbYs6DcizBPu3qFL+jHDnonFvQd6DI+23PvRa01
7FKd/XMl/bohEecMQE/jUyc1gMWuCiFRozUIFl0rVeqYeCf0fuRLxvWtXKoeUb4i
5T+EamDIaSJVf5pHUn5ApGPZ7bOUsOEzPga6x8Ey7pgakBLCDOn9FerIUqfsYhmG
y5L6UtcAf3gYZXWdIv97htooku9ghaJKv3+sVp2Cxg3fwCiYj2w4EuWrrXAau+b3
fDin9vGBQyo6JUg3o4YGO6KOTyk2LnwJYAC4h7a1Omya1+iFm1w9tBSCh1DPsjMl
B3PrWL4WsPf8YzFSEUUIzXr7ptFZQbAaJoQxyiTJOxcf6FtVAPXVmzD93gi5+qAu
ghbWgJbhuojW9vAMUxCMWZQS3tMwVWpuXXch9bVo6DFsoZ2r18SR+WEoLXgUqelO
YGQM3CQwIt+cSwc0AziYiPAdE6M6OAmvufeBdPj6mqXvP2cByvMS/jHFOTXgMGg3
hHO/Q6XiVKA/LOeafvvpq8cxTlwVQSQ7GjjBAlgkuVIK4yujlIeX5rG5M2Fwg4MG
XXmiHEucEO4yk2+BzPx/311+j7WtTitBGeKdsSqIQ9qisWsaljoC/S0xnz5T7gw3
rzFcyLgQn+j8BF2LEAVpDx+xT6MLvCVHpWoy3CJNIvkB4sFm78T/CEFr2h7vur0i
bI/YPavi9qUfIyvEsnFODIVE5MCe84VB4Zsh+1K8TRjPlM8DYaJN5HWnh4hdLAG7
V4x53d5pkVCObXTQk2Rz7MWE2i9BymaXwiiVJpBdA0YjPTGJyyMJPaXJlH0VwX70
BGWsFTiN27G9IqvOwhe3aWGqabWxfhUrWUxpKW1SJBD7wTiGuALE25Qi/A3z2bAx
MeD5anoCedjNCVcw7mmXycKA1J54d0Em6L4EG0vxZGmBGaeTHbpzSEcmTFX/Gzn0
eTnV/bBJWG8V9/6CGPwLKXrF4bU1spSZul1fQyA8fCgtaqLwIjWpG2ORPWj7epel
0JOUHmO8Km0rk5LVHu6kDLj2+dNFNpc32KRSnWwiXHC9goZWObe0VpjsrKudZvFb
17AUFY9vvSAa1QX9k2sEhgMTWtZIj3LwNxBIrBjQrvTPTPhPBfVDEBYCpv89wgeZ
TLumIlh5SuUcniSlfsUgpqwQxhCz8Y0QmkmFJIedkhu9LOBudiSrQ7EeiOaOd7p0
PDgXsQ/sO0zQm60uRy7wah0LH66KUnQW55mTMELBk9DPjYBQWsXomUgdEf1HGtDN
zKawBkELdjZVGXN7p5Xm1UIhj5S93zmXhzM+T6s19mBAdEIO7f1Y/gX6HC/JhR7D
Ba113kDV3TDzE3Vb5k/fsbDAexHxosqg7AaEb6751zRqdbXvBHNJJHgiRiHqh7CH
te9vcTtmYZZ25jYR8rUmjAghmxFs5zwEbvUdt6coKs9Nh7P6LrbSJzxWPMQTHdrG
ciN+0VVXT0WpRu4shkRaF+rxeJmsHfkGIh3bOQds3q3DN4TNJu6U0hTSssfUOByG
2D9mQJ8mT/kmHFlxJiBYQZ5eHXepLvGCE1BasgP/JIhknTBTbcCbaXYdobP4TFpQ
c9nydGbn2Hdt4OazkYQc9fxK+7kPcjyRCeiXFs0MUwH5/zJd0O5Z56pZwkb1YmOM
eENQ2eXXy0LpyznjHYHsQaalnyAHLK0GzodYE3Z4DdQEzH79fZ8LD+3yQ3TEpSI/
JEFRbK/KduQ88C+0429I8JwsjzS3PbLzICaM8axusnAHf97wfDFiritQqdyVABRx
Fco6Js1jOzmhkwFjpK1OfJWN5BvWpcOBSUW4CrhiM35+VsxE9SdJ2tAOIJnN2JRg
YNLGLVMv+QVw+FowcfFt97xNmjVKwqsHVNl8xMfiO/N+jxymOUSAkufuTTJvCCVx
W6zZNf6qxgr85r2mJ2gJ5dv2UNFoEYH/8edC8eHFwQV9Yuy2sNDLoNe0X5Dd8rEb
h9VEdjImtMLrGfksKWgPHWeHA3BxnJGWKwONW93kFyI27lbe4DrOZER9llGPcm9l
bONFPzRoRMKISyZnDqTVToys8ImhoGk4n046KL1PZ5t50MqnAbm9Tl1qZyhRSt/9
lcjUehilMuHkBPjjqgdq7kGiy/99LWLmSFB4hKqCAnheBii5hsaHD6lgydcnei3q
LfAg2m25I4RPMfx36ACfAm+ikhRZ7tILJ/LHQ/JBFj8X+6qSA0+19ZOGu+oI2MJJ
cefWqe6Be8o3mRtiW5/70p7RGaOymq8bQ7i12mQwJzmfgnKVWHYYmeOdbjiTzzzK
MH7ax3lDFaDiRs1bgENFsR5+ctT96UWgsdbQOIS83bkEdUR4iNXwjTSlOUZ1kahF
5+htsx8pdDLhOK0MVgkWoaNr1a2APZOQ4Rt8ra8SU1xio2PLduMc/CPx819GZoF3
pIcCASumBmg0rLih1ZBq3HxIQlxA3vGha9Upb9JYgsHJiGPLvTEI3jIWGseHUkhX
abNP6adYZmnmbjGp8w0Lh0XwN4eNJMjGOQs7NONBN9lj/ZiHQRmPbTowhIFRCwbn
LpI676jhTtXtX98WVLGzimdQb0BlRCmY5XhzC+OX6e8LACZ6/+SASyUzZGrhjLSV
2NizsUfeqohPS0Yp0YA4pRwFjnDYxnNz0Ru6efeOZ7AtDUSMf7c+mpwPBPNpfd4A
FY6Pk5iMMsIRUqf3H2+fy8gqeLnCiWPZ4hXnuJpmQt9TpJkxhObeYJjCmUI/0eea
BFbtuFVCLKpH5BxSKK6lwPJwRgt95bfAwXLbSncsymJv7N7eJScRmvraYOFJUHNd
rHFUx5+XsVUud1fuor0fwArXEcnewCtLFdRdcBqn9RZ9KCkc4ZkhgJs8nyGXEK9M
w0bH7Ygp7K0HYwITrWfB9T7TJAStjgEHl9ac/5ktQCjEm3Oq5JrtArek9O8qpTUM
Om2yba1ioMh6TnporA0Buj9Kgfw/DAQ4N42u+NS8tgP6CECn4W/AygJf5UB2S5lu
m1YdxFtg4miEUYS9zxjeoXG99fh53AGyWkialTLG3yNAVSY7cMNvipdX+xYXgGv0
K966ymZ3+3v1dGxFTw3gSVjurpZzSHNlEF1uLTqKl6VdyZNewMfXL7UkW0eV3DTg
Xzf8cAbns14AOFByDxcP1pKKWTPep2dwXOEv72HU69ZbFzXCNtTr9jP8TEy3SZb2
kiWvNPEUimngFysMrZyq0wBu3X6DuDrzCKIsvXldL38iGrv9q9ErpwItcQMj/OtI
S5/ss+/EW5OmZdxzqdA6sPHwxLDisdD118tG9sWjs6OFWMBvWcb/5uLieY7NRhYj
INdiv4Bm6Lv0OedBbQdN8/QxdFGK47NlT1un8WfDphWLIz2ZguIDrrXD0pt9n9ao
iMtzD+N1KFk/rL0gSrtGDLruGWdsOs+qVFs6/O2ntEtwGQoEoApplDEr5+qgmO3z
OdjujTeGm6ZGSlC4DHuXDLNP3XDkEN8gKKRwMFGc5cRUUU7tYvYgqdVMhDOHsD5w
tnJ3OQLJ9Y4GwxNIWG/8Up6U+jQHLvuYmzbh7nZZL267LbvJw4h7+IV5iaEetHtC
55QlupiosZvsBHM9MfbP3BguQJfHntOtfBrQm2wTrwL1AatHIM3VTAjdbIFjSD07
nhBhXgSVXoUB42HkQsfWsC7FtLNrM4YK5kQE+rHGdDGIR9vRw/gMEp8VUZKcxypZ
0NwMX3I3BxOFSBIhUz4KosUava2pPuFu+/71gFwZ6KXUevOLc3c6dnM0DNRXWHZE
aKN24v4OCJDg0qyrdIT05gjw3IVtOiFAcPioeJVtNjdRahfHd/SZ/zUPfq04tJvc
2eN69GIxVkAr0zqGajiMS1M2egAiN1XpQVKGcCt0P2xXsM4Z/WgBkqXXd71GqNc6
Q/wugRXYiwruS9THRPzQWvy7GE4Q9tOtPys1wcxnIa7CbycGcAEnv7mTxzmknL8j
fQq84WzO/2DVc5f7rJWi0bNGx7phezW8g/i5PZ9TZDLCzyNfwNN9Aq4X3n+3Nc5i
frqi81NrFl2iT+qXBp2+hLvqN2Pzqmnc83FJThisPqblGd3ReLB7ovJ7Qbwq6Kg3
BcW6wIr5GPdpnzXktoXglRgq7m+e1kFATUeQegQ8vErhXM2mdRbxHac3GZpx6nCG
O8c2cMJ7HvMhmXUFQ07ecUsQYP96Ln9vQB+Yngx+UnF7M7ER0kIwM4BEebsI2y4G
EFSQpDPUR07WhCoOgjans/FDb+visaloPAmsLLzzbSpAs4yYcVQK80jBwLCR2uyA
sK/8VKscyEKV21905btnLhb6nEUFCCjhb27SQp469d1WdtFgLVkxvGyHy6bQY8Hm
huGD9XAFoh7GfKmONBvMmDJK745LL+KRg8oaUxqq/UYMoapc4Yy4FW7HtVytL1pm
uYhx8lgKShzxKPCUi44tO16eQZQsxLXETeCRhSLJxySeTPJ6ee9nFGNcAwS7wxKx
e3EfQObv4YsSHkwEiXc1W8Kktzz90DIAAQ4VTwnoj+YFn9+knRw3gmiEW/3uTzjg
f6MeOWHSrSM/KxoYk2xBh9ZvXqGDtV06M4OPFn8E0HI7WXnU1SzwgxnhU2lwHyi7
ZlI1B0gAIB83JLY0rzWKmzM1AwVJHLMOQlLhwRXX3kn+CDSiYOBRNSvwhI8GPylj
UmfnMdboWrXZWXjBf67p5M5/OjGyDQc6t6AR2cc6OFtaTSVQyHyIPKMF1DIgV4nm
t2qBFTU5Uot/Eozh7LeNxhrx/GfQBr52zpjsEV/r3OEe3qEEpx7AO63tdaX6NHRz
cyevUVi5utcHKiuTdCK8YvxsPtTOgh1SGhP7WIV3vc0NvtMB7i1JHf+jcCGzTpiM
c20J6/KDxViOwjFi5NPXiLtAWr9t6xRSZiRIqaS5MebvIl78AMHLlq5fn+3BwbsQ
wZQVc2a8oRjAJAtkyst7LBY7Ud69E2I3f3PkE2DKT7KlRCnOoi6gkv9XPmpRquk6
OOOpCiZsHiqAMIEF/rawWXcYRPagO52l/5Sd992ao7sVwyOXWBm9kmvLO6lsReQv
PThwxieFhGBLsf4zlojfbco/7b/bP/SunTH/Op/G4xPTtEa0enWjI2opXTPcxuGO
tmC8e3JoJgpqQCo46Jlyg7wakU2404b2YcaM63U8iyRcJWK+jtEXkpyTAQA+vH2R
4Eh3sGk7pUxzLMplJMI4XSL976xkjhCt3trNEmX+zykQKjcigGXZH/O1ftSOMh6t
kUQS3UNEYFvogC+ZlFy219Ou+Jt+6h3GGO2+rqdILX4NIZv5cpvmARc6OgD2Y2b4
CEVyOQddruFxjudXQ7L4SQDWXUnY9EnONNYo+w2byBYBE9kMLxI9mBt8WsdFnRDS
j22SQcxHAg0VBdt5hVeBEEQMBumq8ed8bKTktaM6tMR94caKOOTQ7U3+GnD63Zwl
ZQzV3Ggh7CITtQoI8RtSALWG4qFFHsmOV4TbgybupopknUJMP4gMhjAFlv2J02DS
Yrtvwn92wI+SSOHPN4Tblj9d+/AgEtrMaovZR2yASqeZIYlr/4UNUa4w0h5VvSy9
Q8K1w7roSbdLOm81LZ5GF81iQ7PRqtSoWbHfDW0J8PrVxYCovIfpxDKT/tg6XWKY
K/6+5ivo1nCe2lJ0KYrBOh0C78J8O2haDNkbDoHASW9rY//gM9yhWgeiAV78dFfH
MkvspQSUD4SXbwZ4PxlLfSmXRsBtqiKiowWsI7VHBEZ5rq4Xgzk/HNS8jusDPBU+
Hjw5s3xagMlQsUIVeMqW/XCFWpnsOGQddZaDOWW4jnBUfqOeQiTt40RT041GCoNX
6WWeHPIQJ115Kq1gdyH+a2WVwju/xmXO9AQkaGYidQcb5c6IPYdVh9jpRwnxuzV0
cm6m8sYyIj8j39z4vKF7KtZ2y20Rh3cgeRV4AvRaidqBOBX+FjSDuZZK3zTvekHL
i3RbJJMTK/7qX2bIoHLOjmM4IW6/6zg5NJ2MXyYeeZL1+vfOIO4LRvxHoSnzUnrT
w7xaIErCQxOFgdIWQc2sKvBZGYUJQp1W78pthEOGEV1pqUnB/H0v9H3qDYmFrjE9
BZH7GXjMPiZBBP/SCtVYZwJaBwMx1CkjMK6Ls73CmHkc1ZHZsoXB8MckZuQLYftb
v1zkt280h226gqWqZrXz9DLFWiV7iF3o2GQTsacAtKK+DGGeli2zR4WnHiZ9CbuH
HATRkv+g+sZrZ5pFnSx1VpuYg9O3NVDpKoOrgs8cEx3T7F2vVusp9BmbYiPTsvJE
bjHPCmpaKJP/a95S6atmlT1SvYY3xRN6/tACWzgHyg8XB+oRQmHOjJfOFfWrbm5L
Cf7Z3h0G6t0r7D6I/IkaR4UqW7lSuqFnrEZbIiaip9kpj0bPRbeGdC8fQ2+4gshe
VoeRYIRcBVuEaSEOrHHxht/LGVm8ieBBNWN4GVWJo2Vep6Qyqo5zaYFaTKYX1SzO
epD72lY1n+stf2p8ofVdi95ZCPtnzktJjh8a60WNfC2Bd1hh+Z4PfQU8/eljlBhV
5hRPI9VAZfUC4FWWkgF+qIN+i0yVjHPOOqMu+SaOUwIjE0YwqDKaZp2vxoumxLjy
LAbJmTUYLRz5mGgqZRp6CHmDvy1ddjNt1NKc94bsslJd9o58OwlMbRq9lppylwMV
pwBtBqonBW7aVHy4bAV4ja/fqOF4sdgfCTLeREms5pOp3Ghv9IBtzZeNEasorXX9
L4i0j79M2F6Ek5RvciBvcN6BcSic6Sm9W8TL4RpMYmB9jymrZPRaZeAvqeC5r4Le
YuamPksvtBRv97qcxs3OBxBj+8dYfrUU/CedqxmJ+3xSNAQf9wU8q+Bxw7AB/fxd
wXbbAHPAVeMPSHpO/JEJfE26JuAA2H1421LVOv6WRfTLircTo1roHsmnZVMhixwI
j11d9nm9HR8mip8B+utZEAz98LBujiGxRpT+pv5oPrzay+okRxgvr0UrneWlR+pP
cMfqLNhCEAQu6CjbYeogDdGpRYVpnvfqNnKuXqI7WJsItw34U3FBvnTkc10yLIh6
0J+iQu8Gvr6/YVW2wZp6R0/mqTvEGaWROd1FGoLONqRH2TVLPa0CBmCS2Q9av4IE
SLJCeAsJgXFVmNBJbJPcB1mrRVIt+qbluLZdKe7JfKL9C630ia2qRTTq9T1/Yar/
X/LYgPzq5dUNmg/23ahczy6mRgAdVFbiQa6/kQmaRcdr+WxznDD2yS5agVGjXajK
9Abi9wjSC6Wa+ZJ3nOOujuhV5uwlMDNBzAI7j4mZe0gYThdY1wlE9NKnIlNIkHeT
ztcj3acukEEglGNcI2qbu4xv66vCsgT6eZjkdKs6itkWSkbkCe74lnH+7q7r7Re1
YX+c6iQPpiFXpJerl0O+oKIfrKFSD+eP4M+lh71VzmTFFK/StJmnLT1wO8Vb1pkP
tvllZY5Q1YsZu+5t+ti1ZC36dKDXQra1KDkFbPtJFj5xfPgeMJ0W5gVjv3bJdum2
HrtpowBrWnCQWQqfhWaswiZp73/mgE1EWlrXxcr1Ev/7rEEq6USvG0IZhUpVWd45
gXQJJOeCTCa5CwXB0ukpDOTjibfM6jZI4P/cxZgAvPMQ8pmVXDHSLf6lPm0dvemV
Yc1pXZ5WtjfGS6tR4jL1PWgSGgVY5RDcTiqliK3mdkR/Z0Mqfcw0+oA9UtRvyT1P
6k19f1pgbfTo4kLTg7miacHeqCCZtmPXENDf/AuYzlm53wLoJIatiPY+KCOokB29
sQtNYcHc19kqhMWc60hO/mpyE64CCuQyalz3Nwbr+0ldG3vo/107OHfWvrZbI1oD
KiduvGfbGOhq9+cI0q3KDJdisK7H9UN1lk4CJqHjMMXAPtKgXr90G5uZlR3CeAsR
Bn1/drpjs7Ypmgj+2ALtIveUF59DfbFDVA76FR9NTnazcwpbpTXVJA4NEN2rdcli
K6yrI+9135xGCjYdbSypsxTlrL2iAn6vdzmZqwKJDoMffAe4VX0DqZVXRZrjQ+uI
Hb9lqmg2T6eeqmlZHyvgNzHabS0/jRkoWI6NmdS/RZqF5QkW6GZ02qDenLjHYDSN
6aYnEX2O9a/t2P04aamwspBPjIhprhKxmorhAX71OMYPKijKhCj9Gxvk8i50Qv0k
jVwHCNwtSKBjB8p649zW3ZkMvMnOGwAob4saO59X1zFPMmAkPlbt7fplXAzU4xT4
1S9TfrCAChy+Bdp6ZLlt5pzUKnvcNoSem7330ABh0BLJ5t6nTmk9Cf4paTNp4EfS
1p0MKSEUhXwRDUAKJ5rfZDA4ug6/Bor9WdyeT9Ca97jjJzMODTBcObCb+blVCONK
V17cT7vV86GVnVFdbjFt22QUb2pyfjwG4n7S+llLhODKBeAoOgZGKncz/Bmnkp1u
+ncAFXmR33PBDenMz5mnaGDXGAZyGI5T50B5BvFjhd7BFy9WR94JNcUebL41ESsL
o6/LpwLip/agmieDIUWznXywGQ+U92VMt5wQyGN2B8YZ+B22oX0Gc2a9LVYW2iK1
M4KNrQ+frBIOFvZqxmsj3LxjCyZapVEKRnkjEmbqQCxkJp+UOGQRwNYC5EKVGAFK
OxYYcUxSNMfwOaWaVRmYRP3cNIWGxCDOwM7pUH0ziYK/y4pCxPWnBP14N2Td9Ru1
nB7yT+Hf63qn54P77R2MZo9/Uca2H7/9hOCWx9SuJcEw28Fgu5ucUQFi3c30EatT
q4U5awG/Ufc1whm7rQcGASffMWZbMPtIkIkqN/Zj77XCIs/1lK4aqT3zU7BjhOLz
hQ58QlhtHufqh01a2RgY71zJqYkeGLaXo7L3xzfUnulDs1NQCauv6D1oX43xvsti
rK2HZdImVSdON8twkmcchssnTwsg6e+vaRY6Z2dvAXWeQ0bmbA2Ut73Itm6g5K1m
hQ61bp5KPscg6mM4thS3XpZZQPts+Y5UnkCmfXbKe/L/6jU1CsWqrDADE+peDRLX
vdT3vEVe2SULtZEKWK8Yc7/UxE5iubvZ+VgkeQgS3fUOPZWGzlRbnFXm0o1bTMVV
PDxqpZ3IXzNACeMFTR5HCXQkFxxyLFV8LOkCk21eBRzpoO6J3aRjI0KOFayyC3Ft
p71r1JcF9/mk9bj3P+fbPF/knI/KDiTTkAwT0yp1fgrpZTM+ojv9TmRJlqlTZ8FP
u5I45RY4TdJtrJQ5ZhTATTaXKzIZAqqxgqbod/g976QKzBrIci2Uf0I6yt8fuzJR
69lo/V5sx8GDn9K3dwWhl1Jh7AYf2PbFjpZaFCY/jxITKRoa8zoSI+FtdkO4DC9n
djt34biWuYXQHneGaT/FN8sw7G+G54iA7Yjm36QA+MxMFJ2v/OxVpjWgG9B40KHz
zxBMwbBOTzFu0c7sA1j5gR5nlIsSN5BASE6g1zlHmYNmQcDGm/NmbWEGxUy8XnQe
YFpE476dogu7dstD9OAi25KKJfxpRZMg0mKxweiyZB4HhfrmPsNAHxmy6I+0qq3H
LNWrEpJfMecU+EfFEM4f3MPp6VqcH27tlv29aPH62XM7iywJGINEq5zwVQjDMq9J
VTD1QbpCkd7HHaObjWgqXuR38TSuvQPEM0wrCIOrjt0spH6oRmrOo5mO6HpNy11e
eYBiLiarh564cAYFAxr//1eeZoBNRub2UVl0zI0VtbnWsUlfx9EXLo70UT9jcKoq
6QHFGZXfqPhtVis3zex5S3MlU9QHifEFagVP+et4Qlo1GbxjPjnVchtpifliwpxA
fhiJ+14XAjD+bIu19cPs9j/ZJCJuKZOhuVTR1+80o15n1pluChhcZQcYNnfdnfj5
sQS8nwvWmybg01Qx1uWXtKxA4w/D24Qg7HQzZBUkLmHvDp0RIKyIUiJQ2hNgAGZF
8IZAr7J8+mdT8qWI9AGpFBU1S36MAgztPntOKIjlADHusyyFErHcUDPJW9Nlw5md
BZCgYHmXZB2NI3YSFA55wGqFqppvSLzx9QSBE1jf5Orp63LXByA4pmVHpSmFbjEz
iq37KwpmHYDlnAhzKlyxGGw5lwyeaFv2K3y1UFEXRzpBPtPRjuJ4TqiC+zqFkc2I
SaoWBi2FghVj0tJkK7eirixY3QmhcyG2fqpwqfaWYj6+kRBtelydNEFKjXKhiZ9E
U2zaWIN268h7zUI1usk76cmLTulHVurnczVhhWNkeNHTfbsDYZRpSbaKarl78vK3
qsfJF4o3eQIUwWvB6bVKx1OM/yw0PuYyW8YOBoWiSrPhOkZRZCFDExGY5zy3C/R/
BDOtWj8L+aMIZTRxdQ1Eu5+bYTM+4i2suiUoMaZGTOA53frDysAWoafI3FA5Bjf1
qaXKjsEdNw8gRU0bwQ3n/ZXkFI3JIqE3BganG0y9dVhXEYBEag14U0Y72ryV4kqO
lERTxTJFJtulkKOSUNiFX8Q/EG+3o79MwE6py1uXPlqIce66PtNKBenr+0FTjRwG
t0goqubt6e5c8O546quoUapsXI5pZ4oZG/PP55jiUXzmbhFP5QQx39r9yA0SuZ8h
JGJnf0/73jvI/3VDsG36qeARvaownO9lO9g/2C8e7WX0vNHVj83PRKs/TqZnWQhr
DVWzRnCadnscZ9uNSseE9ZQDCvfSA53mQnixQWVnqL23ViksaUhHWGDh1EiKAiw/
EyC+1KaguSwJQJ4P/mVQ1rSYVPXqLA1ZRlHqAIDKMB8QrgwsBsZi7sz3qha6QnYl
0NjHYKhvpafgyQWM5FCZ//Ug69P2+auausk5KdHzdAKms8hSEKpd3kNF5TOs/cSt
852KWdpdrpHLWXhQUqPTVzqbctFrTR3Q7VcVO9d3xRztvVLsgj0Lz9W4psy70YDs
yHWXAbnVz3wKgPzMCIUPJ9rwEE5a2LTG7xduiSy3TRA7zToelHU+YBq0fwi2eY/o
NhGW11obfFTb3Tt1Uz8jC6d+oVplX+QoUYMY1J5nwqVEDw2AaA/Su4Ww5lcZdIZq
W+y3dW4elDFHyqZaQWI4OIfI5BH7Z42Smi8PzPaNDlf7HQekcHBYPTkoDRvajzVG
ivifeS4ZYhKjOhX33GuE4Ydi6GRcgZaj0XJPA56AzL0SoRQT8HgqQPcirnGaiPxA
SJ/GPijxBhLO440UH2G9QyXNCK0+nKw3BHcUdwApSk32fquZHpB4H4Zh7f5hqxyY
pd1fzCjqUJLif6GawzThT6itnQlg/NpBp37pmvMJ7TnBgdh0ylTynY7aqdL+P8v6
GRY8RpTsz2wDc1zJSnFxX4jNtj3Wtx1/Ngg/lxB8pSx5fT1XHQ2NvGh81VFQLSg1
DbGl2nfSy8IM8Omtp17bEeT6H2FRz++a0jE+diM+aUyateT5UITL5A4f0QSvHVWe
RgWN0pWOGMWjgDjYzJaavaBNSG6VO9//OJwt0G8dSi25vR1GWxACfLLrecrMH6Vp
AyPhEViBXG4UC8pRgnxVRXjp7bBpITAbvEhFXX2fwsPt+pS4cgIv9/DroKdkvOkL
qtxrozccY1lr1VMNuRLqD93OTorPiGGQtuxjfLLYNvmTBNTEYYesMYfv5QgY+xW4
gxdO7lJfCyQpJNOZAzA2/PYTIZY3YHJDCHEb7Lu+tRgDA96rphFE4jC53j5J8oTu
RVO4ktU0M2H0R5NrEPe2+cocpbxQ7/HPVNCpJfB4DYqA3lulG2BpVZ/szHPLLw0/
nlfCboCedSfHLDFvSiQrqfor0eheLJzvGTIk4iMDxCHLgGLuMFC6pcrIfFoL4fXs
yE1MLOruzK/tWXqJoS7dFjR86qQghwHHzJZoAL8NDipIuRdmgYQxdMVoSpEXBz+X
NoNpOpNNlffaK1Cs3PpWqvLvShkOrCo1MCoUC6XWCOzHA8RvEUPuga2kGSNBwBeF
cGLvBjQyo7THp+PAays8swd3qx5zFx4X54Ols3EAWQ5tRxMb8l4MwsA9yN8KSxMf
IlC6YjC5rHkTNOaOABTT+3aTJZpdZLj5a1t0sneZ+OjHWTLHxUVBXntHKQ+rgebK
xH4/z/thpF/jNgSt5WX7owPlsN3ai9FVX1QYOraGiqt4mvUy690UbuJHB17AhHpZ
5fLft56UX/UGqNFkMu8hP2M6g3SDXGYshULWeqHaWFjJVadUm3FE5AFSnprqkIQx
4OXp97gomuLfkz3SQ8ViEw3R5V9O58s2Yq/Bkvbm5/BiY4+t7bH3TBPxGJZK/e0m
36TSCEI8gg7+dCvdrEPjU3ZbKBqQVfc2PGGu1Hy/9OfZ8rabM0O8LB5yIIYAzRZL
c1w1hUxgKqD8p4LbrsqdcQzKamVgUSDWBNKlz1KJUxr1ORX9mlNn64DLERf1Z87W
fuSBJnCy0pnuPiSUEtHFRxHcFHShpICbharPymWR//3fuH6cHPjVQ0MGjIN/H0tn
fWfdEmuj62Valnsk58GjMxrR7zFJ9/iSXANcQYVTS8XawgN7/Jz9eUI7DV4/Pz1E
K5CYRNZcZVqQVPMof0a0vXIrj2TDV7J3VHwOGtzA9hlcK0odpz0NG5dWD0tmXrTq
3qESk+ux0m0+7FEKNzCLmVpcpaD6B04u9bnDiHh52JBAK+kl/17cY5OUTJzrPkDh
hthH7FQIyOKLlgXXdESU4pLdv5cwGiIEizPJMMQrIUnmpz1LLvHkMpS6pEjGP4jr
McPaqCGhoSqM3Kshri97U3HYtlU8Z5jRC2M1pGqtG2Dn774xBsM+BBw9IapW/g8o
EEK/cJtv8ryy0BD32TUDJFgRRDnUFemWiu/ChKr872NTPZQWd+nFKiNKVxHstQvS
EfCuJNZ1RUqH/NSI+dMeIcr9aWC7jwTzXpAflypxS5n8SlvaI0QvFEzQr898F3Cs
Ky0l+tYFST9L/K2jCoJUQlYLouNyEvbJeA22kIcE3JIB9EvazDv2mb9T9G24O7BU
eIkg3tBDukd469aVgF30dtR2Q5Ne2yEnO6SGqtL9ieWY/HVWgf93f3P5hPmzWDD+
Mzz46vrBGwadvCWhTnhVK/lB0+aGpnSI89ALEZUuADutRHAaJIxf95WFABUENs6O
XwhpLe7YFujiF485gS549MUL7SiIVY3+Y+E5HG1MXLrXnWTmhQL4jmOzRGHyatO8
eoHoMntjO8In9zzkguzPj9GZACGZz0MwwSFH67uOL8dqT6rLZxigjRrTpVQiEV36
LvBYaLZgkxoc8vigc500hEXPru1miYEK3RkENhcYnkFwXh1QOQekAE7PHgbyIi3n
VmWmaqTS45gLYmQZHPiq1RuZyPFJUa96doZ/BuhXTbREgf338xVd71vhxmdEhBJ+
DFDO32hHCWQM88Tlu/MLWPnoiXh33rpvqPL66cWdS+mQDRYW4bGUtIvF7XMc6kj6
Dl1QRpbWvVdYLdJ8jnmhoaagDSxuao6mdjbrsy9WrJT6x9uZSguVw22KKkYs2Ow5
FlMhaEQZoL689KuGzPKUruQ71qfmxhUEDHlw1Lft4T0qtMtJ1Pr/G3UwZntQ8Sru
fp+YiJCjRV7J/+x8HZD88l7Z8WkTJHb3uO11Lg+5RSqu/oat8jxbHvGJ5qcdQo21
vhNU2GKiL/ITo9YFq4h3ShkcBFsd5+3r08C9Ah1l29mxZoajPQ+hnnJrpPMBX19d
f5n0Tl8nQKxKk/0hiIwzPXRfbJ456O+wGvQIcSBQmCes4YegheCq5T+Yc44hnOOp
Uau93wS5SpmDTkT42gp1suz/catxSp7w0VoiqglzDygNUGb69K6gCv17iFjy/Fui
mp6TSEekLUOERwErHh6fMSSxI87/QoY9DHkk4p2zqTdH/iYmdbAgR7o8KVDRAKVa
iaWVLsPXT7ZcjxF5+4E3z97/HG7r7UCjOSTT7BjnVpZGqHeTSnQNbBnPk7/xRGbQ
xJwlhJk45iVxfXoXZwRINtmGVVCzlvsp1tqmZVBGvfrCX00l2TXUSiHN2jIrpk0l
euIweNJSthpEQGj+bY+SEW3LKhu5iWRK0boUOgP6f+edZ4b/Um8SOog2PVM6DjA0
e2dreFMpuFvYK1Cp/V84dVnqvYkntbjPgLYbXkPil26AixsuNZ2La35X+HKNiN3t
+T3iq2N2Vq53HxVgJagXWnP5fvi0TRWwUn9N0JxVksEEkvSJuORew5pTMJin3pU9
NrCqJNDR7XPjXeRONIyUwd4oAMdZCRfhLcVQNHcBateqLb+4qcvconmClQ6rHfle
zwH0+AXltflFNwkyiwmjPROEeFaCpbofsevs+i9Qf8fvnRThSte0XuoMlsECdjJ6
X9bCvNs01WV/CIjiAvv8o6Q+3bMjYTpU2/nS2gT3OtA0ocLhpoxc69Lj9Qignyap
uj6rgE46aM1RL2QqTy8ztrAqveMPmxc7bk+FdCaCwx30a6RpC2Ov0Dmc7Sjp/g3Q
q8C3PiU8WpdWl132Aq9cevyDW7A9v0O+epKPyfAc0wOwy3i8bkYf3jrlZLawl04M
jeO0bDIsf3LFrPDuz7a08DPO6+MXRSJe0tPHE1FNRg8XRv3ifqmHAH8yl1F+mnE1
V2U+k7eeQXDtfwSfVPV+lUg68laRICq+AUoa/PcBdJKOasm+9K2fk5oNkjEvT21Q
PUiKgPlLEzz+IvAKB0wDCN9tP3EhEIwxhoqFfcXQzg7I2mVUvqz6cPv7+uX78kWC
kZTX9FLC8lA+N+hLyx+J0BgBnWs2nxNR8d8NJyxoRajpJ7hbyzpMoCzJjaHYusIg
+IlzG8nmRdxHKptTJXZsL0n1QtJmOZn5je5j/HgV2TZhiq3Vouy7JPCsHeE0cPHh
sek8Uxx9gwpn5wRzU5b/84f8kPCYa5XFWrhQ1Xf7DM3pP6GMzVgxrcByBvGIxWqq
RF3tbKYxeeW3CMzfxS5AYDXhCYFtwN7E6f8UA68npT+Zd7+tDYeFbfFssTn7co8t
IfIuF61ci0lT0Ifh9ws11BMZmKdpootIo0L4KnyhQ4zrxjGNNxWO5f0hpC1oYsBC
0WRztBRSL8xNaVkW2UyQBjsfcRp8Ka1PubVvG0rFU0YJBGakiMBBgCG40qPrqTlP
n3SaPPyWEpEF7WXRLtxh5lroXj1pLUalJti2Pkb1ZSAsCQ80gxL99oEb61pHOl7F
ROT/Z4l0c3UNuFvtGn8kmUsWDTYAIH9qTiNyiQVfeUTtD9rWmvnc2eTvMeTgVAnM
49PcLzajB1bCvkYj2FSw6KDmrToQYKlKfCiSGk4kNTQc/D98PRSkRo54S18XpwQ8
SMtZJT9CoIMbHYZW/sY62ZdXAnRQduEzQKYilkLRGFqfGQ/4u+qYYS6ZDx+Ctrdn
7/gaK+oaZe8Bu4dZwM7PRjGa8VG/CZKVot628SHmZiSuV8J1X/7aQXax18fNJ121
xVrI9ZeiI1XFDSvpcIEL8C2KETNCORLJ3U2jpnyMzP6oyYHHAqnEkim+3z1qMstY
/St2mFhjW3a/OJ6T4YV6c6JKhPP1N24bT0494M5hve7sjw6w4RsFbeC8xloUGCNY
Ijy0waT986IcKCavjc0ecScMQxqirTukKMmyDkAzEtKbTETP7j0gQbU/nMYDTZ4n
a6wjwi1S8QN47KDvzFCLzW9mH6p5p2o5lV8lOkoEZ12a12H2WcBH37GV/veHQiP3
32VMwywKeEYdCBikiHJCcENKQSzt4qL7ieRymKWSTU6zoDNcuMC+FzN2n0SnPvZp
Z4FXh8FbnNdzWRkFJYL5xjLtg15YI/aOyH1/6kgIXAuOJHvQzfdK8terFrO+MN4p
anrifGJh01dUP5fYQOz+cIlxmyzd2qk5wPxoM/+bucNZdGYpmbo2PJ/Yb6j7hZir
i/cI248W3qY4VLn25sKks/WwaFpfN25uT4gJHgMCIF+sKGQsyF1iDsm916IMB5+3
eczA1XFahnWFTGfS5DeC5ThgDDntsL/WFRQDWhqWmp+z54ajU7mP9StmuFsVF9hb
FZsi3I6LWhlSQo4aBNaO4vpw8lOgUMkjDZMgYG/32B4WA5xHR4+ghEQI/PLuECGq
RXxsJBohU9fkdeDsGThgXCvsj4w5hm8rch7VuBelBpi5og2UxGeQ8PIUg1LIJ+5B
lsS4mtePvzlb6NKrKnKLy9j4GNqPuSnpzUipxChVGQCqKamGNIxzHMdtkwA0Wssc
pWtYUxfiJm5nVpPAz0XJxFumJ5ulo1C6leLVQoNoU0YcREGOVHdhIDPw3b8J4rlN
1bbiKjfTtK+3bTNYmmU11RZmPiWLiJcPfEg0TGci59icFtloLb5p8CxkeoSFjq46
0b7Asvq2gHxXkWWwBH4oiDW9gGUARRRLPpc63ayZL5yk+lEdwdAZEVIAiZ0onpDt
wUML2aTOnq+Lx3g+jUScFMpIdhM63kdP3nUwUpj7wbeWX6+XbRd+UYtzXl3MdAEN
JMwlkWLWuchGv21NhI8njT+E1jDIJUKfsvD3AMeIcwjC/d6kdHdG79GIfCjkvW4+
DPS9AknJWxDkM7Q+JMVv0rF81rxPTm8Y+2gIa6d6ciXfT+9nnIL2939M0ufbdiF/
hlfHq2JwAK0Ov2eUAll5PJ+SvlMeq/xzkp1au0Mz5Ql8vMCs44eppHk1tsQyg13d
6IIS2Eiy1FaW5BAvWXv1IhtEHy2retB0lvTGK4oDdfSx1QVwq5qrTglTF739+voh
/r+98KJbyLsXdEIYIe3e2Mbb+1SdJ8WUQI2dwdvVFx71gdhYLPruDb+o+OwgYdXT
lGPTBZ+H88dMYoc3UTTOgKkdTS9gsVUAUmpahWqahtL1q5Nibp3Pod2k0eGD5T+N
Y5Ebypc1jfK/Mi6DOrnV7Gz4OwNaJO6BCxAj+Tksvm9xAQoMoxHmPVn+CabErJNh
X5EFM1Cq2cjrboVgK1PNvRMYn2KcIYEveakIbkAr8ZzGFSc7ZMnJT+zPQSTLiGHq
2sG/QCSybYUxg6K+/q7zR60tVDagk3/Y2pVStb6YXe2jMxaNb+6AJZ5bHy+6jGPV
zIF3O9syQjoRpM9nhSPLzLDGNtz7IG3nw8NvWvswOTXD4yx9e1gyZtyLBkZ6+IYP
gxzcUBeBSPx2yBNIyOnIRmfhiiBsrUF8ZWnDuIBg/P69XbMKbAaJVpGY3ZA9uBPu
LxpWhcH1OrdL1T/OMT+GHxaVv+kTSzVFJSlSGxIVQCtxICnSwBW2CZPgKnJaubaG
jU/0eWPfTEXqobatPQeRF+iauwiY1IVH/Db8g9RiiOAwJkJ+DcWdMZYkEDKXsb0V
jL/G2tT+nKqZp+AreoH7+zwVCTNiUenOogvpGbBDyMIMQMDPymvatEYZb6YVJ1fC
+TkhfgtkC5bhiG/QDZ2PeIVGODl4S8e1TaW4+GcPHbHSvcuYo+pphNCR87N0xsUh
5/ZmelxID7efveYngXf04yctFKSuHZBuJ6y2LW7d03414BZGuYtu3v81eJJQSK70
29GH5rzx/CyUC1Xu09iFGbtA50Mzr5wMSjoibraQ3rBNV4e5LBCr5He3vxe+fyfr
fPnpqBAGztoFyuu22O2GQGcfZ/AsSgNb/Mp/KYsqDQyEJXHRwJO1/ZFNuq7i8aMp
NyjFA02oI6os9kFhOMFUQmkrLbqBUtXhfaHJvBeafco56PWUbav+KUp1AzoUwu2b
feUjUQY7vjlfn9xWIxBHYUgKVw0Fq+7GAndgHBXQSLhQki5RMDIrYngmjsXx0LNw
CEqq2VRRZhtnHzjufiSqMy9a6xiixkZi11Vd3nGxIeEDmNm7bcIWh/2WVaBbfXJd
+I+0Hh1uQdcF8dLZqDTMmFZjU+DrCGO9HhuCe61Vx4v4lVPzPdmErE2RxvdOiRQq
o2KreJaiXbrYe8v3xl3ndq8aiFjn/zgdMxVXOWVj+ttWLRKat9eTWgMS2ARaoTEx
EQ/nnsAzngUCgtae/BD6Sm/KE8hygQ4Qfk3g48qm9u5bPfRHs1ZWENPIltTnT3Ya
t6zSC5+Rvyp7GJArr01V/gzvlhLrmLEgtS4hnOviHBYmjG6BvJyRtLZQoxilLwEd
qRaBv0c8u+N6hTDMP5FNGi/wDg7ASJjKHbqOAixXK/DGUTpMbVogQwlaHdhfcG2E
P7PiF4nqnXG8Mmyk+INANSQFFgvF4xQkDGFiI0frnmJ5gdi0ukAyUexf9sthnCsi
zRrWT07zFFWJJBDWrQC8aLwgElTsoS+P3oVRIxD5y7M/fPGZaIdNKmRCYDL2nRLF
PIWPd7cbSaJL0aKv/ssvZOdKIdsOzoHIAJCaoZZnSQPY9Lls7gzRhsd3XhJiesKg
uJMRRJGvmdX65lC/XX1BWwPAEx0ohQ0wHPfbUo0XzuQ/Pr5sMb9SoFW+HF15bXnm
+eKDJrS8R8OC8xbFdioHCxc8fonO3YMtQvkrVamTKDfuVhEk3dALRkU1hfQnPvmK
vAAYaknuJNQ6Z22Gw0SIwO0dJO3AYubUHiXVf0FSxHxlSNgjQSBZehilr2WsZNKJ
dVwn1KiHa5znKU3XwzPSyZfTqtjXUACqnOaGvB6nmPytOhCSB7Hbj0SflCFVjy07
asUs4eys+ZOVIPtsascEkrSnPyb1vBIhW04+v7Tv0RVmLCZ6xuXjGLx7KWn01lK1
Q8GhJxWs7MaJ2M/k5ZYvVdZqi+CZ1pSwmM76ukG4lmBxDl2z4IGfc83MVubPuJze
LTdg09NkHaVJVN6HzkI6Gg6rQNvRn6q7+RLg3l6+r1N+NXoD/Kj3RW8GNwc39CAi
xNHqjzrD8sc3VUR7vKEIDLLffCD18dkzJ6iWXTp0W3ImEPV+A0sRUUKlRIZ0DPhq
ygqNLpYpVOJY9CgsMdjsKKY7fmYHxHrI4cJxKPShFp7CcVDtQ9gKjjsRyTMZOoO+
BxCFePMuTExPMJaad5GEUbRulcIaK1cFlOs/sqPNcAFMD502q7pNBjFOux+btLdM
36rqSp85FTFCv4HbpMfu5eFNYSwEdb6IXfsy/N6fCVmKb41LItQj7gDhs4Cc+rGS
Nb9FCVb/AO+vBTAEKd0p+8dP5RO++BWRls6xaRilNNqtzLTN/oRmv2yEcnCSvAUI
0iqJMS3LUqrXFA1AdWoFIn1O+e8cghOb1Bom0nkQf7lYEsKKSz7u1i6AwLhUV1wG
wch4FZThPDfhhd6+8GFtK+OQSQt/3u+Lk6/eyA3MqbpSaYLnTig1bfAp3rrNIjYo
BdOXunJdFP9qwtUc6jel2bZvsygMTGlq0tz6lbGPptcUWtuisou8Oo78zek7QmZM
KqQvdYB+Ns2GMW+ypoQe351UwGbnY3PNyKpA2DjZvDCC701n+zEkW5QSFqV5ARyw
xrFmHzaJwqA/HBOuNQmzsRS4+Ub/Paj5bHCiZ22W48T8ditbyNzxzDH5p1jKceKM
bEhHfe+8D7+6DCN0QA544HGDIk7jvX7f+J6UTlyOKNnZ+nEfFQaDHhPRa+XbACGw
X98+EqXE3ulkl/twvvq/WmhHFkjSMjn1LNSj+3obrzOlii3eoKTg9C0ROKzf/WhT
Q4cHtBrp10wL0CBawVfvS0xpb3zzsw1F3/p6vVkezZ+kIOEJ16RB6Fxa96fxdoOv
rAO62Ei6bDpx24Xw2swBXO4L5M98dykosvkO/LEkavI4kjHtMZbZoXaGVVYkeXG1
E5/LfPrSqnX2yOjvW/8DMMRpb7umbeRWXBIbD2olD5rPQjpURzrOIyRc4KPyWnMD
XMDbH6iNkMOv5Z9fXnXs3gl08nJZtsCNcqhGmLEAfTXMaqUbmOUoSga9xn4x4LLq
P1hyOdNlYe4d9vqGcHVBYXgmS2pOJlXCCVgV46kpbCAs+K6UZZKMrOlMU1UeQ99E
Sj888t0R72Jw1t+4fXUumTfPhP7NGrUrN5ZaMCetiBJy1LWGjlMCfw4dj+sqbHKc
iRry9Tsso2veAvVWGZsMvGUxhmjXNshMAAnwnlatE7m02wFs3YVW9lqVd2aUckbD
xOCN4HUWvMjUErupjnMsKWQHeHwMCNHORbisJHX25uIaVFhiFfCFE9+AYKsdJzmF
hHuRvIQnEN+MI8vi446f2pnsErRk8ERWZ464lfpiYkRnj20Tmedfv59YC5JYyPqC
UOIJakrHLZwhPPQNdIxYtBrGDeX0K2ttu0Qv/0Dt7wEvqVx/AKG5JZh6QYlSXh8v
HNQeZasrVBqy7fe9NXi99VVExgOFmCEJFWtoJuwRlpFt0gGCJnYPBJQu/OVMAzou
ScpQTg+/sBlY8PlEZSBYh7vU/izvlTJdda/jBi6T8DzYy9iToiQsFggRnoT9wCv6
3GlBbVDgjdy/RzNYFuPn0O+MRksSTvCJe4qC7VHR0OihWnp69oScgUGUSjszax/J
KCPvSod4TK9D4+FbVYjnAT/5KJ9ZSCKwj7mcq14RdjtUCYCXRQ4zj+58pbkbj1Fd
2AdVm81Lb2PXVOYFlscJeg7MCfbnwF5Gx6HxcPAc9Mgus17NEJ0w8h/vkZfi5RA9
1L9gGqwmzKVYPON8rHXFoOdIsfRXSId4LP75tc1jM1CHyIzTORqtu+5SHv+lHDGa
MbNuAYFFcUtI8V6zaHSQjYZVF4Heg4wrtNIulNcpWScIBz2ynWJqN3biXNa6D7rh
5at4kLRZ9K1zbMevWiauACaETNEiv/zIdne67aLEB2YRzY1F00KnIpJhZo9OiUOq
JHWiRiQKMWVJ4fyXqGNYfzR15f3VtCHAOJjlMjLMdOZqBd5VHdmeqALl4FInUleq
+daWdky1bE64NCG8rX7Xt6yKadePTr4k7PDbVLsetnKM75TBlI8oSFWAdUUBQ1To
JsJWEyMvE4VQvGjD7suGSiFGuvVfzm7e91HaVpZ9W/BWPyqHgKcJQL50kJErPsa/
pUds6IWjrTnQha0l2SjQafIoZ77jqCXyY/arhf4PteoGDDpWCLwxIuR61XFaey8S
jj2fpjBJKX8/YHfGZ4BHvkZUwXIdeVImTsRaTm2WemG1ZWV/jVhabdCXvWYP3gtW
RePVcMXqyjnTsT+lkxmy6FGGGI+neBd2Nq/v7TJiWD1Mq+f2hzYJHeZvIbSPLD+g
bCNSH7su4hucJFz5KwXYQk3ph5Il5epHL5aRkEQ1R60TrYoxip2hzXABHbVXNGCO
oNxDBTXDGrwkuvHubINMEUmv+qTxTxgneIQahjBcMp3BISoSF4qYverywu5vx55F
Zzjn+Rt4G6pUvSpdAS8KLLRBAGZNKtYL3+o8Z8gSGiyZrtg4UUH/cATQWKVs9L/4
OXin6ElhxEWRJO3F7CzeKYjHU+cvFRRODMdlXAoROST/AQP/OyRrTjhxyF+6PtlZ
DKodq2erZoulnxChUChZ7MlOqYlFJr1OdWo7zmaO2sgR6/wYZZZYF0iL71CL+/np
3kAtrvGCeSq9h+yP8iCN2vFa0Vf1ObMlUcfJ/cJ3n/64v1ocwo5sYd75NdzF+rP8
tpd52p8mm+YjwQi7gniVfEQ70FkZnVXVmEjO4n3oXHSlzrVqqBPALeHaR11wOphr
XgQvvHwfozkOdrr3B9cfPLH9s7+/dNpGXOlH4u8wfoZ5EPhsxF7N2gHIxxzxC55y
LE7v7rMVDQm7BkL47njJXqysm0jaRjx00TU+8DR2aQ6X5fZHuIeLpv/F33i5ZZJp
aGmaYrhiTqkBrJwn4PYv3tZu/3dyZa5hxtQOSqvGzELL+Jr82pkNliYrpQPResiw
edSVLXEaz3Qo5Y4WL3szjotS6FhdtYnP3SZsIHokvT4UBjubA3zvFaeR4dR08m4z
k2zR5zBqOAFuJSXoIqWiA0vn3Q9AC0rr4z5XOns6pNTKQweHyxzZEKdMzXyOI3nn
gKpsM3LtA3vTDg//cEx+sAVL8h+bNRCRUuMJR9QfiMhDYEGOd6DjEoWLsCTFnAF5
qKfVToNJ+MmX0ESOJoKhlvMkEnVv1WFv84Y5DFGPRXXTnWw0N9gzu46+00GqxHtT
Ihmc31kWTkXVphEsUeIgpSZyVwJvh9LMxYlvCWxVZhxeB9Kz1qBLI9jiQ/rXR2Bd
RLj+QnbvqKkrQ1GKjLLNTzU/gWhFm+3uoLaA9VFQoZVIHlLEPUfEKlBDIYSHbeyN
D7aikXGmIKVPo9ryirZCiKX41kGnmZDyLei+X7cmdxTepIMFGlINqGehlXZesBAT
YZmIFqKoyJeXJFzn4jiZG9kEkOjrcrtajvN3YG702P+V+sIAf+Ok9SZwYrGqtZKm
avQAJAFtN+2bZnDBt9Seq+B4qXjOMhguOX4Cn8G9XjOywzhGMJcCCVvE8JARJnrh
IJcWz7NNPsd7v9QYNAYlU9YAmtfBVbv+bl6haPxmwP5tC/6CJMYyk7dQrRAZWlkF
C/rLo+p2UbOhqkFdNhz52kXlfz8Tatxtf7Z6FCnobrPi6/LD90VMbAnguXNQQ1P0
FKQx9/6BE4uonbqUUHRaXj0cdc/1qTz0NJHeZUMl2VSUl64J+sMLPJ0Sd6TrVTqE
uzsOQnocuo/wdxMD+EFzqDlvuGHMNic1kXfA17hg5StfkdmgrpC2PsHW+sJ8VxLp
jtS8SN2oCLJBuhzPN4Uy3YbyszyKnSHqSJCFAAYkOsFXgBPK0pIqO6EFTe9sNDAz
u4wTExOea9QpTDYCSxwEaMkMEh5b3Jkav/dg9I5F/OLuu4o1SMMTQqOKqaz4v/Si
9HzvOHADmSOIYgT4EX8llTFhBMtPtoA93ynUaS9IOTAiyQZAFNjU7UYHLNiFrzsN
lU5p4xqu9z8DhFM2qZ0nqq9C4imSh2jqNdaVehqQT5VUtgCbspMygOJLaZ4i2Hsa
eSTVuolKP2FffQoBPG4FYo2raM8/1ofqjWTawe2G01K70ZwgjeNHcDm8vWVM2MBm
QYRX+m/UnspPuw3+QiSW8L6KLxieg4EqOvF3pJzIBlKLK/dmdBIMaop9jQ2C9eY1
rrsye0G9oYgAxD/SZmYZOXjTgSu8JI9UdIa89JKGTuVSBQg1BwxZSe8NoYBzUTcu
PZLosR1yQjS1Pay2mUixfRsBYiSYgNf89b43XscLzK2Od+WGXrup4Z03CR7UOErU
fti4H8yrYCQJ8H6Gv2v+WXWNtU6oNkQDtuUzl0X933wG1PgMdd3rHLqUNHnd7FYa
SmN1vlwPW34mM9QxnMdxZeYnE63Ece3e2LAoD400gF19Q975ypfzF15CjDGLKCNN
vlAeZNPzbUowLK3pUsrBK4oyiwZG+LspfE0MvcggPyKMbnKdrJV+HUinnngpROuv
/eBkcoqgjW06Lb8qM/zCBXB9Ro9l2vkLBEN29Mnr8mT/KmHE3LIzX8qEDqTF6i8b
DTQmessQZP1wRCMelvP6R4FPag1SJMHkFnbN1oa28Mo1mFTpL4O8dsNTSu52ZFVe
fTKxpRGooysCic5o6myt2xUbePyeZ1t/Ga21CsjdN29ysA5UEBHup6vTP/NsI+Hs
F22g9lunXc1F7Jfng8nPq09y5ig0kZ6RyfOAYx5e9prGvw1TnICMVDwJM2FWSU35
Exu4jS6Jc20oJkkXGG4yyKA77IKddNOPk8OC6lQAKeXvVMPG3hE9O2L/wjPYwyM7
mpP6Qy26J3F5WVfJA9kNs2hoiFvxdyUBQNL9ERS6lIZ2LoG060p1pLQYN1O+knFW
NAlu4hxc1+J/pIxnqMlU2tuUnMJjpdZZDTsETGjNkmeNlP5dpOz79BPxJ3t/6idL
g8ZRY5MWPbKlpix2LUytr2y1Xnd3veN5fQ9C1jAaRUn2jji9R+PUFQoXLfLzp9cl
ZvMbwTSpRTHjerDkmTu2ZEXxsNq6cE3BVrM+qDpeXnR34DoAM02/jqX3t7AKBxji
PUjaNus/sWDuPJCeHJJFrxiPmLZRYtPxSG2ohC/644QibYrX8nMcaTq6l6Gxun3a
r9UJvUVJuLYjdJCjOhSaXdhKxPQk16xLKh+mVQzwlGXc72jeAX5FxIKjsRvbiTSJ
bd1ADNRLXM+0JyOgnGEuGOAAWNSsTtEuXi916kZpuAItazzu96/rqrVfbXMYaNq9
LHzGAnwGGdr4E/vLEiUK+FVIKpE7PLaRUrBXlYuZqBp0QTOoi/i8MhtSC/w0KwN+
HcwigFC17a+ZLrZc9cALIkafgGTlSLNpQ2isGdXj6KniUXQt7hIBPUC0vO+Wsyga
+R62W2DLwo0wSiNdhlDCx70+61RQOuZnmmOmOCsmiZw1o39Fc+1m75+l4vvp6qdZ
ewHYbYkMpJJAMrgC+l5QAJVxO1g66bOhcLpsQNpf98/fpxb76GnpF+e86l7waY/g
exOvK3P3chHHXhYHdKwYBUlEJ22j3dZAWEl+ov39OeigvJKSkPphToJSydJLUYeP
BulzETNg7SRUYIlRSTc4aoq42EHG0UqXvlSxGy/3qlVF5csXgNd8YuunG3miiv/4
JIU1A8iWpVR3zstz+hIoO+TEW4UgJ9v/ksuCWUm8QFja9RRpt4lK2iiC7px7xPTK
NDF/G0IDyrfXItWyKKkefX/9IJ2vEpZjfQn2Yu31reRbwuiJcYW3NOV07kvX2/bC
gbxaN5OukqkieZ/qd3wafbysVfS8mCcHf/CO/w5XoLJK1qNI1WxnxRtiY8O+YVQ5
evltr6Ul0MI8tnK6WypWJSbmZctS9cDXG8DgXtNmUx9kAJEPTuuH0ahQnfYdAjWo
iNnan7WvCjBlSzuoAq9cG711G8/Ps2cbInSy/lMHFcgBg9qO+1CAU6MiFcc2uAof
sug89dDh+jymsePc8IzKnbe1IsNGw4dhz3OM4GqJ1DTZJT6SQJmewZC/clIhSzu7
iXzTmJhbsXdTvIAPc7IMKaNfX8mlZiJ1gKB/DagL44Nspb66LljYuwfTOCF2XxNc
VC3psb6CRqTxHPROTAui87Z4Fjh02EMedcqS++ZHSBUEarbCQ7a29LQxtIFQskVy
8HcLzgnAEnRK46v83uldw23WhR0gguD4CMMlJXlwrVDKtyK++LTfCV0bI4Vo8vpo
40IgMpij2oAP0YwWOfqBWNXxukrs3tybArzATWKkQb5YsjtyGO1wj6+y6zNrUM53
bkj0h9QIRoZ2OeOS3iBBz4ZjBbEK448bNznhMZoZUwC1Gm27LcX/L07lPEHwHODJ
DBD7i+RajuC5nyVyBSsTU5+JIBnym38fqKiTlWNluawOUhiD51Fhb1Qrm9QPDq5b
JTeJRbwW5Xk8TPZS5xTMka+/DWWF0bsxT/IulYXbqOdn+UZKh8qDAEdK2m+INp1u
A2GnDmm1zt+/gqc96EWDhbYYV9ZQYhJNUDpoO3Y8bFd+E5axB4rDrmXk1iEPtvXS
/8DAv70bfBqkzfB5GDI3tIXlk4IAu2iWiYfS4y2nHZyt5hR29J5VLkJ/VxMaO2jP
TqPm+876dqdmCcAiSt6JjzPzS6KNh+/tqshHTAJi+lbu7a9Vjutn0XQk/SnQI3uA
jx4YANTilsEqo48k9h8oFfoCUq7rRcSJNMQzmsQsNTKvgfOgTpszRz4DeY+0jgHF
scB1HSR6Bdzf7CS9KQoew7N1uHrNl2TfU+PTebtZmuHik2x0U7oxKepzE0tDBicI
TeXk/saOJ3EgUnrY5PbP2XyrcjcvesBzGViXSKYl6ncXfSa/Vd56ek+s57xhsLQl
itRLCNm8bFOHtrLPgh+hC3IKbdQZpLl197JtpKDzKOlrQaJJgyHTT48B46+xzl39
oF5/5DQeMrlvYm6Qa/FUJq6dizF7ulBi/lOU/WRrSXB6rk1Cry83OFLV/ROcBjId
LFY00q9l+/3W2sQ5ygelD9ZZpshegrE3FT3DanuoHTbQ+hcgegsXJIJABJxCEFuh
3Tiw0OVjhHKiDMmYFqlaclA8GfTYXtnxQIwuadiQCHGlRd1p2sAkG4m/sQ3UDo7E
W8ccENf/PXCTlIrQGLX2bl8Cgc1J93QcCXDv+GOJzBzpAxm1is4ZizCnyDy4/Wmc
+3u95TRO63jiA/NKRIkdAFgJ6WtRGzHgB3iewBYr5vxt+542dcAEbeN1uYx3hImy
RbqBkxrZmYbNTdFAhPwdDZga+483o4kLrvSIAPRD24Bu8nGtS1UNZfRw++Td+1lR
g8AVeOFcVgzsNZrdtpAErfi23jxAr/hcV0YaRF5tRofv+EvbMTdyvRpYy6ES1AvL
yQtuUvx30OSCulBObHoB3zViUvyxmBzMpgB9FGlNKg8ZEX92QgER//LFJ2AGXsFW
cIBodwBh9Z408Ng9Elah+g9rZL5Y/Lt7LPK5U6410cFek1TEhTg7M2ku4YHmA2NR
0Sg1DPAWrimbDJtS9qi8vEaT7QOsfblnVvpyTuRNCjj0RAoOGC9y5QmYw09dLP9O
DXtrOVawJMSkyu/maWPjrLxNrtI+PgiHKWgheYxDCv6KfEzwvtKqoQ/cGni4w+XX
bzoQ0ZlRWTiErxBWnYn4TRLiBQt2u/EFZxG14bI+LcM73QODw2ogQdrJDVZWnsaZ
vX2lL96btzH1FSBqiXG8D/TW+u4veFPDTcppyoKJ0OIx+FLnwpOXkQWfCB71zCAT
Pll6kWNUYgmYRLNOaqH8AK4uTm5HCzPOZ3qdsKfIGV1KKBaiK7TM5z0PA1lrnpMU
xo+4ufhIrIwyictuUrqAeftHV2NEHIB0xtEmTRm/ihzWEWZmnAYOPgfE5iCc91Ps
iTD10GWF6ffZgeGJrdAPWBsbifF8lRSaus0R2xaq89tbxAjk8zke9hj+SrDZz2wJ
osoj7G7bDtwMhn71skgqBzBQhpe+iH/GhrAqobfKxUnLZgLdx9C9Lra+doNxIRHX
+guKQGNJPAjXinDAyFjaFg==
`protect end_protected