`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
ddtXksX2+yylW5zu6QL2Lhnb2d1sD00763mmSITNX595NcHTEkwn0zB1Dry37fOW
FufOhVzEJp80NC5qZ/+F0Vk7Ik02dIR0elf3clrjeJRK85K4e3Hoo4xn7YbFUIms
l/8VZSb14+JVGURjfswrIyCUotIzlzVYZ6gzoZwDXIi5gQIBf/gI+KxNXPaKV+PQ
Ufys/12rjO6aI/pPlqSm0hCvftmBcnezN2hk1UeXgOIuKZnogjOsf0iJVX2aOOWE
6pD/psybjbnsNB6kH5uFTA5frkzIzkzl5d9+YDm9OyC+k84E83I/7/j+rk4L2dah
QJOvksSIzN867/4Qt8qYTQ==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="MvBXkzurAa5VTw+1JJ70nePUfoQXBvZOku/SMmg4TwQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
oRtzZL4VJ4iwysPsC8SXYCzXS8Fw2gtZTOskLcDV+1B9Nzn1zTyNtlo6lNICRmmK
ZRVu2BmCc2G+fmzynYlNTnSa7C0Cuel6FYpxCBlOuk3OF2tzAmLAuDyOH3Z1Yjzk
a0aHuoCdIRKv7BrZCdALt03JeUmXKPdOmIlkVGFl8yw=
`protect rights_digest_method = "sha256"
`protect end_toolblock="Jn9CQpRhJt4rnzZPRk+dOpzAubz7omckX1MrFd4p81o="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 28016 )
`protect data_block
gD6l00tciPUa6pDNTk/+t0OO0nC/UTtBwLB41d4inuAUA3i/ALrNyoJVcBnAmEQW
ptbcNp5fxEUJjnOxnedyZEuEBxWRieZFQnkRdF269oM0/IE7RVXt0pJmXS94VVOH
FrHpXVTJss6n9q5HEXwYnpIDn9IZfQRxms+IeX/2zKEZUe1y5cN+Cg8ADrX0v0Q9
EQIjsaCCaLKm9z32FFAnIiscVCuDB005dJTanKCfsI2zjk5ii6zG4U040LAD6A+d
si6Ce8y6T2o7/nMlHmxTMGKe7oMNKUa4Bti3FvV0Pedot+SSnlWVY760hhN3/gyH
KOHrTo9x/wyv2F+QI9k17PrYETeMaWAozSg12TpzlRlTB+vnscquqYjWZtHUVedB
ZOdG2Jodc7zyhYGbFyOfj3Rn40WwV5a0YEMzYNYkPlM6X2ciR9nd3J3ZipkxBUL+
csBToILmsNsML2yKTm2UKpmOH4sc6/ykIP/xoQL83HCE6CADVKGJISaKj3VwwLkk
LeU8+DPKHMXik47Lnlai6NeW9+kZW2HX6kU1snw3VVKTD4uNY6OpvdO0M+Qn9puG
wu37HGltD3BY+KOIrOC6hGxr9FCyQGazy7/ZflsptFsNZwQpyotOdr2wI7nE5Akh
yoTDaqLTzK3LRkNsha2Z3HBVUK4KfdUlGyl6tPq9KxJNrDgBEcGmvIuFhIHA83J+
NAiM4UPQyUvQF0pLa/dn1dY49FzyBiXphnE5Zgj6pWP6JSTxMmsIgEucg8zeB0sz
1wnZwbNwifJHV9xeZk3NRWbAAVZcnaCE10Q+8aUl2j7Ya0scErmEyPegoaJdQjXo
TTnzUNUI2SCMmZRoiazXtaOPDgYBwq2TBvCePlywK6gm6aUW094OBgfHUFflhOcp
cCxQlA34QSAczHRY4JZRdJ143ZiSD3BgJf5QXEfay8gIAdQpfwYocCucdf4sJDXa
bAF7eKyWEZIIegCsPwfVAPahzOlpBfec4gay6j/M8ylvNRNBkxoOsvpPA3G7x572
aKPIvas0L2EOnEMtVm4vTv1nPmimm4pqt904b/WtAorV/T3S4ZQKo8Tpgmk+UXmd
GRlDrM1fL4vdUUBHMsawgR87W+PwpZOKs5+tfaRiUrgctodVn0kUxAYGWaJ8jbod
smOtWAqXgV6z6R4Pl4eWRD+93EklDHX6mfCzun8s/xX5sl2IhEIpE5z/zuxMBzHE
bGaRyFZyQWsw2aAhz2OCiBxGAXQZ2YmfQ2jYFtFXp3KU8qQtEAuzg5Jcr1DawBQG
IBKDtAmcj0oys8KYXjF3EHBaq9WIOytDgK19xNncvK5jAW/kkJGDGcjaH2RwJhCf
iBp6+X/TD4/gt28rYrsmC5veb61KAPxdfZbzLqrrBCzj3Y3Qzbsc50G3xYrWEryR
pQx+902WILRcYpJxUdZimpB0ncMr4gFDa5kkSP8HYotsaLvpTXPjcQj0PghIDyru
rpTszq9C7rs3l4EI+7XJ6uaVua7lgxwUL0ndPmt0ln5w0nGLVblDwWZAX2w7/cha
uPicW50P0SlPpozf8lXr8Yd/Sg1XfVfZg5vTTM09dFa1kfZREZJPCQ4bu3dfAGSG
u8Jf/s/X+HfMRutiYIR+bEUuNTix37DSZzDWeneV+SaCoLy/dqryeROq8IcOpodc
9dGB8XkZq6uSWVImImDbNZ05cbfVDDybxkpVAPdcYjhV9seO7IkT+M1JLCVJ+eay
el+GA09OLGi37FCxCYMoc1qnWUXXefko1XeKddAlrFXpA37B9wQo3rrjw6ovi5eI
e9qfbPiWVbeClddJrVGYdt9aUGd4lxL93SIweTKrROy+ZCQFxCHcEoMtY4uTkv+A
Q1uVayoem0evgMeEnLFbP0FjWIrp8avT1Avuw8fGPdI9OdWhYTmSlLXXhAXJcUYm
9DU29iixwlbi0Dk1EL2ObIKy9Pg7twxmkiu7MvYtw77DsKOxCZ1b7OZmVhQx41BE
FTRO7rkDnxvSN4zms1sNx0wabJdPyy39EF+jd85p++QtsFdfyPxLycxUUyhiynog
lTtE0vOdCDtCRPB0kH8iZ+e7HIpTHDhWtqxJiyN8RCQWc+Urf1kZe7w0cfmNmiA1
brD7iMv7pj2h13N+Og4LMJzagbi475oU/Sr1lT94FqfEFfJC/27lH3/t4jc6GWGr
ucXpummLebhEL4w3fZBsgtmICbcr/z0WpXKPnPHQzwQt+J1JbTnlg47J4tN2qbHN
4nVaqskgMgQWaIyFPVjAAERG9q1jhn06ogkJ9fXXIeyYl5kJaUIM7tO0eqEItInh
+IBtnZOcxQYaThcbrKSAYAbeCxRTPEQqaQcimUg2TXi2LwKy3pQIQCYOlCxTqLeh
rDgJIXP2VDv/f+M85sbbYPe9jPVIhmi1U7cy4dIb1w10TG6B6mw2iNasSfdvw7oB
z1PWUK05UEWKSG6mX6q1Z2/n0Hjt5RM/e8wfGPIEIiEQrehmwHTevKbjTHKKsqSK
F9PSposMpuOAbIreJH1BcxksmExu0D4BA66elBiEF7Y85sgYWYOp3mj8KzVNSHh3
vkfDjWG+W7PoaPQP/i8U+2YkAGXAKqKwetqwDeBXiv+pba3XPi30DnDNGm5ExkBV
9VWAsNAjxWH8sGRitD+MUZW/XGF+hYlzQU7H3WO+r6dkEmsSyz3FAdmb227R1Wp3
EA+xHrQ9xJmSMRpZpQI5EsfHeJHWKQkztKUvLDqv7MQeyXsKhge+xDvKVOkoiL0n
Y3Isxb4+3Snb0BJzBMZaFkTRe1fwSuAJ1Em4PEXEZbpumNZ4rwuKGWCfx5azByfp
nKlHa7Hl/w5JS7+Xk/Eb+R8o4WMqwFl9ChIY5lGGZVpkbTfO0owRMGtIZTgBuncn
HlVC88LUkv/Rf8qZ23B+T2qdbg6X/E47VyFNRMjtVukAWotaCXw2r0Nur/1HZAV5
RwcE/BIbpZ43Q3WIuQsm1aY4FYZaJGAmFzGeIGdf46bwu1uAaCvUtS8r1ANVc/+i
j5/Ohg2f9KuA8okwrDEiYAh2SR+FlgfN/spuiheMErJ1zaqVHW1NVGpf7bYpaqP1
xQuLJSeK8jKgP2p1NpB8rpUtJcp8d3YBHlGA0WvUA5fQrtwppnznwh4FRvRVD9As
QIoEVuGVIN+KYFjLyZZe9QZTGqAP1yp5Gd0ZJwGQcsbBQTbQMkhje1untkfgXcnn
3k4gaEaZaXl26Ne35eJqIhA5VVRpynvLF4g3mRf4Hva7RKrqs/xYSQ9NXg6epWwt
KiqjOLcVccnloN5da9Qxu4TFubB25d/ohFXb9IHPctYnbS/bh7CWbaqpsancYotI
h+nfEGe4pa+IPluoWAENlZeuzDMyco4pzMK+t/5pZg3/5J5Jn+q1lWtl5JLZCOdT
T9HRY6ps4sjzfbdx9iLL4ZABEqXR2+CT+GUBJrRz/DRMamRh2zgAVzYPP/9Ctx1O
OrPcsSiUybfXIO309KhEE6vM2yXIFgCvyGJBTpKh4f8FrM9m1owlVR2E2xsOEwHs
DGwiUEuHQo+6wKwqG+EcA2fBs7zMFz6vfHhgYTo7z0ZIAMQgIIfnLj8a6G7vLlt2
VgAHxgtTuY/6XDe5DBCrIgWxFpQZ/c/wjUW+im2gaVn9G0+CTlHn7tkBe08vLwkt
kmatLhwtdQtCrdi1cfLCoYDHcba5iMhT24DCs4iyrKMeBZeCS7GDPiROPmt+kiyR
ld3BUdNLKvKijK/G/ruIbmd5Otmp6Ie7awUk92NCBROYuWSYZqXM+R3d8gtUlRrG
/chDDQwt+4kOxm9UrZws9O1/xin0A712StnqlnQynN4KM6uc8kiMQR6nJtv4+Z7i
LTgZ4CL4AioE1vgd0cZXlwG1ygH55fhNr9xVr51v44fBLNSElnJ+fc8PRWF9DzAI
h+Dv28XpfBmMFfyEVbGkVAZugrMlQDq31d9pfd4nVd3XEk2AfvnglA5f7xkgl1XB
ednMc72L4Y7WkjRVa22zg2X9XzmMsMmaB1rL9r8fiXKJlfTZbGWXKdHxt195yQOb
K9E9AGc3lsnlz9QRXFjhZK994xyhei1pu576dNf2QRImXSsUGhrU9d1LblIL8gmT
fF4BrltxvdH+3zq02mtpfNIkV7TJYwZuhHUAOa4CyzG9xMhS45E4QkDumgwFE2uH
1K2ENHs8lhk3f/qusCOwohZte9sPOY3frNQ810BjUe+1buCyccj4tZJOkYToJNT8
RxJ1F4k7sfxCCixVEYJDLTPHwLn4BSiY7GoqHWepBoXCYVMtV8UZYRUdxfUrrba0
C7VwQo/NWQxzauxNjY+4q9So8mJ0bYEEC+HMiCSC88GjzZFVdeWNkb36aS+ff6og
gP+Zh99o3bW1HzaHZRRGW+FxRPx451nszB/CkepthqGJee/AV86Nq/lzT6JwocKP
3ilgsrdmbUXSTZmiAx89CqxGM+g0GiZYQPoYM1DezpnNLc7+fcRPM9Mpqf0dEZwQ
jd/MrabcyLbCjZ2D4vgGQkEAHHxVEglwqMcN/zb0rPgH5JKCfIkquibMB3kSIZFk
8K+p/C/u8IESUzldo5NJLIQoTA32qU1bio4j8WRR0OWAOVYQ+HOxZZbMM30S8AeN
DqFi547xCFjlyhQtk+u6tKMygw/Z0lysvgYC3jNpAVDL2xs+/78vAFC+FG7Q6STB
jD47Zo6Up8wsyUzaioCn7OCpAn2yz9ZkLV6B5jVVQaoa3YDxip45vIV/OAv+qcmd
Ari9dMmOtCJXM935sxIHMWmuPVKBjadyyrMd3/Kg5cOuViQIogyQoljv8QuZgOAz
gzQdr7H487cewdtRePIFC4pHcXoQLIx9XUqasF0jWqG9V1CesPKvXt2p17l7fCTK
LPWuu4MycKXq2TgK2a5f1Eu9STlbbboYGSgaobtt2LF+0xQvSXYaaC0nOKReZr3K
3m7upzpl+yhNiByY0lV8X5cQlIRo+UxVr/e7NJEyWsW1RkNC3/BXrd91mTrfmN4d
bOS309bQXA2HpfMXW+pKu6tod7ins7+VKRmETUXYkLu5Qq18jkPcfadXc+oATCpq
GAxOJQOS9znenYJhaEq89vD9E7bpiCdaNWCPhtmZjuFpwgzXNBYIKJ8tTn6FhsLy
y2cRVz6/7JWV5Ea7AEZPeuq0rgQUXFWgmJaR9YxOcDutTsxjtyegbtBzLiTcP6Ui
BOgLePV5qN1kbpwvR1Aarb0HXJSc8SwS8jyh+WLnnYipZhVMHmPP3jWJa9O4uHSd
HQ+jimobwHDsIcBlcfZfj8YF24pGAFLSB9h3vsv9lzjsFq5iizgqdsXK+N2qVItI
fLnUezknU36qkJGMBt14d13vTE9NJnObBe1KjWNN2CoY+dFwS1hxkdV1aASppva4
dJ602xXrSN2QmMkfgvJpYMiKJEEvRQhOPIR06fpNPaOSAkK1MMfF3SVMOpa0MHIG
h2VxRyBHHRCkFbVA3OlDFzy28gnSXKnqxUT0kbyxy0+CIU/jQYFgtM1I5SVhs4wc
EmJhbgIpG8fNVo20ct45eYOVwZeIxgpYYW/LTdsz7CQBKoMpSDIgbF6YNxlUWJVN
hJxRU7ImFrvFAfPWLGXCEyPkbZpGYpnqo4nBbqZrMZJ8dmih9xoFXjZ+sXscFAaj
/qi6A2RD0AapXGLSBazb9qw4ucnFCIv3lVNEoon2V3itBQX2p2sCP5dkEXTvfsKU
GhFMJDkn6/R4HnstGw4dBo/PgDUr7xYFmiJqKy5D8R1WItJUdTQyoC0jNlqmT8Dm
XB6dGyRoJb7QKop64kVR1xQzMrmOZ8NkHVf9THRcQl8eKzcyNIuqKBBJcqbur48Y
r1ZVmRNni14Al7Yi5pavRgkzEMNrX5ZIfOgI9dtBc/Rblwk9kj9NeUQua5/hmNrh
tm2/EOUeU6ICzWs8f/lcZS7D571/SyUtu9DqG54xB4xQiaZriyuLSWp9O6GXSSqm
pTDvdLdAjCrgSO+IPo3cBHAyAHSjr13/56Q+02vCIFihYQYEk9CaJHrYbTYqez5Y
iAi9xvPNJbz10Ko5fjL7ECblYXiyDG1FKkVDhWFoJVCbGOEAsLvOYNLzXEyAbpD5
Z4yQnHszLKP8+YtKZfm+FtTqe7dfPeLaQJh9OLTjojWgfMLtta0HUXSAujdPxewD
JrTGkoKKqIMMoeDgl81ywfve99KHh5mUJkpWCy2/AHQBY4L9WoWze+BpIUer44Du
Wnrc8ULdn/ltlSobU/s4Jfc1HdGMoY34No/qcPe22LHq0vTVbkhXN+O0E2nqj7J9
7Okk2qFCppQBCHvoDWZXRkhfEl/+jxmcb+6TWFI+v+QrIFunWPkQhAp3c8GPQQA3
DFa+lZXJGl6GB51bhIqJPFwkzQsyynzBDwTunUCb4MpUagy1gwDUhUr3md/1Azgo
ltLwsTHDxn2SoPxDFwae+3PyENcjWlqqpN6Mc7EFJVWAjcV3muB0EzHcu5SWbVfY
z+n9ukrII9PiMbOVZsWJ/YCvhocWxhuXYeyuStC7BujewQNqYYd99i0hicih9wvS
ZKspJDYBpZcBjJ1o2R3pRaLmiVEolL4SFtOhepHakaAMGqqRC0iWyAf0hYZS5Ok2
c+HslvosHF6ALUmHMhxSMr9FbqZ1lWe7oHHGXOI6tXvyNkpGa8AtuCxvBSBQNXqD
69viWBp//Cl5+p3IllBOB5HHJw+QLgA1Hq2AoaL0cMFmyeKPEcJIRvy9Cvj1fZ0u
NRC0j1Qq3DjsanEGCqXXdE5PJddS6aio7RyRV1FBMPi9kCvpCtuJ6L+8gUEvrouw
mbDU3jbtB10ssIHPf3pEgQLH2x/zydchOY8rFO0reInH9ZoUkcGOsO/MHRQyC0IW
FO9aTaEWvAoluSFdaDl/lGrBSRRAjScDaY8ncT4HYQxagUtEe54KY2vst7gKXNx/
ogCUMwe2qgKa6piDp5z5YiouEXaCn4FWZhNQLVT+mTAXIwtyWWBXD2kIVeRWwVJv
CZMvezk2OvPpxLRGkXMKE722HJ0z4tcNwFp/w7f5dHMx0y24ELHmekzB0efbE2Q2
M3RUDpXIfnZpeLIWGB4O45XUZnUAijGpA0u+peMP5DMkA/FuxEgTE8Zc195Hu9/Y
K7JRizEIUvdCTTsLZX5Ml2gJvwmE/HQQLQz8EC5C3tVoWHBwTgQS1Pho3DkuLW5C
AW1uzPKWYkET7aN0BslZDUjxbW/sbIYZ9Wi+Ox8KJTn1zouPN6EskU3zzuOdSHbX
Z+gYGzJHR3YIqiuzr+2/ZlZXL73Knk3hN9+DXcjdVDwlAFWvZCss4GqqOCzsRiOi
GWhqp3u8shd7WshApEyasLk2jWXtGLgLzdWbmIKlOCVPVn6snAAQK4oYvQXDHpAn
T+1AcP+/Op8wN0M0OrVdI9J/UU4ZCuPN/2BiEtHOq7vu7dTXIJBqNoalMx39uQ3B
wS0n8qIWAHpnak5QbfJxZH+4CIaPrkqUFzgtjkh/2L3I1XDpqS19nFU0h4G+YG3s
xWV5cQQe5u//Buarnm5JoWmXYldAzhZ7vx1pP0rhUVwHxzDI+pAiSsH8gozkIE8w
vYadW4iuEcSa9+MT38YkPrXP6ZFi7hcrjEDhq5oaAbQMKWb2oPsR/FLai+WTT5t+
YYT0AhKjO5egjCL0ZFZ7/D55CETYef3u0kGeNTanR3/0cAEnP3hUZ+2XPU8PKQnI
D+G3W0yjhl84ZC6Eb6Ub/tUZ+1JfvWrllju1xCJr4g+tDjjP7Htzp0iAnN0oCIAa
39qIl08GrBINBgKnP7KrpK0jIazRv9VHICoUYKv9qnVQUj9z5rUH4OpUSHDkTwX+
NMUb5lRLBR7eG9xYpXg5UAovDJLXzvAIZ1cx/iAsmXRD3OdDuDACFjvwJYO/PVJB
b0vc10e2mzxRsAiyT50luQGteU7mqkhlX+hOBShruVH/Ix+hYHVJRzdIsP7afrZx
1Fn3bOaI0Lk1jj+IIQt6hO+9Uu3GieEsjp9HJmKAANgjmXZuMPEQVsM2/PV2Yw9Q
j8Qe9+TORMMFZ+Oyu39f8vWhHEHp7MBktTCwn9Fl9GUUfrPRuk2BzWgRXe2XdkEB
dqDXndD9h9Tdm/KDMn0n0AOsGFSIWInmBQkBMPlCTcpFFhlxhFuipawI7bX8i3qm
jF8zfgDtxVEKlYcieLCkjOKVwMhuqB87nT0KP/nT4rfcz9/YgC6LeT8UQTgdorHd
vrGfiBZyTYskiTZTef5BazsucruActGxGcgLgQe/86v2SCOdMFXFakJNPs8MdPfw
dbPMHM9SKUDNEqWhXqYlKNBG8GY3AufUw7Gp3kqFIFMkIYQkDi1x8+Glrc/btKyt
bAMUepwh5OzeydcgAuZ5lyonQdmXV3X7bSqRXx+G06Bk3YT63Uh6lyFMbHbM0Ai5
Q7kUCmWHjcpQ1cXMrMT8+HASMPOuAAprtwywD4qYty9OkRn9HBE9X3tOkfEA+a46
vjHXvujHGMaqeqoqFzOxCx+/tVlXanXVJLpjvJOZtvs7X6Qfx7qnh2ki7fCuvRBP
L3qhT+vzD5s72H4M9ge95TJ72MFbXJBHE+HI2R7yLDGe/tzD445V0BUEBKVMV4K3
4WuxcjfvGDZVHVT9gHgYH4r5zZl76kb+fhPhth/g50iBK9jMKpWN7nqPMRC5RUab
XObUsgRHzN41hmRJOtsDU2qy9oixD39P17bIWl6yHL6uiqrkphdCdrY9rMHfb5E7
ohB51OGGQrkDf/IO85qMQFL541IgzcqLhgWftc+Eqm5MdFhe9IuO4cP4UU62khI4
zMyUyaSLJZvDZ2l2C9JTXxSSFuBMhY9hExpM1yqSiSLPJiKxB6mBGWFXi7SyPCgw
GzNugxjeIHESKExjXCUcW4fpFgXVcfG41Pr78YpHJ9gGsL4csels23z5VPxijxJz
0RLGFRFk/5dNX8es8GjY5DtUF5tlkYxghSudje6Xklmk0XZORv8Bj+Vo5MOdvYAs
L8EteRE86t5gdzOti8MktQFl7v0dzw5j5Nd6DsyTqB/j0kOQXySDN6U0jlF+8J8U
CWcdVDZeI3hOl4re2p/FgAREYbKkIsiz9+nMuwP/SGWu6vLBiOCaR0B2fU1DKVVO
QWp9zhjXBHGyaLk4022vhw2HSlqRlKGNk+fAaTBMNZDPpscPGpufzmu4bKakvblp
BpDi/jkmoL7T6I6Hxmr387E9Y+qOjum+TRUKF1uBhVME8PQf6cw2dEbUr1mp8SWP
/trcNBLKpavJ8L/zwEjZ1EHGGH+9k6AGTrxqfnz5M1p+DoYhdy+PcDeUHVqI9UfU
ivcxZO9pxXgzZiqk6lv4xI5OTsbxiyCnES/7dgUzpN8kxftHP4HQbF7AMjvGb/Og
tW8Z7miAqAUokpaPRHt0GHsTzbOEoRxTqHqI0bg7BhmnkYt3kAXNK47qdXaNTD2E
4ugPXo+rcaYAAANjwyStymF7X8meeItH2XtHt4IOUTEbRpDO6vQ1HzHRo4z7qVAL
pgrMKQKc+IVTvZgaLFvwT48cWUIkixV/IU6JAf2v0clb16FshRGcFwjJo2x6hElS
dne36QTf4pY+7oIa62BL5fRJAWAkDM5981qF69oaFZrs94EstnX7NA87sOk7a/Lk
DsZiURzMK3H6zaOsVjxUrWUJ4V+sbZg6t4VotgsmraBzdyk2FEInwT4SJfHNiEF+
ooP94LVETA+LbLCCMpYIBJVALF4fNF7wFjtJVd+wpp6c2ieQbRa2Ssbpm/mpKVNl
FB3LOC4kJfDDcHYCOxpfWMIXopUjES61jLYZxztdsvQ9IOIGed+u0CepaaLWOz1G
M5CmFGDAmSekN3IqqjFeJBYiPluar2HWc5zAAc4pLkBxZE9zDUr5Ouc6sePw/skt
qzjX4WdRWNf/GFJ2tIGTOzOSWlskycti0zUCwLhOOZjHRI2PfY+p5wy83QLyCBXV
mE+3fRzCzehxdXTUPiaCZczRIP4yCv7JoHb82wREsKEWOQ81J+I7vuRVlwzzOL0w
atOzvcEXAudiqgiSKwYDaPoh3Lu/sLyC/loY7m8GpbddCfpsUhMlxjcALTXucWV/
ViQjFQdSJDOjAgCBHRiQHFoctZwrZCpdKkH9oSsOkXPak4n2ZJ0aHKW4ODd+ZNuD
HWFjZNnuVxwnMxs4/IexqKqK3Lqfr1M3AUu3mOeAihXrgIiCu302KXs+P3Piggyu
2P5ZCIWi1KXFR/tTQ7hWGnX1NxQiKYOJ3WZUSuQpNyREGYFkiEBclGxevR/KXeem
aJMFF/tWzWHLeI3Vfb7YK/9seeTppePfshDii9ogdpM19YH+Acm9L6CuNiye2tPb
ysN3DwqbXj1EOoHWqb3ukLq7mQ/G59VNSPI+PMj2HN2c/nFdBlNIs2OkRG1K6fjQ
FPn9A//M9wooWTh/d8TLxcF9166dHqfegKZfgIKCgW4f1pKc2MeYr0oyr5CywqrB
x6l5OMhxDAueHDZiOHb6KAp5QI2p8PZT5x4QemnfrNRI0QCyt+QjDbJxJ7+pEUx3
hrW06j+3ZZn2vYdk1KuqNoQKYwG/ECABwbJ6Ws4/88do4mTpa5ENyL9iH+dRHvBZ
mpzifdosZb9Z/yIRPyxwEAQDQCLbwO04sHhUZZH62AhgSj36VtWB7znWkE0HkriE
btwoWFRjsiCfWJtFokzusGbjGfeBDvasz7JQK5lEiNbWQM7cTp+VJwYVvmvP7t2K
7C/LxREV9Tf/8fc4BoGhObDvxAreiUc6LCj1QRZCDTMbkA3mF0ZsfLSbhOuB7wgd
uMMMPuew72lU6mDav9aVDHEgRVxlbSjWwpUREH0PsgndR45wPVe1DwiA4zvovDNp
XR5CBjyDj3Qynhfw9qYD4N8UFj7rNTxrLUjIo00HM9d5uPAm7bVW4qAENRIOPuR4
lv+ifyBVJ6zKJkd39OKFDxZppT42CTjPM62OocONoGPNEjvHXibdQMse6O6P6qIC
VZNUJ3m1YAdk4A1fm3TYISDnKKk7EfIukYS1pOWrB995XuozqfthIFM2kHPTZ/j3
EL80hCSF43b8fmtZ3SIOC0Ksqya8Pb0J7FB061g8mlFNxqFTyYFO8f7IilJpYOG0
vr0X561GsYlRdsWwqFgVu2TgBAJdRMhRJ5dY8pIwiq3w+JpHXN/tG7laf7vapDsk
wkthVKmbvooxC+HBpXtFMQpfHpZwkkuWW377bxNVT9YgJlSh5BeELRiowzUlmtZN
QFUEtEP6U4CviV9JCTG6d2/RkbaRSWdawVCYBM0uveYrhaKSme5MuGLDrHJiFriW
1LQc14FNjop/1kTjSFW0TgXx1bmpT0Q+urV/OJawU3QvRJorntgBHnqWReBYp911
uPhoBDh4is2nav3+tC75Q4Sr/eAd1ZRewFVFcj2cxyMSVblr8VnxdG6Hh0QtMjl6
Z43cim9HJovF78kSE5dd/m/aR+5C2B5pFI6gTtwhh0w9qwzkSrvGtFlKm2z9e4vH
1p9vnbPr/HUiiDwMp0VrT1l4snVw6hJlJBscUFSmjoyrxR/1u+vwfNPq1b59yoV6
PpknKlQ247VdV2TCIpF/ebM1l3wIW2HMDNWdjPHcNgZvtmossNC6q6NrM7KLqJaz
7lau/4/h/rtDEP5uPfrYq0E74NQQCEkCwS0W5bBdu4ca3pYIQrPaWA+TubwC+IXU
SJ96B5Mgh2Ru3B4CyqwTJRsZYKz0cNFBW2D3VWOPuLLQnCbp2oZGWX8a2rxpBhRu
7dRCbd3ONTvmrIxl6Qjrmp0c/VgNZj3Ed4zuOQYJndcIdP44ultgU1rTSIxmYOHR
ceY/8OBxv8DPRvh3sab+VgQAuAY4+FXXKtBEJzNV1h3zG6q7xjJjnd13uDH8cq8O
aw00dPJTu1DRtzfo80IWqjrt5WR1AGMlLIEb2wgyQH0U/UZDG+f2ZYes92DbiOYj
Q51GM/aodjxvkqNIsMn9wzbKrQUq7smbjAj4mnx5NN6BBYa7HFHgDzYbLy9iyFR3
vTPTXPxxNy0A/QkCHO0CKqHpOZRkQ3DRmGYY8GicQ0zXC0jRRs1BnavwiotV1lh4
rT8ouVQVQdXvkXIwQyogvtJGUFBQGhDloJek0yPgPur/Gs7/4xuCFofNw3/zJnUX
O6sMtEW7bbdKbGOmX/nvUfsZRPxFdF4T7FatZRiUvsLHcLupCeyY7ey31EFfJwJH
qR6bojcvEAe0BYoLXB6ll1WCYta4tSzGijp0MjyB7nHhD+S+AvbrKyKjfyrYryw6
m/zB43SeOCSCfOK7aWWKQu6WG/lHpxalMRjz3m/iMxEQpcNFUXdF1bdazvvnVt2k
cBOZXCBPONBTLnXBsGgfJ6sYz1YWb1q4tf3ABKzvdJUkHJelHCGe1ojlrnPgP5pC
ORVL4z23rfOMThcrlwyc6TBs/sePYQyEKE3VH5traZJAGYie/xy3ggIF/NI0BSMo
ERscMthVDYqO7jQgVZw2ZqZIfaJrj2pjO7D/SxvNr04Y3c3xYMBuYnBMSF8H7JIr
hsUMO6jX+OlE7qdoZZ+doxb6mtI2rAcOfvFvSuze3EhX/DPTReWGRwSVr6c05gcf
g0XEqyo8TKSnyDOW3Y6aFFZNo/zE40GZ3JzYoTLmr9SkWoVdi60Q9kIwuB5UNxjE
QOI09PM4ByEUUoAz65aTmmosm0NTNwE0e2UJUCNE9H8ZhNOjbVegWgJtkWyv383g
yC39TN5wXi6LVdTU4HChSUtQ2Be7ov1j2qESeXZ4gXLjZJp4aC8CsO0TpB5CP7mG
UXykHfMs8FCO2O5B7R87nLaCnRrvD3cvw79Bha9mHMz01LJuwjc148sh6s6gFhXX
AklNqVl43+9V0SHGxRHwtcKTrszoseGVYjTKXaR8dzDz7ei/qqmm/aYQgyV5KyRz
TIh93ZG9pggfrNJ+y8bxLDZ38/31NF78NtyQbMsSVH6yq5jiqqsIU4a14Ufwnvm5
gcEvbxKSvc7BVz7H0DbqnyNopRL9D9eeBh4JmubGG/5p4xiWm03GNlZ2yFo56nrz
qOBV7pjN5BqITeBRukTiGLynxocfuy6JiG9frRaBn681Vwj27NbTzYWUJ5MF2MmC
ucish70uI3aMs2+LO2P0nAVrACqmN2DBrAhOKCYEBbSNS5lnH9xckWI+eDnN6U3Y
uIibFgzHIzfJsoNbqwK2wovp/xLamESDKtWcn5rcQ5IPKYECAZ5qqALo+DtngJHd
Ndb2iAyN2AKGFXXAjmrLHZjSIiy1xzbSV0EE70ItU9DBNhngl3PiDNVoQlxReNRK
i3tHK6E9KvYmyhiy1Kmy/8Q9vVjacMfH3ekGkbn5tbyybFSeRnVQj9uXaWNDqAVF
4Se44artRJXOauK6vFTDR5CtVUaIn1NF74o4vSEpT3q52PA2MMA3n4Xt8Krf4YVI
T1ReeGzDyx2Efo2WrPxmXeQuHIuzPB0mzdk8/PwFtsjjkDmTgpMloMiv3TDfGm9H
/tUiH/0Ws6r/dddyJvRDFSV/RaSJ+eb+06ZXVIDj3g0E39wIdzJP6hJrjrMZFz6q
OB8ONwXORKbrkr1oL98if679Rsp6jXM1FHqsJLLxtxc/DPdex61a0hvHv9OKBshM
ss2LLrVftEvtHAQ1jfjneHzSkcvgouwM68Mn/LvkGlXOnJ9ERfoQU4PSrEap6xFL
B4mfr0OpJO77frp3edvyBQI5SR5iO1anhA94vg2p+xNL1pbQo7m8eS3SoOTtLY2M
nc+H+5xnK4a6VWIBsuXBv6TlVzaTh8QKTqUERu4iBzPIsxD+4qnZBnvUqq8jix3u
j3xs7PWj9mIfJQ/w8G1bW9KwaAEV25vPhFcrk0krUg70uWznwRn3cQHynJANZJKJ
SpbHwdWDPyKq6KKRZ/6uCsJv9fluslB0cefMT7bjMt0EP8M4aptE0wEUEtjQGLhx
HBdc+HEffYFrK+EJdOkvBusV67XfhVqxIfgMHy4pNzU34OEDmfti8XmyXPtuZRvN
tm3Wm43oYRIyZTcH1AmuHj/gx3HzThyJEC2rQR3UUrjfJ0ox8SNbhhqI6iXL9ShV
bRoxzFr+ojLsV3FxNqnt93IOphNb6042lLa6eey8DwauvE3/UNxN0T27xuAlWTfH
6meVNN636bXJA1VW7IuO5/qG+6d3+YyqgYrllxaqlMjAdqwaS84030Xsjz/dH6VI
pkTvG2O9xcAGCXJzl2H1Q8xj3IXVSNYXNGDV6rSM/YIXjPOeA3juzNmve1xB/a7O
8xi+Uotrf+v9SC88NapGC8TZLvY7kKQ7GUsx+55kOMBD9VxUM1xeUzOkmd1CTx13
zo8wPcCJJxpy1YQr3HB8oKz5YthSXBOpsh2sbCjOLdXB3fOaN2PE5XNxPJmrM8bK
Shk2gfay7UUsdBrUsZG+cij4Yed6sJ412C/XnbcgPzH4/guzCiMfNzyI5N527g7J
o1kaVLer7QJJFI/Q82m61pjLvywFvp0316kwxhPklAN+wOb4HFdcLv9p0JEn2qgX
K4K9nd0ot0jp4rFPNlrsPPyybG+bwUkLanSDfriUV8prJNqSJLpHbSZnre/iNlCc
gns+K90KbByK+G0X1LjzFlcQeJvpngJLEADnYufp6FqqqwnWcuScfZnl/+HrhIqF
JAWs91ikT5pegZg7jK9UurQX+wN/xRW7vN+eYOWNizJH0fp6vsSq/QFj0JBhdYVz
xaiDKQqkmDsAFXq7w6EWnfLlz0RwjhDoS++undMSmBxA+IEGBGflFxeVoJDR91ep
bYiYm9FoQhGsxX7OYiTeD1GRXwzSUTUehAwnYs2gm3pklmQrRuN5KR49cXMcLHnu
hyZBnDWQ0URZp15zJ+hyMSRl7wveyz5l9s+ptJo2KS5lhAdwZwcLToDtfOr+l3PV
WTUhcOmiz17PhjzBdPoPCujXhLPa5/4g3fAmMh3d+SMuhi4EQ5cEItJ+VKFqnrpz
sNAgvDgH9Y7MFEoLmbDco9vQ/a5S8n8ZITlp25U+Da4bm1VN/xe4fhzZ8SiUdNaU
4XGs0yF5F3rOqg+ECcsph0mo62EcJ6I4i1f5qeKk/8dtryFRDiZQqk1L+linyfSx
3Mnn14BohilLCEHkmsPW6W0J0LXabJkNPg9w2njNXq4z2FOd+vDojGGMwff86CUe
9mYYJDFlnLjPYdizgdav4WaMmP6LLF66KUUJI/dwtbU4qj7CxmNMS/NV8OJ6nxxB
T1a6AE0uKDWDabplmwRz+3zZtuu14+JJZzVvm09ldWiffRRAty4SH5gSdZP1cU8W
aY5hubB9BfSqMX61YvrjmgiIg2GjUGPOFOG/rXKKwIZDsSw1fsBAeBcuWKnY91gG
VksbzLAC7pxSsUtHwG5G5cT3MwkjX894R1BkthCJ8pSPmKdAASU43J78Wp0/D7DA
Wigfk9Fgx3rftE+Og2VWm2q7Ke9U2hLcWRg+dguyRQVXFXNA+O/MJY7RsvYVxLbj
iKNsb64kyH6SABcRbx2+vVnLmo07pIvkOjuDOP/HrKFLzncY2saQAwanaELyTZlg
kZ2c20P+Mi5fbrU/KKv5yGtNzOsEdUxaqZRqzCPI7Ih5CNh92m8PpanlfU9Bb6v+
FK5NQIvb68499JJ9EN2qADtYdTi5c8YxpCkvpNhJz4SLCLxE5ei22PxSYKxaQcpI
W0DxvMlksY4gBqgE8ux6FNKLEJIZYxUD+ey7LwyMtGcJxaB0CMcJI7Lh3z0j25Qs
CZVMz+N06zSfbnNpGxq8j+jISa+aOm92QGWebqHrKgubZtJSQmNl8dCuM0oqRlo1
r5+xwCiD4JbJWP5+Ie65FBS8Qjc9K9LjU8HGmH4vtg54pUNcHgPzrnv/IrKhX1Wu
xYo6fiSftfIknLuXSUnqpfES1Cya03pZCZb4Q4DoSOeLnVZS175l89blL5HCqoUv
u6oELWc9gh9C1KQtPh+LOCBclKBa5ltA3dr//DZe/8+Mk04BJ0Gk06By3aJrWd+O
IJ8CdGB34pIE79JGalkBYUFZNisqKkgGC/sU1GnOv/yCR0jQmrlZuU8z2/FK100R
pvh6L3q1e7h/q1/Iuyjj4IJ32tkSt9JMW1GAkXBtnrwgyIJ35Kq8nAaFJTjXTTdo
KmTNXkw8fywwzjAfmrUav0eRWjalm+t/hfKwf1Tsx7xFD6xDHLmV+3/ucRD8KRvu
SNYFUcdylDyJpSzoqYybBx7Mrof6GVqxnNR3buOnag57dmt3o3UHh2YtYCMZdEIj
+ZLCr4wApYd0I06udGX7Oumpio/Z9JYqmhcpgcyUxYFOX/kZBf/eKvZ/UzQ141NA
7ofbkxdSGIp8v3xwLm1OSc6h88Al326Bt29AjccVt82o79L8/Zvau9kumAAl3r0h
b45Mz7yMGcek1/kY/mphqkIlDIDmb8fXWnBb8T4hlfvNw3AAtyRmsv5pNdk/eQva
SdXKyhluXfifpyeoDT6PGqGoXINnxm+enzEJ4t3Hr929fgYOqlng/FegIEnKF06Z
ORm3mXqp7CwbcHv8vVCcW1oWPmTn4SztfUYQnZKLxu0niJNjMCi8ByUXAZCiNE5h
3Uw3P8IFp/Ncf8/blWShCPddHQBAp+RrMVMzumdlRi9D4bKI9g9kUnDLMwhB6xDf
8VpICv5TNA8zgxv0obrvjsLwE/KxD8p5DKBt1El1WSXxBq+GvxjUq/r/YRwjJYUw
ZBvfJXzFvdu5tAOqxojDSkTeitu1bN34GogzrLnBM935TEqxpTb5D4EXxTVoug40
FjAKedcUXTmyVhuhcjSKmGLTmpS+75PL9ACMkKbHK6HDfyI2AMiw87pS8BxNTHJS
kCdgBJ6QUAflMi+OBHU/MGV0xNT4r6XfaM0e1+2LqiX2A+GkTdHkVEiaj/p5VNKp
GmqYy2HSQQ5Q1s7seAqiHBZrWE5JgPE3Zcso3YRmVn6YT2oDZgexzIUIQnBhSlo9
7qeT7YGV3fK5uPmLOy4a1/ztkarKR3GBsCo0QgKPFvDMsSOX/8Ucldtt+ipizG6o
sw9QXko470916/KHOg1os0vU/jtpVVrESJykOUkscR/+9cyRjSAjaW9znsk4vFID
3WESVZfw0D1TAxXoS/5tx6p5Yr4HxkA2ONU4VbMrowxaLxX2vlzGjdkitpHycjOp
4Fclas66s71GlE2wGd7f9N6n1ZZvXe5ymkeTba/EzNq0iVAqQaZvLT2wYR6CYXmc
4d8I8rfB43VWx6Mc14NLJTBNt6AVVu/p+4+uqTKTWGBcOViMaqkiBwj8CO45asmS
AIqdX3JfHgdfZLVkK9Qq572u7EGNBBMMp6Z0pW74bw0ygN7HlONtIBl0OaKpkp7y
Df1QX+rgHEKmq4GujRQts3UwKZg8dpHMQHdyz38cUptpWVuGlSfXhNKfvtRMtr9w
GLUYwIM+lKzwdeRvYCXoPYR0Wl3t0MYkWSfU1cV5r2aT67YBMQCCJ5BaD+OxY1Id
q+5LmG5K3RGZ+pHV039UI8+f9JUxKkdZVbD3A+RrGy7b5lIpxpaOfJfVPYP+MUL/
xgBaNafITdeKjqHvVRcGGuRYYvzmOl8K4ilCnyiDsgnItguMZVROMHzETqNv2j3Y
ScUCU3BvSghWrqi83ppAzhBvyoiQMjhr4eGfOA75qjsgUWmW1wm8DqXMJfU4EBWp
/MjgedaEyV3QEKKPT5oMj/uwsBMpWDCy1faS9rbUd8TQzv7kM4F6C58rpUOupu0C
W57o76SPsRv/BY9xZPmqMpp2hue8PeRH3tvpVojlZxl2N0sMt9T/xqIL86J3i11d
kfenLB3iGSYhloQ1POM+G0x84YkjhxBYW6WKr53X+lSsUr+xEb8k0rhB1zzmk2GX
tADHVAjvrr2d6U3QBKPwfUAnoxttJqtXdwY+5Dd0F2yVK+h8C5Jmydn6MMNfubK4
4Y7prv1nR2gKMgax0qv2kTo3ZxbHKYH4uZ0oqhUO8xYXdKUTdL80oactAWDnV0h7
YyCV9CtWdYP2CPAQCmc48yY6RCSOvTajFV3pz0sd0MxRZ56KafiB8JsISUniWocQ
m6hVYEl2Vt+H/upC/KXzKun3qbpsRWSNl8ZpPERh/yzuCyqmYXssfsNGUrgq5CDQ
3uaa89TbU+8rXw02DCECB38G39snwLbyHAaAN+kf08I0MKVW8WG8dm4YBtaP6r7m
0g/fC2cOpLpLR1TZqSUx4AbWWtMgj2ukGAS+YH/qki8Gycsr5/Vl/l7B7k/uZHFq
vidPZCSvWfmlRJ8bHo1FOmriB0GPwZTySj+JnvX6tHSNQxKp67Yf2+aeVklMhP2u
iWGqYJVBegMikgBqposi6isJof/3SoSaRh77SMzIAGl9MAGRwEZh1MuVvkUBaWfB
CL+qPtrwiXGD5ATWVLm+I7AAsy2Sni1WoylyKXZcCfT7aFvOO+/czaD50HalyokB
fe/nbaQtT/nbpCzNVkrB5317V/IS4opT7j2hxG3MFFeB3iPm+CF6GrPXxUPd8AEz
/roImZl2aOCLKkS1je5S6Z6oy8tooWXx9nxOPhKJ4gFIOhHOQcGTzYsRNxCNboLw
qnTo9K3F4xdUhSaW+Wfy8LkB6o7JETlfzHOP4Ghils9uyEUGR9iABbXL+HK0IoHL
IhrHhgXu+btjbCa7YhwxYZ5doFRfLjTSQNNo3mUFL+ucF6CwugtLWdG7yOLCpAXS
GfuISNCrGXxtuwJHNB9C8srJMHxDp1iyBJ3BHJ4zoKcQca++oR3AcxpupMkO8SSD
BsK9T/4ezhw+R8TvHZgCsOU6jvCgz3xrmqDDXEELL3S99SzYoWffzH8EwFIAHPcb
pjkETY1TpLA7QKyOcKuvo+sIHnq3tHYmLdPJYz47h+6xxDDB/PcTHpyr3WfFGPQy
dJOeRiFKlGdXNGDF7KuHGKTYVjZZROreCnDkMPpI3wnAvJawGZF0y+1bI9qZVNJ5
varXj8LCEbgMw0S/FBW0QN3sZsUhUsAUfNacNjnUNkiUrgwUqfXrxyuk8UPlWuk/
2qBhXHFOE0+UaXIZ25jfRqJP32+ccxafNuDtqbWKwl/bC/3u3ERhp37hoDehui0n
G+zfqyf2DA90nBISlaGTNKtpjHtrBt2marvqsZ8rWqlbauwXBVyQUaK++5SXLcO+
grXYDuVEvk5cgFV0dQ5l8C85ZBLnLtHFBVF9P7phUiV1yX5o52BBVc4ZNsMZFJMx
21b09K6/y8OZHtH6lOml0krnKnC48092LbFTivjNIZ39c0ATodfLYq5CSZtPg+Nr
a32BC5PrSOhYIWLBtsLOb6wMqy5Pq45VKH0geGDmu48jae0vBkHxmJ0HmgMcXWf4
UVNYGy0cSueQpmpeI0kZMvquvtS3/1nEJZF/4mmF0R6P4QSFtffINMUhcV2gkE5p
5lIGbAZ10MkbKddXv2SjfUHoQhnrmlRKtP6wg59PIaTIm8ejdwIiUgKfysjvNs+v
8m3b6p6QQephwNDW7M8bn/6VLEkDCgWzCLvraHRL9UudrduDV7fsXBycAemDB7Ta
1kZYfkisM0IsjI7MdQIq+C5bZxqr+Al1O17spmigLVynHGYPwJ5cuVvNJshfOhb6
1H6zwAFHZ9jtfKhc816WwxuD9Fok2uld0IksJoKA78a8Vk5TIu3jm7emNcyPEyi/
LfEO4+WxAfBrHhagHGHPQElK3WJLkjmo0vue73p9pN80vOuzvvsLy3H4pNDEKnNp
gw2wHr3Ej/h+P/jR2ZVv+xi9ZaP7DXc2LZwVPdmXddnP1YVt57A4Kes+4+mEGTgM
zP8hA37YUwx6FYX81nFCHJVeowMe5o5mBR8VF1qC57jWYH6AWVl+aQ5QkDZZMaa5
bQK5cmwhINlmEfquCMC67cRJAQNxkiGYSx1VaSDh6CDmiqo7m5fjCav2i2n5xmXY
2dNqO0PIlfvARPg4e6V5L6WGhe4WTvqcYc/knokSqgTE7GWOCGnQelKcZwWrj1gP
cyUaorYIxuIT3DAP4Nx1uUKSJuHoAR0fG0Ith1O6l3n4/EH+B8MNhIGMzSCQMduL
4KDdwIMcODkHkwN54wDG5z3xg0XRJ9ZViT0vG02xsO/wLA9vRvYS2knLcxhJY0k6
zNjwfUOKOPVBwzLschCaqLyeTNpDkeNjtY7mN88d1t6LkN6dtNAHg3nIBi0EbCNK
Sr7rLqAJ8U7a4EPKp8vMn92NpbhqwOvQk+WTOscZuxwYkeKPGmElr0U5oFV5+HRu
p9QBHt/+f9ngQ0VaZ4JWeXAEzWa/x/5NCAbSAOUj0fsnpsY71QdpjjYWXuL25cHZ
p7/GKYrbDDiwhAu/NRjwXgrBjqI2AOuuX03UQN1I5UAZPaK8e1h7hXsxfPZCl9mN
R71mo2SD+pw5Flla4nteNxgZUZHA0aY8/Uj3Y3WoPVWhlEBobkmANP+/YVw7XEfX
PsfuXV2lY2ulMJJ7Z2XxLBO0ROSFwzVM6HEXJOv8gr34JZZxiudyWbIyQYLjLcqa
6BBfe9RQ3kyRJiIqcH56CrNgKPqKFpkUqRQswkBUrsJ2oWyyuydka8hTbp+oUErI
jsiYmysXenVICSv8NC32r/wxmmuL37aj/IyuVsVB/GhbzlCOdkIJuOlu3n1tl7Fh
RVq4R3Sl4r+1t2CrthdyAooDFZlwSluL7CeBILtT0jDxkSaZc4kA4TqZcxj8Zhad
oQaVxLISr8VGViSeIhqSpUtx3ko8BFJTMKpT4M2ScxHBPkPgyi+CxWlHREksx3JM
ZiZSlTJXcPBQTzmDOIgby0am0q31LuBFTlIJfvKVTYVromHENWjcdudIs5PHZgdp
rWJBOOCCu/qDqPKClxlJbvB8Y1y4YUi70qeU0VIMCfvHg5AdY8uA/U9asd96TiYr
2StXDyw1PjLiLu4NBTCbfNHwiGGrd92iFqoq4xKqQy5Z8kgap6fFeildT3FiCJZ+
ft4NnOANEMv1RPjqNera6Hw7N9IURdyiF0ccrb26TiKQfuAbmTx0YYCRXbzxnSmV
crKgCt6bNOub4SlsfmLgV4iUSZE/HjWQCIMrHAUV+DUn2XaRP3pFWp1Jbpi7lglD
zTtlXR+dd81nAwg58hilRAfK4HbRTuvmQ3pl0MZeWGby0tc7jMI4wLn48/bD/ETS
i+XFBVHao6NC1UCB+unNXzenozsOTHN1Q4D1bjkp3K9JYuEeVpRV01z7hUqNCuRP
OkHyInnfy2Kz0KS7A20lGbc+i2OWhOjxVTPUyUtwnoYAEJfWlROb6mkC6BYG9kjV
JTdfT84Bwy6FtQxrzlCEpGuNrSPyuVeOSKTzpOJcEtwe0A2a7a/nzgBoVYq6j7Av
Sg4G2eVb6NSOgoDk0rS06yJuEA+tBOddyDlr+3oXB2iHD9qO5vaV7lfPez1jULX1
XL5yd3d94/gu5NRzTKF5TamCAV3+lq4u6OzYwXRgZF5KfB5BFih9xJYKxqSgeciK
8T0FZL2UhcpFr02t5An0+2G/ye7ptw9Z/zmkiGTqFfIeVMS/c9QrFNAYRwaLE9I9
cclkWod7cQeFSwNtVogNDsddxoNHPycnkUgVJ3ZZoLggAKH/VNYTMqYpy1NpPDWn
93wK+w7fqIsSH+8QngsdUJV4EVdrmy5tXbu/cKBSM+VFAVI11Y9NjKzi5mw96Jr4
wxkzHo62zfzeQkhgD7VWdA6XrR3PVVby9vG5c4H/k16cHyEGtPM0COEiUem85KGX
iM7HFhvfpfnX65raT+PZDTu33/NkenSK+OKH6myYabf/btCYA+dimGWQ9iV1Wgch
BZQjSyi11FiWkgw+Ge6Qlu8sdN5isG4BkEX8C/1IdHRodCjCWbve3QLIhq/9OKHw
VXBohPcAEhYdn0sJBkm/KX7Khbc1iUt4o4+gt60Mlgy6+moISukIpQUu8gaJHXxY
3U0P+IMukjmURTPyU6zrwSf31XAMVvyPtvwZIhntzpZdlyy2PdY22OQXYcf/epkx
ni/uvQpIpv9R4Ft8rwOIT3svCmzniNIJpV/NzUNV8nTo5yzDdmcGEOV8qCJFVn6Z
+Xzt/avo/YJ3fHQBqOgDzIzhCmNydFCuBf70w96uuCOSTfyAIwETIyVGD6wAGWDO
cX+eVswU9o8odvVKec32oqB9D34ijUltlE+S41i65RoeJoy3pOMK2Na7n1ds6CHy
ZD7UDQnwK7cqM/vU2Rum0L5ufdRTopS1pDAIbXEhKTVCrWQygaOrzzo8/8JxXAZz
D99W4r6vqpC9micION5iq10uXnloRbjrdc/LrsXjp+u5Rypl2QjT1rCwJ4mwrNMt
qKvQoY7mj8i0wrUXBzIz7t/OlxhF9hSNVbbCJqIep9CZUJ3beEtyJ23D6Fs+5vbS
bRabq6wNGBgeVzlY1D3Cw0tpZnR5rGOQP5FwFjzhSevLBI0iYeRqsx5+GUT+0QMN
rp7fPSm4ijf+v8VHbyuMS+qksE707u+wWuwHfqzi3r90BRDHfpl2uNRsakeoI8YS
r7kDuWUaTMzOujHBXQf8nPnsEljGl5J9L+7sHfU2up8rPBMqe280p+HsfY6kqthW
4hGI/fb3b1wltZlZPASNfuSJUlACxvHZ76xgG5NtSOVmcQs1AKXQdvAUnB9S2XMS
vHg0J6YPa0M7zQrBgUHy+PXVH0wtcDzfTMTptVTALFHLbVcLLUZWeh4+7HZ1S75I
OW5AfXU1UYKIWUWGlBCLtUNgFKmv3J7wtTuWFQ19Fz7MX14izzBr66F21IhFgX7X
XS3qngahs/P5shblvsu12j5yxb6CQFhw1CJgwBSKZ6axK6OTGM2R8VBQ9VhfM1Xc
UKhvI0khToEZ3mvbxfiil8THiyIDiloSmsPoYy+juJmjlHJDvQVKNCP4o5h1ze3Z
mkBYiZ/Z1vWw/nEtQ6EKqRxSYyFLpOdrlSh1EVytxbkSEM4mie7Fe4ghVNaIFE6n
Rm9XMIlvuwglszBbikCFXwXHtI0HuF9E0LI7ntF8YdjqcJSGRjt1/deYHzx0XX4I
/ejNiQvfg48CFXcgARTe5SoAKQklHhvrmIJSbvziaEsJpCP5Qc02rqP3k0A2hmkh
gDBWc5Yw5Rm0W5sMl/7Bif3gr8tiULWMPOyr5LQenkeA2fl5C5IuIsRDNL1Lvfk4
PGlu0h9hgKjLgipiHa1yEkVFwdqG1pEx7wYAY+IdA2x6KScH13ebGf3s3vijNgcx
8q6ouC7Ti8soMdoRxFpqRlOPNXEKSI5zBFhY2ZG66VN2NKWDu3N3Ygi6Wa+tKtKn
xAg36s3k+4cFdHYKZNah2gwV4WAAr2x3+Oh6W1ONQLoE6JGVBp+KQ+AoXHQt5Vbd
BcJ/9ClzFWAVl0/b6P74+XqxW4qSNhiS4Chmr93mjnVK3hVAjLM8a5AaJPlFiJnR
ELjllDp5/FBz+UoK2X1tT+l+zosRwjFUY98R1J8r9WNsh2NdsYyHw2nEFcBJespb
S7pMFg/qSy/VOx9ft+JceZVKYtnjmacjzAi8YvMSqnuVYS6HCBVtq+5CuxkzyuDi
3wI6/5iEPbb9MhyR4o/xVtfVwDFSoVzhSiISw39QTduTtNCqbTee2Ng+jWtUTfRH
YboS8RWfOvygoygsiBIVH9b7eeETbXq3ZsbG817RBcDvrW4qD6Jvst7ROsRkdcxq
ZU6a9TfKDVC6GQ5MC4+qynNH1XhI3KgmZiTu92uUnXeiP4s6TFAr+aIkykx0JNM6
bbrkBy9YdPUPdjekLczxvYIqQZbdaPVqbsmcHooNUL8pMRR+l98EiP22vy0J1SBg
C6gU+mim6ry/0EjmUUP9LNtkBu5imI1e4B3XOsdv3MkB0kSnsiR4dyLJrj+B+H3v
vC3N4N+y7sxAagH3KSJO3iHQdUIDl3sMSAWTjrjQXS7XdiwH26Y821zCgpDP7I/G
BZscDJRO8oIRZ9NwjoEpW1sXFgvZlXo3p331192jWfl/P2AgxgtZj0vCi7LAmlWc
wZhJEkuc/zYDemVQEvAhE9Ikdqz3eR6tc4Nj23zILa62tEaWoSY/gQz75VRc1ue3
fkS0X9iyCV64VUVMzbnhqCTSvDZdIi4m+PdcCF1rgIB37AXe0OCVoFCeHHssPqo5
8gzfJfkb7aDzXArlEfM7hyv1XlmetRrEGRIy8DqNjvAdkCNKEyPQjVGK3Ev7o236
AnL3NR7QqXxMMzN0ps5fLoUYyQAbFB4rlwSRE8DuGJ0iIdcALKMxPQvidjafMWXp
ARrfex+nXXWD1WIlVZPWWPNXHMW0VaoQjObTeWRrU+qof7dEPBxq0yNw3oGMnqBy
zUaYV5Ww1H3IEBxn2rqd7/5DhgocSzTHxFrT6lU5J7Jfc3y3J5FmnL84kHhAlUzf
6z6gLklrB7lY/cqF/CgaAzdxntcnJ85PkOxPAAPB72JSuImGhJQj5ZU5Ybzl3bZA
r5eR3+JKEyZhQQZUo7clduduq+hvEYbA61/6COdigKTXsakEa98T8IRUjg+AbHKv
qKcP+byErun/qmIL01ZD772liabdJAU0ems14k/UGF92A5/bLE/OQheGCXfvmE4J
aho45pFZTBzHaKmP/OV/0ruYoYArqRVXC4dldUWVB9rKhj7MieUx43kQUgfPiKT7
gFw6mHNdz6E26tIpGkOHKOZx3q5BEpSpUEpldzrbB8ke7XSUH3J15nzKL+5HXvCV
hifc5qQW9GFcd0UJQ8115fO/Sfx2qdg3kKQXceHNo4INcOgT0CgpIX5/e/dxJIXu
txY/oGb5OkSWUOtFacpoTQ0QvDmtjKAkVhbdFXolVof1yQoNeH/oxzn7L1BxQU/n
hCfjom8iP+YEvgKFTV1CtAv3zmOIpe+MkwE94aT27uxQyXunPZf0ZGGePPjteiKU
vy7zScj45eqMo4C6B7lNy4FPf1R6DJeDMG1ikVJ2BUyJ5LOCgHzMQM7Q+JDi1gWu
5ZrEIybthlSvytxmAn4xUB4iDkELPYh/JIVlvSG7mafE8QMecBCleEFjk2QBN7c+
EaCl+8qjvB8wU67ph4KTqypL9peg/D/UW8SB/B62zaD13P+7k5oHV71A4fKy4nie
p4p0hLKQuIzZGEn5iR2i8Oh5VKBq837TzeP+5BnOZP4rm5iiUTdcmJXtK8foEz1Y
67E8nupN+n/ZgUMQt8akAhYrH5yAljWk3opS6o0LLaowYojb6igNThyLqC1Lgi8B
Jx9OIRZAEcGZlcgcnLGCnaeCGIlxRWmtGZRv7tttNwjfE1++2rVJLi+Q9aOemf5D
59UPkCUXQ2SLCtTyqsWbYHb5jZWa8DhzWn+gaUtbKkTmjtt/sI62aFTTc847PbWA
qnZCw/jiYiL0FzAjqGf2HJs9bIU0wOuYMbPTm99r0hfxrMZQ4XAkpWF8ApI4zrV2
22Ryqd1vefE1NLFTgtlzERWlxj+hIjpfvU/MwQc+zWNfXHFmnaYgdKI6eIEHrsZv
dKa/xwJNmPKgPUCP04vfv/VhPjOMYnjkKA8+7Vtr3iUgc6FmXbnSRV58oE5HuSo7
vdk5BEMShlkvTZ6VBrWjOOeaDmW6pCV+ejcUpC3eupHc7yHoNZDnbnYe3H90GQcQ
Wrcvj9/J3OG/90GpswsiZGieMjhUbPr6RVbG0rBv4fYcs74G2FytU57CeDPrjtI/
MZ22CzZluRsyn5kAveDVS2j/WmiHQU63sdrYgCknEpPQpRgJnJzbZQvqStOprsKg
fn4KrgCscbaW8+pTIytKaBx1AuRv2Zfq9T52blBfSDuxC5Ak9xAcW+MIsiL0uz52
vm/bmoPIFKNlr+52O5QWSI3Rw/gWaSUWrIvaGufb3GiQ5bYyJ0VGM5ZGOsXl8O/l
vCnns7vYkde2mje/9huxKZ7UvtxaBdq/KEr8bkcRpfXJbBEdPNc0CLrnkcrlRH0j
FrUes6FDOqcpbmzCqKvXbv4PLoRqi6SHm8UKs2JrYhY4IHemFv6iZQdDmZkHIHKf
EZluUyG83HSXop6wvghN9U6VNhNgA0o4iOePSYzrX1Jo5zmBUSyXeJYHfUSWYfU3
4r9jI0HxQz/nhQ5cLWbO7xfGl9X4WhAMHadPLqRHRycBP/dwUeltwLyHADLy8rj4
D8jocu+yj9WVsWPCoz71Oy3RVpv5KHpApSzVtAHtqU1O2TgUcREyu0l7p6xDZi6s
jusueSJT/+A1ea0gpXXnDByAf50QRROx8jM8wYyBCtS3K8WQGCGJy+qMmfnXLk2S
99PUzw8z3RQD3tc7lV5+tLvR9eCo9qd8vUH58PpzDRFrphy6C7usjjPeUoHUbVhu
q4S9MlGyDOjuBZ0zkLKebNJB1qwqlYKJwYnUTZtbQ8s0Vd/ckgUdtjOhzADo5aEi
PZruEpBc7a+Uu3cLBQ41rR5S48gqAF0OZn+fmoXGitS7upqgkCG7Ou9i/FWsIIRB
6bRN3rCizMEYDhUBuBcoJ6wVyZgD8ECcoA9VEy/dGo4oha4XwFGpecUdhK9wSikN
UI/eVmbBKf3yX7kM+jYN4gNDTBiDzFl+ysXqM51Ko+gkzIZUDDqUgnyJqswPEDo0
9MxI4bBc6XwKhWR9sW2v0uX6HEG2Us+oMQPiwiWYCLfqM5C3cfTZmKjazXtJMwf/
7/mX9G+7jjCwg31vOrh9GkXCBTEU5iPWa33C7k5dMcxuiMJQcH81ZkLNgsdptKnP
Hxje7wjIiH1koebp14mdRzvOrPQHUXJGwC0DHb2QXc6SBjcLidc1/191sVcPV9hk
W1P/1SHMzBLQ8/3/K1BcpCL4OWwCviCxmTTM1+2Bc96wZMyQGqxIH004kw/c3l+E
PyAoyq712v800xQmW86Hyt7jvhmFXYaD7kGA9uzuS7V9Ds5Kl8Bt1AqFvjk5mCNK
T722cv708xxPjy4O1aKMpXk6hDysJXfv3Q1Ahhnuu70rKeNhfQxhGQPcsmPf2TY6
CHRZPra73uoRmzIKpDzs40JVDnVa3ykFIOBLniNjRC+5M9FE5obkLG/8hvbgYUye
8WdyLWAHNF4V4FAUs1zldakKllwRyoWdwrmFWx8r9oCylT6+24aSvF44TiU4EYuB
E6aKYSxcgBeJK49v4seqUGk5bbO1BfUe/QE1+UWN1p3TJLW+zmGzP1xUPl2IyoNA
zLB3tuPKQ2578z6f1M1tr0iw6fQOmsL7lSp18s9XkVIhEUbTrx0xUK/1wycB6la9
L6G+oCaXqR7c4HlnH+l8rRCp8qNes5VPKUAv1OI5BY3zYBy1wP7oOlnpUJS2//lL
fNbEAhhPhIvbbKt1l54sKk3odOZfRDq52SiaIj6lWz1+wqEznVE6ZZ9ALD7zRvZG
+5FKmMUiOczIWMTTV52Cc49bWSUoraKv9gpsxiUt1ZK3//ho5DVKNmpkOUixZJds
PFSi6o6OnEuEamhJQVsifOnPpgJpub086SU29ioluLoOUj8d7hJidL++fiLNc2XO
w0mBAzYLEFG5Q20SkuqULHd3AvDG65apv2MvLriJc0MSsIsteRm6y55x/QDyuive
uvOJ0g4qePLymMq1L89YYRpMUhn6hLVEh8AYJ8L+cf3eSEcNOT068U8K8KFTnzeW
I4PB1y1zLpqZCkOxsaJcoOtKN/AxsoMLFtK0EdJa+SjFwkwt7hp5ThU1s1FooWsB
QG6mmJ2rojc6pCZWQqsEjaWtKzGV+YbEzuNOsDvOHkWnedqkJHAVPd3mRfGRx9VA
nX4DOjsrl0jN90hiBZNWZm4WV+rn3lF5lYqUylxYxqeFJwTma0l80+hZWn40RCzD
YbmPqFzLFfrPd/f2KymDdzUL0v+DkeReXAB6w9IEXgNhg424B0cvLF9kg7GkXh08
lte0thr7F6HxH2PP8isz7LU4N0fJsaFwIuVpaL/8qrVozHpDtHjk97bfq82i+G8/
JR3Q4vriNkEWPnD19BOmqfL8MW/QFhHJtOuY5dMRrkvtRZfi10JEQnAe9k0e7D51
+J5Cawkw3AUmv2xyLfP5nijkIWvJhb1ERxWnlF/H61tG55rI26dhPaMl1Vg2Ixb6
Pd4j5UP6qoDBXtTAkf0TFZEWuOco6LGXHk9O36P8avrWum9nJTMWzXtDCfVb9OQr
AzJZSvDjy9KQNN3vJixzykw49DrB8Y8KSRT6vwN/ZNnWeayy2ktJEzwvSE28wxlG
b5WroKd2CUWCP3XxyVi15fSlQeMl8+UOwrhoOTkSlYZggnrK3RB2W0tcaMUkbGdo
YxXQS4bm0bviYa7X26ewXGXaKm8mPQIHkFvvhIcOI44QR3GSnGGIfPQ795mcoHRr
vSdpnj4RaEdM9EVZ6M0Df6LbcEIySnD4QyOrnIWuWUy93/IpeQLmll02NrRYMI/K
BFTaJ1qEI/KLb5OUG1hWVgxvldqCXJwjzcLmqgYl2ug7nGXjy2/Gm+QExXy3z83p
IHhE79zzSwMd6EGuXbu5qMiJVCy2NCArZJJw1RO1kYMFLJfIFloOX3RWOhEQU+Iq
6iXZdFoQCYoC3n6klcHeZTYO9Ln+fajYMBIVWmaHtUatOcvYUnW4Dlt4B7ppmTvp
wwuPzIpXBu8psbT1jULwqggs0DmFmLpxNCq9a4zPfFXZ22l/RDn/fvEJGhZN6QRy
bkAMU6mmr50DBT94HDcmLUZ7cGysZA5Bey2fhglBOKiw7dPg891JCWdjUuOJKWyU
VUGxlWpYCdB1hQ6xaynJZdPns3ui3e7NwCubLPi0YWFaKfqRWmqYaXcukIvP35Hg
0cjJP1B2kAQZPbhlCqh1zZlSnpwtYiNaFq23Eqv3w+RLTvLtEvfiVl+bA5B8BJuw
8tAyubUs6rQq245a6ueHAD7E7fNCy8uhLg6lLLD7x0CzDhdjrNYj5zzjAxg1anQR
OpNe/oApzTc0PbBpwu948WxoDXl5UyETsqwDWR9Z7z09bJDzllCxx8PxMxWLT6UZ
FN8HHIG0BbAYVCZ3SlqFYvfe7Vz9Bg9t37OCKCVLqW5kG/YLvsoZ6LkEwh+wVLMg
6A82SPCz5tpytSfwIem6hl59iCTO04tSipD/TmWCk5wqu+abMPLgGbZ2swBMh07d
Th9xxr6tcdnQz9dIWK0Iv6sWKR4aw9QDg2kgfpj6vS2nkxIaevsgCJN8ZzsnVZqx
/oWdIEp9JRjNglpo1aXwodQ6P3e1YPNjLP/PkaubvV6BUyJfbaY6sGVz7VJbCFkI
P7sfXu/jI1WHU8TmvkywlIy1W1k0aEAjfq4dtKrdx1DJ8u+Jdeszw+oZoxvr91Xf
CeMLNs+RUC1UIcmWsTzCKXimOaY73ZMbappwB1Ivd90EjRJvjV1ZTB5tKLZ2TnEI
Wbfj20qoK/PYRbDK+Ejnry/SoqnN9bOpYqlTsiUWSLZmM2p1P5TsikKe1tdyf/Un
Y+Atj8B1eUp7ZZ42DS/34SoHayU7xY3FImOB3qbc6OFqpjCbXhBm4gQZ6IpctZaE
UEnGcK3BxfMP08wJoaAEHJR7EVrTt9yvvtf84ZUAoDAHq/pmfY86H8j6h+MR7aL2
V3AACinMwA5UcxAob7Rnnh1b0CdAsrZCBdL1ainqJEFaf0AyapC3SO6yl/qJ8stP
ydH7yHkXCxcxhgzD1RkveY6D6jfDKonxu1lwRmbsgN9z8GTanazTqvpjd0q6532w
Du+7HnlM5h3KsoOV5AvUQ4it/KAcZHWG6XQkmcl8OoTYzlGO4p3P4JWs6QQ1tn7t
brpbW4TFn/p3E74oxoEj/LGazEbygWuhc5PnyBwliTKILZxTiIrz5ROvKPn3G43s
ew++LNyAwEoJ+n5xz1LV/mzF1bEVow+1asAsbqVrfKAehxLjYEADeWopsK/YTZAs
es15LZJbV7BEZMHTEy2eHU5vUWMaaKFVhZst1X/evt6yHSzFH+oURkefs37sSTaK
3SctXMYlhqL71XxlcdKV7LyJF6Lo87mkNeT5nYHEQHhaRrqMpbX+x/bk9hUfd3p0
qzuH8S6fZo0UW6OtuDmF9AdaMpGucrIiSlSc5lfsm1Rz6CPSRA7UHKKIJ+F5oSNu
s11J1D2/G4KbGXPoxGD0bM3+Zhth5OZCBDs06J4Pd+uTb+aDbNv4u1a4Gmwpluwx
1SOfShv8xQ12ju+aUxuxeFz8rSFqbwE0u5bvdmdL6hgG9n+rXjzbl7J5QwULRROI
onCglwn0SlDHaxnyueksu3Evuwy6M6McvTCYvniEnAGn50TS1RyRjHW2adfX6wAQ
AbcNsUjAPPppeswZrU2d25aQFdWZ0Ho5zs5A+kV6iJ81YFUtRklM7i+IwT6IHthv
VYVoUFegMkPGh/nr6IDwWnOqYeJ3DArBQ3NRyajwIte1gdQCY5NGXET2gFc97dNJ
bWKWJ8tWZ8utznsp9kfG+dpq4frNniFd1IGtK5OkbKC7IN9y2YUHuSxB8kFIeREo
TxKiWBOZ6e0oFguYP/hjNvTEfFQuFakFZEe4mm60RnNDzH4itbovt02xNOjR8UcH
G/LC7Mu8483HI5XRxVoNKBr4FjwmK1NaypZetnc1MisnX0VCNA106yqjQdtolnFZ
LqxIzwzUemX3qjKsOMJytcWUYb5RC61EoxQ6mZyA9u0TXtVQzOGiiQbmT2woWenI
//6wJD9Sog8YCmDoQcEeE2aJaw3kGpuUoyTKucJvo08JCtyb8EItkD+GqfAoAlaX
iSiYQZMjHLtDn5Ptqn+ftEwj/iKNlxxOz4DkG1Gr/SpoPj3kAuzwuzM8vaeM30rA
ZG2MjTgA51eDsNwF1ggmbJPxVuhh21R8V4vj2j+QZ9IpSA/zfr6g3xF1jN0wz/m/
elNZMM8MtwvDKhoB9egGgMFyavkWca+FuRHem2pRPWeijl/OdBreSmoz48UHjN94
XPvv1xW40NTKP1KfK5vysLblaiY9Xr/WZwHEge7WfHcdjo3sbwoioWjHLvKo9JGU
rRorWWqEH0nFghhYN60f0NOyPqKAgAS5L/BtzT+fhqkVDGvON/qiWwTZzVZ22XsD
3LjvBTAoy3l7I+In1s8VSPG3++Tx89as/WqQGXw0ElgnEefspxhSDBRsIxVbHW9U
UFv0P7z6pOfECtvhKLI/FLsx1tTutoewPeGQXfXg4hfnpG19Lkoc3m6K+SjuafeY
DhaflfNJ/MTlRPi/UPh7w4mV6M2FCr0tbk08rHJ6z7GaUh0enTdRzNqbWsmZjblC
WbcRfe63mPoFYwjpXZWFYMl4wos/l1IVF78+GKR/aaTKtG0s0DHVMHFQ7c5Wy56L
bX7UZLQNceG1BaUZNupg1NJ1HRMUg0sJ8FMrZJbv/O3U6CqhQ+Az3+AlM4Lvvbyh
fjlswbfrqZUOsUXopzBss1/R+1sbyUKCMGKaYi4YyTBX+iBxDoHQPuyySqIx5niQ
ZzfULtaltN1yxGkAotUtOv/66ShBHykgbyblCaQtaiuBSOkUSj5al6knx5a9Nf1X
NDcnTqfUnCsysXVHE6r1/1CUEG/OSO7FpvXCFkMZ0APKoQRyUEi5gtI8+kNsUieH
en0pmCRMcEthRwHsXlR/oOH2nqgWVOIKWrHyXABxd0VJSm8nGpDOvLQi15syBKPW
aMUQtBxGyE+S9Rfi1g0TJIQoDHsvZeAYs0eaNEjSjp5lwJBsUCzpbhRCHqnxq0/A
KqDGidgL3LMx3d1ydtjBMZjvxC0CAnKfskip29m+s0MGGhzjnAZ9l5oHWHPo0x0J
puT07EmrlyT6GGA5DB2E2rQfysWZuiXK97mmD6mwSuIV7txhddkY32T3W1Pp95SZ
XT88sKcgSP0w3sOXHx0Pv3UJkwhu1+QRXzUWJcGk6pKGbn0UgVt8qlts9/DLlSqu
riyePkIKEBxkSlVGPAp+8qMzuKKFNSxDEGMnTCur0LEMRrI2isCVusFr6HzAFv/X
HtmuAIrzwHQMrCFy5vRJ9tD4sxYmAm4FntF0NQdc3+1L83WYKX+ozst6ET0cvd49
T2oPJc3zKgKjslzJ4011LRJxpOSmnUiZ8sW81jTW5blz5exCkixIcOp0e9ZVyQmS
0meJIY1kKRJs+gudmkPnqWC0cqX2cxQTLGntPX6vSId+Ba8olOgGwF9wrtG9kpxA
0X6x0Vb5nTyGYliFm3oQR0nPCUyj474l+9ZWGXPuHnYueFuI/xtdZEBOUtzCCQii
p4LaYiTkOqEUU1oyz2BzGccQnU7YZXxWydOqVmdrxKWzQSljxcFtj7vgOZkMWaef
5OQ66G2mtxmFMSdRcrm6L4RBTyKlPYn0ComO0CYjE5UzmF7gidST4HznxP/l1NRb
Jg+qKM7hs8QQZyuaVTtvMUMRfuEAp6IMIgK70LFMo0grgvJ+jdZUuYRHnH9DriML
lxMbZEqyfY7HRHL/EZAFBL8obq2ciLUbzDO+q4W8q5OQd7t84SNjG9p4PSKY/r8n
lCjQhjGnzrLP5pkq2yH1/+gL+9lanV2r5aguu+Nb0k37cwNrPHsuiNK+Jr2P+w5M
CitN59sALwLO7EX23KrqDTANGeAxQcp1uGRZ5rt9pqIS74UBapo5XToznCjJOOMC
t5ykmpPuppx3qDzGJ8W71Z4Ib2LV4gpL7KkW5fCRm+Dpa5NcxVc3qvFS3pxoyGY3
jyTwos4G4wTwzxtAlrIAjWsH3n6ggX7tShHSmfQoiXaDZpFmTP7/bbXXZx5f7FJh
7KbEscNmXf0NjNcg3F7VAjlx4ngXVOiK/AXKWmucFNbHi9LbGfXDpGXT0pBk8b7F
zStL6ydy0mSIhxdMtPbF3RhNmos6LSSfsJEGucVKCKjkwxbx1pLhlfIoEQPvVv1Y
pFoTF0QEIKExJKwHJzD4e5/H/atMDnVyWeHph/mkHI5hKdNQ9mgfmaCiwj7ANVl8
RGZ6Ztdspk3fY9w878tfsvTJZR11Eo/4cK1GC/nCc74mtkhFxv/PImGktAbIh4r2
ssqeEiwpbn9Po7puzo4MAVJ5nb8rIALXf554zYIwzHO3Jwk1D9R8UBAuN6Qid9Ma
DAL9qRpeLJfXKAEK7EC+VSnizDBs6QraXkCow3XscW20kW+myHJqRhbwjkAdD9x4
L9FVpLzLMJIVKKetUcGakVaWT5yAXbujGgathSFZMExJMX6D1sXzpEsdg7pkTmFJ
0o2wMPZZ35hnMEF0a31IEKvAwGZ/7egqXVIYrD1dB88A+AWn9MXDx45i/CtUUrMH
/BLV1vD1R73abok6TsMWjJN45+aoZvVV9FgA0FkF2ICZ4jOmaTU6FRHs8Ey12FCR
/k0I+3esKlzJWla1FUaQVExYlVXrJz+6xoODSPXyHtKBK5bTsRJWviZqgXchOJcy
Du5zgrUcrV5y15QNVMFzKAvTJgdOck4q7D3vy/0UvT+3/7o/+ThQzIWKa0it/jZF
y6Em7gdCYhMpRUQ8+vNpFY6RnRp/Wg7n3+jKQOK/qEyTPCkzzcyVhNCHjsPGq0qw
mxyawmmmnyP3yuLRKa4IgQ4RrxW1MHJ9pTmACkHCggp9NSI8ANYgYnGRUGHbdDyl
6Zn/+/MtMOWAsb8fepWgFfPWbWAflkfgzvmzE/x3icSiUhafzZgTL3YfOvh8z1Nx
xG0u2dYF3VuRxLW/twxYH9ax6blPNmreaUu4yAkWkY2eqEo1zO7Jp/c7j0L44Sip
qAcRgygmB5KVJUDfnq/vWRvgfRXkYUeFm+Vo3ktv+HaXGoPyIhyMSN7Ieb8daRUP
YOAmsQYwELPn8XW63OKi47byUB8bgNDOBrsR/L1N4XwEUAnqpPEJvn/p/e2cj0Xr
2WckV/56gzgdz6XoIqecLm/g29J3EDsS0A/5fPMim7Hs6WuKyJ+x6tkgzwlF8gSO
jI+P353ee1hrcfefuLYkoJ479Dt4ZoE2gXiNC60z0FJJYW7HvuVNLFAWUKNCsPi8
37V4eJlsl8WahWaFfUinwzY/mXbisxmp5A4A9GCwBM908ECKY6+EH7GmcwwMKQXu
20T4hzek1gd4oSKfGm+N3+imjYbE8yImVvkk8MZEGSpUe5qybU7ppp8r7ilCiMm3
LRhPYY/rG9iM8h+CU/FLf2M4Xgjjqie1B6G5LUOQYJLgwa1LTIuPMVhaISqSBFQi
cW5PcrH/fimtxIaRPVoRylpOPe3CiM/JQBnz/s9CX/6jSby8C6kmvKByOaTNdgQH
slhk640jbXV6VAbP0nhI10GRlW5H3nDJbOEEhKKuf+bbYpX7b4OcK/AikVJTXLOB
3uXkBT0X++4UM/9o+XvPYHZ8jhGkTBUs/Incdl4AQ1wFFpg2Dynentp+BFJ66cHa
5qbfqD7Fl+QQxEaanPkBxkUkFUGKQqgVV/no7Z8FbbmMxhJEkEnWT8bs6UT43kJ2
/2v2NinFrpkqsU08mCDslwN16u/PMNvUqfr0m13yh5HOwdXG0DDKoFUwDu63OwyM
ewUhFf+A4FEVjDB7GASwPbrJSgfcebj+KmG1vT3HVdhzxSh/1I60zclW0V26Zgc8
sAsXE/yYIjeZDctIWZ/mm0M66iL8mEEjrmqr3iLVzB3+u6RE4p7xL0m6mhRyXRGS
GIMis3/+nTjQeZJ+Do70d6aRUbtukEAdOUkq+Elu8EfgGob9unD82U3kMQV5c86s
a6TwmPk75S2oLU5X4tePchC2IuMXzRgclI20yHx6aCPmJFnrZy0cq9iugEMdoGw+
tvIXz+jdZCYjuGXBvFH00jMiVSXWxHXcHZdH16NoI4k8zxOdUUCPuKdWMdAUFjKv
Ud+TV0FR8rM/u7fhDLdygemDqap6DGHJMyDNB/w0KkGITK8UVfCc0VQS/jaRO5sU
oB40dLZ1/z96eGKVUSbCsAUf5mfmV24+AMExOLHA8etq4pM1eX21ycoVuky4iJ0o
UsaZvW47M74lVjmJB+3jADFjYdSksc2qx8AhkOgJ7xdifX23EhH9ppOEGRl+axON
uXX9VHcqYyOjSP4yOjHPJrQiaN9O9lU2dP8pzzQSSP89aRNFN51UGM1q2Ge1hl1q
BlSKpM6aN+aqWK1fAro1FEvoPD0l62BL4hnvL8XBhZITELsRBOc+IQaarL7rVOue
5oUFJouIMjDt7s7fby9WUuH8wgHjJobHZXf9VKisg6pCny8HpJUmEwlon2qov5jw
O5gSUpu53aIXYtiDdnTcBo/kjGDE4B5eGQ3KY0jgdYULcAe6xznagTD+IuuW2kpD
C4BxA7znuSYhGDh2oui8b1fWIfKMRK3WMaAFMwW9Ft0JWUnspu0/vTB7Goyj2W79
bFEkQ+Mk1/lp4mXvgSvpwSrUaQebzdjbJ8oBbxYq7/Oc5mzkl6szrn0tuLKjaTm0
B+9zEzEZk/roq3KIkPkp1hpPNYTyfwj9roCMSfOwqIoSOD1AE9Fe3LSMCkm+mWcp
BYWrzZllxI3BYQ7XigM5OyQPXfpcPgOhA4+aV7bLGEH5aFmo6sXPjf/lq5X750Q/
BQsi/UjiyS4OeYpLeXyRR06zewR+MQ+t+i9CxGJ1260GYr+1KYB/10bcp3ykGzZN
akZq8+zYZV6KXIwQVplgKUeE6MKKpFMmd0WR1QVyQFDZsXy5zT2yGrs3FBaHZpOO
GLIcY0HLUSi24KTMzZbNUQTyP1SNrAVseUmFROFJAkwQHIRe7YClN5oqIFxLWed8
73RAnabHRg7zttsHT7hJmCIMuOkNKVZ3gZamyBRD8Q21k3oLz09qr0FzxHCta/62
9ctrvyo6dWTQ0x8CqNmWJAD0Dq64tFkFvnoCmhrXQAn0Z72KjwoSqMklvIlC+DFX
4UN2tF9WmznY8v2J+pWfY7GSyab2zNLPnFJP44Nl4Q5z7SeomBSUNnnZ0ghqBHKF
OM8nfLps4bqPnsL5T+QhR8KUJc2uC4/doQg5aMHIWy3+U7dnEvesm/nnBN8nilC4
Z4PezlwmdKmhCyOqNbnqsKkEztqAIZir3brZ7P9DORjC4mjHOW+HuGugJCMQDEND
S4l14g1cIsGViG/hQ850zXUMuuN5v1k5cPKZnwyvE8CE6x3sZnyr8Yg4wod0nMeH
aSnPL9E/4TWIkRtlJZ5lKevyANl6ChLF2la17GFVDj0gbIdCuO+rpHu+b6u3vB0j
kFCCLEcDvGKCBSSrWhMVk5wuDRWhAzaT35doalRwf0k5JK11wMJ6SKMG/yIP3EOq
YdBLMDLiJVT5OuHoVHFJZeBTuqCgIglsPGgkKHgJ3Id3gK0mC4Cg8nMYZEwf3Awo
aIn8l4PFriLybFQ2C9ThqDwiRu0vh3kPvhZz5UJboRngUxbH0mIG5BkDXG11E1KT
m74+8uxKM+QDjeyFewPnOYDZgjgKvKdCp8JshQyPluUsUFthhyH3+0/tsF99bF2W
q+prtkqeTfY3JzUAh/XEuTYaM3HC+qSiRztT28Nj97uS+7biI1QkKgR2lrFdResc
YrNIGQ/MnyXBKq4kr8wzMFPOiB/Zq/7Ib8rfGlCjnbjvLh2l/7k0wznQzGSSfbCr
7UPdoe7/bxVNFCwniyoqMdtR/DYnRhVDARwPEWDkuGu0iis4xzKOdKYk+yIE1uyf
CATh5WKWNMcPjRgeiXSiN/ur/Rog012odK0mFqETTSLrVItLml60qRCsbKqKrEUc
k0tyXkEr4L7s34DjPvN5mkTV2VerUwGX8p30TLC/6TyjcFrRkakT/JHjO4cF26bg
BJKm+LvcBWAAc8De0IQ5PtUjP939q684Ql+PVQCrbqeRHByQX8KJs8MC74Rw5W95
V96+urVJz9RHdBVsi2DrwzIZXxgKalpm8clHS/jEMVmiCqj0QtXfIoVFzP1yPkJy
q7wHP9Y1s6YrWQBq6wc3ug7iDkRmk25HV7GTadP0ENWClQLxyNWxmbYpDFnLOvHu
400OqR3YnI1nTiBM+dti18CSMzewfLlUOgN0kn8P4jbye0ys5zAhd9rWdAbNG8G/
NnHBy7NzjllkylZ05GgPzFustf3TVgUOLL66H3f28DGrkIISAziHF3A9fPHcszBb
Iv6ikbFe3iy2UvVjOSiRA6vcVAR2lac8/mFUntxaCmWsqxnOMx1yuxYLexajyvSO
o1t1kGDrmY/GT66potc467GuhWlCusYdTupVJrViCZoVvlNtt1P0+NYpqtwDHmu2
kExTy3/uuPQddn1rEPW5kGg1fP/zNBR0ziBQUtagY+2M/1STEyhKzwBXlwqpF8dG
qiBTGIaio5uaN69vGn/Oi/DAa9bHcZ9UGkmC99xbWKT/JCBejVqol4nn3Z8iU869
IcBJOV5pm5oLXDdVnvHJDa1SYf9HImBZzIwOER1QkwXL3KuD+PDNjG0uzDiMnazT
3tzqbF0U7daWSrYrQOQXyFA8pBwajsI1a4DeScg789LbKKala8DnGEjTMP/lyY1N
ng6Iqfok9u/DQu9ZZBNeS32unY5PsrtwVX3JY+rA5FakQXK951OrViKCntNO23oy
KqyGjry+zOY/ECFS5BypIiGVdWMQAQ+Roc2/Jsf8/xwgPcCMxMNAq4vLYaDmV6Vu
cEgoBn4M+4Rwwici9/Ns5Qi1jM5snCA2rZuByCX3Qns=
`protect end_protected