`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
ddtXksX2+yylW5zu6QL2Lhnb2d1sD00763mmSITNX595NcHTEkwn0zB1Dry37fOW
FufOhVzEJp80NC5qZ/+F0Vk7Ik02dIR0elf3clrjeJRK85K4e3Hoo4xn7YbFUIms
l/8VZSb14+JVGURjfswrIyCUotIzlzVYZ6gzoZwDXIi5gQIBf/gI+KxNXPaKV+PQ
Ufys/12rjO6aI/pPlqSm0hCvftmBcnezN2hk1UeXgOIuKZnogjOsf0iJVX2aOOWE
6pD/psybjbnsNB6kH5uFTA5frkzIzkzl5d9+YDm9OyC+k84E83I/7/j+rk4L2dah
QJOvksSIzN867/4Qt8qYTQ==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="MvBXkzurAa5VTw+1JJ70nePUfoQXBvZOku/SMmg4TwQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
oRtzZL4VJ4iwysPsC8SXYCzXS8Fw2gtZTOskLcDV+1B9Nzn1zTyNtlo6lNICRmmK
ZRVu2BmCc2G+fmzynYlNTnSa7C0Cuel6FYpxCBlOuk3OF2tzAmLAuDyOH3Z1Yjzk
a0aHuoCdIRKv7BrZCdALt03JeUmXKPdOmIlkVGFl8yw=
`protect rights_digest_method = "sha256"
`protect end_toolblock="Jn9CQpRhJt4rnzZPRk+dOpzAubz7omckX1MrFd4p81o="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 9808 )
`protect data_block
gD6l00tciPUa6pDNTk/+tzLxvdHE2s3DQL3/JqqujQBC/Ei+vcAB8wM3doqg5vTg
mdfn9XB1bLOis2CVSfu295W2DNwHfMSTc/8BhCDRnTlLIX0UCJs9Za0+LoM0rMrV
T7EjVWppbP+Em6PkVKCwlmIQ7JKaifJ+Y+kjw9HCGboYo5074hY+K/CBbfsBQY86
akxgwqRomai4n3Z3sbNPjn3fD2OVbbr/GfEPlBofsA2KZpoCT4j6ZoPFT72P25Wx
Jqn6rhQwHss6B3/548DGmvXLz+xvsiYCosH2xiaIztjavh6ZaFNP5f6jV+YxSZD3
Bo+jZKjXds5KW4HPsImADIo2JuobDEv3Hp9eoxieW4i0O7exQyre+IPaDiJB0VLe
dhxOWEJFd27iSeYMYNxBSzRtX4tIqzYA4Kxu3Z5Pk0bTUspaOOq3s2E0LT90B8dD
ChhtGGYyFMMPwMZOetaOOn4Gi+eYjImkQyUD9vts75fHPOBMDsQ8sn+i5HuptVOI
9pd9phbhwbNUq10cd6qzBMbCl4VWdnckEBWY7ZNqKREhGJbjHN5rUuEpuA3YC5QT
7kUKKzeo7AEIAlQhE+ITp+r0J0sJVGtu/nnhKb0Y8lsxd6V2miQ/iYXyZCB/4sqD
wpomCKrhwXjVHy5+gck07nIWXEmm1JxEsFClx1rr4qnivVNQ/Htl9g3A7b8FCA5H
/tL1JUG5iCNQciV+zM4Pi6IcAfi3bF9eEdSuOvkj2ck54UTZEiinKPInk57xg8IB
O4FaTi6P5P5jn2B7ElzWtUvcn4ROj16Q0B4IW9bgb5/hHlccBMk0wvsELQn0jcDx
pthS+WrKlyWXAB7YZ1uMlcypweyGvpDozVb3ZNwrDjfElWXBdbZHygWODZZ4DT1Z
ql7RUoceTluvAv+knXeJMZh8ZiggNHp5zSBBgcngHMCX61qTUI4Dqz6NCHgf6JuB
LnqfIahf7DDCNnu6OufK6HFsswGRFRHZ4/KFpOseoGe3UTGnejmh2QOOb622xiWp
rnpefGoYRhLn2kbtD4HSlCJKNdMuxg9fwKOh6qmDkIGyV+p1Y1Uw9TODmDY7zuz7
tbCJoXkq5kQmcqmeOHbcICay/xxCoPUYHRonWqMeDkpCq8sRmXEqW7WivwhoX7B0
BdSc4q/wIvqJf8+ZUd9tcaJfREmx0HKPRXYxfM9ouEKbnyLl3b+PIPogWKNOXgUC
adfyJMk5ew3A3Yp/NITFxDB0gXn7gpRoV5A34knGnILIZiDEj4wOHPUWg9bLqy2D
tJYARTHUhb2e8aOH7KCnktEDoSaquJHKOZe2iJ12mLBf0X6CdV1dV7wJMhzuiSX+
tSp6hjrcenZN9cFm6Dop/6SLfLqx7ndD4s2RXWAhUgce89znZtt1VstWywHpSOYA
UQifjKxcSMpmKeRvKAqd3DKBQmRUyJrvvtdzoK3yss1fdLrhaeBcSNtpZpkuji4s
IP5lf80b+ITo+Efgioa7U0+VI1Aqp9Ne+RGVKFkQWZiawiW6AtLudWL96Ffa0ryO
JNk9g4pUHKt1raZcwK1sV7pLNA+nKAUKLHyQxpivCX/yUE4v3/RdKl1ztAsNGNyu
Vmdt5HKvmyypR2MBsRxoHBuhJXiXzo7VAXSuXbiT3JjE/45U9d+nyrUSyCAt1tmH
qKqWE9tTRkBgKDlDYNhSoeyadcbSALMS+UN7QNdEl8xFH+YmSzNKdzm1qOZJmqS3
DCgSPj3pg3fwqVxMMjTbBAddumoBBn6cWpdu5tbjU6O8mZESrckmkMAZ29SY58Cz
cZGJZyJoJlyXGfDp5iGz0F6OeCETVcN4ZIe0tDqVoY1NK2fT6pDSMs0jltQBVCOv
Xe3tt4E70G3CEiMiROvL4IB7Z12usFpWl2R4qM4Vv7iEbvzG4OysAHobYH1ltpoi
yq76n03YNHA920SIrkzYaS2CBQEYQp+yjGmEUVuuW7g6A4pWzu36xRDFUprMZZo/
5YxcBSNQCnEcDujZqlTtkgTz6zaae8eVjmASZuTWgdGkVNl17cdN1ogn76wuY6kk
Mb7U4T286N6CfuCqKznlcsgI0Y91Tb1fi5h1sV4a8qabd0SLz1l30FPqCt6h/M/9
34qXInlMYuTtDPwq08TdT9r4I11Bezbhx2KHlVNA/Cf/TIWauAAOhDHfX6QgJ9T/
5efVnr8MFpqU/AgGq/0CDZ5yjGzSXk3CRAEmLUplyc3XO7XyzJTus5MPIygjqwJj
4sts6wA78chKt1CdvgCX2d9XmY2I9SvdW0Wn3TjIbOBRLqalalNYRQk9AWnYfYaS
uuscLwngKwGhNVeidP/DlxnK5Fo2e44EglWsAV0bih3+HpGc1hzcR8782Db4sDLL
kc6Spxwx50nzEnTVct9YrzyydEo9NfsJx6ztc32rb9AFC5JZSNYV8Ph7zaftdY0k
8nXc1atMTOZ9qh5lrYcbLGiPA9avDQigJ/1yUF18zy76lTlJW4MhO1KyE60XNNLg
e8P77qK/0snU7Ywv0NwYd5A/Lt+nREHwkhJLNfx/ENE43P2m7LAtw81/Nk4/Xz6Y
laRrRGAX/BYYUCWeCh/DQJRk5kt5ZwvQIShes2NVzSvTsZ6cRgFfa1yBkvdto9SW
5RmgovR75zR+hj17NMMMjyWS7J/ZmVHEhxRJ2UlkNjdxrdYSNMukYtrQGIQpGUoI
MgytZn58YA8GdrChenpzXzCnBzucZ4S8+BAldLw5xyhRBbt5K9nHves1vsJkAYBY
XSvd1gkUxZ/rrzQsOYOZbNNlqtK2bPFzcTWLd5cm0AFvQxBQgQsUO9k36OljSgat
xczBGZMJNXZz81TUvFwOnXFaVLoLYQ52VCaTotAoYRkCzCLCJuc1J11YfYMVckwO
olh0KHq0/zYe6X9CpxjwrZQLMOWolXyImalef+WRBWXU0EsCAVZiss3ZrMPjG6D7
AW2D9E/nmqUij0P0+4dEhk88IMI7wjE/45HE70sEDnq5IhaTO451h4Vp8YMOJbgj
P0xZZ2s9EB3k5BgQJ/JOh38EKe9Cp7MVLnEdaGDYW+YX/APYuQVRWRlfF/8uLDFl
hFAmtez7pdufq+Tgldz29oS9ztJBmudjr40+1joml91Vq494+Y3eKDatlVEY5P1v
36yEOuWtAe0LDgeCHDgLwvM35C4ZBsJXAgeI+gvFU7s54rxF/xLHjV9NWSNmDpzB
8utPacEK5iDf2gR8IErrYA4bnix8H3fRQqndxHVGkfSblhWFkRI61zL1LY8aqT4h
sWbm9u7l0LSHUZiwHBx2SvJO28Cn3IxdpGSAnQ1a3I1TYdtQOcjL8kEYD9yIQdSf
PuKDHFOdfhEE5ZOAK6Ov0a2WsKQEH5L1HAuJs3DsIAN0B1Au1FoxRb5+OS+HzY7v
KYgIgJDSchy6GYUTA0UX6A7/UQOM1dXHc6wUzRXWyJk5SoMTjlurrlh/HNibL0fL
d9TO73lKn3esh9yIscGiQoZI9jLQ/W1gzBXXnTG5W9eYdQ/sLhQVyvexkwuB1XKN
Juq/n64h+CZjanzhNLVFG0pKFnjZyf7+aO44ed5LWKie7HmuYS/cJdU/cDlFAWSN
Cuvoh/zAyZBgXbBnPsX1Ah4PWS2cbivvM3dQUAPJhAg8XSYiMoHYc80uVdU8wlYD
y8HqtctMP1ORUSoZGzjknJ01sRwuqZ3jDrcCfyeOsiouxmQeE4H47bQpCtRPnL6z
CIjtMVwOjFPP5gMc+7SXNzbnuKiuWMKqvpEFTnkWLsHIPtRFMwDG5qj2wpX/bfRG
EBRp8IuerXX/mesGXumHF6dmMbba36zaic7wb+NvZdGevL5fyan20tnXsoAFTZHJ
dNA0bkEuiCEC1mH5LNOtnG8OJzdhGyI/nUnwfkx6+H3MjLwPt1ufTK23gaIwSzLT
5ePuQciJTloSOw8+W/MiL35zbgOXX5YwCO8EB5K7U7E6NifeBfavsfy7dOpEuvhc
ipPMPmB5V7rfLl36jgBGdO9qSPjDiDO6KJYNOMQFXfZMQIRkHbLQC8yPPqaN8Iz9
gx1P1HZjSfTanEf0qQmGwBpMMsWJp2rY8S6I8L3jyYxVY4wM41uJAJjI+MUjMwkg
WfWQlSSlEqjQ+dnmoNZjop3Go9hatQd3FFGOGE6x6OcXNOL01GEnUFWTlTckkjhs
CC8yLclJu5Hc6zUEcJCu7qbkb0Y6uzNTzqvIj4SAqW9lXsppDNypDHb7n65ADYct
At1sXhbh+2jmktw5JmqxOZXAgQ4xL9m/nXK/3nGO+6ctfagcszsXy/85iNRp9ipu
pN/nCfgHw7JgEInrxsoxZMPlpYmiyjMBEl/SrGu+nqpBbB1SpOtnCO4blQPjG7QU
afEYe2zI4Otlyr30AHCrngYADZJ1XA+EfsGGzT8ll9f6rNpRknKc4rDjGPnTbZIQ
4/2kQg4YROsGUBnsvjdxq2D0H2PWNj0GHZSau7DCB7Gw0uUbsbGxObk7bwdD4/Vk
rbMu6d/HyHdKxpbDpHRK2jzaDzufqx78fGMWuYa5dpVeBXt4TNy7EvWePh2m8Ro4
uHnf56Mgk2xEi9L15EMJG5iZdptoS2SDTe1QZmZ3nwEjnkSXWj0yUmmNxouEuaEo
bxef1aga/RXEz2nJluE+jjk3pQX1fi0a3W+23CHI39ek9eJkXEIFwbAjjdxQF3TE
qiOHGyLkbTH3jgxWBGodvbOCz1X9F8JKzHUdVlrUxuF+J6nphwK1svRTRyvh5QbX
yABLj7sygMgM/zandhYAKM168XgxOTfoqAIbWLY9vOEBJ7I3f3roKRstBS1aNSUH
lv25BOk+uwIATbQy64rdyA4hjjgRDpjfPMWtTmfJ9VSupriguKb6APwKq47egT1Z
imVALX/Wvtq7okLPYQBlkQxFzNnDTRYWIR/Pi+axyLCYBuE71Yy2lQjQyVCdTShc
prqJO01H/3lINkr7Xl9GdKIi74g4nSLoKoVxd9LhIp/g7Le09ACmP0UF4OkNP+re
eAav79gkkgTGyhNqHLFOz7+Ea0oWlD9dvjrAMA0sSNaSPAlgnP142N9uPkAfNdZG
BWl3GiVTsQEOwj6chSxetBr4spn4i5lA/dd3vjoPmkf1TTjxLpJq1hUckf9mbfq/
AvsTiYpnwyIfKS8+wpHiExIqGqVV07/Pb2QTkWa6xkdLpspKKK42ADJJ0+VCeRCr
a6IR3vHn2vbzKq75plW6EcRiOBNpK5c0XySL9bDuKkC5k8QN2C9fwXitWPI3/0lJ
kcqFF/CNEsqGpVN19MYaPrDZAAvGiQjmxh+uvm0RKhZJzhKrHsjJ0k4Raypu20CW
ALMOrE2e84zx3xs0bR1E+SDh48I+Xc8qGARfzkdnZJt7uToKD78Z5wgVtsgTGsvy
UEEw5uGEJL5UYMG9xKGosDV2U/nka7fhyDi79B1BPb/SxVEp5YhKuY6TsSnJgF5B
+ZnleUtUMVCJt3GcQIQHpJ8AmuBWNiNHeOww9iKPCHO90LaPNwqBc4S132EbtTGO
uCdAglExXnwqV52KR6lzCMc1NbkQsyIrXVL9dzIomb5Y2bP0PiRScESr1w9qeDYZ
aOlb/jUXN/vwTt32RnFwOEGZDBbzoTzQFu3SFisOJDlk0mz9H5aOJ+HadQ6wpdw3
S7XUIzlkjgSMFT3CnWQl/OrrWfGBNcOH5uw4tytJ9GfPSvURJEOzS83dXD9Y6AbK
0iYE2OjjkZL9Q0HsyuneWCvWnT17PtP66jUCxSFVRmk2sIzuhZciVoXKmtxfweTe
ePxDsPhk7h8lHW4xRDGlO7Qve+3EgN6DJGikdhoAojfgiwR+yS3ZhH0MLlp57hUL
cllrCiyMDt1md9SA0B/tqtooKLeJaoo/uLgvh9UiLeF7xi1K0QOTyGOxiezuL8FY
U7fiibypqXXahDirFN4fjmXiDScYfMt2BZ4wclNOiaOeMQg3XTsPtDrQrPptzONj
0eFgIqaEWZO6wKG1dzHe6MyS7Ls38isDjGO0viBzGvnAjDzyAYUKu/APQtApMIeh
eYSVOH7haTu1aeU+BL6QmI0IMWdbfQVRkHmnXOEF2pttYRVF0pivgP2rSsrykrR8
c9H93UrvtVB5G0rgCYu2Zq3wsl2pFScJgdjpUQvtMSqD6mlAx4TT1h7bZzRMd7mK
FrvAJPIhM2mJglPaMhPLnhVd3x7B+nTMCB1KmC9CGq3O/gtPqPopAq8AA3cXKv+m
D3aX1j2+rQHFCGXMrUjtt2etbmT6kFNwT1bE3aGGuA/zd9zHtr1+H0ncBWWm8YGe
kiVAlEx2hgtUqT426l48y8z9XOmOCIgrssNgoSNHRbTW08YLMnLGkZpGY50ug/GI
DSfCqhui4MrhKiDy8EJRcglFLeiE08VRqHjNhT3pEgOeabXIZY5GqTLbH6nBUrYM
bdywH/64s8NQgmIgZfJ6FJa7JgAmOUod8Xfh7c9V5Bz1r9XEDO9hMbM6HQKEAr9T
HD0Ollh1i4kesfOSeZhbULtSieMvnjQcveTsKB/UqvxrW6TgyeguOmzFUJE0dCWV
0U6K4esjXl4pE1RyKgsqSjUAkLWrXLarNRrj3c/x3aetvCb2KvAdz4KzMMwNMvIF
unvgSYF1a+/slPxX2j2JLHo4juyrplXXGg10DtKAM3VHh2+2DmCDfoYQ0jyoeNcx
9cfjjV0F37hcnE4QlOeh4q3KOWWJsp1kwR9Inz7lzjy4RQTQECMNiZe8bcXz6hzZ
nfnjhhSN+dephnmybmhOL6jn72fKxA6/2l1kf11534VXIccLYLL2iM8eONm94ajt
Y2DmDwBk6TwgMeDikjgCh3vjdVlP7mljtox0ymUm5FJiwFZbEHcO1JWCVArx+0az
Rs/df3nih6RXAfbTv2sLuoBCerz6/d2ViODtn3sQC3/YT5YJRZGk4oYJfsncgvuM
tWO0gzGKwE+ArpcdEuksuEhuuuSfT9vOjP00nFkokXuMkjH6R77AA/ww7DugGERb
rJk8NjJ3TD+CohB9bbp3vVspVd6PLuqylW/SOXZZ/FBIP699cmc1WAt6a4wUyPST
VttzWKZG1Z1Aecx1WAZ/G2Bxrp+IvswHzpko9YVzxy42Zc/j0BF7iuERo2EC7h7h
g4op6E2KzwpMdCt5/uzAT14hm5waHrJtnXMVs9bjpiyrpj/j+Xte5sBgW+SfXsQ6
EZFhr6RGi4lpRKihk8xrX2rHPYwo92XWvNQRZhYhq1B26CTxV1UQcw7xFPTMW2hS
zr5F9O1qOst7cv+Lrh7WKevL/aFkWPU7PxKeXUcqGkvNtHnnfjvMO4ixHZw6utXF
81euV0sX8NcfonHY+4ye23G6pdV4xh528OFt2/h+71kzIe4Glp99gsc9B/NBrOyp
PvA18qx2AxTxfWv5RZewJho4P6vMGwLBXA2y/8GJhCv4clCs9yomTeGpC8pqMhbH
qyPHtvXYpHrTru/dSCkfQiTTQfr8Qf5mkwgX3VBNttGgRj63nA7AQOIS80b02+ed
xi2fmRipBKTS61dae41u0L7HRPE+mnO12bX04sOgbBRZ/KMK3JH2DBP9zdp+nbd0
4w6RPTabIF48MRtJVnNSkNKw8LCi011aryiwFHzlxAD2wHQBbHTLumKKCWgH7+v2
hSuuAQZlxD2o3ft5Nh4yDc59PhDTTn0k0ZdLdilGTejEXz5q3TQBjZNxnpnwaUld
5OU2bVagZ6SDot8rqqX1YetTW1t93n1FuiY2vEKxO3nbK8t4a91S3XA7wkzRzCrZ
r1sau6rDsOQx5wvmrZqb6V9T8Om5QYAf+YhsJmxgp1bYBj0WMBL7aiKpTfi8mwzz
ptiyCUafNonGeeuHX6IUSV+qGFDWZqnyTNDNYpLesc5EC/B2W5r2OVl0nSlm5z6S
Jrdog9U2mqsvcJuN+HVkAScsf3aICOiXJuebRlcwMhIPf9yqk4FTjzhiOAZmFpfW
B4TivbiP4HQW98F/EPU9oJ0ILoKchvaRAryyLx8lO66XcSlaXFuQEE/EBwq26lxB
afFpu7tlNTfMZ8QjgnjnHwFIVnOiUeYEv5QQNrd6nVQIhUO8KiqwVwSg6tQsUhmn
aLzUTS/T4LODfPnx5+q27Nm6AQblsFKPJS0PuInMQiQEQ86zICXEf/Gu8/ZM6Pro
LQSVrV9s57ODk84o4zNrsvFxujBo10yY/AAlf6J56t6sY7XXP2yNGBnblX2WZ3rt
svIlLBsdR2qO3cUoaZ9jYuFpn6fn1FBiG8/cfhXoovv7kLxpTStvE6IjYAu7mn82
psXZUP5+z1Xet3SgDUfL0KxJg10l2a4L0DcMRFlZkewsG6K8IGk+irqJMTFHWWTo
ae7IqjD80+lKxK6Ios+ykL9MrmiSgIs6hAUxQmR+xZw9+yByu+nXHQJgiPR3rgp9
HRBeptSTq8JA0M58ynO2EfL5o25BRtoQNNalHnBQcjS86gVNhFhklMI9AZ9XNYIv
hR8N3XyKHuWsepJkxnwGWFl9KhjJACVDT31as5cTSUCOvI+eTUMg07rfCPLT4QSA
RoUMeh97F5SFurFB3gKr1mkKMJbqoWwGkPlzEzHwzrlZtMp89WMBMG70pQMjGY+Y
NwetJI7Lk8nil2HW9a22QHVeeX9rBRNCqLYqZXFm5yDj6ryhB9KeAzXrhG355vB1
PTUstYIlWYu3XvBMWq2zDCyRdQLmMo0/je/51Qc74P9ljESzUSoLHkkpfmhutDMg
HoHEcbek2r+c4O3bdCMz6yO5P8daWV764FTfHZSYKyNqWX2sFfU2hL9pdA/Z5qBW
KQVgRtVXBiyuL0ZqqFv/eXBpKfM/VnIqorQr4lbrsJBOF3lCuk3m6ElDW0KpXANL
+/NT18hMy83Ul7gmTMM2Q3RkNMjwSOoZOsiJ/09+3Z6j8s3q0Ak35pRr4mKPayoZ
IaO0jIMEQdCcVzVY+a11WVcLCd5NvMVI5wrLNdSXHJQ008ucH1dOXidR6cijkBKn
Ktqqt7tNsFIBvjpkOKulBbT+z3hggEZbgZGfFjGxmnq3tabKwsnFL7Ph49Su8FBB
GaQKVxawJlchZeQJ0InfEbPdLel+l7dzF2G2OEordc6+G+6cwqkkuAdpJUjb4mxq
6XtOw8RtgtA+E9CHQC9y9Zm0NNsCpt636L/eeJ2vs4ZaMfuPYY7VH2RSIxDrDnbc
K1eCHBDz+TQBpCoDNHOs6pF137OpgJrZwNc3syUPd4VAyEWn/zFbYLwHRa4Tu7Wq
iFkfclDHatCVenmLwCFWgdFU6o0cYxyE82uEsJJ3SGNvyNnW6rb86Mdd+22AW63j
oSa9ZFDO5yuVDirPG7S5s0ZDV7ITZy8Sj1da49F9M/yCUtrM01PWL0iw2JL230kb
UkhIei+K7u5z8Rhr1uIhtT40Kkj3GdQKh+w5a5cQpPnNrgrr8jtXVQbJlTxc5QvX
qNvrx2u1HUaliUlEEx3D1Ar5bo/Fpu5f6N2xdeLMd8/xJ0aMmRJx920xzRPkgbBB
qyWybnWEtLjMEhXPIiWP4GWz0cGoWqXDBUi7tUnBE8aJ+fJEnXAMse/mXOA7edyE
ulAZBd0S80EBBmqaHheWdjjfvhSRB9vNuY+qO3foszCHSaZE0Eap3kN+5bDy/4Jb
XC5W+00qpQmdTLl9qEx6FL/mVg/L639hLP4GaDej1Oh7+FtrGe0Nrzvfm28nYd3q
KF+SaYfHvvq6D24EiD2jbhv9Y6BUR8+McibUj3BGk+9r1TZMTvF2Vy/PmarTIGk6
djh/KwVOqUNcjFXJsGJ9b3g5CsIFuhPA3E+orDtOtt++a8XY/e7p9ROS5LypUoqu
JUwxJPtdzzslmrJcUaSHTp78KcSB7+pnz2d1GsXwlVfkfj/2xeXALhjx/s1vaWyT
q7425rrauhDZzWBhmjA5lTnpmVmVtVdtu30gyHJkOFRYFudUJdcxc7Dx56Fho69O
DmLLpPPKJazJN8h9gZf8GvP2WRQCZ/BlTCg4fAloFAFsaXTFJK+2SphgrJamIQMh
Cd+g7j47eauxsxm3xGTR55wXRZqEFLal6QyrqvuWSwrI2AhWZEetJs/k3+nVGAue
ySFwVu/2G5IBGN69kOqAMxBRDpmOPKSa7c4BYqQCBSpuPMavp7vexQqInnDAnjcs
gOH2m/Wou0M06VEHku4kT+3qPtopuzY9sNW98saAugIXB2+Ag/Ex+2n5lm/CXnkU
ARc/GXOIP9jSEmtCj7DVHfA2LMLTYbwfLJVbhNUpXOTBEavnpQ0JLuhyfNtnjtQe
DYKQRTbPipDnSIDi1YlSahmNqXIK0omVBTbmYF6RMMUFHSvLdbwuznsbOnPHhD3X
tSl2a3tphhNrd+7BvfASbdLdT1yrMtpeUX1gKLcdA4pZfJ6jOtNxA5Ai0Rk7SPOV
eCR63AT303cSLHG0b+8hGrGOeo4crURlkRMjpUTlFBwSFCYDdR+h5yASxV8tg3lw
gDZBcK8lEra0eYkEYuOz/b3coBbJHRT+lvB45f9vMLlivzkrXX3cI2hTBGFgdmlQ
6P1VwOO/4n8ny3zRyI1pPVCtp9e+wOtrmQsf9cyrgHnKPT7IRvxthhochmo9N8eU
K7babCVfVADLxV7fp+kJDsIyG2BILvQtxsWtahhFlK9SpxCcRx/+hEsh8TjZ9rcn
voMz6+rwksVpnMry8gBEn3nxVOO0YLF4NG0FeCAGVOB3iScZtYT9EZyxtBqMp3sp
uv4HpIaEylhM93AOK0Z5Q1fBkteLQz1n615mGrhoO50agd7ezeKDT2lFWWX37Q2I
3LtIq12bDisa1KuAwNxwreJxtMEa/8TYZ5F9FluQsCEeWLz3ktNrYrxFziw9fWMP
TOayOvwCEvsaYhqUtRld4ZgHOq/sudv19PuMUHDYwdp8tnTwpOflpr7tKD0lrIEX
1XJHKRaT13EZ9FfNve3pcDIhFkptWYnRBQhUeA8giVKwr8hTy2bVYzPuPt/DSjoB
1lfvCLX4Xn7p31JLRW0gmmPZ4qxrMKifdGLp0/zqmSH11g/lrmBSBuH3mhq4NBcc
ff9JBlcgCj7zI8w+6LAowzCOd4ECVNrcy0PN8vjTLAOvA2a65x7wp6CGTN5TRUZI
ErW2pey414/5bun+uOi4Ur0W10QQwJ9Qhkp2h9YFswD1xFZ8B07j6kUyLfZx+fPk
jfxBOUDRrBBbPF0h0f6ngBMYyW7L1VaEOX97anJK8cMdoYG58tYCXxgPLgWTzuJ0
w1GjttZyGPl6qhiBabGN6bBn5TpPJd+iyhB6LSB3q7FPyClZgalM2vjwAmAE3IHU
+uBiHEYRmfkZoaCNfsZmLc82baVYnslaf6OoM6mUghAQH8PB9JIK3Hoy03WBaycA
76mT/0mxi4nC6o7m30sLYHzoCPmKuNDmyCJr0IhdpDtcnzBytZ31BRTLCaGv39Ry
x7r4igXWWAosHCk9iPVbbvMwtIxEOmjRtOQM+LRcGFsodW4vkOI3aRkib040bpK+
SqokhzfJ7G1OiPM5kA8LLeV3h3I9jNJQ1otDzsm+uOw903UGq88ZotuKzF6WcYrm
S32uVYdguMl+4JkTKRunYZzlalZEZ3Nuv3F5Xo/hCjs8x4XVXrMaoAhTe3aCPzQP
ff+4LUxCmuacCa8BHnra12ENZurFFi/QKY7zvNagos8KFRF+if3xJHGznf2ot9Ur
o72mYpC6WXM8uJJAE2PsCu5Me3DKvqpiaJ4aN1ImBz++cQmeOrXjd2HHG/R6+ng5
5LxiBKB6pPXrKHpLhd7qxr1qs5P1RXPqFNnG2cWlZpsRcfEe0vY1KHbcQK8tWFA+
2XCnSrzjohnppfo1V7yqGcw7hSIWhNp/TPFyFhlWZ0ELV8WXAWKGWdK/mvPAPoUh
r+5ZVapDXci1wsba8n0NQvR/yff6yOMhn8plrrbiHe1cDoG/iWrd0N72F3yzDFSs
TEBkVIftAYZ44cTYq/Uemlm4IZwgL/btL3mj7bz94xbFExyzMSTJyRrSXX4HVL9T
CP2OnfhdVPQd9qoUkkMB+HqamHfVg/8ZacrlGEc64iaSUKSLQRcjDTTaR6M+0q2K
E9D5hLHG/WsLQiwC7bCkOjJf0erN4KR/zUnK/+lSrzjrzDGBlw6287baFyh8yj07
Ei4QjLGYy9XpVBHhltRkBUzzkOhiH6igHeeYGzN9pJbEAwO/sXPDSbqFVf7zPuLY
U3KfW7tRC1MN9PNyBoolZKAcALq5T3tOs74eimyFHLuJaCVkc8Jq+A3JiV8FsUth
EDicLjjspxF0TfhJW4LihHxnwONP2d/pkprg7VjJt02A4ZWt/to0C/b1X2+fT9UB
ZSQ8+k1pYfjU0HstpypNa6hQcM3g1/RJTENXzKHLsKLwtVYMKDnUp/BfJc9AUaao
hVLM99G4QIXRRhapO7s/zMB0F5tVoxFWN+ltQzFVhbbDUWcsIrMX/X7TH/YuFF5M
n1u4zO2myIFgcATG+13FdjO2+INhPrkRaPjWZhoafKJs516sw6AAi1GI2r2j/VTS
al2o4rQxZArFpq9bzzxnbOS7RIhhan92/3fWlEIBMI+mXWCb3JjG03rTGXocEDvt
vK3NXZiUYkBWsuNWLCEZRtoT3Ak7Ocn6s686q+PJiTrJeJwHTES4nTmVbp/vx43J
M7L0fOaUgElqA/uhhrYnpfLkNvxgeF8ph9/xgnRDusQx+QLzFnptSc9abURmglnT
cO6gq6gauEO6olbvI7xh0NYAteSC8VPCMRASGSQNUQ6XyE3uoMZscNzVyHyaic9N
j/SyjCu69T64Eo61U8QdkKg9OnrmOEHU440NLEU3lhr5QpSPvxdr+mT9O3lmk3Lj
nnKzRKsKo7fcaPR4dnSuKVuvQrbSfdBPTr2AChoEzWN83QdmPyhlEEZuC/hbyEoX
kfnkCAI+EdT4yorBgl0DagRu1rSHXbrkAWOMRrO4dNLlhcxprUsU+JLN0apiIqFy
LM4Aj1Ns0aoQxworS+PAZjsemphJ+j3R1NqoWaE9jdevCU4b94R5g7nusoOa2e94
QXgYekKiph5WB7dxKoOdgBKOJ1ao4e99sYXmvDXVzXGYNludbTxCbe/pYQ7LJPLZ
IS/vGZ12tT0ff8IgnqPNHw==
`protect end_protected