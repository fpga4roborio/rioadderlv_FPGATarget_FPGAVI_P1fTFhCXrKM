`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
ddtXksX2+yylW5zu6QL2Lhnb2d1sD00763mmSITNX595NcHTEkwn0zB1Dry37fOW
FufOhVzEJp80NC5qZ/+F0Vk7Ik02dIR0elf3clrjeJRK85K4e3Hoo4xn7YbFUIms
l/8VZSb14+JVGURjfswrIyCUotIzlzVYZ6gzoZwDXIi5gQIBf/gI+KxNXPaKV+PQ
Ufys/12rjO6aI/pPlqSm0hCvftmBcnezN2hk1UeXgOIuKZnogjOsf0iJVX2aOOWE
6pD/psybjbnsNB6kH5uFTA5frkzIzkzl5d9+YDm9OyC+k84E83I/7/j+rk4L2dah
QJOvksSIzN867/4Qt8qYTQ==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="MvBXkzurAa5VTw+1JJ70nePUfoQXBvZOku/SMmg4TwQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
oRtzZL4VJ4iwysPsC8SXYCzXS8Fw2gtZTOskLcDV+1B9Nzn1zTyNtlo6lNICRmmK
ZRVu2BmCc2G+fmzynYlNTnSa7C0Cuel6FYpxCBlOuk3OF2tzAmLAuDyOH3Z1Yjzk
a0aHuoCdIRKv7BrZCdALt03JeUmXKPdOmIlkVGFl8yw=
`protect rights_digest_method = "sha256"
`protect end_toolblock="Jn9CQpRhJt4rnzZPRk+dOpzAubz7omckX1MrFd4p81o="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 5216 )
`protect data_block
gD6l00tciPUa6pDNTk/+t0OO0nC/UTtBwLB41d4inuAUA3i/ALrNyoJVcBnAmEQW
ptbcNp5fxEUJjnOxnedyZEuEBxWRieZFQnkRdF269oMgUfmURdWbVfXAn14WR8Uo
U6ofnMPARL0jOem8b82wqVfVmgKXmV9zpj+CM08GnFNQU5svZjg5dRo8i31z+liI
7ZVc1l228TIDi8AXbXSRCQTvSndPwdPorUWLWVVeF+mBQd2dCluzk5U7iKMG6bBu
CCQM7TN8EaEvMexMTBMXukqse3Gwmuq3BS1U0V8c8OfluKoJWj4zkd7TtpoN6Go3
4idAMe/TziwYoxtq1z7TIa4XM/rWwCJiHi5hSV+vDL2bAAiQ4fHgyg/+S/fJxOO/
rwOVj8+0QKhTMA6hmoKtwc/Z/6sa12QQgGyfC+euHS2vUc6Vb3FN2L/mS9LKHGr/
MN9aV1fhg1Q6mLEtHTpp+SAuMrbVIjpIZA2CYcZQL85k6Mjv6aG5uZ4HOdYYbDEC
UpRb50Ecd6C2jKy1gZYsl09/rEU77GAgAtLPD2wlfaT6gU0dYrA1FUBOD4tclT/I
XBMZu2WNMWLGMoazUPTgCArXZVcelgkB2yR7yg+oqrHvZRCXdfBDaue4wQ5z+qwD
pZmARltDHs5rLdxPtsBErIKrZwU04c3QCYzX8bVOPHn7FfVXDUCzW3P1/TUmlRZC
xvql3J+EqbKlzrSbLuNqZXDcQpultTdA6NRz3HA5Ox3OZoehl6MU+Fayu2XQoyBN
uIuLL5dHilnCtjpc8g91bzDE4h9t5aqzp6zqIzMECF+5Up9jW7eF7ZqbqMYIFACJ
emWH3sP/AIAuPLCyOl1QS0C/couwF3SoIipF6MTzrxjKJPpLIBIevDhb5aIgpJ9C
turVmsAYGJC7vAWxF7f8iIEkU7on+KY43NPsazqTTFAsAexQDtXyZvJsFbjbQ+Od
5MXL8pdLcmgJJrbUF7kiR2VMupE0DxZIlDQu+swn9PDj6d85GKynRxtOO7+Xm8SN
6yE+ZbHqXbWJGMDtwJkBqnND8u7Z4Ljgj8mThKoUl3lxgHMRsfpbICOq6Mnf9VeK
n46iid7DC4qBA3sCjNIUvO7Xca3U0tv3+/5qrHpbW8dnb9KaOYhvGnh5yapWgyts
nQlnDPHG1imX9gqHOpDtk1wQ00HGWQG12WA25sueVoL/04Q2Jowl4brCQs9zElrK
NmsE1OQ1XAUColySj+vzucmbQnNjaWm0t5IajunJbtbew0g3AsloQovVLVCpDCZY
KB0Gjh8uVyTy1lOXgw8lVUipTSo1nVfaFd3x/zq5hS/Kw5amBU6IaYW2GA07yI+m
x85ULjOgorVk5ypYFBP2B1SfvvueADJvdRUbloqg15u3WGYG+/T9VN9XKbuNEANj
Huwx9GWpPAJGLQFc/HEICvpK1nB0CacsJ2M0g3iAUBE+DWdN4yz9hjyvTJKi5WQs
YvWZFi+n9OTo4axiaqh4AZIrrA8Zm01xQQm9Ei86IsWJ4hZgFSNVkaKqcAyOG01I
4Q6kA99kiTPWPZXcocvZejqPFDjwyRVHhyqLN0GvhTZ8D8kBEQ9njDZVItSZG7BH
jlK0Tg54fzWfUYVA4CwaWj1VFbaAwPdHJFjE9Er/qHhNfy/gWU1Ey5g7o8EplEc6
yEBUC5VZ4y4KOLFLlQrfohpy4qOBnOBvqwctnch0XDnDmLsBbNCmHzBaCUf+y3aX
lg8At3KtlHlF5wTwA8/+LXixb2Eg6+2ltsqvNA+hZpaKgJsj5umRvSUhK0VzzaQ2
JjKojF0uXsdSUm7E/nnWRHlFKlSzXupMsVOYv9YCrc2cbM8EZIw3vtMdemta0DNM
t8/76RayIokhlP3sM/Yi7fposyw5fa+wKfQ0Bpc1RSvWpcdGwYB+K4OhjkPhHIWI
imhrt4yPDisoa+zQF5YjoM6+qLSqSTC4mxpgsXh49kjdvlF5eAbTzEgSC8wJD75N
NgXNOFVn0Dy4jZwNidojAIacZmD3TEV/zAu2YmeAckQhhQHRFs4cEqU5kOGmNhIY
GZ9zFsLSVBzLabWx5NZh5GcFAaYGuH+QJWlbrPgJMT3Vqa3e1E/Zw0N1bJcqCqn4
bIKr8o5SGEi5k2s/ZmLM3hNZMJ/FO27fOkhi4XNAP2RDGt6QZ3vbLrTFr9wq4DvL
f9gH/H/0x5w+ra111JxJqMkIQvBQUBhGr0U2MGfkQR0YgMFlquWpCQTDRzj7M7aX
kBY2V92WsrnOus7clmobm+gTwxqjNmIWDwUQp+R66OdzOofNbGe9TrdZlC0HxNg+
Aw+fIdIAgT0abWHRQqYnLxNE3oa4xNHfUTUpYT6gaDpXEcw0/t2cu96g2LHzxewS
EuKa/iFgDi7hf6vFeL8FwN+1kZn5TuiJDZb98sULdaCQXaFGJbmOjqE7K0uSm48E
TCRwqxzjrepqSZJg48nTgaIEtinIILGhQqKIhg+/wr5uzDcKoG0Cj/CumUIYPmLx
Ba3t88WMFDuArSPUAmeH7paSjMU458PDJfPlvtgErsxDzMXwlJHO78SF98vgk+Qq
aCVUq4eSvpvFLOV/tTGbWNu9FD0pg5O647dxnwhh2m5ekJIJf/x4ek38z9HwxDdn
t2cqOBmPy7Il3kTCHCjGoVDl2TDDbkU5OQ9VtUMWq+KXdAHmaNLcVYruEze6ekVr
vglFlHsjkmgPmUuLWZ4y7RRzOnmonyx1GjIIZEyJc7lUJSE9s6l1aVaxqSobUoF+
silAkdXP0XcvLUgyuJBla/nA/EIsxXeQKUMNpXVK0AkYKkS2stqLSGAaSXCBceoo
tJsv3mt7WtPzPHL2SrxV2cwCw9Pd0ig9su8ZrABe/S/ouJaO4mHrSXhgzjDz7q3H
4DNTlbq4PPdzUlCt6f36NC9rfLTAvwqxQuZADCoEbwT/inUinLTnY29tC+zSFq80
eXo30YzlQskYNquWg6+cqZvsZHHoMu+ICTyPnL+OHIrQdavImKaVrTFEGFN4b2H7
dPpIn0ZvKHJ2vtQh5RcRsK2tNiLXB0TbxEHzjtY6ssr6g3TomZMJhK7S7C0jJbkf
netUf3dnec34j/kBmBKxM2GtvO0N8t5RU8u4Rijm3Objntzx6RKJOPGgRdWD0R6+
yn0ny7S0ENPzurwjkCk+rPDUtGx8H0GhSSNxa4X+RYIWuDbPb1JuZDVB1UoU3sDZ
9DU1V/mxwdwznB3/4aGtQuI4RWyqJaVocCpWvJrwifESVJoXTkICQbHLzrqxNQzl
0jqg/TzGl2ZJitsQ9hT1+a4KSnfezlww2RDG41regM42oGK/Om+CRe3d90K4dyvH
DfHH41uojvsaGg2krVUiOCzNFISiHR7xh5ypip769soRZi3LRIFMkp70+kf8uzoW
VQkQ7s8L7bXYKI2K60DJoRIxAwLXFInGH4gSkPG/5P3WAw+kTfemBgTQMHzZi0My
RBDOjHA9aMcroBBG0EUxSYyQSV4/8Zz8t/NpWqWruYM2eYD/Pv5iBzAy8c10Efyi
dqGfKjG/YhJkjGo4xdgmmFESEsnCXozRuxd4lzwjeP7YnmLvvihb/DGAslATt+M/
ZPkYSV5Qp+LXucVNa33YtQYVpM3GzXmUjIdrTW2mt5swkdX+AwQWXTNRyWrREv4A
yBssUnCtsUOzZgwjoliTuhekxhIg00LakV91VRf83JP1/cU+AIMbb3aLipeXntjr
0moQ8Y0w5cTlkd1BFIBtqahZIuxz4krCAh/GiYxrfWShAJ6LAmkh65Iw/xH/l7GE
hVuiE0yDXjtzjuImn7FZuL30wCQXMxqVZkQ48pD3ufGa14Ccf9TUJL1oXnZb9u6C
ma4yCMzs3weLj1izvRrDFAjPhaUMBl7mWLYP8mDAfmTiIC9N9DU0QD0gwZswBC86
zBMK6CmGpo2/Ewc+0WnpdmxtcS5PKYcM9qq6El3fYVq5iiPI0/OxVv3VK31T9NSL
0WUbfSofH/mqZVwESsjChLL6gpXpTlNl4DGGoDOj65TxfXYvf6Df84IunPxbcugC
6jrOpA+X7u+6SDL/nZubAW9q1ew1Rt+tbfwONskibhXXbahWEMtSQBcqVQRH27XJ
qELDRfRXgrzwBgWVWUEhoRFJLY4GNmL5WzhEZiFV+cUO3vls8j+3YKY1eWzwsVSK
2Cuh+ds33yKxfoCbe9CTwte4QlLWEpHk6aDcxcEBj6EiACuQ08xguAZYe6XBY7S6
WNWquICq/EfaT25YtKn3oUptrYSu6q2yq6n4PF3u80xd1cqiknIJHh2SX7XkIXVH
niZmttw0XUIS4bQULZLPx9XkMQzEVn2XBn5pKJTHxmKL6BmSGzeF3FuhESAJDAfh
HWcjmITQIQpHWxwMAbtlIk/CPEpuTOG8mj76TYZnTFmpGn9Fra+MuqyLa2xzi0My
KU6+hFaB+jUC7OlnWEqwqrsZsePP0lpBwaLuwKpkT1G7di7euJMfFI/Ml1hh/45K
zfp0cwQa5peGeTcoefXpRCPhbHAFjzONuA4mHHrJhwfhWXHeG/WFZdBJTjmTJLDU
2dwcdP4bQVPR2xQnioNxdyL+i+C9Woj5mjZw7h/PP4JWxIBk7aqyiOD0oZmMdNaQ
Cxp832RvWqATFFqwegvvJNNLBgLZ4so/cKmLq+L0hGSUikeUzSMzSe+29FcBiBK/
Enznnb8XNAQv5B+JIVDw1Tfq7YCJn8wpLMLEzBncZLgFxJVa3Pje7aLTa+7VLNKo
eUijhGd+k4y8N0hqEh1xbIi4bUI9FOXW00+WAgXqf8MVcz6HQgDU6pSkyLCY5Bhn
/lMCC+if2+wcKfQuxWu83DBeVzozw8zlPw9gPA+qhYO3hAdw+R0CVQGAj/eIOKjC
csGkQ1uyE3uIq2EL34aAjTWx3iJY6yfXnzHT8MQqRKixIbtdavqWEmDf/dpPmh9B
IpPQaYh/Ft6D6aLYi3nAoSPYyScjxo0r13pUCmnUHY4KDcm0UhTJBI8xCWCfxRGq
Ss3vH5pwED8Bnxx6gs3BiH/W+SnNwxobTKfaKmhUKcVRL9SzIjS2vAklIwmpCfb1
wh5KdI8DlpLBdCQ+xgFJUdtn1/NEzCFivQJQ05CcChzeASFkR2nU+BMAMFRiyK0H
PgW6pv6zjborCA0vFNon6PyjMzQ3Htg8qT+5ERYiWI+Ji7D//Eu8nmytjS50xeVB
ELjcSf7KSpRTeE2Es1t7KOH5uWKIjGI+sE1mcHMH9137zxKGs6s1ilnls9i8Apm1
+394WYLXUML/5IbT3oYvOr6tMr6ggTMq56cCKY77P3iJZCI4CODxkukoMClGVQzk
tN5KeLCEN8TAUByuKRuTd93nbIH/6voCG/LcBrs9qKuUcw0Y+3sd5kbbe7YmlLJ7
c0DSGFeGm5qkhWZK6d7KBHSqQNWZebZplErAEZfNyOepfIGWM07MAblxQvXMirXG
F/DtkDzpIuBNlLI9bSNkz76RdFKS3W2cA6npXMuXQm02calUnkG2/lk0jLdVXTLc
u/jZajJ0QrkK160Z9k4fnpqbZbVcdlb8g4GmTa7oDFYwxZVgV5mv9Q3EEUkzTT9v
s7Wap5arPm//nTiVw4bxFwOn2RIUsvlcWYAvmL3J7kPVET3an9k+rA0Gu3i8tqDw
mYL9NLVbzD/N167KZ6TiYO/uTvaixK6ycHtlcKBTF4Q9QmFkCzRI0+B1+MWLX+gq
CR7Dymy1jzmWHhZhT63hS/Lj4v7pZKLVkxuMa/754UMHnat6aMRfBkmIIpy3ufgI
tccsZCpFKwA9t+rZ4ptJ/rEIm7wBwK0rAmVaSEN8iVha6bBwh3/O82nMQaZ0i5oU
EpIRUYd/vWojoPdTgHqK4tp1oLp3g/aFhnaKiPW9FbCpIEQ5lWoiHX1WagNuP0wJ
+Xc93+q9HZOPLefzKgTfvlRtmuMqe8uwU/xaQaHoyJZTgUnsMG0zpxjjDiQVb28z
AsSgpHAi4b+D/ljZZUY/s1cJb1iPak/c7JUljaoq5I2vl3u56mtiBjMyg+4jQytm
orkj60z0ZfMrGqUsTO59MlMqZGXx3OVBNjo8E/bf64wOpNtKCf+zuEQIgAu0S81I
jbSj47TrfegB+n+ux0RftK4uVcpKgOMjPIFw9GsHcAgIGixzovY3LHdHKVv5qyPM
sTamIXjBdwjYqt7a3qBoWmBh3FQ4EsTW33783n4BQWz55qaUursr69mzcIuTa3wE
E7b8W/EvwbCLWwyirhoxUvK8y36cGFGqYH600rChg5pF8ngsy0Aa9v2xjXUiLXyk
uxe85a3Dez0VSe8TD7kWlVK7h4dalpqK574Q+gt8oBQpQeLqDUZtSJShhZ1Qc+rZ
Z+v6StwugI7ta6mAqSvaBsv9iOAw5m6pMQkGh6jhCnDxfKrmVcBTI7/BHiSUNw/6
PQDHd42KlQxaarl/vYJA6iv52+wOAwI8CvhH6KbZ22qjNUmK2GaMXFY7GKYHusZO
JUzYS0gyewauW9cNri5M5PqQlBSZraK2D4K/IX/4z/AQczf5S6LhwD3OvBuHq5Uq
4g7Eb4qhJv7EWXE2XxN5tgFcGgQ9WAYA2C0d/wNc27qszOhmPS3P3v88SiB7tBSv
8bLA7lIMMSsVG0LstBgtCod+YBmaoDe4k/E5rYJWHSc6b5D1qULNYwdtz+ROuOFA
6JwnzGKHLlxVmZCySh92fb/nPLjuzRpgWVI7P8QtlkQ91u2h7J6KJU8Qk+UALRh6
lF0ixO+zC/LQtO1sGsH2vHJKjlqAhqPK17I+TU28hPcYml6ikLUl5+FyyvS1EB4t
uNM8apkj+HtZ+ism8MhJuwwjYENPoplwu8t3Ff15PH2ZNDAGU83JvApEPuBLdqmT
L+5DM3/dE43QX/MbVxnFkv13DlHAE9NLiVjcPMzbTqC+1GybGu91y12AoIdL0vqC
03AjWWN9Vh3UhQcYQRY300DzVyOte/JI0Dl793hkkdg=
`protect end_protected