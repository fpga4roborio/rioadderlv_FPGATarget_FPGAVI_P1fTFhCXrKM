`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
ddtXksX2+yylW5zu6QL2Lhnb2d1sD00763mmSITNX595NcHTEkwn0zB1Dry37fOW
FufOhVzEJp80NC5qZ/+F0Vk7Ik02dIR0elf3clrjeJRK85K4e3Hoo4xn7YbFUIms
l/8VZSb14+JVGURjfswrIyCUotIzlzVYZ6gzoZwDXIi5gQIBf/gI+KxNXPaKV+PQ
Ufys/12rjO6aI/pPlqSm0hCvftmBcnezN2hk1UeXgOIuKZnogjOsf0iJVX2aOOWE
6pD/psybjbnsNB6kH5uFTA5frkzIzkzl5d9+YDm9OyC+k84E83I/7/j+rk4L2dah
QJOvksSIzN867/4Qt8qYTQ==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="MvBXkzurAa5VTw+1JJ70nePUfoQXBvZOku/SMmg4TwQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
oRtzZL4VJ4iwysPsC8SXYCzXS8Fw2gtZTOskLcDV+1B9Nzn1zTyNtlo6lNICRmmK
ZRVu2BmCc2G+fmzynYlNTnSa7C0Cuel6FYpxCBlOuk3OF2tzAmLAuDyOH3Z1Yjzk
a0aHuoCdIRKv7BrZCdALt03JeUmXKPdOmIlkVGFl8yw=
`protect rights_digest_method = "sha256"
`protect end_toolblock="Jn9CQpRhJt4rnzZPRk+dOpzAubz7omckX1MrFd4p81o="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 5792 )
`protect data_block
gD6l00tciPUa6pDNTk/+tzLxvdHE2s3DQL3/JqqujQBC/Ei+vcAB8wM3doqg5vTg
mdfn9XB1bLOis2CVSfu295W2DNwHfMSTc/8BhCDRnTlLIX0UCJs9Za0+LoM0rMrV
T7EjVWppbP+Em6PkVKCwlmIQ7JKaifJ+Y+kjw9HCGboYo5074hY+K/CBbfsBQY86
AyoN0MKhsIx+eViNgnWjA1/QcH9yxb5NDX3k9oAK6bTLHYByTU74ABPyULkvp6zB
4vM754ayi0DX4XqlPZuFXbfxWprfSUZUMAcvVAQa56mU4FjWM9XR4Wxv37V8tJ0c
LsmjZmYZzhErpOiHD+Hts+LMl4tgQ8ObRnvavKxiO782iMC9aM3KmEuCSlZmqT3x
Kgkj7etMFgCW5Zew4/u09wBJP5Y/diAVwYWCK413GHvrvNArGIa65WWx9ais5A3t
rfAB6Xyf02YNxQyXl3slpe78x4dtWnaUQqTI4yWWFT8v0E/bwe1YYC2dLwAN9wEo
sgyenrjsZzCDGQRsVZnY79YCLPweyUdzOJRaRbMP+ZTZXrIXsKaYK82X6aVf4iJb
cwahjkM7PahhFDppEolgAYXQ5V4g3u9mstGk+2LSq08e54/4r9aRSGHdNxxhD+a7
4UDEVgNj68N4f5wFPzKm7VRfcW96d3eyprW2oUWXcd0H8SWJl0WyaS5KxzkaxZHs
ZuEk+zd1EAhb2czjG8q4WJtFHjdw5ftkL1byqu0bUaRyMoQObwG2yfObBl7gyziM
WzU+ucYvVlso8qqUblyOdjfNnXlyAFAwuCkQsTFhcKtZlTnDX91p+ad/36lmIIvt
Lfd/zWne8ArxYkrPExMOfUa0ZqhVw258mWOsmtXhOa07xa6qAj6ffBv2lrewlZhi
xkA4Q5D6AQc0TtAkqtgTeuN/v3EBvWMiWZob33HLsftalV1Z2N3bb6Ep+5Bf1M1P
MQsx7s8AE6n39/Y8IjLXtrSf1ItQaZkIY4my1V7mDPD2QH1DU/GiBcZUtkKcyvp9
HxU3J1ig/dKryMGYdBSFHUxibJU59PLUmjMXlUOk4J+LLGqfVahWygS0r21bO6jB
PQXccgzfu9P5yazacF7vyjlfqbOQhDZODF8S7vrstUMN8LmDYJuLlKSlASIlCg6S
OqHaMA+u0GqjTNNMQSqQ+iRazQNVBg5UBA0vs/6aS0Z4dAn/9k++sEzWntdx5eYJ
0RxG2ZZph29j/p3sAmog497++IOTm3ASm3ruZAS3E5YQBGQXGzM8zZfKqwQhlrNS
FRiQoCIXNWLTcu5ylkew7k+NHc3+HnHh1HKksS+kJwSgcgYzQVtW1EWOCCImWJXG
pUnCGdCTp5Zt8lZLKtVd5Xqk8FweP4/RDYAgX2KbzoX+p281JH7oGz9CylN5IAA/
eqoX04Anf8yvj20y+KnuZMStIbalP7MfZwyiG2+QpVmkq9/5DiuW2voVqLoE3QQT
V3pQFlkFQ00JkhVqODAyIaymllQCcqx5vPKDEeFnRF3GgeGd57mOpj9F+ck20JUL
ni2VoXDHuv5X200uk642HQ+H6MerVxVpc+zhSwUAMgmXEwd3Ail7Vp8wVqd7C0Km
Weqz4Vdq/FvQ2ylRW/f8PGu6qGvdFN8rLa5pbapvNyYv7YqRpV5WlXobtTCeilPw
WeGscI6rQHBaWfdtDlAxK/hwAiQmnQrTm1ffuuLiuTHUSNHzR0sd0m6r86NjFeyp
nEbLxwNiMVbFFfz5RNMv9vJ0Jz00+E4O1kI0qX5DoZK9G/dTuOLsPxGIVotVfV4d
CrGLIcLEZJp93rqLcau/j3CKMdLT1xMEh4dULATOpNn7JrjqCS2W3sk3TBsrfGSV
DSDi5ftWq2uokxRbXCYq1zTJKHdXqy3rnGwK1IA1yDUYHQY5WZ+d0F7/DVCK/tlw
BRZ6A5kbFT3VscdLH+c7pq7BoW9lhwjoSzaHL8i89t92z69KP5VFm1PXXbMocQH8
Ab5xIf0fDBHl6Pcea0ILzqb4DRjfIhDqn8hFOF/2Fvz5VJ/6k0dZkWWp6JmmP1GA
nj2Z/gQNNnwB2ELxF40okj44srfOJZOFALr7xtW9RqB5j65RO/Wn3eTJvLaYqKq2
hB/VNR5qqPRqpIl/sWY4fkL+lFzSeG3Hzn/9crZZqc+qAeq6IWc1AVTnn9+G7gS6
UAtksCpA+ufw/9F6/kmPFZdiSkkgzRSGClUj6q11xoVny2l8eA6MYD0TXBYEqXqC
xOI90iezGNDgfhyhVCVSf16RGujsv1mjQAkuv2/+57tP3yzfTblccQDWj6jxQyzZ
65/1uOXe037x82jr7LIbpReJjTUcFXZbBYlH1y85mzzL/PPjsH/LquPK/ILrnNDk
jpS8AjZoutbUgmgg70nFS3okozWGVhfJ/P4Ficuy14Cz7nikIeC+xuzKGyKwtvuo
Nj4xkhmjyAGcxOsszRA04iCnJDAP3o+kM9ofNA/3N7YEBAssYr3LyafkYhDRI1Nj
akAcBaIGfKHsk/1FmNeoksyc2LxMRhy1VxWl6+M/EgJbwXyIf5cmjV+jkHxa6xQ2
/ou8mdY0/zdRP5Y0fKxafuIecNnVJo52b8LOtQc5yjESXlzm1K1gE3VGDzxNgPx4
IcnrmCKQ+f6+D9hQn5rXKeecYB/vJdOJALyje/lVB2D+U2hZ4TIvBNloGhnVtnNG
axKM4QQZxYi7A2+11kJGgE2kjDAYkXAUEMx7Zvu9FavDtdvasSPirgOH1EtTJJwD
6U4srdiI9ZIf6YVSOp75Eo+Nx5McWIt9ZPBY/4A0joXZLIMZspy7Qqa/LmJaMti2
mBk6/q1F34aFW3k7kZm7Z174AKxVvm6k7LDJcTmCAGbvTf0+XKeLjha6DjNP9cRr
l8iTIyOeiydOjglKmc8w6bgyhBBVg01kx3gFZFoaNdL0s0IUf3PI3kFEHmx+jJiW
Gifn5wQAm8xvLFcKT7/GoCnlAxuXn0vGKI2Ynt2y74QZuRfJPOH4Ii9OxPrbzevj
fCrR46RpyJ8f6DK/+YsmNiIFdCH9bd5Hd3VkbZkWWH7tKoNJ1S8YlclrojU/rVUw
PBY8YNGvWWeaofjQYV7EhcswDEGn6U6lhh8FgcGpukjh+F7VvuvXnFDisGxF1woG
D4mhbLBC3Ew3alResjaahayC3NN+hclxGS6AyKKrF4EZK9mSyiUBxJhXd9lFQm7N
vJSs8u0Fw4QD7XrxxGeupOTIvuCOcTlK9wJRvhwALB2nKLNBw6napLnhshS/wNEo
xitDgRKnFJ33cV3vh5pEIb3DrXNAWDUN6dXWHE9hgJwRQQ5RV+3RcgAPPl3lgsc3
U8PY0y0syUH9cwfPhzI05PTo+9sAIKQNyjD0WITgjIJObtm867uESQ7ZpRkRggea
Zu1HgirBi5pmatr2MPd8738+OFfSEB3f499NkZidG6TynkhsyaNC8JhbwJnx/WjL
+ySkl/gmD+/g9ztjHKcBEjTOZHW5VoUxZ9hwNGUzp3NDrikDiR47yT4fQolYWYZ8
cJWLBB0fh9yCmCIYRRKThWwWxXgEc648JyoGWNukiPezzn0Bo7bX/uIUyAe58FWE
1tQeOoLBb+Ey37lwbDWARVCgHAscMzDydaccUAqjFDCzc7V5JRTcqUptYKrRpzQ2
ONlZkOT+4vpAccESxqFpAhhoGqdAg1u3F5qmER7kXCYgt5xwEmE3LMRcjqBo5bOT
f3IOh8LNbIKGuVAUmpr/HqPbQt7kjga/r0tp4gfHAd6zyUbAxydR61biMyNoQl6o
2ANgcI8RC91/PhSBZuzLLuJl/N6AB8uZLHrZo0K82tyNhCP+iKK71OTQKmDKfpoM
EmkQBzD8dYz3iZ83JgnDcIgGOPcp+zDOQ/zCINlRBcrUCTnSdBFOwtB99BE7/yr9
+9wlOp9BDOopz7HXCH8mGWVLnimF2iAxYDP/uvqjQ3B+MGHUoMGiAMPqTQLGFYrb
bmdCxsK2dsy/0PMkt6+yplSzolS52AhbDaCKbI5I0xRAR2eH6JHqLbEhUy29CPo5
ZegL53yFoSBjRUXUOu1ccjzaop6ZG0XkB3F8E4N96aiwGUNn91ygd9u78ykYDrON
YLC+YZYqRpQMB//YmxBCatkgZLUzk1Y82SXuCn/LR6r4FtC3P0WVRTGcdif+AskU
yPBjURag0XqXjlUr1+eag986rckJ9FVgD0e3wuXlJ3V5+T7fBa9vqB6wf2A2wUa2
Ijc3vGvwBBJmfjhEZ6Y01mcfOUzz8mk/EEx/tts2KhOKaTqBPJKOUJy3EIZPCD1v
8ldzssPSQ65/riQophBXbFu9MZEbS05he3liZLbqBL6PGtC3DugQWAjA0Jl3rF4t
o6bjkT4hog2+Ej3RiY3/72GBxNJqPfIzdhUEBdeZiPLY/PYZK7W7K7j9Si6onpUa
FYqbt42r0EuHq3BspD2ViOZNlIdxhZ45OItP+KfaotW4EbpsJGrGCtaupVmZsMU8
Mi0OLe2OFtvw3NFK7IGjEIQPio0tbOvipOyeZfIILwOpFFtZrQRd0pMnfefOmXf+
t/g+mjYus8l/3DAvyn4a074iHIMEU527b72iWRLrDdzlSz6434LQS0/w12VIsB6G
cVjsitu69Z/VyGiMeI6wQ9Pe+szH/jHjJrbQ0hmZvqTD6ojMzsCqeDzq94wFFch2
KpQ7fS/eyq6X8EZIoMkDgmFPzDlsQHQyxCz85EDQ9pH4TbHxgz0/yybRq3QVUg0u
CehH7Zi3gK5IXeYDoNQgpAU4vEHXdhypHsvHeI70AHOndlcLAsPltL5ZZsObflkZ
3EvVRIL6KxXQNWD8Iw6I9CzgCfk3PKE3tkY0i3mPGvFnQuExTcqHTLgLkRxmf8i/
o0nFgl1hlYh8NE3ZeX2S1zw42LxQe0nbtbidprdLXjn8S8RPxpMDGZZwCKbqwvAm
Wf7FK69N0eMRdqm/Zyuer/bhwMW8kGekJoZOTb9eYsqJ1u13lFMjU4GUAUgpM/hK
vpWAR8M3xTilE/J1XeN/Wu1R+unS1mRXOYiHOjDKzsLYx0zblBUgjxFehjwIiONp
WSyAJvBh2KypykcD8jDrJv8dycL9qVDy40a5tdcxMdNNrdVPEAhZkBXLH/86dakh
U9M9n73NWWF1hHIL/bPeEZ6/E8+84CHZe+JLLYVO9m/A3G2P8WzhFtEETwckbvTL
niKYH51QE7kfDd2WOsiuEAbdNthnVNsVv/J2brLrLu5OESt5FJXsbyp7hJ73qNDo
NbOEQlMnBXGWOlFqVqA2Mn473tWNiIhUQ6P204+zOdJ/wfBaocI+tQBBUJyOZLUm
vaNWxwkaCzQPZCrZWLumd+F2HpUdq3mFfvd+eYe+DBLp5yRrMcOsynKF4JwfPLos
IPk5HLrzWwkgWG9+HWZuzBzPk3zpbVKFeheGtUSiwYSPQTYKibawYedxdogg8A6x
RZCzjirrSFjyjVqOqp/IwtqNGOoyO9N1VLMQEYGFtKH5vEdFvTaep2JjOaNb963I
e9N2hKf0i6iWh1NQ2FXgZ6QamNII8NZkWvN+TOoqC/YjdeLM21yY8Qm8ABANHPcU
/vnVg0ZEuMAykzbA8QtHOsg9bTy3ZCQqDSc1H9/XBBSRg/UepmX4gZ2gCyY7I8Bz
g5Y5NTk4y9XjBOrM/wnlrgb5ZhcrnJECGjh7/eh9B2NaFQEmb0bYMcxCbUAQ5e0C
oMWK/KLdWMmyeqE2W93RzANOfO6+PPfjl4a6XJQwGz1ySXZHEO8H/KToXfJ1FR1d
/NB363TqZBKKlrnDGnUzZ7PVNm0JIi66OFcOvBakRLDTVefJZ8isY7FOP7YCnOf0
xCN5+BUIYUpKEo/9twO0vdDwABre7bSRUrQoWhbpHCA2olh2H59ltfTGL93NEuL5
g3MTCwX2+a3wlyrREuFXZHW5+0vaQs245y+mAxWrAxAyUy3UpKt/ss7LFGG1rSa3
CbMPfV+CIsUZ+CBcJebwdvOoAyINwBE/pXBRyu20gmGRaGsjJ9HvS1cpovrZgAn3
NIV+gN+39BJh0MwNDS8TwxOwKPIoVlEBw87qD0pF45rvbmSPYB4fjDwEqrq61YFX
8RrrIa0YZ9Sr+XnOP5H/gk/gDjR5Tu7TR8G3UJB3/5rbxHKTdl44y44HZj5Y2UN0
TaZwvcf4Ueb3BPfzaJIC76YoLn4mvjFwWQkkZdXNb9vqbFVt9yReYKRAoROwVXdr
cwKZroI+eYlu3RlE/FG14p+tjYfQFX44k3V0WUoKfWucoOYL4aLPESNPui5usoQ8
DhvZLEa3zXAEcdOeaKkf8m6jfpmORc5ERV3npNkN5PSZHsd2P5PErl7u3+elJkZx
zRuMRn6q0XyHFHFdB/+azx4Yl4KtlVB6h3k8hIrckGM1U98xYbYo3muA77OpRSDd
DkXZ9mh5Yd99tt9FCQIgGoBm7vKdq7TTCyvWiHfG430a3YnzSDCDQsFYl+WHwU3N
I9lmlFOcYv38O4GHzpXVPJzPPq8goo6Yshk/AvkROFsMudMHsN/fla5Uv+yCN97J
O6TvfNX6xwxxd1gthGjWOmdbHq/I8kei31nanYGVZ3AjVt5KZ/IZfazsiWfPIEMx
/xQ+eI2WkgCBa9qCdKW1tpr5A7IIiHQ0zs434bO5AG0+XJ7dyNoB/gh7QGRGC3yw
yGObXQPsv+t12NhrW/YE7U8b/DRIqyGsB76AwEYWUlKt6g679t/5eZWafUoLUan9
KHyYGh2By/pqY0D8TYhMlkwe63JEDi49ko7E5LnKV60JlDj6mdIsACCU5yerLk92
WerTC0dlim7u251pqHHMqPgaAUohwcZBZhh5SxnNdFtJVdY04D+J13rvXXI1imdS
5TnXlas5PT4d/vcMhUvKQla3qAMtdlVSkvxM1K+DFczfq54zrzD1dT69s89FpvLN
QyOlWi+S2Go2F7B8Qg5sQqGnTzsBqJR2lhazWBbH3oN61gCIGoh4m7ujMPaOP65e
xhVgtV3F/b1Pcvi7In6TzLSukbOgv76Bv62l92IH1hra6RFKgOeRkgCp8zjAaGnF
vAc/WbC7IsfplFPKVrdg3QHlniDYhYUL1TRT2nB+txUE7LBaKH1LXMdKzAleEMhE
u53v3fg/Oz6Jre4YH5GMMmJnRCQy+JMAxaeX0kYJz/Zyn896tnqjxuiAtMOZzFSP
ZqXx4GSMC/sV/rWt+wHzsu45rQw/hUbmeeC7cFjFMmAe7P38lEe37EAN+LJ+wHg8
ptGVEONhYUn9O9c+60r4heFflMrv/3eWucTxUeyD6f87fEUuc3UXKErFHre5NtJG
S+z+il0h33s+hetGmj7JSDC6/eMHn4XH+oGxH+FWYYLO5fTKYJYgp1OcZoVIEbKT
ZqLpDvtOJNIF/8NvNekzYwS9aGz+Y7V+25r0/R14SvtpBxZr1SyfzJtkmmHvzwvU
VR+XA+vxxcKre0apZ2Kwnovg6IyzCSMxIOIsFTDgGf4eBGYfjaq/gFPtKhPe5d/b
YJDNUwB/JNFRJEvOn34VrK3FqIyzGF++z5ruNrviZrHJH0O6gSSOAykiNcOD69Fb
RaoNSC0QqkFTO18nP6BsEXAWUkdD+RWWM6kdk0nx4vuQbHpdhcV1HvIxwIpvFBfH
+3QOQmqDe//gkBBp6Dc0tX+v24bM8OKRLfgmoX9GE+PvJUQBUnssDXyy7DuMyelD
v8S+kEbYZxJ3p3300CNIrnvfZlB04f3OkRZpBHs17lY=
`protect end_protected