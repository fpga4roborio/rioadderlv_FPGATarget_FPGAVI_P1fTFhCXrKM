`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
ddtXksX2+yylW5zu6QL2Lhnb2d1sD00763mmSITNX595NcHTEkwn0zB1Dry37fOW
FufOhVzEJp80NC5qZ/+F0Vk7Ik02dIR0elf3clrjeJRK85K4e3Hoo4xn7YbFUIms
l/8VZSb14+JVGURjfswrIyCUotIzlzVYZ6gzoZwDXIi5gQIBf/gI+KxNXPaKV+PQ
Ufys/12rjO6aI/pPlqSm0hCvftmBcnezN2hk1UeXgOIuKZnogjOsf0iJVX2aOOWE
6pD/psybjbnsNB6kH5uFTA5frkzIzkzl5d9+YDm9OyC+k84E83I/7/j+rk4L2dah
QJOvksSIzN867/4Qt8qYTQ==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="MvBXkzurAa5VTw+1JJ70nePUfoQXBvZOku/SMmg4TwQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
oRtzZL4VJ4iwysPsC8SXYCzXS8Fw2gtZTOskLcDV+1B9Nzn1zTyNtlo6lNICRmmK
ZRVu2BmCc2G+fmzynYlNTnSa7C0Cuel6FYpxCBlOuk3OF2tzAmLAuDyOH3Z1Yjzk
a0aHuoCdIRKv7BrZCdALt03JeUmXKPdOmIlkVGFl8yw=
`protect rights_digest_method = "sha256"
`protect end_toolblock="Jn9CQpRhJt4rnzZPRk+dOpzAubz7omckX1MrFd4p81o="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 7168 )
`protect data_block
gD6l00tciPUa6pDNTk/+t0OO0nC/UTtBwLB41d4inuAUA3i/ALrNyoJVcBnAmEQW
ptbcNp5fxEUJjnOxnedyZEuEBxWRieZFQnkRdF269oOvEbEWFjTJI8OIXaAzBL/l
vXZzIKlqgYJHxZFv/GOuhbcrJLRip7rVtUe+3hlSfPOPLtabqVmdv4mCbjaoNwAu
iE13rXtGtYbkdwy8CRU5s7nrmywGNdBEssvUE2OfjIKpPSV/1BDpB/Br8Cx3ZfMG
wgCeWCn30OeNF4f4lcRzHGHQFAVleBB0+KWcpJB0+LJep3srhoumD6Y8X9lBoxym
x8C0cPdY63JoAzfCyw9+eD/dpqCg83pgnkdV9utRX7WVs9N9NFv2xbgZCZapMZ8O
+sE7BmlzXQxvbPhVcrYZmgmZisPQEXNT1CymFDLMsHfEWuVI0cL3FL3dfkF4scfn
H0uPwmRCU0S0H/0Ih/X1GGx8Au5qO2LYsAMKOF91Vr6wFLFb4q60dNuqeUWOsuND
abzuYdUORYRr86IAI5OYL2kNwDWG6WtEIRzPkE8tUIvLmkBHj456DSA6KJAyWKVB
0GUKydIRfERYee1giyG+y30H4M0SLwyjgSRSqbpBvR7qyVpVMcDyLJH873Wo8pHa
Tcr+mZeMvMuX3mn2JeH6QSCUP+wSifAYgycWrQf3PcujKIvO6uw1JFajq7M+GYih
Mq0GYq43K31zcfO1XaZmUbgdVAV3rUOlvhUKUIWR9YaLqs4V7WHCss2SYUEFWQUb
3OxQUjdUYsOVUWumKmNi5MDbaRF2jHLuBJ/GnLzvqMpkcJg4Ddohc/KIic4ASDej
NcZ5eqGn6vWvUZNm9d7Imows5a9bClU3Jr0wlMLb8X8N2IuFBTe3S44ccC6Smy7a
bHViXV0ihL6lVPb/OIqSTIeEvK1l1rit5M4+FsN4Ugx8v5VsU0m/enVyhzMyohGv
drg7MKIrhspbTJju2wx4FPKBAMZhuQ121FB+pSi41RKFEUYlUGmIOxsaeyrW4fb+
sm5Y5GOcfqRNZLfzorFSIyARpOE0sqq+6URlrCNu/hRZcbsDrJN1xg0o/XY5meRK
V9KMA7YC43aYPr9gnohzOomXvuiDWt17IQzrzW+nGxfeu+2gj7pqb5V/z8ynRb3O
ShOJOo1jcXyADagrI+FG7hIGc3Q+GxRk/4yAoYNcbDxJQU9xOjFqXL9FXFbpn75P
dIbQ8fWQuzDFKWyLy3tdi3yFjKS+x/Y7sAiY4YkWcSgQ7HCu7PJkzdQoWeAU+lnL
mCRR5k1s0c4I+v6+uW5D+jWmnEBCZTQYNaNCUDKRAZcRHKnshB3tKU+H0XeWXfUR
ijrcvtrq+vF16AZPDO4KgsYtdnC4NSZwwZM9Qm1MIgK7H7DmF4qgHMjxXYgzLJj5
jvihPs9wI6+4XRO1nLSJjHQMktF1IV6B7a48HREcat1lAMP2AGzK0xngFrx3NRra
YTnBLmKb/RGnRy7zvEwjJNov434eGsOhJwVEoUMLkNbnE7c3cjlqPQt20JMofQ2Z
ieL00MELw6SF/MAH0bgWDG3Z7XcG7u9YKNzdFspzNUMAg4j7x7DADNfLdbT6G1jI
ROaDLQ3vqNAfml6W+EW8g5Zx88sZjyvsQGQjODE2idK2ElMUjRFVIx6tjA2bzM2z
ec3QHxgHwtdz7ajPe91pMU+bzTjX4JBbwShSz9dsvReeJgmk/irR3RwjMjTAj5ra
+dnU377SxFBfJO5GsHQM3lWRrp43uee6lYmU1tYuEjRD2RFMiacd0e9RK2Ck71ns
HUAw7bxwK5KPkvHWKfV2LeFEIQfxA5BmaL3+BEtZksV+VLZpsqQE2vK16U7wFUjO
T+J+tWQI6YgOIulwhKIhkhHUTBRWR8mv5+zO3uAEUsPLuwecBGvLc6SXnpnPiTKj
4MWDvpkG6BAdSTU0Ri6bGpPhUSm2ERCS0diVnE790apMncG7+7FTBpnGELrrs1cK
bKk8ZJGxw/U7JuTmpgd+2NcuHo0t6p5/bqrQirhptrNiaN6e88B7aCmIEPR9TQnv
ZeBZx7z+MDS6TUQQuxL92ez0DlzQkuOlnKrla1h+bLpk77ShoVwCaApuWn0rW8cg
ygxb8vTc4HeNwcnLpIxonyofqOF6PCbh4Oakz94b6VTxmeWf6iEfObFvUv+5Gc3a
rFWQKW+c2vdk2nPaN3dLNG7UnnG8y2EfkTUiQnGGZkWh7pA+nobcvyBhaDlS5LHz
BxXWF38AA1+XVkS9qVDWQf1O2txoU4K3APqN9UOFHFp3qGt7lhyPx3TKPzfKnex5
BtnK1ZBCqH/enFJIz1MWAmPOEuAUd4O9uDrCVVzQBh/8dgIuOCx2vk0cYmIEoaMi
41NS03axk+a8iyQ0W4wc9lsTjFyEAHth2hbYIOu8m7tjfvmseDdQxGIPbX3HU8vb
fN13GlyBhGH2cqIlrcw5WshPhL2ecUYB6Z9NQdzHbC5QqmgLGncVBHzq6lJDKg3Y
xcSveT0sb9v4YjSJWIedVXjWqrMCXcppRlFTLSfitUX2yKb3ZDojiJxK+oxpAeWc
kvUmMkjbA02NLKheaGEcq40NScvQKx+DFCmeGc3I9+fOmoiN64u5/WRorWkst5jm
veHLJaXx3V5IZTMOD664C5V4bK9yTCuwnAaBNLhhlIjY+kfJcKz3C5VOXb6uw7Qc
r2ksJDQL2NtStJ8yh8YwXwprfh3z2zMQWOC+1SbmRT6fwNGS82gY2Y3PgsLeJCGO
3vUGwbdUwn15FBbZbYZrqCNVin86RpO88249SGDzV+kHqPw9145n8tzoeZjolDmW
SqUk/NSr9US0unt+AjrlNqgRNheATb+/ovAnj0NFYjvkf3SRkdGwgzZEi8RIj5h3
mRNdPGN1mLoZTvP9/jNELzfaKzPGmuegPWvQPdRDaZmh4BpeSdHpMhiU/+pm0oNy
2zxpja13sEJl0/mI3D+Il9emVXrIayG2DVp5D5C0pCTd8c/HYMm+jC1iUyHfdRca
MXo3A6bWaJR4VGyGWT6jPDaVmdxP4aXnR3lsIlXD0gDURuIS3aOTDUdRrWQV3gfk
kvv8MxvGydCCMuajxnWFJF1/gYPpkK1x3eE9CyUQe1DCS6UP8ujtebaFk+w1Y870
3EuXyZNC5VnH67GuHl3ptveCfcSx64SAOoqAeJGtPkZ4KErREChpRPnVe/x2GWpy
WK6IE90uAM5cCaKPr3QtszHrHcbBe7Q+20fUP2jMFMbP8OeZLxtP4eIoDuSNkisU
AlmTP+Y4rj1UpTol45+vs19U3+W/87dI+1dvxtUFCi1jmpHyWRbPK82jKW9k/VaV
A7TwWKF49LfoHEOcCufIP/egU316HvLndh9whCXinMmZEaeo3INq3yRlmydom3sr
EkIR1nprfmb0PLtqpORYromsFTHUNTXoc9PHoFgDxXxbZ7dgNltDD2t1SaKeIiVQ
GCgz3GIWjN1dBLfS+xZvCVgsB+sMWkzyKHlGIdjEaGfv1Eo+0f9MLR/v/Km+tbWI
6CTQm1nx3g3XI7DDgFkMgWs+tnJ3QcP05H60hCXII8XcOAV6DjBnQyrIH/enNjNJ
S5lcoImgyLJg5SERLcm+yjD8y2+Kn41ufLrYYNRMIf31WEhYUKkWMmxUEG+Vru3F
4TPHc3U4/aY55teLhG4r4aFYMllXO+dkkAo/096+Sg/bud5+GBnitmqGc0IWrj7G
IAbEA+5Qt8JJ2Fb0CFQYlgsoRtY2M7Dl+x/mDWt7qAJ7c4pnYVpmeUuY+tzXBL0e
A2zyTrqxnpXWDjuPi6ZZ/N1psD6sktTgo85Ear10Bo3CLPaz55U39vWuDUmjB13c
esNgFSvLa4oHSdGlYojbdHQM5eQy01Cu9W7mAmC/xzs0a4Q6EEn2SPDCsW4U8J9V
Vj0u1dvOOvC7XyBA8HZmZwzDmeOCGc6NCSTbw2Y+/+DCklZC7HEeHAg0zJylhaeH
L6adPvDNdLmmF6uNJ+XWx2Uv0EcxmFKtjhzqLbetlkiEeaDx+OW1X52nUmyIo+Wa
+cVUCEwkrfQQ97Rsb0iBkcAQn+mWj+I0JcwLVqr0rMymvrSf/pi3BogwqFuProbl
puN8dFISQUt7n0W4mMDdiQ0ZOLR/2DF64E50qRf4mZEHToGFf/42fpVBCxrhJ7EL
P6o4uUWm2GNMR+JOtc7Tl0Pl37IgnSI4Gj3w7PV3LiKK0dlnXFOdylQXNOKxN4QL
d7IFegmI+abDfDcz6bU1NU/y3eS51N3SA8zcAvKk3+Qb/whM9u7vsnDg704aC8lY
ZPSWNGbygfK0y7WIZi5N/u4SjqkNSAAQIpOhatM5U7/leA+HdGAehQqB194rMXpS
rIdIUl+XhJ1MWo2TQS5cJ4mJ57pXIScX7Q55xNMgWDlObRirWq1sdVAh7pqkuLkJ
Rwb+7AAlVsylDNlhUWKqsSWDRhkGfWjrpPClQkL6jyYae6SBrzLHAdyCHUFXDaFS
+G2/anEZBMlHdn/kPa0XGN5bfldGIHcBIlZji9AzIWeN5hgx47qE3B/T8KDbVXIT
xbo6KL9+tK1QJzR24bGP/rjdbHwp2JOWdMEKUychoxDQAJc7QTgtzfeG1hvFYpbJ
P1UvY/n4dyNb1mip+xVmJspc5eLV3pflBSBxNomuYrtAvL0j5BTLR/hubkCIzotI
Iv4HgjDPbWIRCVnxMYr7/ig0ia2bShj1Y3qdPO9G83/OgXT0RUboEjoLy3G6n7zF
4R4CIbJtg5NGdo81m6LQF7+xCnPw7WB7HMOhmvGAawTbjvD+h1EDjx/k/0KAGXLy
XX33xCXfEwYgnwTqxfE7aqo9JCnNc7jrJbpFGVFhHqPAAZXbuGm1rqHHrtaPKDWi
sF5a05r4LeG74SCZx+wVEaug8jVJ3IKWbqmtDS2uqNskf4N9a8+HbTfOBrBeZXEj
iJcgZdtZ0zR86vfaZHoQplBYhybrYT1iPuG4zGjvZF6ygTrqVcdM6mKmOz58D0m4
o301na7qgA9W1olJt1E9ReRUPaiWpNn1XMe96z54BdQKjUiiWX2fm5xABvNWMPm2
dGO3//y0cV1v3NnJWB5yDUZaVGzKvlt4rSey1wVYnmNI5g3W6AImTm9wHGqeqY1t
GTaET7hcQWwXf+LmbmTciPcxE7Ej/+FoE2DoXQbwgM6Cp12nimDrYtoPDKB5B+IN
wnu0dWGZnXSDZG13l0MUtUmip/4CQ+frrndfOQ9iNCrILeEimly+ZFJqcK7UzQnj
TPiSt56KTxZQ7BaUXdOgrWyhfWGPpgUkXE7HsWHQ9B+BmxHs+/TA2J4GJMnDz10q
LtoQgZOasSCk36X1vtecG0ZES4wMs1hY5SKURqyFRcrBuaBNzvRcY7Ckd+6Rr480
QG9xYHO53Ui1HV8/5Ga7a9njsD0Zd1wB7/JdmD2IC3THNVjOKdYiWM08rG5KJFPe
HYjAaZ452TBiavnM9PY1WcAoy/50WCF+WGDBWAtJcT02Upi/uv27xv7GDEtDIkLw
kAIhcdKRim7s4tNlEnBcoXYJ4RSmJX0qpHt53PiPMbDQ1XL6Nj4TJ/F3zuqgMXzG
w6ZOXHZ7JJG3ZOQnm/8eEGefoQe5PwbRxzkxHfK9mmcm12/z6/+psFnKvQORAkmF
Zbh34T3dcLJz2cycd5oGcS8u0FKaUAcLEJ7YNobF09PExniyq8Yk5wsFEqnHIDIK
Wp8oXtzK2CnJ8YGopEj9excLqU8Fw+3CTy8XmTQ9KP5jAZpCQmKGa6fi8o5zDrgt
eZvZ22T0l+XbDQAI090B0uIbSOPBwRpIoru7xFTKwFtiemH+9nSwHdEKGtn4DZU/
foLsG/rp3GKdWa67V0QG6phbd610e1sWh69QIa9pcZYeTkwj/902snF8zmpY1QUT
TxX1tGOIHw00yoc+GWJujtVvLdxzeNgSOcxr+7yoYKwFrmJMMtWZYCx3VujJmQI9
SLMku2/97T1V3M2VMqJHhF/ehtsnGDwfmaxlnjT07CtDjb3jaGGfe2wwUYCMwgWe
/4EZ+KoXHVf17xVFyxEOVQ99AnJUJLUgw3ICcpy+wEWCq+qkcIaILWhZw+kVh97m
WBOiCFLX8QuYPZxEtBiUFA9ih744lEfSDadsW5ApaXxMBrNh7GY9K/n200GYD8Kd
eniVsNAi3lE3Sdx+zS3rIQzyL06HhayyBqZe0+drST5CQhF1KJ1Q6sPEyKRMCsGo
FZ+NWVGgkE4XUERNwKVCmlI2iPwDAwxQVG2fPUDV+TVju/hpSfzjwfG7bTDEh1HS
rM/ES6RcBfG5kV0lITv+Mvb81UTa2Jk/p3AAOGM5ea5VPXIurH9FeJsneDbMo+Fi
1BpnAt9JB6kBUhHOJrCv5EWzOBSuKSAsuTiWuGrMRMWwZb0fpC1SmFq8gaL20R0d
iBbncCJWTH19nLTmt99NXmeq71VrJAb2RoSvqKsX8PZ556RuYP5CLxlmvDUCxEuX
foRTObNvFDhuDJuJUOcxkPBYLL4kfN5xLSfX+rzUg7/upmHHxg/enuVPAO+GPHkT
Jz8Bx25q/N6IvTSKfMpb8Djp/AMZECYoT2KZaIwkM6mtL8HoGkGShD5igGc6ajpi
oHvMMqOPLc2RmgZivXbdyTPXqmWYBwft0jtMHFSuMqVS4eZwiNKcvbQe7PjlIbQZ
cxl8hZnaMgDYGL2ukgZWYE8aX62e4qzqJi6wReD2lELVCi8ELRSzOTrazZ32z1h/
fpWoKPxvW22q6dAr+ZeJZ0q4py8IgMxriwGIUl83wWb/VuuqQpa4bNaKFAsduKge
dBbwpiyi7JKrx1ZKHiIKOncobZQ8auJSOzJM34dYSS1twnk9B66bQPuqTo+Jy2D6
xLSM7Ns9efaLtk1hqOESf65OEitk37k6pvBUK9q+oovee4CghJgsa8dvYS/EoEW/
Y6bdeASxrkrYPuYsL43cOOevfDkuTaGkR2+rAnYqRp1iCpBu+2B2sujk1N4Vt2ta
PdKwn8NTeUUxYjmKPJS2Thv/n/WVaxz84ULkbvJN1bFU4s1D0bvQumtmdRyCS4wR
/Y1m7yI+D6PFn9wWTYAJ51zn83cVuCNyo9szUu8ZQq23i30snxqkocz68/d5CfPP
rQXsZwi/aT56Hc/fVHjVZBu6xEUqAB3ET+o86EXSgkkoJSqB2bmnC+V/9YPknxpw
cyF2VzhW/7ZtipsJjgWlNVVtwllZ6cAGAk2J/+w/EvBv/RkhcfiLqFMGTokh3ZNg
dH2a6CTzPOQT9YkZOTZPzdzQp0uT4alffASu/cn7gc6PG/CvzeDe2SED7G0GBCeq
MVzETHWpzz+1bzT7jm5lOXyBEV6ZkscCFV9DmZqcjwKUbBtPPDhYqDv0MplEIOeR
8mGLiOmnPW8etG/oOtl4Qnx6zJj3VfU91z2gQmwoXHy4Pfy3RHovwsTUAH/ZYvMv
idBOTowD+DWSTCZYCYizo3IwhEyAj4WdORSDKu3a0DiEG49YcMoGI0VBE6M46TGY
fOlWzWDpIAVRw3eP0uHzzrzOzQdr8qbJyf+H5XodViHho8TzGu5iRA9VSEgsJZwv
vxRyO09AVOX/bslQxpk6qy7LNl+lBJknkU8Haca4Ls2IXMN0g9byFG5cs2wZatuH
vaWDccjQDYlpw/fxC4vmYvBr1WhZXkkCMbEN0xskesw+F9/PwA02ukWDkV7uVIkq
6p5vs07Yo/z72hKLGzFrbZU1s3KZbFJmWwnKU1dIeEB47avxb5qP/q0yJEUQaA/h
YZ9yW4tIFL9l5ZKln7QVr7U7Ci02GLnOjXC6IzQTFwTKslyqPWRZ+5D5Ig3LBc+f
tTphbl/MRYRc5G+hC+my55EhyPNSsWowIvvNZSOLKxkQfW+kawWPNSg2PYKSX+AV
TEKL/G6fdrNxnFc+vnmbmozZvI2gsckPjdQPqGARcuWezr2mgjnIZne97kYJQZQG
Lv8K+dcfLJTb3yERMHJkkSGYkdWPmA37CQRZxEmr40e9386rHMv18h+KlN298sRd
crb1VE6VYpmMRXIhzLYqicz1jANulNH8WGb3cG8yEnZYqvLcdhRGSFiaZfSqpdLB
kgYTnNS5JEilZUJRANrCXa+ZDRYG3d9ZaS4AhXaJRi4D0Cxj/XfAYmuKaTsjMTac
CsV9R6HchMGnEkEz0Dr38JYTercmKVG9FWsl6gGP3PfqnhfjCpjIpJ3DhcuK5BVL
YAVF9TY41P0Spiotp54AOFY+UECP33Y4AQH+dhqjfZvvWm4g65xiHAe2//zfV7Zd
8+o5aCiWaIbN827cA99RSZzjM+QiIBM7CzPn8QtaXyzmdjzEtmOUcqHrwEhKtDlO
vwSb9pAMVWzKvvVSGtRbw0UTbr++X8fAvTUxt281BqyqoO+n/tDbJjvM29O0oruB
1uod7fi/5nYmLVGiqAnOzwl4lEgn+siEVnNoZNZ+t1kxnG2xQIWIunEhgkP/Zl3h
cvdfOhvp2qSLh55kmHTO9KBVgDgq8LR/0sAX+TP0GRoVVkbbzkxcugdXnfFSB0Ql
R73Oxd7dUc7UcySq7iyyIEhJDDw29GixLP0XMeR1l06snAb4WaeahS7VDOBZeDcn
+zQT6EZQ0pbsVV1GtoDBAzDaob6+l6zqlXB/OILHWHUw78GoWzl0EsRUgn2crjYs
CLht69mm6KHWDw+xy6pMR4zzxg95bgkCNT9NkhsC06Qdw3r/d4vQ2gUiIY+LARHm
58b9dTttfHkfUe5tXFrdgtBhEMkjetqt4yxeX5+Q2i1C8gZcI8kRVcTB11WBukk/
WkqZebK+WU704CsKdIJLakknFuvLdlSdVoPsGXlAyVPknuPHNQZS/oYxZVgY/94M
4/0ia/Efh4JdLPHlfOFOQM6/Z9jsWodKuPz0pRWtTq813Z50DW+5GI5XhC25aEjE
pu/cbteDBzhHpWQbTKxVj86tM/iT3s8684e2KYDH3M4/2VNAcqySEDX0tmk+hzNf
MDi4SFQO2hMJTEH8K2xeoz65Vum/vtudtyfLb53uDTaWIF57fnRJAVJhXQEZpbW2
ljFLN6P42vpzayQrHhUgflMs6cBtr5BfU1rJzDp6fq3otvwEMLs6OPxQeyKAOyDw
gmK+zEwADK0avR/RaDMVpW1zYKbfWXCFgl7M2UML2wXhZKJflc+l7FWrb/TH5IwU
nYXSnSIeHKy2c9vpOwFm8Tn5fpJlYhAfSwDaFi+kEQM+8dnMP3LZ0mzp/GFE5S4M
yaCh+Dw7Ua4sBEO+lKuE7qaeRwgVh9yRGqTQkYr5GtdJRDLo0Oc+M0ytxg2X6Jq8
OPVaI8ODizhXX67V9Yp3M55NBYtYsPUdPcJo7icPY6TLdfiZg1g2gkX8bjbYLvNJ
l7apyOHjxW+61ZNI8l4puAiAchHkn8eWXgRmbm3XDaKoDp77ieiYKNJkh7gfoMbo
3H0sEln6dsJA7pW2HZNfu2VeLaSTtx8ilCmxEQSIVuB6IN+yU8m3QwBWI3/BbapL
+V0p46hju2sY3lwXt7bUtmvek7l84VCWsou8neN238KmbzGKKl0gJ8RBYLQs9COT
XFLm9d3Sc0rSt7q7+dwJUQ==
`protect end_protected