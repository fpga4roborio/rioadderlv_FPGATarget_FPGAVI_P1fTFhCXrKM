`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
ddtXksX2+yylW5zu6QL2Lhnb2d1sD00763mmSITNX595NcHTEkwn0zB1Dry37fOW
FufOhVzEJp80NC5qZ/+F0Vk7Ik02dIR0elf3clrjeJRK85K4e3Hoo4xn7YbFUIms
l/8VZSb14+JVGURjfswrIyCUotIzlzVYZ6gzoZwDXIi5gQIBf/gI+KxNXPaKV+PQ
Ufys/12rjO6aI/pPlqSm0hCvftmBcnezN2hk1UeXgOIuKZnogjOsf0iJVX2aOOWE
6pD/psybjbnsNB6kH5uFTA5frkzIzkzl5d9+YDm9OyC+k84E83I/7/j+rk4L2dah
QJOvksSIzN867/4Qt8qYTQ==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="MvBXkzurAa5VTw+1JJ70nePUfoQXBvZOku/SMmg4TwQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
oRtzZL4VJ4iwysPsC8SXYCzXS8Fw2gtZTOskLcDV+1B9Nzn1zTyNtlo6lNICRmmK
ZRVu2BmCc2G+fmzynYlNTnSa7C0Cuel6FYpxCBlOuk3OF2tzAmLAuDyOH3Z1Yjzk
a0aHuoCdIRKv7BrZCdALt03JeUmXKPdOmIlkVGFl8yw=
`protect rights_digest_method = "sha256"
`protect end_toolblock="Jn9CQpRhJt4rnzZPRk+dOpzAubz7omckX1MrFd4p81o="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 15200 )
`protect data_block
gD6l00tciPUa6pDNTk/+t0OO0nC/UTtBwLB41d4inuAUA3i/ALrNyoJVcBnAmEQW
ptbcNp5fxEUJjnOxnedyZEuEBxWRieZFQnkRdF269oNzUphiVxv79PGfwjY8FR65
+THWBmy//q/5wJVPY0/teghTU4kP786wXR2et3JhqKy2aW1GO72bf7VuTpTH1E02
tkQOjCi8OubbHdEXSNe+6+wzWSXDMrfDyMaRRMufm5Ju5zKGOhtmpHcZXklnNHSz
/HM74903+OddD7wzsTtdRTrRm1mCox287Y7x64PykHuKkPqt1fYRV8Z2a4qrVa+T
/lR5ULaHj9MYL+Ve5wBk/gozeSG8n5KgH9K6YTitb2ovIUh+XyVsDUyjc1r+WPTA
67+m/uQCIIPmEc6vAq88DgkOwMGjpRZftzSF/xn0El96/MhPqpoccBEXvDSQoQyD
hYlcffboqhuJB49gT/0WWs+kcwoDwybnev7DhLQInDS/9GxSQSORI3aSkVIIaTCx
k3tpFuwoU3UZcmdxH0Bz63UNVjiKGxSJHjlnMN3SElc0Dcee8p1RsctaFS1MvkYM
z6eb85SyonB6FuqJ5tDmAkabIMlsVYL8CoChMYMwWBe+QhZ8scKygw8Z91gs/CyD
5bMbCVWTA85+3WMCmwPg2Qu1r+ixovkwTIEcCfW71N/545OySoh497mAosQWLeEF
1kKQ4RyUawQnmoRMY1GiimftCDLKg2runX9YFYBU4yx/sdrNgG/Jx9U4KFJl4VSl
Ffv+8BSWc+5NCUd0bQw+TVXPNpLS0pXVKt4JTHrDSpywiu5/iyt+j/RChRscR+iJ
4sg7jd7x56hbXJ74ng13bAnEfqIFsZU/WApr3OjPv7+PEd6jH9NsnXpTG85XhRh/
C+4+073s9XMO9Cw9GQ0MQ1bZhKoD88YR5d7Pl441MqyCgsjIyA271X7EwrZbRFTJ
pEJfEftI8uk8lGuNM/VfO5QeDtj3oDVKpSN4CM11+yCsXyJciZKI4/oRblEOsQ5j
/S2CH8SHRuw3WxXCCDC5HD/u6aYcrvGhQV+RXV/6Na1wNW3UbLp8CCgLHN9KMAiK
8li16qrLnDsT2QFULI+KNesSDEGz3+mvEn2YZmC1t92zXREICtoCdsI/8IGYETl3
LG67q80WfUh7HVjz89QWs1Js38YVeXZ/piVQkuTfpJNWF9qR7iZBv5xkWu6r6q6u
AZzK1xBgcRZrtYlvs5LqPOyaqmnLa0VjnInSeyIYThVKoz/kCd8MXu5XWq0Mh+Ug
LESBIVVRuV3JMWYklUdaua0h616tUShVW+4wstV2h9aBg5jLBDuE2FONHk0md9EM
GvqQaoHOL/dkJlt3fefq1ibIovcA640BqNPFmbMjK4QlYGk6bP4RsuDhYiNQGuou
aEFwczdIoF/eI8IRAMD9bqe1mZG/2hxXDznlrV2QvmX/cvhX4A445ES9e5gyqNxK
H6CIII8FyhIcXllBz541rSTRAYL4v1geFxcUvoG0APZznt2vA9k0KL/u4AS4H9bT
yMLXk0a159IH01w4jn3WVOu3YXZAIHnvBdeFsdVB8ummpQJNspVQwWzDPUh78MfO
Rok/TqlUeReAb1ZKj4EhGX5rKx52jxdN+1W1iEBvx2H0swcXUrzjzdwKP3+eVNTj
63dg6gpsdRe8XYpx3PgrBXpSmVJxMX3FRZAndABzcvRxpi9luvK4tepZ2CjrRajO
YQCC2zqHycdhLnViyB4Vog+hSOl31E/9StMkTD6tUGkEUF9vgBLq/rHopiQcRp5N
qcCz1KysxNJ85OIKLO9K15IwP3vtEDmYrUYtCxVx1BN+XEAxdGEfA7+Ftd/U1C5L
aaH9XFhUdYz11dtftklswy5y852dwWfdjwz34v0v5GKMN0ZK1bUJGYUT02lMGow2
k805g3UyJ2hni4mzVwgcaR2xk5Co+O/iJTGOGzq6TctIVmwDJQFw3/otgL1F3Kwd
3HOCMFTwMslVzwv/U95YyDjQ+8lbOoVrLBYshreD18kG17lm91Quo9dR7W5891lj
wWuM5bHApA8tCGWyjpkit5cVwzh4LxvQKDiF3b/tA82pVxlZRSejBkQbZdsXlU/8
W7tF2/RUTZBh3PA+b81lM7hQTLHi/GotMsM/2ZHvkct8baoRmBWjJ7aP1Q8Zfeae
4qfpoLxv94ECYu7x92HuubazNuWSTAfA8R+vLiYa+euN98z5Jf/qpj0gIJW9qOsF
hO+bXR4B6d6U0I0EF0g9h8xw/rhc5U3FkOelTu52VI7lISWnqU+ANkD2dxphhrvt
DXWz4rAfJrIdBGucOOt4tQJlLL1hVYADNRPh71j7UfDys3HXTWStegx3CHYUh+FN
l5ZskEoACGelr6a+rOQW3ME7i4uRZL8I/7Ffftu6RLtNiVCIYggs3RUN1VSLyDQi
vp8JR9Y+dWxtsKnnyeicm74cgXe7mz6/sQk83pjUSt+XLbJNX/NDnCDDzaV2lIZO
z86KRq9JwwQ/vaXLTRcG/h6TsKLmzEmp23RmKjuO+mRdbsekjFa2PLUHIVr7hfUS
eNCFVnpL3ORaLWRJ0HEEal41RvyH8KmDehMV0x0p2EKtgxK7FyOiqYcnpEt7rBFi
AGZrAxp7ZvYNC8FxvbCilS6Sh50zJWjKrPo5SMR/w5/SDLCrBcnOmJsUIiCFBShT
sIxMmQIkPLF61SkQwqxxfoMhk9M3EHOuG7f9pgy/PVvkPP7R5q721uvKLrbHxjNT
UpHI+18d8iVh7lT8sdJ0f3OJ59yPiausBEDV72bTFDs2pt1frzGyMwES4VczhmB5
s5l/Mz63+rC/Zn4skxWf2aXz5UA3T/iHvExuLqW+OkaGkHMUrerEoI0KFGA3mtwx
axTkkn7UoB/UtNRMSaGAhI5D55dHbdVaUMKU9ns5zsgPcchZImHE4I46lkwAU9cf
oBb4aPQ/mX7CHXVAP2esCOi2UBUVXFfaFOr+AjpcVkj2G50N5DGEuV1qoMVYr1nS
joz2Ph46TZmiWNbOU8YOcwwdYvEPuEY1qYDz+JYjmbETHvH5Pc+UZkq7R+tlU+Vj
gcoCI1/ZqD3PPAHRcJ1o/iW5W7wx4ngSn46BS3rce1LCdZ8lEQLUneO1i4YUY5wR
FOMCFiaGlN/S9w1abKhxnPNa0hiGCiD+vhYZpRzrSSz49HjQRnpAfcALf91OeDDh
35oei3xYkTE/FWTm/PyFp9cVE9k2QkFJlgSeUqBQgN1eXBEQr4u/0uqsN1yJ4tpW
zKzcovhEXmSSMoZtAXqiwTxXJ0O0Dp7Ck4Y6v8vEq1G7LWtE3TEyO4fDZ0qbyBGk
dpvk1qbvShXSegEDDUyQZkgbE0yLDRzgstdYwScTZhHJo+RdJZayYUrz/rc0YUT8
wE3ygnLaQfgumZGld9yhtK7ZN1ySxSUmKgkkHnsLKJKSLDZ47TPBdmi3h2CrYRKR
z6BjVUT/NLKJIC3xIUf7XY7/3NJ+FwsQqUWTdkv+Zz7anS6y/tp0hQ0833nNTtCZ
kvKKSuzLqXk2TkpYCVPyANi9XeSLIGwlPYnisl1/Gj5iAXd9AqlYnsu/gsRhpAtb
Hnx003nGkAxr6/kJoOP9aqXB4nu+WTFi0PamxDS9AcMCfhlgjLpT3kNQt+GZuFpV
6wZnOT0yPeXrsKtMR1VjWUMR6VseyJYZgELPiVejBP0akjP7f6jtgIvlUZ1uDOHl
mUzTtcHHXQeWqPpsV2M5MNCgN4ejqqHJJH6RhJUEVzf3x+HCTGAgxf9QlL0/m2D2
1qZVKs7jUxsO4L4NMuiDmshUD5AC1vuG8sLxu7pzRa66klNr+kKBGgEqelzQlVZV
Tj/mi4QZbWE/2Ba0Kq69rIDG64tgKrlVNwzrEygQTGrhOnO7wpkcSFyCGXUHHHRU
UC7wmBk0dtdpjxd4QfLo1Ea68BfLgSgisiOFgp3yOTsK4Dh2H/HiYOtXUI6BjeVW
ZpBka/Yx+1j/mXoSiwqlCfFeTn8IZsRrnQhOKzjC4qKqCvO/ylWNAWwU30KHmk0f
LUGngnym0zMI9JLM0unlki9p79BqDPa06FhaLIgMrBO9EDdUz8WbmP1yuVGow6zh
drXTpRcFLln6bWEQCUXd1E3C7rDhjMjwjAdGfC4MCcRb1g7PTvfHs8gZG3dl/Kez
3tYdP/+ptQ1uHz+P8bbV9xkKP54ZjDD4lBphStDR3wmeycI30D7MEng9H2zbMyA4
lkuXb3OQkQOdViztXsNy6iRXawaZ+oYdczZPtoyXnM93PKFxds4oFEBRRFkmvaio
aprpwegSxXtkMQruBfSuPyHlVBWFDUulq8lqeW2qppby1ag1LHTN2OZ++IoR/0mk
rsOKS0gdy64exQpFgeNLRn/GqomGLZb2ILyqaRSBn3PsT7Yr7Pv+RxBwoS3q8FXC
JTAiHeuKs1py/2gUmYRq4QydYGhESbAU/o6sGzks0qe4a6ZrP1UBjXC2lg0i8CIV
188oCkVMv4yItypjPk8i6Vzg5KRa39wl3ZolDRs9Invd+nSKEOh9liT5dQhthlez
9uCVHKFaK2nAwYj2CI6IANwtTaF9MvmFA0PgBqC5peC+v3KE+AzKFU7mdTAd368J
EeFuIjC2bR37lRww1xK6oyxNIA1x91CuDwU6r+R+a1GXjV5ftlcdA1DBeAzn4g4C
+adnSBEZBNq07cn1WRsD0YK2xAchwhicEqEIlz8kkAtA2hTt0EcdxLDRifrebh4F
VrBdIIqoPy45Vtzo2ULg7bzgY7yYfEdT8Qm+116peovJKavkaxkycxLXuh7Oxp1k
Sts3oD+RTc+TDf5EAxPplDxznvLmZBlV0syPMuEIBNmM2hHtNuizk5IDsKNY9Opc
vDAPr8hsZCx7TTjFmzNGSQk/gHCpDs/Vjzq+F8GKom8YJMMzUE4bzEhMe2whiAKi
7DI56Dq/gXqdh7cBE5J63Pb6yPYrqbWwb/oW/vdpo31+PS4RSeZ83weQ1+1SFS1T
qTHs9sM82hy4hd4ob3X5/gAzxTPI748ZkCXnMjuIqWqOJ0FzT/rsOZaUhJGruXkK
A1qBi8jTthryMxn+hhGnEr0fYk+8bJ0KaGmytMLeFeAptUCJixJgskxFf+eHkqWm
e8RjG4U5ULtznGuqMFzy1SpZQWOp5Q6ntxudRHrLTXv7oZW8B3iiJmodaVpV2x+l
un2yKUxlZUsc4R9H0CJGn9RPnpCVGEuLT7QVdtc9u5ABjV5pFsvksvewyDJY0FVL
OkAcQ8ZAyzS3mRjIxrJBP2yaX5ZKhBxkQgf2FRLlnzHzqHmLBR8F5wmNpzcuBP69
pRQlI2NQgHhyNgf7X6dEiffxFWPEvqjlEu2b1T8jYC7VbklqX4D1XTwOGNvhJDnJ
yaUK9D9lL3OCD13Uue4wKdMw+DRHn48EB8G08lx9OGH/idelbMsEteUMmSBrIGMg
1AFYep+/dMISucxXDqwXwEY7ahyoK1gpuZ355y9Ar3C9/VhOyi6ExDNCi84DV/bV
77PHimdEErvsUA+boxfiVxoWNrHBlozEDD4/8t+1BUIZBNW4o1Nl/ZsoiV/zMx1e
XRlGUia3hNIuuXV3LJgyxgwLN4Bc2toOOD7JEet7LJwsfIDCS09Lg08mVeIp6usB
lZI8/2wjdLr2WkPauey3culb/LJBZg7FUJwYxpPp2Q3kG38evJK8NegaxVRFUmCx
pNVb7J6gGLfhD0ie1WuveFBSYpv6cTYIFWZc/VbQgdwvA7w9DSiGT5kwDzH3Oo5H
0WOOQrBpKIkAbxK8CVxXzSbsJkJlPm8B0Qf0T9GTY7VCSqdZpEs33R2COn4T+Nlb
2RgkbVvyCAQlDvFCsATRuM8i+j+bqm2uRkwj5wZNnhUAZY1rnFGgKQUjdLKIc2De
mvdsY+FNJDnpOoW/Yt3+1NpbQesTDQN/vYfJo8KsfVmIu18ZCffq3FH8rmHyz3HY
5DDpdRj4hj/g2tiKS4/jevCNbjJfloWljKyeGAhXN592iO1duXl3/pSmdvT6c0qk
C8cOTFwHOaMFzNVdII3D3Gd1woCtQUymuDOEO1zrn1I+KJ9oURLcHnidufZB/IYu
QIQu+vAktKtiuCYETllN0JVT1odH9T5vWWAqZ0o82DYRF2QmnPtVOIdFM2ob4I44
nEZA2utiJofkIAVex8U0pPI5IA8jlk5g+/69DM7k2JCiuew1mceWpWtcEltmwaN3
OVqPXXHqybYH6jKE8CXBzeoss1Gtp6ac5V0/cr7aCtyK7yzR5fbutv16Wd4qU8iU
gVG5P35+YmvrAexYDDZ5hMSWuejoBj9H5C3eIdSGlRz71BhH4HgpZ/vxoxbZd5Qe
Ua9mnWxDlHTAontfy/Vf6U6j8ip2ivNKAc3dWKUpPe7OHGwzvRAHAhx5qnSCuveC
cdRSthCfVMnaxYXl87/ukWhdFo08jbvhWUHf/vmKkV0jJXhRYY4AA8is4EHpuC+q
wrlfJ9fGOI2gIEiQM0Ac2xornetieev5tmSQLKj6Wp1FZE8wQhrtU91sHg+sJELw
AYzu0A9PN1qPHFr8zXchLxkLO3QL5iKL03xXeaNw1fZ5cTJBP6cT793LiSnHAckH
V9k1QDO8Vrq6FfWPFp0F/40huboMvJ+scLjhdV4tbtQuADXExSq3EdMO3JgMperY
6gMKkgSsdsNHt3QbsoRIGa6I60b6c3dIpyakB6wmCwBX0AoBmpG8sSEWewrJnCgm
S6x17f0AzhoJlLuiCFRuC3AP+KWYFkGN4DEaeZ95gCjVMV+tauK9qV8pg4K2vxhs
JMxCLAP415ijHyRMxCOQ+PZtjxYrUK6M25ITqo+DI1Fi4fpW86SDHvqejoZN1bMW
UuiP+HwzLvBRKSovRFz0d1jYkZyBhQVHGitAWIjCFoha2o/Bi0hED1Hp3miq1gbm
WWI+NJL94Ied5tbMwRmzLuGYILKACFaE5lZXbF0n5Y9FBs/l1Tf0mg7F5wwzT+Zn
chcwnq7fsyWXhgUfg7fBl4EBaEPZKIUso9OyQXbePqMIqYY35D5utLMXXtH/3lpS
/loxn4TpQvDmeArjQtmaRENAE/BxGG8JaUt5jmS8XWADjUZmErf1ioxAjDg9XA/M
fjG1G+AzgPRJ0RMCVNGvUMr1c9KvLz+GjcwYGsBc1emcnFF/BhtoDaO9n1cwiXGn
toMTxY5gsmwz9ZYPwOAt7lwmiH9XZp11yeCz88kLzXfzDclUxJzsoBz8hD0Zny4D
Let+jg2tKI+g2XX9U+7QM1MH86Ofg3e8SuLZh6GQ0yB0Wwg1tJPhxGbXYXnyO7mv
abP5zICWbnnjAr79LrYl0hZFNp97LvpsB2ooxd36vBcM21H8X7kfeUy0sKLwZTsA
FYw72crFAM3XLSBDTfKVmBzIF5BpwjZtAHxySCEKubEHmhua4xye/7boTikrit3M
w7VzQsJxH1+5OLPRfWOjODSu4G8IMeOnnJY0zHilL+tVReTVuXUI2OWc+3+oFQQH
rSfyZj2bBXj/Lm+WMYSYJhrhdbsduIVVd+F9KuAXgJahFo1Fm0QSTgVXDN1ag+i3
dUMwvnSvwuVkpbFRbuh5OLZJ0E5Csex58UbgLXaKj70/BWnSryE3JraSikU2PSo2
3s1g+FRAs8dJKjR5MQmKYZFKXmt5riIoIiSbEIXwz7jNKakyUwOr+DSFCRccIc9V
GqTwmLXivpg/tcdOtJSZsVRt+5scDWiha9RTPNWmicaNwkIrWWeut3JEx64qj2uz
N/shh/pNlx1JFeM8WOuBNZzduQVSYi9dqb4C8kHubSX2kHcmACdUbMuesBc34I2B
BTORBjdXauUKDapbeV0qim/OZgJSljv0fHJlpDV6ABjPIwVXqPMXo1QLrwhahKGx
vg4YFc7O70jSdT2FkZTl2eqHPOmOJ3vSxvfzH+gcEHE8Y6F3IwEbVkyHncWulPNu
lf+8oXc1wN6oe4vyGFOKSj2HNr95tItyqlq0/IdM6SDZdw+GYaerfbY3hKwePsqD
mLDuqjL4uTw9/dDEIn6emWpXeQpeiJT6IjRj9ZP+Xn6j8XEIA2xvIGmTL+NdHhHP
XLdgf5NjCsBhtdAQgAv8T33g/sWh3BFPZsTSLwjAUR0+sp5+X4MsvWJL3OSGREoW
2HlZClCX6Q5SWrcS08SXstdYY3CIFT0X57gxJi+gKn7UPJ1MzM1219WYNUQrS77l
G3Ls32uj9gqZXVF2xwPN/lqPac1Imxf/TzFGQW6UuG5FgkbeVggYmqjO4hYTNpD1
stSwSnelZxBVJ1yXB8+231iqoq7KeUfEjfAlTwoAqfzsmYXeK2os+/hp+Gzx6UBW
b1CPlAkF5mA9M+umYZyzoLuYvtzMZIYpZmFAuvuvSj4RHkfBb+O5HdI7o+AYuqB1
wMq9Bdr+IC1C82ikL9n2P+rONO8YxLdNwchuQJ2SCyfrPa6Lfc3jBYG9lC+hPQj5
3p15Wb85csG2rqdoXN8lwXfBnYMXZo9qNhQzafryNmbwdv8sYsGP9QR2IxQ7tsFb
7mYwRCBnMNd8zIiFanvRTTTfxdNM6/VxyXQvV6I0T8twWchpMO45fFUL6o9JQSOW
DQv4TBhUCoBavLL6F9zzhObWQBbu9HJclJP+2EAMiQeGUnGgAgRlK1aqTtlZz3Ca
ECJUzDNBGIG9GKPabDsd3Uwythv+5yqEneB4U72BAHoflVV5TLwYvQc9duSqCEC1
+RTGj1Ml7eagFnERFzquaKY2U5sQ5UCJWUKQcwhZkA50LA+p066Jaa7M5p3nld6L
xcHXmDmf6MkmZCHqL/k0xG/U8YokA32cq+9I0dYer/W8VQmCUcouvbXI/VwbQkhX
m0tbopmX1gV6jeoU5iVLeP1SAOGpPjrXwIUBREQ9gZoGTbk/5upG4lvxbU6nCIe+
KUzIWl9//h58pRhlCrTomQxBN5mlYP6aEuTn10wGmJj3/aZ7NI+hu9PEobpeIiTK
kTkc26biD1ZynOwlpZ1EmfXNmqGPG+iNenlZS6fNGA5xGAy+aqVzDPC4WlawiHFv
1UxYBVbf9loxGTwq4xyXw8giiFxw2vwRPHAJQ03/p1tEshRHiAK/awgJaTqIZyXV
M8SqF/TqMAcbvj3GiEshVZH1YHTHhuHugYF1FSliPAIG/2zyl90wSKjynpQGPBx/
sCcgxz8ZeruspDsPXpzgieTKebIjXuRZqI+CCJbwAd6BwVvoJ8X3IZHC/7dFL/ki
FCZEwNYmu7EbD5J9QSXU/4vqmZXNiDRNvmJYzd4VUw8R4Q0hBvZUpg8ovQlbZ24G
s3gA0DBfcJvXbh7EK///sGPgXtmGo1qUHwgYU4S0xrVcYAE7vgsOcJaDVfwRkYsp
Pq6JyXmWWdpRTe2NGvu0dNkLrfqwUk/w0y7MjZX6A6fqw9sFkM4jEa3/YEf4EGD1
7itGzyxuq7mpf33MJdU06KzT1Svn2iYXjJfNnwfLcouCoNV9m0vi3sm5/Hzt6czs
Uf2RtLMuyZbZuqDKgvcDJ9mLNcCSpEgacLv78m/56PwxGmfBuj9C5gNQbj9ujL35
fYfL2EmNduJ7We1OYNcVmI4OZT/njWdmOFOOXVg+/t+OXKli+Rq2lCYbg5bSHWGf
S0hJUUTjB67Xc+a2GayOXt8SzaRzEqyDX9IEcTHqhzBaCMw9uCpL3B3QEcN++JOd
NUxxHX3z5fvDkKwlDQROHBGgA60Rcn+UfyUagonTLKZkP7i6GkQTQQEEDyogH5rp
p8Q7O1Q1xfGyClxsIay/1CzLACd8soOPPY7nXdAHbMbc/hTFYUthTE3ad5IfW32e
oBL8mvMjJnD2DVUPdgmMak0snG4IptMBw2aduQoS5+4+pkS3Pk7VdK/gQGB+WPHW
fh8J0D4gT7ESDiy2BuPAAgPErg9KgvwgIy5BUNCs+K+vLYFryIdRy0x/sczpEeCq
Qaladb5+47KM0zdD9duvmSJ/RuAVfU7Mp5lBxia1AHNGFkF+QbZ00fggJquuzCjW
5zTeHLr9ove5wUWxuXlj7nIAiBwZblBC88oSqiokcUbk6pZIiMB6ZJ6s64LB0bzw
BfV1kjoauN51en29lqco5vm1VWOp5+3w88ewKqbBCouZNwx1WpkxW8ZienjuFxYc
iSX6k+QWVTjKwA4wW7vvP6YwLEIspKQt0OhEu9BtruhO2xANw3JJDXXEJ816yF/D
+s6ISepCr00l6NZitWczoMnUddcrB4HpBOPofqgIi3fbTQ5KL6PqVYV4nsIpqwNT
u8X5fEMgnl0HvZuYs9koJb6suqFw5xypvEkQiB2duj/PVBmN9hs5Uza+5NH8+si6
vXjktG63ITpbtj2a4ItT40b2z7Jg/SP7xSmwOKNN/Tyiod6AEA3xlwmoM1V8+Ttd
TrjPy4aQF5t6n/WwACppXJWcLSRE9xQaCp/3lXPGTdUgYJ15qf05/RNiWkGTfp4n
dHfCHbGuEZEBUEjnGeRjgRFtdW+DJ5WgHotshX8iafY9XC7hRVCGEIefblJDtpEd
Hf3LdPZnrk3SRSk7lPJBlKpHH5rC/lXaMrnieo/kBFCwgkT1z+qyV0BBSCjtiXE3
tps0hG0fdjPhet9JDwRWZNXO+KXsgxxiiEkM0V/LhtYgM5JwmQefesaVRIUjn3Uw
QOHEhuNOrZPqekGy+/lMCLVAB+J4fcbcfUOc1X7BtPGEqnr39Mio9ZjXyCviVcjx
GU+AhBF0zcW2OHv9XpdXY+xh6uiXWgQYMCtMFCVuDMztkz+Ujnv7YCmV5767r5Ny
UGJSYShpNA6YbhpBShm/FTTlCetNG+4orL5DhbXjSdxSINur0GdAcN17pBs0uzN8
zBimHKGy7l72UrQ5N3/dlfggAEL2/hRNzfvoDaW3yC5JF1zShrdE6Xn2pdh5sCte
GEjbnSW7nvzTbh4/ydQV8OdQe5ECLZdnyMB+KL9zTq2Rd1WdyQ363jJmSxeKgZJI
FF5B6KVnYmsgWxQKAXDJhiZjr9u3IzAkT/hhhTCSwxNjTgYF+EnpKZBegEpRvfkP
sbaHZ0bOWbN+WVKKfJcWWYjs5or6RwV9Dj4bkMGrPCbGv8mGgs4wM1ZTOv6ay3dK
80/bipkyKZec9sA0HMiSmM/4M5XAAQFlH22Fikq+hrBRI3ZgULraOentehW8Oy57
Zh8TYQic8Ia5q4v0HylGWYWzbIXIOylVhICWZHMpR7V1smOws9lpcuINfIw5dEMk
yXnEoY0GAnZ4BUJO9AxoDb5dkf3IbErXGnbNfF7RGVnRsmw7IanIyN9AnQiu6on6
eU7xNJlCIQaIFJxs/eK/QjDy+CtGuPi/0w1Yy3e86A6Nyqho/IugEBowGJM+9ijU
2RQP+wV2Ni8w5//E86tFQazK57e1m/aBE0FyAOpDN95BFHFTQhXe8A9eOodruPBx
chiIHLJOhMXjvCwzMMYKtSlOSicIfOYtMSS6mHCkqx4aIgK89QojdpAAk3ppc7ie
dydSemLr5D8OaKVZdh+Via5V1rN9pngJqst8B9B/JxX4/MsdxGaAeWQU/4N5tmDR
+dXrzkGn79IJVyDyrOzzl/rtT7vYII4Z0Nn/li/IHJs8rjFMEiu0SfOye3aQmSvg
MaOI8kib1sUfrOrkmVbyiTFmUUiLrMjkFUUmqUH2cxtbq4Hvb+YZo4/04zRx7sqI
XxEEScgyH4L9CQ0YoJ+Gxd9PKJ7KLxUtfbzhN2F07v4OM6E6veHnCLX/VOX8Zc5D
4EV7Rqi9ASimhXtMm0MvVxON8JYFS6gqTlOEWc4kEECLL324BE8Ekn922RtcxfXf
lnT6lqhSV6d1jBsTNMJrPoOkhy2eQcn9Oprh+zUwzVMieahp1j2SlrQ7ZDj5ooZM
H/BMQrwrbtYpC+MIGalxtAnMsT8vln0olGspjKgyszhKX154On3jlJc95+AMnMX0
++PmP5ZCmW8QcXPRFVwUGWfbyD2dpCtCcXk0EopLwc8zioFsLxjub4eH/edre9zl
qLOzSYH+DTBtBDxGbYQQm6ug3hHRSSs65mahmzaq4zHMiWD03IwydVIWQsuXTi5I
gbwJg4CPVBjkkuFLHdfkZuj2pwpKX7kwdJSBBfU0vEOry0MqZE0lJ18TKP3kCY42
TMUf+A+JSVVPhRyEpyPQvGGM1AaaQQ+581YIVj9uPhNUdXKopSN9OfNQuqe7Fqqp
NSi1rN1FVWKtt2qJ244dyaKe+J9kZIACj5wy7rfjTZzHuTI2IEgJii0Uhy3+jMHT
Aofw6gMunc6rFwlVVmNeXzLLBmUwl0BjNsRTMYtFOFM2s+0xlPtdufqgoaKTsYun
hwBVS3h+JDQdTA2qrNp0jBd+imsGtgxfJnw8h3KK2r5aLWkUd0jHbXcxZJAhAlRV
tdYmW0lDVB7+76UA5m8sjZpFow9jwvvkidFvQJ7dpw0eCxS0I5NJJG6u+4LV+ZQy
+OLYJt2y1QjgAmf0sdXBsyw8RIeHRs7krmhhjkvfg3VvM44H3ov1vs9PH9Lch9Ll
GPLyoUpiZwYTr+1tL44EJzAE5K+svDNtL8bkkslRV7T70i48oSlMubYFOoAY39QG
yob8ms+r7FSlGrm3Vysq32shxCDj2BG7KlV5CazqQn+3W40mLmDiOnDU5Vxrc1lZ
g7weL9z6u1qReAB0bhpTBCXkdIkmraCld8TN6aVOBwu06Vb7MsUonD5RpSwq4dt2
fYXQoM94iJKizBLTLVCzA72PhrzwKN8HZnwdTn+Dts3+69ML/hIphaxdgmKTsEM8
qDuEVvroQZO6u20Tg7G6MnbBUBYlaX1DKJXwBhrldSolb6+9OggmTSATDYHKyTS5
nBGzxxkY64ZjyCKZTHeHFnwvPRzLg3accpp2gqtGMhKDkIdaXLeJRaA525CwGAdM
tOND2R+QhAW011/J+3YYO5MvseAeQoQaMs2GZvDGrckf2XbBOqFygFNAhwNkShcn
FumPSThNcYHcTjebVOmGTAjfOReRaeJDixU6kcj84/oI8M7ll0LtbDcPgXGhxVCT
+QbAP/CSvbq2JCD6SE6DwIpC6INj5J3q1dnqlbJdOcnZkgOoz9tsxkes9+CQulaM
Dm3SRLuUaJqTSCy+sx/PfLFIKjR85Zt/0r75qcCI6tXgVxVZo6ouPXDFpTld2XF7
lRg62sNMoCngSUSqCZ3IJfOvQzgWiIT8hAlj0j31jGo77za54dDT/483keSMdj7B
6VynKIBCETHbB6PoFrcYTmUlCHKr9+Cweg7RBYiD3BMwxYfmOgRi+Ce/uYlUJvuL
W5gaxLA35ZpPj1bW7cCRVf+ZZx0hBH6c2NgaE06FhZcTskJbiZ1918WOk1t1DzS6
Kx879JuIvVcdX9b3NWYy+JZcyRwZsAFZ5uBhd5MX+SScu8rp6pi4FQY0l5SYEAWB
tfZr+MUUp0hHQCOg0jxFZ5VrUK0Gd0nS/Li4ODgGulgAZlABf4KfUX/8/cApqgGT
I8F0P1ToWf515LpiSpieBy9GkefHuA9UMiDfKSyuHtZcJmKTlmXgzOheuZP/QvyG
nUlQ6kQdhfEMKiGIsEOpSf06SHnmlecN91dLLb4UFLygyjkxVkZjFIOwyOyeE3g7
qq4h2JwEyziSpodGkXlOcc/CgAAvdk9OSY5Me2y1nPB180wf5L0ZALGVjrH50fpG
b7ATKVRmeABhxHusigCU1HC78QQWSY7g1Xmfx+OU/Uk2nuJ7pL4fdeVe82xoAtYZ
Hc/dt4jvhrRgLHTcgo066OAEWwoKnYjttzXQ/b+m+IbAT6zLkcD9DGt6J0mqTSG6
gNN1sp1iBZ2lS09AsBf4Qvxb75FO2vkdgNEQjsneieXFH8BVJno4re5gHckaKqBG
jHOoxU4Hz74MhswAYGsLQzHRD9/f/91SL+Jjh/9Wgv8YmFAGKFeUDprqluXiQKOg
5a/c0yNghGog8abVWMod60DSLXfOVxE0M05uwOKVJmUNSMKH+2xhEtxdGMvS/YIo
Gydom0FwsT473DItlXCgiEsh/EBuYopVQPvei+WhgpfuwoC9jP+NZCiu5t2JFmp4
z5jyk9vZ36KkPYmwvTOp8I83FaWPHUtIG7u8bQM0Y16t6YpQW1DW4Whq9Is/NMQp
DrRvo67PU5RA1kxM302Jn1ujQG1txwCjotDjFcFfAJud6fdiORTxiqb12tQZRTFC
a3UtbrVdlO5cl/jzeIqoKZl0jf1Rmq6F3DHvvNSMm+PEjlGGkumCoo2c/23b/N2e
g24a/XWSwNKZI+NNeoyxaNBw+QKjt++yYeWzmJM9mFUqxtHu4mvriTP/ocftJg55
8xMBYCcYwWH9tT4aqdadWEXSl6ZQHkzCq59ELmfAnF49VM7cCBgKJ6vWKhIK6ja9
wlPaY+hmFytFDVEIsOulLtJRRjJ7e7BGnn5AkTbyCiJUahgJQiCa+fUSIdeSfP0r
/ABLPd/paawOAQH5qVqKJkkHhbZ+uiHWGSM3BwudqTCvk4tdS98nDxK9J+8EDOV5
oBCXFOMALYUC+Xg3LPGa/BAAiDIEmNo4Lh2t3FIT1QnZyqJ3L3RBr2279wu+kO8K
hWrYbPYal/2sigQVjuEt1oTUa2T8LMCxeGpnD/1Ywsgl4No+oGaHsGTL7FzPGP8Q
V9n1G+n4icYxUsNoP3Yiyv1KgRff/B6uomNiKWQc3x++bAiSdooQXGFgUBwNOkJw
AgVFg5CIie2c5+yHr7AGm/W1CNvlM+PkfAHUqPHjB9MYIgSgMzD9MSXFxEQcsqYu
rLsucsRVNbcDHuE+iQpYY+LK1VhA1KlxqaG5DtPGnN7/nHXm1q04XDOHnI3UJeSl
5iteaL314RGtxVAeCO9hmAcUqEh1BNytdixpj3FwvNAZblAE01vEzR4+0jt546NL
a2j1fgf0k9osjIqycPFSWZJRCfyBkPekYIsnSf4t9JftCJCMllA/b81Wxbaz9BIU
HtmVWU9b41cFgkzqxzC99t76MgWTARyZkgIy0/w3rtIwfoju12bgFfr8kggkDgbR
DAFf6VejAwTWRbIfK5FzaHAPLVO6rRQHsYdxU98O9TwQcYPwQPU+e5I4EjXVw20q
tjOK2lrIN+lru1IuP0GZi09E4C2ZbithW9aK7CprCv+P/Z4NLGvxUVhIzNWIUjK2
3sJW1/GhkECjGv0u9VF+N41LUbm8NdWakett5kVpmXuvdAVl5RdaX3HP16EhIjgo
pa9dYy3/7SmRwIMF+YIk2BepbqQQKiaGQ3j/tWcWRTmSHIlKqTBk3+ZGHHdjakl5
+ClEqZz0aSUBo/PwSJkDOKFSjqkYKHRG5uviHNIGS29LIf4hnaVAT6o6QVQ1LiYA
aQ3gbidVLQr7n8FvND0d27Dwf9Ub8l9QrjJvqcF7Fxsi2L3XCZsO+rJUjm0zSIdQ
asN9rLXUuka5ay0h/kzQ3W/ciP+YquotsdJt1fc8XUDtwuqqIL+3cwGW/6mbQyxK
LmhwSn040uoKv3ww3cf7+bIdgXLeFSOKKiwIZBoI5fuIPttPcjneVhJu09DziNL9
reaYnDCkcUydSof3cTT/C26rf4TrTH7g3DYv1364q3sRv24KKKR7KHChrkVOppG7
e5gnXqzltcQp1iFtsw+7iNsI/6hKC3BPUdusB3QHXSuXlV2BNVXblPJKcuI4e2Xm
5GCiqqxxbG9nN8VEHBKencMxJyvT5/IhC+IbY1yCqtUBVu1424ywQ3vZPbjxqg0Q
Zvgc8vkcaE8ui+1Us9mB13kEYhAKKBejI9JWjmxDSiTT+flBFue+VA561QmylWK8
yuNF8jz+iOgVKOURzRPM2VYyue1ck6e+O5DHhVhvnlMIwO8qopfiKht9OBXWQ7Wb
l3DTNlcXdEGZPAagK1CYCWRge2dwrPGM9kgVwb/1arCWzxYnIcpIYhUwFcz8Pakl
xRPdhBF5nqLZo4LATVlj2dnTpMl+ZeVEw49d1OROliNvCyo6XDpEEq+C+a7qAAxO
plTnGBHXqAPuAaD/kttlFMZJM0NA1c3IEDaRm4ZsXJXAlQnTHea1IuG/iohfxvE+
nWTCo7pYBkg6wCWlA4xB0bqfuVz1vQRHYDCwiLXl8Hxt5SUEJLzGmR4qhTJ6YoYZ
OD49GQl9QT2gheNj+qmkMFw3kzjqqzgM6VBiWmIkJd3QbtfATWWmGzmqWvGjZoz3
z0H/CdwFciCEEIzraKVAMOqoii/Ah29C5qwojxpEa6pse20obdgtFp3A/Kor9BHx
HNc/ksFC34dyt8tzr/2QPm4VVU6kXyUpDpYqrYk9cqtUZVJZRMtQSvyOiO1QGuqK
oOUU5Aq6Mv8fo+JWVuRwM+DkqbupJNyUe+E1HpfF92L6lfNrMpB1kMIqEwN3ehau
85Lbh+qBkr5BMSDJIYg2ZabRLqfgHhsMBWXlTNSoWtJD3/DP/70SLci3CB30HXOx
uuz4Curythb00bFkxlbTY0d2ep/10upL/W5EqrnnNB97frLtnYSip/5hZhz0GSSg
JJwUrytThlB5HF0SWxewX/QrWn8tOJv3Y/xlfa47DPj4fwQHRQdVBfzT/GRakyhb
ZyTD4GLUVK4tNijK3iCg0HpfiXek6cSfJJJbiyCw8r2dK6WKLwJhoFoGwNjRS0+I
anPp5u1Cw2MQp0r4i23twLXL2w8h+LOTiGdmZgsvV619VSEH+1msfNTlH9dSe08g
JGaba+XyWALMR6uHN5LE5sc/AnLgc9BKlueYZd7imgC0F5wfiBXuWYJ5ZiAT9MbH
xTsfBL7VS5HBgSFW0CJ4RDWEP+o064muiVDo4e2UNKQdYtP4Xid/xwV7LqsT8PAa
AHu2e5FGLeK5xoU8uyix8xCDS6z7gJ5L3pMJJTc+Z3q156SOQ2agf9waxJKxVR7C
DzIZO9/RGzFzlc+qb8T62eWRCvNjudvbaQnPLsaUE1p3iddXAvRmicKmsm3Rc3UD
zjHDE9u/AcxgegWwd3rgscgk2QpeOSU7uREmKpletVyu/+mLg3FlX2nNSzjYBT+b
YogPn36V2NI8M0kdQD5bX9ibjFtq6Fikl2D1MkAmkfs6EOP8o/Jv8r1tX1MAFLJD
0bhKY8UWdKZ9Igbs7OmiKaZc2o133RKRmt0A/rm9LoZ/d5lsUtg4jUDv+4bKtNDQ
PhPI8Ca6zFjfJZZCR35dAhWCxNRsZ0E1vH72a1QrFAlC+3HEIpdZGqo3wog68m2Z
LjgBw1/YfO9CdzVwh7pUFOEUeZNggD7SJawXKKIyAPHgfTSgpGjt/OJEDoJSZP2B
rG6uE7nJK53izQNcovfaUuzWSgLx8ARtAwnfNyWRcYtOq8BuDi8LF2jiKAe38N2i
pFqP6gHHAdJ5fcvTobHqI2VLQEvk4pkbvwNeNv4c5le0Wz3Iz+U5cxBr6QleZRFP
wk07afeI4Fgu6pdOjx6YSpTRTIz6kFEkooHianFJXEVm0V42uMvNu/1dYT3tS689
6DKzMCQ34pBguy6eZcNW4pvk3S+2c0MmrovinwtnOhgVNszgfN4gwuca09Z87r2T
GtNTRrm1aPVoLcRG3rYf/WzSasIUBEoU/v+EeTi9E++5H5RjPC/cMRC4beBUaiA8
rRlmQmgy7ou3Hx2kH6wOTOmT4U69WGwmy9usvY4ssrO5x/95oPDgyNP84lwAHaPB
ObRFGsbD1G2sogRsVBGb7BURAh+ee1WxFP7fKfJAGTRGVcCmWyJ76EW1CFRQbtcN
1m5SnmQRddfC6KKoO2al/43yDbJclaku09pXMKAkJcbUzrUOoAtDGFxTFncSJbYh
++2fTAF77pA9ezeVIM4yGwmGHiin7bVBQFHrzDVxpO1rqANvJDyNG/7fdq4H0wEF
vIIVuNyM8V6xu6CiUShUuPHnAy1TiKFkgrQL4Y9B6r5AtlfxKSMCaGgMlNBhswTx
DbhAVIyRUW5h5h6WzY2l5cwCCAZDwrFd3alr6d0fNo6jAhcYwL64CEMnyY89YzDZ
MoTzzkXQF8ldS3PiKm3kv1u50SzLdFDeR9TR2SAUCz5wZ9UU7BODU/0KHVKFG8Ws
LEgYM3M7hAyXRRShpxBrJQy/yHUbVMRBbeefVBeIqkaNZNkf7wSN8didRG5xpCZE
RJe3xQqXQgyImRluoyrT2tFCR9T3i9ZTqwLKRTQBysnrJGLPTjjOL0bJeQSqey2l
AwlXgPV9C+PUzNB99Nc4gBMGF3OvPDsMm9hFxWkF1uHjnsPLlpIoZ5I6OZIqKPgF
oykzOXFZD1wL7NpRsIuUZLZwPwyNc6gclxAqCdZRZ7r2u8bb5zKBu6iogvFah+6R
uRMwhHUyc1WR/L+JnKX+wBU8MTxZE7TJNEwId6jajC3+DnkSY93fH4CUFBV0+cww
E/2yTxm4+Kgwnop31QzLNpeb2Khuk7Ks1xY9iBmjRLmPOn4CTC84dZywvRZQxe/f
T/IxjcuG3mNFdKlOCI0D2Q934Z9/BuK3MXwZuumPr0Xv9jkywvY9xYpKGp+FOZ8A
yPfmPXZkaFByLZESjhrReNuI3BrvcpsS2yJHecLat+D2BEMoJDc+ltCuxfdLPBuj
T1A491Gsf/i//bGXI8/a9v57EUawMMkGJeHJWTmuhS/0L7bmFMZlVOd7UgRRMVtu
T06LB2w0mGtFZho3zhhzAYlTXmHnmfBgN3oqxvHgh1md5WD6MdfOEf/ormkchOqy
EJ9vQ7X58hjc6xg/9WVunjEcxpqEptlGwQQCIRqclAhethVsdJPcrtUqetTwvzZf
WAomhi7beOHsXIt7MjMFdfeZO9zMCataBMd0oclI6X4ZJ7oAOzSC4V72nY/69Mqs
jJuOo3zjLzqiB62SKxdHodzLPhcGFRhOg/0f37kB9TXP5cFBYayLjPK6xr/Dk/CZ
v5Dqd8p5LJVfoPjh329KX1/porlVLFPukmOMPeksNh1DVHMq97Biq5muhJFmU/X4
w+aGB9aKYgboq4eDpkcxvuj10oairDQbuu4Mt2RLfVuhapVP76JaGl2X2RlT2Z86
x7ax7Gul+AIZBaNnDnLazknIoqDLsJMxBtEsz9kpc+IfV4vTILMZf+8QU9GGkz/I
awSzjApZPOobcpE0KTEPeabqsaxk/fwLB9DebeWrokY/8NbdZeeBenH4eedUsSx0
QCBn5NSpjhl+z26j9Z5Ika4B0eLRUb0BwvpzR0nU1DNeDSRMHquUhwH0NbPiNXw/
yCJWg01g9fB27YtGlRxKTLhn/6A5KZhbt6108yh8l6TLVXgMiZMeNfXd6sWnGpYZ
/d+Lg+lVkDphzNbfcVc2D2jwDkg4nckxgQxyIYG+x4veYEL3deDNbcR0qf3A1R9W
NydrBxUwzRia27+vWwhUkHuZtF9NTDgxHHsWR2+CjZb2O4s438ZfKuOXYgb/v3Ce
xAt/kAUG1DS7psJVdv+q1G7TMXBgaWb7Fp8zNEuTIz5r55KWBVsLuisbnzZETiQj
n3weBxDFiNtycgTxpWROU4J1NxtiiHyMmP7e9r6B6TMRUj6HGLAKtcQHdzq5Q0+8
43ciry4Uk/kZnGFC8skGp/KVCARnHj78Lyhw4l3CL3cpe48e6W1JTu/bp0lFBtCw
brDM/KNuHMuhcqGIZpGqXAmJD09/L64So3vN4llRJkDXkSPbChUuKXh++JLsy1Fq
yFVwKMeohhg9STAbyxjFWDgmUM+SBBtiRJ3wHBAFBK76QaPbc+N0kh20EJ0QF5cA
akipsK1htEPtLwiegDJcUT7PqloehxPy+1PZ27z6OirfD7FRITyz2RqivVVTgTYV
8NOM2e70zCXqfsqlw31WXgayq7jx6o0NZzPeVw7X5W9r6Gundow6EZh+WqwKM+bM
R4dP3KoCpYmOzkNiJ8YJlJaH4S1TJWH53XZX3BuPAfdt+O6/LdKw+pGzLzSbj9cY
XTcHBQ0rQ/aieJuh1MQeXMC3HI692vhjFKl6gr0Zh/TSXpiPSJFTqpXBqDJtIBfS
M836yZuO8CaDqTb3nP4JyNmvx4EtNUk1dcDoO43nLm56jAHzZGwjgGePjw1jYi8J
ngBQoFl74QHQ/Oo10on9fNss8J+UcmHhYqnXgKlm3JkgV4ODNzbCO6uZYNzmUaNF
88jASu/KH18miU5QQtiEbZKijV1w5LYNIMR+p1XAidKcaox7IFJvyVW+GcCOZTVk
XRKQXbzR7KnY9kONPvfksq/3nyGRz7enGXQ6S6nLJtTUuSEqZ99vwma6vq97BrAL
xyW85Gn4B3LL8udy2DdPg3QvqU5WHy/aApW+o0aR/z2dLQwiRQPduzB9XKYEC2bD
cpSFlqRzG9BPX20R/PwrsGcZnML35IFDFaZ2KUayS5Q=
`protect end_protected